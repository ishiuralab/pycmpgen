module compressor2_1_64_12_shiftregister(input clk, input in_data0, input in_data1, input in_data2, input in_data3, input in_data4, input in_data5, input in_data6, input in_data7, input in_data8, input in_data9, input in_data10, input in_data11, input in_data12, input in_data13, input in_data14, input in_data15, input in_data16, input in_data17, input in_data18, input in_data19, input in_data20, input in_data21, input in_data22, input in_data23, input in_data24, input in_data25, input in_data26, input in_data27, input in_data28, input in_data29, input in_data30, input in_data31, input in_data32, input in_data33, input in_data34, input in_data35, input in_data36, input in_data37, input in_data38, input in_data39, input in_data40, input in_data41, input in_data42, input in_data43, input in_data44, input in_data45, input in_data46, input in_data47, input in_data48, input in_data49, input in_data50, input in_data51, input in_data52, input in_data53, input in_data54, input in_data55, input in_data56, input in_data57, input in_data58, input in_data59, input in_data60, input in_data61, input in_data62, input in_data63, output [17:0]dst);
    reg [11:0] src0;
    reg [11:0] src1;
    reg [11:0] src2;
    reg [11:0] src3;
    reg [11:0] src4;
    reg [11:0] src5;
    reg [11:0] src6;
    reg [11:0] src7;
    reg [11:0] src8;
    reg [11:0] src9;
    reg [11:0] src10;
    reg [11:0] src11;
    reg [11:0] src12;
    reg [11:0] src13;
    reg [11:0] src14;
    reg [11:0] src15;
    reg [11:0] src16;
    reg [11:0] src17;
    reg [11:0] src18;
    reg [11:0] src19;
    reg [11:0] src20;
    reg [11:0] src21;
    reg [11:0] src22;
    reg [11:0] src23;
    reg [11:0] src24;
    reg [11:0] src25;
    reg [11:0] src26;
    reg [11:0] src27;
    reg [11:0] src28;
    reg [11:0] src29;
    reg [11:0] src30;
    reg [11:0] src31;
    reg [11:0] src32;
    reg [11:0] src33;
    reg [11:0] src34;
    reg [11:0] src35;
    reg [11:0] src36;
    reg [11:0] src37;
    reg [11:0] src38;
    reg [11:0] src39;
    reg [11:0] src40;
    reg [11:0] src41;
    reg [11:0] src42;
    reg [11:0] src43;
    reg [11:0] src44;
    reg [11:0] src45;
    reg [11:0] src46;
    reg [11:0] src47;
    reg [11:0] src48;
    reg [11:0] src49;
    reg [11:0] src50;
    reg [11:0] src51;
    reg [11:0] src52;
    reg [11:0] src53;
    reg [11:0] src54;
    reg [11:0] src55;
    reg [11:0] src56;
    reg [11:0] src57;
    reg [11:0] src58;
    reg [11:0] src59;
    reg [11:0] src60;
    reg [11:0] src61;
    reg [11:0] src62;
    reg [11:0] src63;
    compressor2_1_64_12 compressor2_1_64_12(.src0(src0), .src1(src1), .src2(src2), .src3(src3), .src4(src4), .src5(src5), .src6(src6), .src7(src7), .src8(src8), .src9(src9), .src10(src10), .src11(src11), .src12(src12), .src13(src13), .src14(src14), .src15(src15), .src16(src16), .src17(src17), .src18(src18), .src19(src19), .src20(src20), .src21(src21), .src22(src22), .src23(src23), .src24(src24), .src25(src25), .src26(src26), .src27(src27), .src28(src28), .src29(src29), .src30(src30), .src31(src31), .src32(src32), .src33(src33), .src34(src34), .src35(src35), .src36(src36), .src37(src37), .src38(src38), .src39(src39), .src40(src40), .src41(src41), .src42(src42), .src43(src43), .src44(src44), .src45(src45), .src46(src46), .src47(src47), .src48(src48), .src49(src49), .src50(src50), .src51(src51), .src52(src52), .src53(src53), .src54(src54), .src55(src55), .src56(src56), .src57(src57), .src58(src58), .src59(src59), .src60(src60), .src61(src61), .src62(src62), .src63(src63), .dst(dst));
    initial begin
        src0 <= 0;
        src1 <= 0;
        src2 <= 0;
        src3 <= 0;
        src4 <= 0;
        src5 <= 0;
        src6 <= 0;
        src7 <= 0;
        src8 <= 0;
        src9 <= 0;
        src10 <= 0;
        src11 <= 0;
        src12 <= 0;
        src13 <= 0;
        src14 <= 0;
        src15 <= 0;
        src16 <= 0;
        src17 <= 0;
        src18 <= 0;
        src19 <= 0;
        src20 <= 0;
        src21 <= 0;
        src22 <= 0;
        src23 <= 0;
        src24 <= 0;
        src25 <= 0;
        src26 <= 0;
        src27 <= 0;
        src28 <= 0;
        src29 <= 0;
        src30 <= 0;
        src31 <= 0;
        src32 <= 0;
        src33 <= 0;
        src34 <= 0;
        src35 <= 0;
        src36 <= 0;
        src37 <= 0;
        src38 <= 0;
        src39 <= 0;
        src40 <= 0;
        src41 <= 0;
        src42 <= 0;
        src43 <= 0;
        src44 <= 0;
        src45 <= 0;
        src46 <= 0;
        src47 <= 0;
        src48 <= 0;
        src49 <= 0;
        src50 <= 0;
        src51 <= 0;
        src52 <= 0;
        src53 <= 0;
        src54 <= 0;
        src55 <= 0;
        src56 <= 0;
        src57 <= 0;
        src58 <= 0;
        src59 <= 0;
        src60 <= 0;
        src61 <= 0;
        src62 <= 0;
        src63 <= 0;
    end
    always @(posedge clk) begin
        src0 <= {src0[10:0], in_data0};
        src1 <= {src1[10:0], in_data1};
        src2 <= {src2[10:0], in_data2};
        src3 <= {src3[10:0], in_data3};
        src4 <= {src4[10:0], in_data4};
        src5 <= {src5[10:0], in_data5};
        src6 <= {src6[10:0], in_data6};
        src7 <= {src7[10:0], in_data7};
        src8 <= {src8[10:0], in_data8};
        src9 <= {src9[10:0], in_data9};
        src10 <= {src10[10:0], in_data10};
        src11 <= {src11[10:0], in_data11};
        src12 <= {src12[10:0], in_data12};
        src13 <= {src13[10:0], in_data13};
        src14 <= {src14[10:0], in_data14};
        src15 <= {src15[10:0], in_data15};
        src16 <= {src16[10:0], in_data16};
        src17 <= {src17[10:0], in_data17};
        src18 <= {src18[10:0], in_data18};
        src19 <= {src19[10:0], in_data19};
        src20 <= {src20[10:0], in_data20};
        src21 <= {src21[10:0], in_data21};
        src22 <= {src22[10:0], in_data22};
        src23 <= {src23[10:0], in_data23};
        src24 <= {src24[10:0], in_data24};
        src25 <= {src25[10:0], in_data25};
        src26 <= {src26[10:0], in_data26};
        src27 <= {src27[10:0], in_data27};
        src28 <= {src28[10:0], in_data28};
        src29 <= {src29[10:0], in_data29};
        src30 <= {src30[10:0], in_data30};
        src31 <= {src31[10:0], in_data31};
        src32 <= {src32[10:0], in_data32};
        src33 <= {src33[10:0], in_data33};
        src34 <= {src34[10:0], in_data34};
        src35 <= {src35[10:0], in_data35};
        src36 <= {src36[10:0], in_data36};
        src37 <= {src37[10:0], in_data37};
        src38 <= {src38[10:0], in_data38};
        src39 <= {src39[10:0], in_data39};
        src40 <= {src40[10:0], in_data40};
        src41 <= {src41[10:0], in_data41};
        src42 <= {src42[10:0], in_data42};
        src43 <= {src43[10:0], in_data43};
        src44 <= {src44[10:0], in_data44};
        src45 <= {src45[10:0], in_data45};
        src46 <= {src46[10:0], in_data46};
        src47 <= {src47[10:0], in_data47};
        src48 <= {src48[10:0], in_data48};
        src49 <= {src49[10:0], in_data49};
        src50 <= {src50[10:0], in_data50};
        src51 <= {src51[10:0], in_data51};
        src52 <= {src52[10:0], in_data52};
        src53 <= {src53[10:0], in_data53};
        src54 <= {src54[10:0], in_data54};
        src55 <= {src55[10:0], in_data55};
        src56 <= {src56[10:0], in_data56};
        src57 <= {src57[10:0], in_data57};
        src58 <= {src58[10:0], in_data58};
        src59 <= {src59[10:0], in_data59};
        src60 <= {src60[10:0], in_data60};
        src61 <= {src61[10:0], in_data61};
        src62 <= {src62[10:0], in_data62};
        src63 <= {src63[10:0], in_data63};
    end
endmodule

module compressor2_1_64_12(
    input [11:0]src0,
    input [11:0]src1,
    input [11:0]src2,
    input [11:0]src3,
    input [11:0]src4,
    input [11:0]src5,
    input [11:0]src6,
    input [11:0]src7,
    input [11:0]src8,
    input [11:0]src9,
    input [11:0]src10,
    input [11:0]src11,
    input [11:0]src12,
    input [11:0]src13,
    input [11:0]src14,
    input [11:0]src15,
    input [11:0]src16,
    input [11:0]src17,
    input [11:0]src18,
    input [11:0]src19,
    input [11:0]src20,
    input [11:0]src21,
    input [11:0]src22,
    input [11:0]src23,
    input [11:0]src24,
    input [11:0]src25,
    input [11:0]src26,
    input [11:0]src27,
    input [11:0]src28,
    input [11:0]src29,
    input [11:0]src30,
    input [11:0]src31,
    input [11:0]src32,
    input [11:0]src33,
    input [11:0]src34,
    input [11:0]src35,
    input [11:0]src36,
    input [11:0]src37,
    input [11:0]src38,
    input [11:0]src39,
    input [11:0]src40,
    input [11:0]src41,
    input [11:0]src42,
    input [11:0]src43,
    input [11:0]src44,
    input [11:0]src45,
    input [11:0]src46,
    input [11:0]src47,
    input [11:0]src48,
    input [11:0]src49,
    input [11:0]src50,
    input [11:0]src51,
    input [11:0]src52,
    input [11:0]src53,
    input [11:0]src54,
    input [11:0]src55,
    input [11:0]src56,
    input [11:0]src57,
    input [11:0]src58,
    input [11:0]src59,
    input [11:0]src60,
    input [11:0]src61,
    input [11:0]src62,
    input [11:0]src63,
    output [17:0]dst);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [0:0] comp_out17;
    wire [18:0] out;
    compressor compressor_inst(
        .src0({src63[0], src62[0], src61[0], src60[0], src59[0], src58[0], src57[0], src56[0], src55[0], src54[0], src53[0], src52[0], src51[0], src50[0], src49[0], src48[0], src47[0], src46[0], src45[0], src44[0], src43[0], src42[0], src41[0], src40[0], src39[0], src38[0], src37[0], src36[0], src35[0], src34[0], src33[0], src32[0], src31[0], src30[0], src29[0], src28[0], src27[0], src26[0], src25[0], src24[0], src23[0], src22[0], src21[0], src20[0], src19[0], src18[0], src17[0], src16[0], src15[0], src14[0], src13[0], src12[0], src11[0], src10[0], src9[0], src8[0], src7[0], src6[0], src5[0], src4[0], src3[0], src2[0], src1[0], src0[0]}),
        .src1({src63[1], src62[1], src61[1], src60[1], src59[1], src58[1], src57[1], src56[1], src55[1], src54[1], src53[1], src52[1], src51[1], src50[1], src49[1], src48[1], src47[1], src46[1], src45[1], src44[1], src43[1], src42[1], src41[1], src40[1], src39[1], src38[1], src37[1], src36[1], src35[1], src34[1], src33[1], src32[1], src31[1], src30[1], src29[1], src28[1], src27[1], src26[1], src25[1], src24[1], src23[1], src22[1], src21[1], src20[1], src19[1], src18[1], src17[1], src16[1], src15[1], src14[1], src13[1], src12[1], src11[1], src10[1], src9[1], src8[1], src7[1], src6[1], src5[1], src4[1], src3[1], src2[1], src1[1], src0[1]}),
        .src2({src63[2], src62[2], src61[2], src60[2], src59[2], src58[2], src57[2], src56[2], src55[2], src54[2], src53[2], src52[2], src51[2], src50[2], src49[2], src48[2], src47[2], src46[2], src45[2], src44[2], src43[2], src42[2], src41[2], src40[2], src39[2], src38[2], src37[2], src36[2], src35[2], src34[2], src33[2], src32[2], src31[2], src30[2], src29[2], src28[2], src27[2], src26[2], src25[2], src24[2], src23[2], src22[2], src21[2], src20[2], src19[2], src18[2], src17[2], src16[2], src15[2], src14[2], src13[2], src12[2], src11[2], src10[2], src9[2], src8[2], src7[2], src6[2], src5[2], src4[2], src3[2], src2[2], src1[2], src0[2]}),
        .src3({src63[3], src62[3], src61[3], src60[3], src59[3], src58[3], src57[3], src56[3], src55[3], src54[3], src53[3], src52[3], src51[3], src50[3], src49[3], src48[3], src47[3], src46[3], src45[3], src44[3], src43[3], src42[3], src41[3], src40[3], src39[3], src38[3], src37[3], src36[3], src35[3], src34[3], src33[3], src32[3], src31[3], src30[3], src29[3], src28[3], src27[3], src26[3], src25[3], src24[3], src23[3], src22[3], src21[3], src20[3], src19[3], src18[3], src17[3], src16[3], src15[3], src14[3], src13[3], src12[3], src11[3], src10[3], src9[3], src8[3], src7[3], src6[3], src5[3], src4[3], src3[3], src2[3], src1[3], src0[3]}),
        .src4({src63[4], src62[4], src61[4], src60[4], src59[4], src58[4], src57[4], src56[4], src55[4], src54[4], src53[4], src52[4], src51[4], src50[4], src49[4], src48[4], src47[4], src46[4], src45[4], src44[4], src43[4], src42[4], src41[4], src40[4], src39[4], src38[4], src37[4], src36[4], src35[4], src34[4], src33[4], src32[4], src31[4], src30[4], src29[4], src28[4], src27[4], src26[4], src25[4], src24[4], src23[4], src22[4], src21[4], src20[4], src19[4], src18[4], src17[4], src16[4], src15[4], src14[4], src13[4], src12[4], src11[4], src10[4], src9[4], src8[4], src7[4], src6[4], src5[4], src4[4], src3[4], src2[4], src1[4], src0[4]}),
        .src5({src63[5], src62[5], src61[5], src60[5], src59[5], src58[5], src57[5], src56[5], src55[5], src54[5], src53[5], src52[5], src51[5], src50[5], src49[5], src48[5], src47[5], src46[5], src45[5], src44[5], src43[5], src42[5], src41[5], src40[5], src39[5], src38[5], src37[5], src36[5], src35[5], src34[5], src33[5], src32[5], src31[5], src30[5], src29[5], src28[5], src27[5], src26[5], src25[5], src24[5], src23[5], src22[5], src21[5], src20[5], src19[5], src18[5], src17[5], src16[5], src15[5], src14[5], src13[5], src12[5], src11[5], src10[5], src9[5], src8[5], src7[5], src6[5], src5[5], src4[5], src3[5], src2[5], src1[5], src0[5]}),
        .src6({src63[6], src62[6], src61[6], src60[6], src59[6], src58[6], src57[6], src56[6], src55[6], src54[6], src53[6], src52[6], src51[6], src50[6], src49[6], src48[6], src47[6], src46[6], src45[6], src44[6], src43[6], src42[6], src41[6], src40[6], src39[6], src38[6], src37[6], src36[6], src35[6], src34[6], src33[6], src32[6], src31[6], src30[6], src29[6], src28[6], src27[6], src26[6], src25[6], src24[6], src23[6], src22[6], src21[6], src20[6], src19[6], src18[6], src17[6], src16[6], src15[6], src14[6], src13[6], src12[6], src11[6], src10[6], src9[6], src8[6], src7[6], src6[6], src5[6], src4[6], src3[6], src2[6], src1[6], src0[6]}),
        .src7({src63[7], src62[7], src61[7], src60[7], src59[7], src58[7], src57[7], src56[7], src55[7], src54[7], src53[7], src52[7], src51[7], src50[7], src49[7], src48[7], src47[7], src46[7], src45[7], src44[7], src43[7], src42[7], src41[7], src40[7], src39[7], src38[7], src37[7], src36[7], src35[7], src34[7], src33[7], src32[7], src31[7], src30[7], src29[7], src28[7], src27[7], src26[7], src25[7], src24[7], src23[7], src22[7], src21[7], src20[7], src19[7], src18[7], src17[7], src16[7], src15[7], src14[7], src13[7], src12[7], src11[7], src10[7], src9[7], src8[7], src7[7], src6[7], src5[7], src4[7], src3[7], src2[7], src1[7], src0[7]}),
        .src8({src63[8], src62[8], src61[8], src60[8], src59[8], src58[8], src57[8], src56[8], src55[8], src54[8], src53[8], src52[8], src51[8], src50[8], src49[8], src48[8], src47[8], src46[8], src45[8], src44[8], src43[8], src42[8], src41[8], src40[8], src39[8], src38[8], src37[8], src36[8], src35[8], src34[8], src33[8], src32[8], src31[8], src30[8], src29[8], src28[8], src27[8], src26[8], src25[8], src24[8], src23[8], src22[8], src21[8], src20[8], src19[8], src18[8], src17[8], src16[8], src15[8], src14[8], src13[8], src12[8], src11[8], src10[8], src9[8], src8[8], src7[8], src6[8], src5[8], src4[8], src3[8], src2[8], src1[8], src0[8]}),
        .src9({src63[9], src62[9], src61[9], src60[9], src59[9], src58[9], src57[9], src56[9], src55[9], src54[9], src53[9], src52[9], src51[9], src50[9], src49[9], src48[9], src47[9], src46[9], src45[9], src44[9], src43[9], src42[9], src41[9], src40[9], src39[9], src38[9], src37[9], src36[9], src35[9], src34[9], src33[9], src32[9], src31[9], src30[9], src29[9], src28[9], src27[9], src26[9], src25[9], src24[9], src23[9], src22[9], src21[9], src20[9], src19[9], src18[9], src17[9], src16[9], src15[9], src14[9], src13[9], src12[9], src11[9], src10[9], src9[9], src8[9], src7[9], src6[9], src5[9], src4[9], src3[9], src2[9], src1[9], src0[9]}),
        .src10({src63[10], src62[10], src61[10], src60[10], src59[10], src58[10], src57[10], src56[10], src55[10], src54[10], src53[10], src52[10], src51[10], src50[10], src49[10], src48[10], src47[10], src46[10], src45[10], src44[10], src43[10], src42[10], src41[10], src40[10], src39[10], src38[10], src37[10], src36[10], src35[10], src34[10], src33[10], src32[10], src31[10], src30[10], src29[10], src28[10], src27[10], src26[10], src25[10], src24[10], src23[10], src22[10], src21[10], src20[10], src19[10], src18[10], src17[10], src16[10], src15[10], src14[10], src13[10], src12[10], src11[10], src10[10], src9[10], src8[10], src7[10], src6[10], src5[10], src4[10], src3[10], src2[10], src1[10], src0[10]}),
        .src11({src63[11], src62[11], src61[11], src60[11], src59[11], src58[11], src57[11], src56[11], src55[11], src54[11], src53[11], src52[11], src51[11], src50[11], src49[11], src48[11], src47[11], src46[11], src45[11], src44[11], src43[11], src42[11], src41[11], src40[11], src39[11], src38[11], src37[11], src36[11], src35[11], src34[11], src33[11], src32[11], src31[11], src30[11], src29[11], src28[11], src27[11], src26[11], src25[11], src24[11], src23[11], src22[11], src21[11], src20[11], src19[11], src18[11], src17[11], src16[11], src15[11], src14[11], src13[11], src12[11], src11[11], src10[11], src9[11], src8[11], src7[11], src6[11], src5[11], src4[11], src3[11], src2[11], src1[11], src0[11]}),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17)
    );
    rowadder2_1_18 rowadder2_1inst(
        .src0({comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst0(out)
    );
    assign dst = out[17:0];
endmodule
module compressor (
      input wire [63:0] src0,
      input wire [63:0] src1,
      input wire [63:0] src2,
      input wire [63:0] src3,
      input wire [63:0] src4,
      input wire [63:0] src5,
      input wire [63:0] src6,
      input wire [63:0] src7,
      input wire [63:0] src8,
      input wire [63:0] src9,
      input wire [63:0] src10,
      input wire [63:0] src11,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [0:0] dst17);

   wire [63:0] stage0_0;
   wire [63:0] stage0_1;
   wire [63:0] stage0_2;
   wire [63:0] stage0_3;
   wire [63:0] stage0_4;
   wire [63:0] stage0_5;
   wire [63:0] stage0_6;
   wire [63:0] stage0_7;
   wire [63:0] stage0_8;
   wire [63:0] stage0_9;
   wire [63:0] stage0_10;
   wire [63:0] stage0_11;
   wire [11:0] stage1_0;
   wire [19:0] stage1_1;
   wire [23:0] stage1_2;
   wire [24:0] stage1_3;
   wire [27:0] stage1_4;
   wire [30:0] stage1_5;
   wire [23:0] stage1_6;
   wire [21:0] stage1_7;
   wire [28:0] stage1_8;
   wire [30:0] stage1_9;
   wire [25:0] stage1_10;
   wire [21:0] stage1_11;
   wire [18:0] stage1_12;
   wire [11:0] stage1_13;
   wire [3:0] stage2_0;
   wire [4:0] stage2_1;
   wire [7:0] stage2_2;
   wire [9:0] stage2_3;
   wire [11:0] stage2_4;
   wire [11:0] stage2_5;
   wire [12:0] stage2_6;
   wire [9:0] stage2_7;
   wire [7:0] stage2_8;
   wire [11:0] stage2_9;
   wire [12:0] stage2_10;
   wire [10:0] stage2_11;
   wire [9:0] stage2_12;
   wire [5:0] stage2_13;
   wire [5:0] stage2_14;
   wire [1:0] stage2_15;
   wire [3:0] stage3_0;
   wire [4:0] stage3_1;
   wire [7:0] stage3_2;
   wire [1:0] stage3_3;
   wire [3:0] stage3_4;
   wire [3:0] stage3_5;
   wire [3:0] stage3_6;
   wire [5:0] stage3_7;
   wire [4:0] stage3_8;
   wire [2:0] stage3_9;
   wire [3:0] stage3_10;
   wire [5:0] stage3_11;
   wire [5:0] stage3_12;
   wire [2:0] stage3_13;
   wire [2:0] stage3_14;
   wire [3:0] stage3_15;
   wire [0:0] stage3_16;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [1:0] stage4_5;
   wire [1:0] stage4_6;
   wire [1:0] stage4_7;
   wire [1:0] stage4_8;
   wire [1:0] stage4_9;
   wire [1:0] stage4_10;
   wire [1:0] stage4_11;
   wire [1:0] stage4_12;
   wire [1:0] stage4_13;
   wire [1:0] stage4_14;
   wire [1:0] stage4_15;
   wire [1:0] stage4_16;
   wire [0:0] stage4_17;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage4_0;
   assign dst1 = stage4_1;
   assign dst2 = stage4_2;
   assign dst3 = stage4_3;
   assign dst4 = stage4_4;
   assign dst5 = stage4_5;
   assign dst6 = stage4_6;
   assign dst7 = stage4_7;
   assign dst8 = stage4_8;
   assign dst9 = stage4_9;
   assign dst10 = stage4_10;
   assign dst11 = stage4_11;
   assign dst12 = stage4_12;
   assign dst13 = stage4_13;
   assign dst14 = stage4_14;
   assign dst15 = stage4_15;
   assign dst16 = stage4_16;
   assign dst17 = stage4_17;

   gpc135_4 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc117_4 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11]},
      {stage0_1[3]},
      {stage0_2[1]},
      {stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc117_4 gpc2 (
      {stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18]},
      {stage0_1[4]},
      {stage0_2[2]},
      {stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc117_4 gpc3 (
      {stage0_0[19], stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25]},
      {stage0_1[5]},
      {stage0_2[3]},
      {stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc117_4 gpc4 (
      {stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32]},
      {stage0_1[6]},
      {stage0_2[4]},
      {stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc615_5 gpc5 (
      {stage0_0[33], stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37]},
      {stage0_1[7]},
      {stage0_2[5], stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10]},
      {stage1_4[0],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc615_5 gpc6 (
      {stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42]},
      {stage0_1[8]},
      {stage0_2[11], stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16]},
      {stage1_4[1],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc615_5 gpc7 (
      {stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47]},
      {stage0_1[9]},
      {stage0_2[17], stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22]},
      {stage1_4[2],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc615_5 gpc8 (
      {stage0_0[48], stage0_0[49], stage0_0[50], stage0_0[51], stage0_0[52]},
      {stage0_1[10]},
      {stage0_2[23], stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28]},
      {stage1_4[3],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc615_5 gpc9 (
      {stage0_0[53], stage0_0[54], stage0_0[55], stage0_0[56], stage0_0[57]},
      {stage0_1[11]},
      {stage0_2[29], stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34]},
      {stage1_4[4],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc615_5 gpc10 (
      {stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_1[12]},
      {stage0_2[35], stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40]},
      {stage1_4[5],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc606_5 gpc11 (
      {stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5]},
      {stage1_5[0],stage1_4[6],stage1_3[11],stage1_2[11],stage1_1[11]}
   );
   gpc606_5 gpc12 (
      {stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24]},
      {stage0_3[6], stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11]},
      {stage1_5[1],stage1_4[7],stage1_3[12],stage1_2[12],stage1_1[12]}
   );
   gpc606_5 gpc13 (
      {stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30]},
      {stage0_3[12], stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17]},
      {stage1_5[2],stage1_4[8],stage1_3[13],stage1_2[13],stage1_1[13]}
   );
   gpc606_5 gpc14 (
      {stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36]},
      {stage0_3[18], stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23]},
      {stage1_5[3],stage1_4[9],stage1_3[14],stage1_2[14],stage1_1[14]}
   );
   gpc606_5 gpc15 (
      {stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42]},
      {stage0_3[24], stage0_3[25], stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29]},
      {stage1_5[4],stage1_4[10],stage1_3[15],stage1_2[15],stage1_1[15]}
   );
   gpc606_5 gpc16 (
      {stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48]},
      {stage0_3[30], stage0_3[31], stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35]},
      {stage1_5[5],stage1_4[11],stage1_3[16],stage1_2[16],stage1_1[16]}
   );
   gpc615_5 gpc17 (
      {stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_2[41]},
      {stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41]},
      {stage1_5[6],stage1_4[12],stage1_3[17],stage1_2[17],stage1_1[17]}
   );
   gpc615_5 gpc18 (
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58]},
      {stage0_2[42]},
      {stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47]},
      {stage1_5[7],stage1_4[13],stage1_3[18],stage1_2[18],stage1_1[18]}
   );
   gpc615_5 gpc19 (
      {stage0_1[59], stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63]},
      {stage0_2[43]},
      {stage0_3[48], stage0_3[49], stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53]},
      {stage1_5[8],stage1_4[14],stage1_3[19],stage1_2[19],stage1_1[19]}
   );
   gpc615_5 gpc20 (
      {stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48]},
      {stage0_3[54]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[9],stage1_4[15],stage1_3[20],stage1_2[20]}
   );
   gpc615_5 gpc21 (
      {stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53]},
      {stage0_3[55]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[10],stage1_4[16],stage1_3[21],stage1_2[21]}
   );
   gpc615_5 gpc22 (
      {stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58]},
      {stage0_3[56]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[11],stage1_4[17],stage1_3[22],stage1_2[22]}
   );
   gpc615_5 gpc23 (
      {stage0_2[59], stage0_2[60], stage0_2[61], stage0_2[62], stage0_2[63]},
      {stage0_3[57]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[12],stage1_4[18],stage1_3[23],stage1_2[23]}
   );
   gpc606_5 gpc24 (
      {stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62], stage0_3[63]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[4],stage1_5[13],stage1_4[19],stage1_3[24]}
   );
   gpc615_5 gpc25 (
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28]},
      {stage0_5[6]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[1],stage1_6[5],stage1_5[14],stage1_4[20]}
   );
   gpc615_5 gpc26 (
      {stage0_4[29], stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33]},
      {stage0_5[7]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[2],stage1_6[6],stage1_5[15],stage1_4[21]}
   );
   gpc615_5 gpc27 (
      {stage0_4[34], stage0_4[35], stage0_4[36], stage0_4[37], stage0_4[38]},
      {stage0_5[8]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[3],stage1_6[7],stage1_5[16],stage1_4[22]}
   );
   gpc615_5 gpc28 (
      {stage0_4[39], stage0_4[40], stage0_4[41], stage0_4[42], stage0_4[43]},
      {stage0_5[9]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[4],stage1_6[8],stage1_5[17],stage1_4[23]}
   );
   gpc615_5 gpc29 (
      {stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47], stage0_4[48]},
      {stage0_5[10]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[5],stage1_6[9],stage1_5[18],stage1_4[24]}
   );
   gpc615_5 gpc30 (
      {stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage0_5[11]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[6],stage1_6[10],stage1_5[19],stage1_4[25]}
   );
   gpc615_5 gpc31 (
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58]},
      {stage0_5[12]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[7],stage1_6[11],stage1_5[20],stage1_4[26]}
   );
   gpc615_5 gpc32 (
      {stage0_4[59], stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63]},
      {stage0_5[13]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[8],stage1_6[12],stage1_5[21],stage1_4[27]}
   );
   gpc606_5 gpc33 (
      {stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17], stage0_5[18], stage0_5[19]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[8],stage1_7[9],stage1_6[13],stage1_5[22]}
   );
   gpc606_5 gpc34 (
      {stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23], stage0_5[24], stage0_5[25]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[9],stage1_7[10],stage1_6[14],stage1_5[23]}
   );
   gpc606_5 gpc35 (
      {stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29], stage0_5[30], stage0_5[31]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[10],stage1_7[11],stage1_6[15],stage1_5[24]}
   );
   gpc606_5 gpc36 (
      {stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35], stage0_5[36], stage0_5[37]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[11],stage1_7[12],stage1_6[16],stage1_5[25]}
   );
   gpc606_5 gpc37 (
      {stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41], stage0_5[42], stage0_5[43]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[12],stage1_7[13],stage1_6[17],stage1_5[26]}
   );
   gpc615_5 gpc38 (
      {stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47], stage0_5[48]},
      {stage0_6[48]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[13],stage1_7[14],stage1_6[18],stage1_5[27]}
   );
   gpc615_5 gpc39 (
      {stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_6[49]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[14],stage1_7[15],stage1_6[19],stage1_5[28]}
   );
   gpc615_5 gpc40 (
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58]},
      {stage0_6[50]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[15],stage1_7[16],stage1_6[20],stage1_5[29]}
   );
   gpc615_5 gpc41 (
      {stage0_5[59], stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63]},
      {stage0_6[51]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[16],stage1_7[17],stage1_6[21],stage1_5[30]}
   );
   gpc606_5 gpc42 (
      {stage0_6[52], stage0_6[53], stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[9],stage1_8[17],stage1_7[18],stage1_6[22]}
   );
   gpc606_5 gpc43 (
      {stage0_6[58], stage0_6[59], stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[10],stage1_8[18],stage1_7[19],stage1_6[23]}
   );
   gpc2135_5 gpc44 (
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58]},
      {stage0_8[12], stage0_8[13], stage0_8[14]},
      {stage0_9[0]},
      {stage0_10[0], stage0_10[1]},
      {stage1_11[0],stage1_10[2],stage1_9[11],stage1_8[19],stage1_7[20]}
   );
   gpc615_5 gpc45 (
      {stage0_7[59], stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63]},
      {stage0_8[15]},
      {stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5], stage0_9[6]},
      {stage1_11[1],stage1_10[3],stage1_9[12],stage1_8[20],stage1_7[21]}
   );
   gpc207_4 gpc46 (
      {stage0_8[16], stage0_8[17], stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22]},
      {stage0_10[2], stage0_10[3]},
      {stage1_11[2],stage1_10[4],stage1_9[13],stage1_8[21]}
   );
   gpc606_5 gpc47 (
      {stage0_8[23], stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28]},
      {stage0_10[4], stage0_10[5], stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9]},
      {stage1_12[0],stage1_11[3],stage1_10[5],stage1_9[14],stage1_8[22]}
   );
   gpc606_5 gpc48 (
      {stage0_8[29], stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34]},
      {stage0_10[10], stage0_10[11], stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15]},
      {stage1_12[1],stage1_11[4],stage1_10[6],stage1_9[15],stage1_8[23]}
   );
   gpc606_5 gpc49 (
      {stage0_8[35], stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40]},
      {stage0_10[16], stage0_10[17], stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21]},
      {stage1_12[2],stage1_11[5],stage1_10[7],stage1_9[16],stage1_8[24]}
   );
   gpc606_5 gpc50 (
      {stage0_8[41], stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46]},
      {stage0_10[22], stage0_10[23], stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27]},
      {stage1_12[3],stage1_11[6],stage1_10[8],stage1_9[17],stage1_8[25]}
   );
   gpc606_5 gpc51 (
      {stage0_8[47], stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52]},
      {stage0_10[28], stage0_10[29], stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33]},
      {stage1_12[4],stage1_11[7],stage1_10[9],stage1_9[18],stage1_8[26]}
   );
   gpc606_5 gpc52 (
      {stage0_8[53], stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58]},
      {stage0_10[34], stage0_10[35], stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39]},
      {stage1_12[5],stage1_11[8],stage1_10[10],stage1_9[19],stage1_8[27]}
   );
   gpc615_5 gpc53 (
      {stage0_8[59], stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63]},
      {stage0_9[7]},
      {stage0_10[40], stage0_10[41], stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45]},
      {stage1_12[6],stage1_11[9],stage1_10[11],stage1_9[20],stage1_8[28]}
   );
   gpc606_5 gpc54 (
      {stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11], stage0_9[12], stage0_9[13]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[7],stage1_11[10],stage1_10[12],stage1_9[21]}
   );
   gpc606_5 gpc55 (
      {stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17], stage0_9[18], stage0_9[19]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[8],stage1_11[11],stage1_10[13],stage1_9[22]}
   );
   gpc606_5 gpc56 (
      {stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[9],stage1_11[12],stage1_10[14],stage1_9[23]}
   );
   gpc606_5 gpc57 (
      {stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[10],stage1_11[13],stage1_10[15],stage1_9[24]}
   );
   gpc606_5 gpc58 (
      {stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35], stage0_9[36], stage0_9[37]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[11],stage1_11[14],stage1_10[16],stage1_9[25]}
   );
   gpc606_5 gpc59 (
      {stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[12],stage1_11[15],stage1_10[17],stage1_9[26]}
   );
   gpc615_5 gpc60 (
      {stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47], stage0_9[48]},
      {stage0_10[46]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[13],stage1_11[16],stage1_10[18],stage1_9[27]}
   );
   gpc615_5 gpc61 (
      {stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage0_10[47]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[14],stage1_11[17],stage1_10[19],stage1_9[28]}
   );
   gpc615_5 gpc62 (
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58]},
      {stage0_10[48]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[15],stage1_11[18],stage1_10[20],stage1_9[29]}
   );
   gpc615_5 gpc63 (
      {stage0_9[59], stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63]},
      {stage0_10[49]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[16],stage1_11[19],stage1_10[21],stage1_9[30]}
   );
   gpc135_4 gpc64 (
      {stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53], stage0_10[54]},
      {stage0_11[60], stage0_11[61], stage0_11[62]},
      {1'b0},
      {stage1_13[10],stage1_12[17],stage1_11[20],stage1_10[22]}
   );
   gpc117_4 gpc65 (
      {stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59], stage0_10[60], stage0_10[61]},
      {stage0_11[63]},
      {1'b0},
      {stage1_13[11],stage1_12[18],stage1_11[21],stage1_10[23]}
   );
   gpc1_1 gpc66 (
      {stage0_0[63]},
      {stage1_0[11]}
   );
   gpc1_1 gpc67 (
      {stage0_10[62]},
      {stage1_10[24]}
   );
   gpc1_1 gpc68 (
      {stage0_10[63]},
      {stage1_10[25]}
   );
   gpc2135_5 gpc69 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4]},
      {stage1_1[0], stage1_1[1], stage1_1[2]},
      {stage1_2[0]},
      {stage1_3[0], stage1_3[1]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc615_5 gpc70 (
      {stage1_0[5], stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9]},
      {stage1_1[3]},
      {stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc2135_5 gpc71 (
      {stage1_1[4], stage1_1[5], stage1_1[6], stage1_1[7], stage1_1[8]},
      {stage1_2[7], stage1_2[8], stage1_2[9]},
      {stage1_3[2]},
      {stage1_4[0], stage1_4[1]},
      {stage2_5[0],stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2]}
   );
   gpc2135_5 gpc72 (
      {stage1_1[9], stage1_1[10], stage1_1[11], stage1_1[12], stage1_1[13]},
      {stage1_2[10], stage1_2[11], stage1_2[12]},
      {stage1_3[3]},
      {stage1_4[2], stage1_4[3]},
      {stage2_5[1],stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3]}
   );
   gpc1406_5 gpc73 (
      {stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17], stage1_1[18], stage1_1[19]},
      {stage1_3[4], stage1_3[5], stage1_3[6], stage1_3[7]},
      {stage1_4[4]},
      {stage2_5[2],stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4]}
   );
   gpc615_5 gpc74 (
      {stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17]},
      {stage1_3[8]},
      {stage1_4[5], stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10]},
      {stage2_6[0],stage2_5[3],stage2_4[5],stage2_3[5],stage2_2[5]}
   );
   gpc615_5 gpc75 (
      {stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22]},
      {stage1_3[9]},
      {stage1_4[11], stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16]},
      {stage2_6[1],stage2_5[4],stage2_4[6],stage2_3[6],stage2_2[6]}
   );
   gpc615_5 gpc76 (
      {stage1_3[10], stage1_3[11], stage1_3[12], stage1_3[13], stage1_3[14]},
      {stage1_4[17]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[2],stage2_5[5],stage2_4[7],stage2_3[7]}
   );
   gpc615_5 gpc77 (
      {stage1_3[15], stage1_3[16], stage1_3[17], stage1_3[18], stage1_3[19]},
      {stage1_4[18]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[3],stage2_5[6],stage2_4[8],stage2_3[8]}
   );
   gpc615_5 gpc78 (
      {stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23], stage1_3[24]},
      {stage1_4[19]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[4],stage2_5[7],stage2_4[9],stage2_3[9]}
   );
   gpc7_3 gpc79 (
      {stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23], stage1_4[24], stage1_4[25], stage1_4[26]},
      {stage2_6[5],stage2_5[8],stage2_4[10]}
   );
   gpc615_5 gpc80 (
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22]},
      {stage1_6[0]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[0],stage2_7[3],stage2_6[6],stage2_5[9]}
   );
   gpc615_5 gpc81 (
      {stage1_5[23], stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27]},
      {stage1_6[1]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[1],stage2_7[4],stage2_6[7],stage2_5[10]}
   );
   gpc623_5 gpc82 (
      {stage1_5[28], stage1_5[29], stage1_5[30]},
      {stage1_6[2], stage1_6[3]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[2],stage2_7[5],stage2_6[8],stage2_5[11]}
   );
   gpc615_5 gpc83 (
      {stage1_6[4], stage1_6[5], stage1_6[6], stage1_6[7], stage1_6[8]},
      {stage1_7[18]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[3],stage2_8[3],stage2_7[6],stage2_6[9]}
   );
   gpc615_5 gpc84 (
      {stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12], stage1_6[13]},
      {stage1_7[19]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[4],stage2_8[4],stage2_7[7],stage2_6[10]}
   );
   gpc615_5 gpc85 (
      {stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17], stage1_6[18]},
      {stage1_7[20]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[5],stage2_8[5],stage2_7[8],stage2_6[11]}
   );
   gpc615_5 gpc86 (
      {stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage1_7[21]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[6],stage2_8[6],stage2_7[9],stage2_6[12]}
   );
   gpc135_4 gpc87 (
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28]},
      {stage1_9[0], stage1_9[1], stage1_9[2]},
      {stage1_10[0]},
      {stage2_11[0],stage2_10[4],stage2_9[7],stage2_8[7]}
   );
   gpc117_4 gpc88 (
      {stage1_9[3], stage1_9[4], stage1_9[5], stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9]},
      {stage1_10[1]},
      {stage1_11[0]},
      {stage2_12[0],stage2_11[1],stage2_10[5],stage2_9[8]}
   );
   gpc117_4 gpc89 (
      {stage1_9[10], stage1_9[11], stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16]},
      {stage1_10[2]},
      {stage1_11[1]},
      {stage2_12[1],stage2_11[2],stage2_10[6],stage2_9[9]}
   );
   gpc117_4 gpc90 (
      {stage1_9[17], stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage1_10[3]},
      {stage1_11[2]},
      {stage2_12[2],stage2_11[3],stage2_10[7],stage2_9[10]}
   );
   gpc117_4 gpc91 (
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29], stage1_9[30]},
      {stage1_10[4]},
      {stage1_11[3]},
      {stage2_12[3],stage2_11[4],stage2_10[8],stage2_9[11]}
   );
   gpc1163_5 gpc92 (
      {stage1_10[5], stage1_10[6], stage1_10[7]},
      {stage1_11[4], stage1_11[5], stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9]},
      {stage1_12[0]},
      {stage1_13[0]},
      {stage2_14[0],stage2_13[0],stage2_12[4],stage2_11[5],stage2_10[9]}
   );
   gpc606_5 gpc93 (
      {stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11], stage1_10[12], stage1_10[13]},
      {stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5], stage1_12[6]},
      {stage2_14[1],stage2_13[1],stage2_12[5],stage2_11[6],stage2_10[10]}
   );
   gpc606_5 gpc94 (
      {stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17], stage1_10[18], stage1_10[19]},
      {stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11], stage1_12[12]},
      {stage2_14[2],stage2_13[2],stage2_12[6],stage2_11[7],stage2_10[11]}
   );
   gpc606_5 gpc95 (
      {stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23], stage1_10[24], stage1_10[25]},
      {stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17], stage1_12[18]},
      {stage2_14[3],stage2_13[3],stage2_12[7],stage2_11[8],stage2_10[12]}
   );
   gpc606_5 gpc96 (
      {stage1_11[10], stage1_11[11], stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15]},
      {stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5], stage1_13[6]},
      {stage2_15[0],stage2_14[4],stage2_13[4],stage2_12[8],stage2_11[9]}
   );
   gpc606_5 gpc97 (
      {stage1_11[16], stage1_11[17], stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21]},
      {stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11], 1'b0},
      {stage2_15[1],stage2_14[5],stage2_13[5],stage2_12[9],stage2_11[10]}
   );
   gpc1_1 gpc98 (
      {stage1_0[10]},
      {stage2_0[2]}
   );
   gpc1_1 gpc99 (
      {stage1_0[11]},
      {stage2_0[3]}
   );
   gpc1_1 gpc100 (
      {stage1_2[23]},
      {stage2_2[7]}
   );
   gpc1_1 gpc101 (
      {stage1_4[27]},
      {stage2_4[11]}
   );
   gpc1415_5 gpc102 (
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4]},
      {stage2_4[0]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3]},
      {stage2_6[0]},
      {stage3_7[0],stage3_6[0],stage3_5[0],stage3_4[0],stage3_3[0]}
   );
   gpc615_5 gpc103 (
      {stage2_3[5], stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9]},
      {stage2_4[1]},
      {stage2_5[4], stage2_5[5], stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9]},
      {stage3_7[1],stage3_6[1],stage3_5[1],stage3_4[1],stage3_3[1]}
   );
   gpc615_5 gpc104 (
      {stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5], stage2_4[6]},
      {stage2_5[10]},
      {stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5], stage2_6[6]},
      {stage3_8[0],stage3_7[2],stage3_6[2],stage3_5[2],stage3_4[2]}
   );
   gpc615_5 gpc105 (
      {stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage2_5[11]},
      {stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11], stage2_6[12]},
      {stage3_8[1],stage3_7[3],stage3_6[3],stage3_5[3],stage3_4[3]}
   );
   gpc615_5 gpc106 (
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4]},
      {stage2_8[0]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[0],stage3_9[0],stage3_8[2],stage3_7[4]}
   );
   gpc615_5 gpc107 (
      {stage2_7[5], stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9]},
      {stage2_8[1]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[1],stage3_9[1],stage3_8[3],stage3_7[5]}
   );
   gpc606_5 gpc108 (
      {stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5], stage2_8[6], stage2_8[7]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[2],stage3_10[2],stage3_9[2],stage3_8[4]}
   );
   gpc7_3 gpc109 (
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11], stage2_10[12]},
      {stage3_12[1],stage3_11[3],stage3_10[3]}
   );
   gpc135_4 gpc110 (
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4]},
      {stage2_12[0], stage2_12[1], stage2_12[2]},
      {stage2_13[0]},
      {stage3_14[0],stage3_13[0],stage3_12[2],stage3_11[4]}
   );
   gpc606_5 gpc111 (
      {stage2_11[5], stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10]},
      {stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5], 1'b0},
      {stage3_15[0],stage3_14[1],stage3_13[1],stage3_12[3],stage3_11[5]}
   );
   gpc606_5 gpc112 (
      {stage2_12[3], stage2_12[4], stage2_12[5], stage2_12[6], stage2_12[7], stage2_12[8]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[1],stage3_14[2],stage3_13[2],stage3_12[4]}
   );
   gpc1_1 gpc113 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc114 (
      {stage2_0[1]},
      {stage3_0[1]}
   );
   gpc1_1 gpc115 (
      {stage2_0[2]},
      {stage3_0[2]}
   );
   gpc1_1 gpc116 (
      {stage2_0[3]},
      {stage3_0[3]}
   );
   gpc1_1 gpc117 (
      {stage2_1[0]},
      {stage3_1[0]}
   );
   gpc1_1 gpc118 (
      {stage2_1[1]},
      {stage3_1[1]}
   );
   gpc1_1 gpc119 (
      {stage2_1[2]},
      {stage3_1[2]}
   );
   gpc1_1 gpc120 (
      {stage2_1[3]},
      {stage3_1[3]}
   );
   gpc1_1 gpc121 (
      {stage2_1[4]},
      {stage3_1[4]}
   );
   gpc1_1 gpc122 (
      {stage2_2[0]},
      {stage3_2[0]}
   );
   gpc1_1 gpc123 (
      {stage2_2[1]},
      {stage3_2[1]}
   );
   gpc1_1 gpc124 (
      {stage2_2[2]},
      {stage3_2[2]}
   );
   gpc1_1 gpc125 (
      {stage2_2[3]},
      {stage3_2[3]}
   );
   gpc1_1 gpc126 (
      {stage2_2[4]},
      {stage3_2[4]}
   );
   gpc1_1 gpc127 (
      {stage2_2[5]},
      {stage3_2[5]}
   );
   gpc1_1 gpc128 (
      {stage2_2[6]},
      {stage3_2[6]}
   );
   gpc1_1 gpc129 (
      {stage2_2[7]},
      {stage3_2[7]}
   );
   gpc1_1 gpc130 (
      {stage2_12[9]},
      {stage3_12[5]}
   );
   gpc1_1 gpc131 (
      {stage2_15[0]},
      {stage3_15[2]}
   );
   gpc1_1 gpc132 (
      {stage2_15[1]},
      {stage3_15[3]}
   );
   gpc1343_5 gpc133 (
      {stage3_0[0], stage3_0[1], stage3_0[2]},
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3]},
      {stage3_2[0], stage3_2[1], stage3_2[2]},
      {stage3_3[0]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc1415_5 gpc134 (
      {stage3_2[3], stage3_2[4], stage3_2[5], stage3_2[6], stage3_2[7]},
      {stage3_3[1]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3]},
      {stage3_5[0]},
      {stage4_6[0],stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1]}
   );
   gpc1343_5 gpc135 (
      {stage3_5[1], stage3_5[2], stage3_5[3]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3]},
      {stage3_7[0], stage3_7[1], stage3_7[2]},
      {stage3_8[0]},
      {stage4_9[0],stage4_8[0],stage4_7[0],stage4_6[1],stage4_5[1]}
   );
   gpc1343_5 gpc136 (
      {stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4]},
      {stage3_9[0], stage3_9[1], stage3_9[2]},
      {stage3_10[0]},
      {stage4_11[0],stage4_10[0],stage4_9[1],stage4_8[1],stage4_7[1]}
   );
   gpc1163_5 gpc137 (
      {stage3_10[1], stage3_10[2], stage3_10[3]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage3_12[0]},
      {stage3_13[0]},
      {stage4_14[0],stage4_13[0],stage4_12[0],stage4_11[1],stage4_10[1]}
   );
   gpc1325_5 gpc138 (
      {stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage3_13[1], stage3_13[2]},
      {stage3_14[0], stage3_14[1], stage3_14[2]},
      {stage3_15[0]},
      {stage4_16[0],stage4_15[0],stage4_14[1],stage4_13[1],stage4_12[1]}
   );
   gpc117_4 gpc139 (
      {stage3_15[1], stage3_15[2], stage3_15[3], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage3_16[0]},
      {1'b0},
      {stage4_17[0],stage4_16[1],stage4_15[1]}
   );
   gpc1_1 gpc140 (
      {stage3_0[3]},
      {stage4_0[1]}
   );
   gpc1_1 gpc141 (
      {stage3_1[4]},
      {stage4_1[1]}
   );
endmodule
module rowadder2_1_18(input [17:0] src0, input [17:0] src1, output [18:0] dst0);
    wire [17:0] gene;
    wire [17:0] prop;
    wire [19:0] out;
    wire [19:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI({2'h0, gene[17:16]}),
        .S({2'h0, prop[17:16]})
    );
    assign dst0 = {carryout[17], out[17:0]};
endmodule


module comp2_1test_64_12();
    reg [11:0] src0;
    reg [11:0] src1;
    reg [11:0] src2;
    reg [11:0] src3;
    reg [11:0] src4;
    reg [11:0] src5;
    reg [11:0] src6;
    reg [11:0] src7;
    reg [11:0] src8;
    reg [11:0] src9;
    reg [11:0] src10;
    reg [11:0] src11;
    reg [11:0] src12;
    reg [11:0] src13;
    reg [11:0] src14;
    reg [11:0] src15;
    reg [11:0] src16;
    reg [11:0] src17;
    reg [11:0] src18;
    reg [11:0] src19;
    reg [11:0] src20;
    reg [11:0] src21;
    reg [11:0] src22;
    reg [11:0] src23;
    reg [11:0] src24;
    reg [11:0] src25;
    reg [11:0] src26;
    reg [11:0] src27;
    reg [11:0] src28;
    reg [11:0] src29;
    reg [11:0] src30;
    reg [11:0] src31;
    reg [11:0] src32;
    reg [11:0] src33;
    reg [11:0] src34;
    reg [11:0] src35;
    reg [11:0] src36;
    reg [11:0] src37;
    reg [11:0] src38;
    reg [11:0] src39;
    reg [11:0] src40;
    reg [11:0] src41;
    reg [11:0] src42;
    reg [11:0] src43;
    reg [11:0] src44;
    reg [11:0] src45;
    reg [11:0] src46;
    reg [11:0] src47;
    reg [11:0] src48;
    reg [11:0] src49;
    reg [11:0] src50;
    reg [11:0] src51;
    reg [11:0] src52;
    reg [11:0] src53;
    reg [11:0] src54;
    reg [11:0] src55;
    reg [11:0] src56;
    reg [11:0] src57;
    reg [11:0] src58;
    reg [11:0] src59;
    reg [11:0] src60;
    reg [11:0] src61;
    reg [11:0] src62;
    reg [11:0] src63;
    reg [17:0] exp;
    wire [17:0] dst;
    assign test = dst == exp;
    compressor2_1_64_12 compressor2_1_64_12_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst(dst)
    );
    initial begin
        $monitor("0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x %x", src0, src1, src2, src3, src4, src5, src6, src7, src8, src9, src10, src11, src12, src13, src14, src15, src16, src17, src18, src19, src20, src21, src22, src23, src24, src25, src26, src27, src28, src29, src30, src31, src32, src33, src34, src35, src36, src37, src38, src39, src40, src41, src42, src43, src44, src45, src46, src47, src48, src49, src50, src51, src52, src53, src54, src55, src56, src57, src58, src59, src60, src61, src62, src63, dst, exp, test);
        src0 <= 12'hfa6;
        src1 <= 12'h599;
        src2 <= 12'h4c4;
        src3 <= 12'h86b;
        src4 <= 12'h918;
        src5 <= 12'h58d;
        src6 <= 12'h52d;
        src7 <= 12'hc01;
        src8 <= 12'h508;
        src9 <= 12'hc4c;
        src10 <= 12'h69d;
        src11 <= 12'hadf;
        src12 <= 12'hd27;
        src13 <= 12'he97;
        src14 <= 12'ha7a;
        src15 <= 12'h660;
        src16 <= 12'hc13;
        src17 <= 12'h7d;
        src18 <= 12'h7bc;
        src19 <= 12'hcfa;
        src20 <= 12'h774;
        src21 <= 12'h4db;
        src22 <= 12'h968;
        src23 <= 12'h46c;
        src24 <= 12'hba3;
        src25 <= 12'hcfb;
        src26 <= 12'hbde;
        src27 <= 12'h269;
        src28 <= 12'h77f;
        src29 <= 12'he2f;
        src30 <= 12'habd;
        src31 <= 12'h5e0;
        src32 <= 12'ha4c;
        src33 <= 12'ha98;
        src34 <= 12'h2d5;
        src35 <= 12'h7c4;
        src36 <= 12'h759;
        src37 <= 12'h8f1;
        src38 <= 12'h8a9;
        src39 <= 12'hcbc;
        src40 <= 12'h5f4;
        src41 <= 12'ha9b;
        src42 <= 12'hdb2;
        src43 <= 12'h2cd;
        src44 <= 12'h5ea;
        src45 <= 12'h6a3;
        src46 <= 12'h453;
        src47 <= 12'h496;
        src48 <= 12'hb14;
        src49 <= 12'he7;
        src50 <= 12'h446;
        src51 <= 12'h54a;
        src52 <= 12'h962;
        src53 <= 12'h7fa;
        src54 <= 12'h3b2;
        src55 <= 12'he7;
        src56 <= 12'ha45;
        src57 <= 12'hca9;
        src58 <= 12'h45c;
        src59 <= 12'h443;
        src60 <= 12'hd3d;
        src61 <= 12'h4af;
        src62 <= 12'h76;
        src63 <= 12'h49;
        exp <= 18'h1f3aa;
        #1
        src0 <= 12'hde9;
        src1 <= 12'h771;
        src2 <= 12'hd2b;
        src3 <= 12'h964;
        src4 <= 12'h85e;
        src5 <= 12'he64;
        src6 <= 12'h925;
        src7 <= 12'h6a5;
        src8 <= 12'hcb1;
        src9 <= 12'h13e;
        src10 <= 12'hec1;
        src11 <= 12'h38;
        src12 <= 12'hfd5;
        src13 <= 12'h5c7;
        src14 <= 12'h4ab;
        src15 <= 12'hdc2;
        src16 <= 12'h882;
        src17 <= 12'h72f;
        src18 <= 12'hc55;
        src19 <= 12'hfda;
        src20 <= 12'hcfb;
        src21 <= 12'h4f5;
        src22 <= 12'hb8f;
        src23 <= 12'hc97;
        src24 <= 12'h207;
        src25 <= 12'h3e6;
        src26 <= 12'hd40;
        src27 <= 12'hae6;
        src28 <= 12'hf76;
        src29 <= 12'hb6b;
        src30 <= 12'h896;
        src31 <= 12'he66;
        src32 <= 12'hdd7;
        src33 <= 12'h3d0;
        src34 <= 12'h3a1;
        src35 <= 12'h899;
        src36 <= 12'hcdb;
        src37 <= 12'h145;
        src38 <= 12'heb5;
        src39 <= 12'hd2d;
        src40 <= 12'h6db;
        src41 <= 12'hbc2;
        src42 <= 12'h5fe;
        src43 <= 12'h3a3;
        src44 <= 12'h32;
        src45 <= 12'h2d5;
        src46 <= 12'h278;
        src47 <= 12'h60c;
        src48 <= 12'hb5e;
        src49 <= 12'he8b;
        src50 <= 12'hc9b;
        src51 <= 12'h9ee;
        src52 <= 12'h598;
        src53 <= 12'h4c3;
        src54 <= 12'h850;
        src55 <= 12'hb25;
        src56 <= 12'hf84;
        src57 <= 12'hd71;
        src58 <= 12'hd2c;
        src59 <= 12'hae8;
        src60 <= 12'h61a;
        src61 <= 12'hc12;
        src62 <= 12'h89b;
        src63 <= 12'h6bd;
        exp <= 18'h251c7;
        #1
        src0 <= 12'h114;
        src1 <= 12'h4fb;
        src2 <= 12'hb21;
        src3 <= 12'h530;
        src4 <= 12'h8c;
        src5 <= 12'hf5f;
        src6 <= 12'h246;
        src7 <= 12'h222;
        src8 <= 12'h404;
        src9 <= 12'hc6;
        src10 <= 12'h518;
        src11 <= 12'h6ad;
        src12 <= 12'hedf;
        src13 <= 12'h92c;
        src14 <= 12'h7cb;
        src15 <= 12'h8ca;
        src16 <= 12'hd99;
        src17 <= 12'h1f5;
        src18 <= 12'hbfb;
        src19 <= 12'h2d7;
        src20 <= 12'he85;
        src21 <= 12'h720;
        src22 <= 12'hb05;
        src23 <= 12'h5cd;
        src24 <= 12'h8bc;
        src25 <= 12'h35;
        src26 <= 12'h1c5;
        src27 <= 12'hb85;
        src28 <= 12'h70c;
        src29 <= 12'hee1;
        src30 <= 12'hc96;
        src31 <= 12'h66b;
        src32 <= 12'h842;
        src33 <= 12'ha40;
        src34 <= 12'hd15;
        src35 <= 12'h42c;
        src36 <= 12'ha8c;
        src37 <= 12'h37c;
        src38 <= 12'h39d;
        src39 <= 12'h6e9;
        src40 <= 12'hf5b;
        src41 <= 12'h59c;
        src42 <= 12'hba0;
        src43 <= 12'h6d6;
        src44 <= 12'h686;
        src45 <= 12'hf11;
        src46 <= 12'h589;
        src47 <= 12'he1d;
        src48 <= 12'hf96;
        src49 <= 12'h342;
        src50 <= 12'h586;
        src51 <= 12'h40a;
        src52 <= 12'h8b8;
        src53 <= 12'h321;
        src54 <= 12'h4bf;
        src55 <= 12'h974;
        src56 <= 12'hb3c;
        src57 <= 12'h114;
        src58 <= 12'h9;
        src59 <= 12'h334;
        src60 <= 12'hf2f;
        src61 <= 12'h293;
        src62 <= 12'h948;
        src63 <= 12'h70e;
        exp <= 18'h1dcf6;
        #1
        src0 <= 12'h540;
        src1 <= 12'h8ed;
        src2 <= 12'h9fe;
        src3 <= 12'h735;
        src4 <= 12'h2dd;
        src5 <= 12'h592;
        src6 <= 12'hdef;
        src7 <= 12'habf;
        src8 <= 12'hb58;
        src9 <= 12'hf8f;
        src10 <= 12'h64e;
        src11 <= 12'hb08;
        src12 <= 12'h3fe;
        src13 <= 12'h443;
        src14 <= 12'h873;
        src15 <= 12'hc5d;
        src16 <= 12'h55f;
        src17 <= 12'hf17;
        src18 <= 12'hce6;
        src19 <= 12'hf6;
        src20 <= 12'hfbf;
        src21 <= 12'h62b;
        src22 <= 12'h458;
        src23 <= 12'h7f0;
        src24 <= 12'hd9c;
        src25 <= 12'hbb3;
        src26 <= 12'h278;
        src27 <= 12'h5ec;
        src28 <= 12'h77f;
        src29 <= 12'h1d9;
        src30 <= 12'hb93;
        src31 <= 12'h995;
        src32 <= 12'hee5;
        src33 <= 12'hdb;
        src34 <= 12'h951;
        src35 <= 12'hacf;
        src36 <= 12'hf4d;
        src37 <= 12'h4ac;
        src38 <= 12'h570;
        src39 <= 12'h455;
        src40 <= 12'h7db;
        src41 <= 12'h203;
        src42 <= 12'hbb0;
        src43 <= 12'hd85;
        src44 <= 12'h76b;
        src45 <= 12'heb8;
        src46 <= 12'h4bc;
        src47 <= 12'h620;
        src48 <= 12'h1de;
        src49 <= 12'hbfb;
        src50 <= 12'hd34;
        src51 <= 12'h6c5;
        src52 <= 12'h721;
        src53 <= 12'hcf6;
        src54 <= 12'h214;
        src55 <= 12'h7b1;
        src56 <= 12'h210;
        src57 <= 12'he2f;
        src58 <= 12'h708;
        src59 <= 12'hd74;
        src60 <= 12'hce4;
        src61 <= 12'h6e2;
        src62 <= 12'hed0;
        src63 <= 12'h901;
        exp <= 18'h22432;
        #1
        src0 <= 12'he69;
        src1 <= 12'h64a;
        src2 <= 12'h772;
        src3 <= 12'h95f;
        src4 <= 12'haee;
        src5 <= 12'h1be;
        src6 <= 12'h327;
        src7 <= 12'h925;
        src8 <= 12'h654;
        src9 <= 12'h3c5;
        src10 <= 12'h16e;
        src11 <= 12'h292;
        src12 <= 12'h2a9;
        src13 <= 12'h790;
        src14 <= 12'h1a8;
        src15 <= 12'h65a;
        src16 <= 12'h2b;
        src17 <= 12'h46c;
        src18 <= 12'hfad;
        src19 <= 12'ha31;
        src20 <= 12'he6a;
        src21 <= 12'hfd7;
        src22 <= 12'h24;
        src23 <= 12'h456;
        src24 <= 12'h83a;
        src25 <= 12'h23e;
        src26 <= 12'h779;
        src27 <= 12'h481;
        src28 <= 12'h800;
        src29 <= 12'h3a1;
        src30 <= 12'he5a;
        src31 <= 12'h8dd;
        src32 <= 12'he48;
        src33 <= 12'hbdf;
        src34 <= 12'hd2c;
        src35 <= 12'h922;
        src36 <= 12'hd61;
        src37 <= 12'hdc6;
        src38 <= 12'hd5;
        src39 <= 12'h4c0;
        src40 <= 12'hd06;
        src41 <= 12'h4e3;
        src42 <= 12'ha25;
        src43 <= 12'h13;
        src44 <= 12'hc6d;
        src45 <= 12'hd5d;
        src46 <= 12'hc06;
        src47 <= 12'h1f2;
        src48 <= 12'h94f;
        src49 <= 12'h272;
        src50 <= 12'h4b7;
        src51 <= 12'h4e5;
        src52 <= 12'h99e;
        src53 <= 12'h345;
        src54 <= 12'he20;
        src55 <= 12'h625;
        src56 <= 12'ha52;
        src57 <= 12'ha41;
        src58 <= 12'h226;
        src59 <= 12'h5d6;
        src60 <= 12'h59c;
        src61 <= 12'hd15;
        src62 <= 12'h892;
        src63 <= 12'h85d;
        exp <= 18'h1e512;
        #1
        src0 <= 12'he62;
        src1 <= 12'hf5f;
        src2 <= 12'hb14;
        src3 <= 12'h24e;
        src4 <= 12'he48;
        src5 <= 12'h3b5;
        src6 <= 12'h1a7;
        src7 <= 12'h9ae;
        src8 <= 12'h705;
        src9 <= 12'h252;
        src10 <= 12'h221;
        src11 <= 12'h7d9;
        src12 <= 12'h630;
        src13 <= 12'hf33;
        src14 <= 12'h524;
        src15 <= 12'hbf5;
        src16 <= 12'h972;
        src17 <= 12'h559;
        src18 <= 12'h44;
        src19 <= 12'h2d0;
        src20 <= 12'h451;
        src21 <= 12'hcc8;
        src22 <= 12'h5e6;
        src23 <= 12'hd75;
        src24 <= 12'h58;
        src25 <= 12'h30e;
        src26 <= 12'hce1;
        src27 <= 12'h8db;
        src28 <= 12'h18d;
        src29 <= 12'hfca;
        src30 <= 12'h8df;
        src31 <= 12'hf66;
        src32 <= 12'hf40;
        src33 <= 12'h364;
        src34 <= 12'hb1b;
        src35 <= 12'h730;
        src36 <= 12'h48c;
        src37 <= 12'hf9f;
        src38 <= 12'h83c;
        src39 <= 12'hc07;
        src40 <= 12'h643;
        src41 <= 12'h38c;
        src42 <= 12'hd16;
        src43 <= 12'h5e2;
        src44 <= 12'h8f5;
        src45 <= 12'hc2;
        src46 <= 12'hce4;
        src47 <= 12'hfb4;
        src48 <= 12'h4a;
        src49 <= 12'hff3;
        src50 <= 12'hb7f;
        src51 <= 12'h6b;
        src52 <= 12'h540;
        src53 <= 12'hffd;
        src54 <= 12'hbe1;
        src55 <= 12'hdb6;
        src56 <= 12'ha94;
        src57 <= 12'hd1f;
        src58 <= 12'h6fc;
        src59 <= 12'haff;
        src60 <= 12'h7c3;
        src61 <= 12'hb13;
        src62 <= 12'h7a3;
        src63 <= 12'h808;
        exp <= 18'h222f0;
        #1
        src0 <= 12'h27f;
        src1 <= 12'hbfb;
        src2 <= 12'h637;
        src3 <= 12'h43a;
        src4 <= 12'h9e0;
        src5 <= 12'hd87;
        src6 <= 12'h456;
        src7 <= 12'h98d;
        src8 <= 12'h3f5;
        src9 <= 12'h198;
        src10 <= 12'h99f;
        src11 <= 12'h3fe;
        src12 <= 12'hdce;
        src13 <= 12'h4c6;
        src14 <= 12'h69f;
        src15 <= 12'hd55;
        src16 <= 12'he7e;
        src17 <= 12'h266;
        src18 <= 12'h6a7;
        src19 <= 12'h504;
        src20 <= 12'h9f5;
        src21 <= 12'h532;
        src22 <= 12'h156;
        src23 <= 12'h359;
        src24 <= 12'h676;
        src25 <= 12'h49c;
        src26 <= 12'h467;
        src27 <= 12'hea4;
        src28 <= 12'hfcb;
        src29 <= 12'hf41;
        src30 <= 12'h4d9;
        src31 <= 12'hc6d;
        src32 <= 12'h9dc;
        src33 <= 12'he0c;
        src34 <= 12'hea2;
        src35 <= 12'h8a8;
        src36 <= 12'h5c0;
        src37 <= 12'h534;
        src38 <= 12'h906;
        src39 <= 12'ha62;
        src40 <= 12'hcfe;
        src41 <= 12'h7c2;
        src42 <= 12'h9d9;
        src43 <= 12'hce4;
        src44 <= 12'hb87;
        src45 <= 12'hf6a;
        src46 <= 12'h45c;
        src47 <= 12'h980;
        src48 <= 12'h133;
        src49 <= 12'h2fd;
        src50 <= 12'hb07;
        src51 <= 12'h509;
        src52 <= 12'h149;
        src53 <= 12'h5da;
        src54 <= 12'hccf;
        src55 <= 12'h8a2;
        src56 <= 12'hf37;
        src57 <= 12'h924;
        src58 <= 12'h343;
        src59 <= 12'h2a0;
        src60 <= 12'h1a7;
        src61 <= 12'hcf8;
        src62 <= 12'h56a;
        src63 <= 12'hbe0;
        exp <= 18'h2078e;
        #1
        src0 <= 12'hc6d;
        src1 <= 12'h70c;
        src2 <= 12'h2b;
        src3 <= 12'h8;
        src4 <= 12'h30;
        src5 <= 12'h99f;
        src6 <= 12'h55f;
        src7 <= 12'h7d7;
        src8 <= 12'hd7d;
        src9 <= 12'h714;
        src10 <= 12'h69d;
        src11 <= 12'h6ee;
        src12 <= 12'hdd7;
        src13 <= 12'h4e5;
        src14 <= 12'h157;
        src15 <= 12'h20b;
        src16 <= 12'h45b;
        src17 <= 12'h126;
        src18 <= 12'h1dd;
        src19 <= 12'h891;
        src20 <= 12'h9e9;
        src21 <= 12'h787;
        src22 <= 12'hbaa;
        src23 <= 12'h721;
        src24 <= 12'h26b;
        src25 <= 12'h365;
        src26 <= 12'h60c;
        src27 <= 12'hee1;
        src28 <= 12'h346;
        src29 <= 12'h2a0;
        src30 <= 12'hd72;
        src31 <= 12'ha7e;
        src32 <= 12'ha5e;
        src33 <= 12'hcbc;
        src34 <= 12'h4c4;
        src35 <= 12'h216;
        src36 <= 12'h7b4;
        src37 <= 12'h6b6;
        src38 <= 12'hd6;
        src39 <= 12'hfe1;
        src40 <= 12'h54e;
        src41 <= 12'h66;
        src42 <= 12'h129;
        src43 <= 12'h518;
        src44 <= 12'ha66;
        src45 <= 12'he3d;
        src46 <= 12'hf81;
        src47 <= 12'heb2;
        src48 <= 12'hc99;
        src49 <= 12'h601;
        src50 <= 12'hd35;
        src51 <= 12'hd75;
        src52 <= 12'h432;
        src53 <= 12'h9cc;
        src54 <= 12'h70;
        src55 <= 12'h2b8;
        src56 <= 12'hfba;
        src57 <= 12'hccc;
        src58 <= 12'hc2;
        src59 <= 12'h6c4;
        src60 <= 12'hf9f;
        src61 <= 12'h48f;
        src62 <= 12'h9f;
        src63 <= 12'h743;
        exp <= 18'h1ce0e;
        #1
        src0 <= 12'h96f;
        src1 <= 12'h7d1;
        src2 <= 12'h967;
        src3 <= 12'h46c;
        src4 <= 12'ha64;
        src5 <= 12'h277;
        src6 <= 12'hb94;
        src7 <= 12'h799;
        src8 <= 12'hc69;
        src9 <= 12'h5bc;
        src10 <= 12'had1;
        src11 <= 12'h583;
        src12 <= 12'h45e;
        src13 <= 12'h9d9;
        src14 <= 12'hff1;
        src15 <= 12'h8ec;
        src16 <= 12'h7c8;
        src17 <= 12'h75d;
        src18 <= 12'h643;
        src19 <= 12'h4d9;
        src20 <= 12'h2ca;
        src21 <= 12'hc8d;
        src22 <= 12'h16d;
        src23 <= 12'h72;
        src24 <= 12'he45;
        src25 <= 12'hf9e;
        src26 <= 12'h712;
        src27 <= 12'h8e1;
        src28 <= 12'h272;
        src29 <= 12'h368;
        src30 <= 12'ha3b;
        src31 <= 12'h361;
        src32 <= 12'h977;
        src33 <= 12'hccc;
        src34 <= 12'h329;
        src35 <= 12'h5fb;
        src36 <= 12'h24f;
        src37 <= 12'h4c5;
        src38 <= 12'hce6;
        src39 <= 12'hd2f;
        src40 <= 12'ha49;
        src41 <= 12'h4c7;
        src42 <= 12'h38e;
        src43 <= 12'hfd1;
        src44 <= 12'hbcb;
        src45 <= 12'ha4f;
        src46 <= 12'hb5a;
        src47 <= 12'h9b6;
        src48 <= 12'h60e;
        src49 <= 12'h7d2;
        src50 <= 12'ha66;
        src51 <= 12'h57;
        src52 <= 12'hc93;
        src53 <= 12'hf39;
        src54 <= 12'hf5f;
        src55 <= 12'hda6;
        src56 <= 12'he59;
        src57 <= 12'hcf0;
        src58 <= 12'h24f;
        src59 <= 12'h822;
        src60 <= 12'h50c;
        src61 <= 12'ha69;
        src62 <= 12'hc2a;
        src63 <= 12'hd0;
        exp <= 18'h2172b;
        #1
        src0 <= 12'h4e9;
        src1 <= 12'h4b0;
        src2 <= 12'hb3d;
        src3 <= 12'h5d7;
        src4 <= 12'hf6d;
        src5 <= 12'hefd;
        src6 <= 12'hf07;
        src7 <= 12'ha32;
        src8 <= 12'h9d9;
        src9 <= 12'h1ee;
        src10 <= 12'h55;
        src11 <= 12'he48;
        src12 <= 12'h12e;
        src13 <= 12'hd6;
        src14 <= 12'hd94;
        src15 <= 12'h86a;
        src16 <= 12'hc01;
        src17 <= 12'hc04;
        src18 <= 12'hd2e;
        src19 <= 12'hf61;
        src20 <= 12'h602;
        src21 <= 12'h304;
        src22 <= 12'hab9;
        src23 <= 12'h845;
        src24 <= 12'h512;
        src25 <= 12'h445;
        src26 <= 12'h642;
        src27 <= 12'hd2d;
        src28 <= 12'hc4e;
        src29 <= 12'h50b;
        src30 <= 12'h3dc;
        src31 <= 12'hdaa;
        src32 <= 12'h562;
        src33 <= 12'h5f3;
        src34 <= 12'hdb5;
        src35 <= 12'hec;
        src36 <= 12'hee0;
        src37 <= 12'h2c7;
        src38 <= 12'h147;
        src39 <= 12'hd82;
        src40 <= 12'h799;
        src41 <= 12'h9f6;
        src42 <= 12'hb22;
        src43 <= 12'hb1e;
        src44 <= 12'ha9c;
        src45 <= 12'h7ee;
        src46 <= 12'hfcd;
        src47 <= 12'hecf;
        src48 <= 12'hb98;
        src49 <= 12'h62c;
        src50 <= 12'h8e7;
        src51 <= 12'h1dd;
        src52 <= 12'ha5a;
        src53 <= 12'hc3e;
        src54 <= 12'h975;
        src55 <= 12'hd3;
        src56 <= 12'h4bf;
        src57 <= 12'h68b;
        src58 <= 12'h302;
        src59 <= 12'h3e9;
        src60 <= 12'h700;
        src61 <= 12'h132;
        src62 <= 12'h843;
        src63 <= 12'h31e;
        exp <= 18'h20b7e;
        #1
        src0 <= 12'hdba;
        src1 <= 12'h7cb;
        src2 <= 12'h51;
        src3 <= 12'h21c;
        src4 <= 12'h6f1;
        src5 <= 12'ha8b;
        src6 <= 12'hdea;
        src7 <= 12'h289;
        src8 <= 12'h8fe;
        src9 <= 12'hede;
        src10 <= 12'h685;
        src11 <= 12'h653;
        src12 <= 12'h112;
        src13 <= 12'h428;
        src14 <= 12'h1e7;
        src15 <= 12'hd18;
        src16 <= 12'hdd2;
        src17 <= 12'hd4f;
        src18 <= 12'h9d;
        src19 <= 12'hf9f;
        src20 <= 12'he92;
        src21 <= 12'hc29;
        src22 <= 12'hda6;
        src23 <= 12'h6de;
        src24 <= 12'h7d4;
        src25 <= 12'h88;
        src26 <= 12'h7b6;
        src27 <= 12'h7a6;
        src28 <= 12'h2dc;
        src29 <= 12'hbed;
        src30 <= 12'haa6;
        src31 <= 12'hb0e;
        src32 <= 12'h964;
        src33 <= 12'h2db;
        src34 <= 12'hcba;
        src35 <= 12'hd7e;
        src36 <= 12'hdb0;
        src37 <= 12'hf97;
        src38 <= 12'he46;
        src39 <= 12'h9ca;
        src40 <= 12'h57e;
        src41 <= 12'hb59;
        src42 <= 12'h889;
        src43 <= 12'hf49;
        src44 <= 12'h235;
        src45 <= 12'h99a;
        src46 <= 12'hb38;
        src47 <= 12'hdb;
        src48 <= 12'h577;
        src49 <= 12'haca;
        src50 <= 12'haf;
        src51 <= 12'h1a6;
        src52 <= 12'hd23;
        src53 <= 12'h31b;
        src54 <= 12'h622;
        src55 <= 12'hf4a;
        src56 <= 12'h2a4;
        src57 <= 12'he98;
        src58 <= 12'hc9b;
        src59 <= 12'h168;
        src60 <= 12'he68;
        src61 <= 12'ha1c;
        src62 <= 12'h239;
        src63 <= 12'h7da;
        exp <= 18'h2200e;
        #1
        src0 <= 12'hd81;
        src1 <= 12'h49c;
        src2 <= 12'h6ff;
        src3 <= 12'he7f;
        src4 <= 12'he4f;
        src5 <= 12'hbff;
        src6 <= 12'h3b5;
        src7 <= 12'hfbf;
        src8 <= 12'h1d2;
        src9 <= 12'h78d;
        src10 <= 12'ha43;
        src11 <= 12'habb;
        src12 <= 12'hc5;
        src13 <= 12'hc47;
        src14 <= 12'hb34;
        src15 <= 12'hb14;
        src16 <= 12'h225;
        src17 <= 12'ha;
        src18 <= 12'h37f;
        src19 <= 12'hbb1;
        src20 <= 12'hfc7;
        src21 <= 12'h8f9;
        src22 <= 12'h89d;
        src23 <= 12'hf54;
        src24 <= 12'hbb6;
        src25 <= 12'hb8c;
        src26 <= 12'h1f6;
        src27 <= 12'h875;
        src28 <= 12'h17c;
        src29 <= 12'h62e;
        src30 <= 12'h51f;
        src31 <= 12'h715;
        src32 <= 12'h18d;
        src33 <= 12'hef0;
        src34 <= 12'h775;
        src35 <= 12'ha2a;
        src36 <= 12'h2fe;
        src37 <= 12'h3c0;
        src38 <= 12'h5fd;
        src39 <= 12'h49;
        src40 <= 12'hbe2;
        src41 <= 12'hb05;
        src42 <= 12'hff9;
        src43 <= 12'he44;
        src44 <= 12'h5;
        src45 <= 12'hd0;
        src46 <= 12'h38a;
        src47 <= 12'h444;
        src48 <= 12'h9f4;
        src49 <= 12'h20b;
        src50 <= 12'h290;
        src51 <= 12'hf84;
        src52 <= 12'h565;
        src53 <= 12'h9eb;
        src54 <= 12'h765;
        src55 <= 12'ha7f;
        src56 <= 12'h77c;
        src57 <= 12'h20c;
        src58 <= 12'h7e9;
        src59 <= 12'hdb;
        src60 <= 12'h53d;
        src61 <= 12'h47c;
        src62 <= 12'ha2;
        src63 <= 12'hfdf;
        exp <= 18'h1e75d;
        #1
        src0 <= 12'h79d;
        src1 <= 12'hbaa;
        src2 <= 12'he6;
        src3 <= 12'h4ee;
        src4 <= 12'he85;
        src5 <= 12'h1d3;
        src6 <= 12'h90d;
        src7 <= 12'ha8c;
        src8 <= 12'h8f5;
        src9 <= 12'hb83;
        src10 <= 12'h92a;
        src11 <= 12'h766;
        src12 <= 12'h514;
        src13 <= 12'hca6;
        src14 <= 12'h7ee;
        src15 <= 12'h8db;
        src16 <= 12'ha06;
        src17 <= 12'hc06;
        src18 <= 12'h73a;
        src19 <= 12'he8;
        src20 <= 12'h5af;
        src21 <= 12'h177;
        src22 <= 12'h2f2;
        src23 <= 12'hf34;
        src24 <= 12'h7b6;
        src25 <= 12'h94b;
        src26 <= 12'hdbb;
        src27 <= 12'hdb0;
        src28 <= 12'ha6;
        src29 <= 12'h83a;
        src30 <= 12'h7bc;
        src31 <= 12'he87;
        src32 <= 12'hf99;
        src33 <= 12'hfdf;
        src34 <= 12'h988;
        src35 <= 12'h827;
        src36 <= 12'hf3e;
        src37 <= 12'h377;
        src38 <= 12'h622;
        src39 <= 12'hdd8;
        src40 <= 12'h2df;
        src41 <= 12'h721;
        src42 <= 12'h776;
        src43 <= 12'h5af;
        src44 <= 12'hc3d;
        src45 <= 12'hfec;
        src46 <= 12'h66d;
        src47 <= 12'h54f;
        src48 <= 12'hf0d;
        src49 <= 12'hfae;
        src50 <= 12'hfc7;
        src51 <= 12'he71;
        src52 <= 12'hb6d;
        src53 <= 12'h510;
        src54 <= 12'he02;
        src55 <= 12'hb06;
        src56 <= 12'h83e;
        src57 <= 12'h6e3;
        src58 <= 12'hdc1;
        src59 <= 12'h725;
        src60 <= 12'hbdb;
        src61 <= 12'h93d;
        src62 <= 12'h9e0;
        src63 <= 12'hd2d;
        exp <= 18'h25524;
        #1
        src0 <= 12'hdd7;
        src1 <= 12'h380;
        src2 <= 12'h2b;
        src3 <= 12'h2ea;
        src4 <= 12'h828;
        src5 <= 12'hf65;
        src6 <= 12'he0;
        src7 <= 12'h221;
        src8 <= 12'h1cb;
        src9 <= 12'h646;
        src10 <= 12'h22b;
        src11 <= 12'h8c0;
        src12 <= 12'hc4d;
        src13 <= 12'h5f0;
        src14 <= 12'ha78;
        src15 <= 12'hdd2;
        src16 <= 12'h621;
        src17 <= 12'h226;
        src18 <= 12'h694;
        src19 <= 12'h2;
        src20 <= 12'h380;
        src21 <= 12'h5c4;
        src22 <= 12'h28d;
        src23 <= 12'h466;
        src24 <= 12'h8aa;
        src25 <= 12'hcbe;
        src26 <= 12'hb81;
        src27 <= 12'hee0;
        src28 <= 12'h31b;
        src29 <= 12'hcc8;
        src30 <= 12'hb90;
        src31 <= 12'h2ba;
        src32 <= 12'hfc7;
        src33 <= 12'h4b;
        src34 <= 12'h2a2;
        src35 <= 12'h11f;
        src36 <= 12'he01;
        src37 <= 12'hddc;
        src38 <= 12'hd4a;
        src39 <= 12'hd20;
        src40 <= 12'h6d3;
        src41 <= 12'h969;
        src42 <= 12'h131;
        src43 <= 12'he8f;
        src44 <= 12'hb7b;
        src45 <= 12'h2cb;
        src46 <= 12'h67d;
        src47 <= 12'h5c2;
        src48 <= 12'h789;
        src49 <= 12'he78;
        src50 <= 12'hcec;
        src51 <= 12'h18e;
        src52 <= 12'h612;
        src53 <= 12'ha0d;
        src54 <= 12'hd7b;
        src55 <= 12'hdf9;
        src56 <= 12'hef6;
        src57 <= 12'hd3d;
        src58 <= 12'h8d3;
        src59 <= 12'h1a8;
        src60 <= 12'hd1b;
        src61 <= 12'h3d4;
        src62 <= 12'hd67;
        src63 <= 12'h511;
        exp <= 18'h1f845;
        #1
        src0 <= 12'hcbd;
        src1 <= 12'h90c;
        src2 <= 12'he43;
        src3 <= 12'h4e3;
        src4 <= 12'h981;
        src5 <= 12'hf;
        src6 <= 12'hb18;
        src7 <= 12'h803;
        src8 <= 12'h20;
        src9 <= 12'h9f8;
        src10 <= 12'h8ce;
        src11 <= 12'h10a;
        src12 <= 12'hd73;
        src13 <= 12'h17e;
        src14 <= 12'h9ec;
        src15 <= 12'h59b;
        src16 <= 12'hf6e;
        src17 <= 12'ha5d;
        src18 <= 12'h430;
        src19 <= 12'h538;
        src20 <= 12'h743;
        src21 <= 12'hdb3;
        src22 <= 12'h24b;
        src23 <= 12'haf1;
        src24 <= 12'h5ec;
        src25 <= 12'h9b0;
        src26 <= 12'hdcd;
        src27 <= 12'hc07;
        src28 <= 12'h880;
        src29 <= 12'h445;
        src30 <= 12'hbab;
        src31 <= 12'h12e;
        src32 <= 12'ha37;
        src33 <= 12'hb60;
        src34 <= 12'h4f7;
        src35 <= 12'haae;
        src36 <= 12'he63;
        src37 <= 12'hb91;
        src38 <= 12'h515;
        src39 <= 12'hf3d;
        src40 <= 12'h890;
        src41 <= 12'h3;
        src42 <= 12'h9c9;
        src43 <= 12'h5e6;
        src44 <= 12'h562;
        src45 <= 12'h706;
        src46 <= 12'h702;
        src47 <= 12'h4c6;
        src48 <= 12'h915;
        src49 <= 12'h7da;
        src50 <= 12'h738;
        src51 <= 12'h273;
        src52 <= 12'h95e;
        src53 <= 12'hb72;
        src54 <= 12'h32d;
        src55 <= 12'h4a9;
        src56 <= 12'h43b;
        src57 <= 12'h937;
        src58 <= 12'h2ce;
        src59 <= 12'h190;
        src60 <= 12'he2b;
        src61 <= 12'h64f;
        src62 <= 12'h676;
        src63 <= 12'h519;
        exp <= 18'h1ed82;
        #1
        src0 <= 12'hf47;
        src1 <= 12'h97d;
        src2 <= 12'haad;
        src3 <= 12'h3e0;
        src4 <= 12'h757;
        src5 <= 12'h58b;
        src6 <= 12'h9d8;
        src7 <= 12'hcb7;
        src8 <= 12'h461;
        src9 <= 12'h879;
        src10 <= 12'h624;
        src11 <= 12'h3ce;
        src12 <= 12'h5db;
        src13 <= 12'h9a8;
        src14 <= 12'hbd8;
        src15 <= 12'h8d2;
        src16 <= 12'hb36;
        src17 <= 12'hb0a;
        src18 <= 12'h116;
        src19 <= 12'hf53;
        src20 <= 12'h78d;
        src21 <= 12'h228;
        src22 <= 12'h506;
        src23 <= 12'h4;
        src24 <= 12'hb15;
        src25 <= 12'h1ac;
        src26 <= 12'hcdc;
        src27 <= 12'h419;
        src28 <= 12'hff1;
        src29 <= 12'h63;
        src30 <= 12'h5bf;
        src31 <= 12'h39b;
        src32 <= 12'h6a8;
        src33 <= 12'h5b8;
        src34 <= 12'hc4e;
        src35 <= 12'h318;
        src36 <= 12'hf41;
        src37 <= 12'hda7;
        src38 <= 12'hf47;
        src39 <= 12'h262;
        src40 <= 12'hcc0;
        src41 <= 12'h734;
        src42 <= 12'h463;
        src43 <= 12'h3ae;
        src44 <= 12'h430;
        src45 <= 12'h843;
        src46 <= 12'h46d;
        src47 <= 12'hdbf;
        src48 <= 12'h3cc;
        src49 <= 12'hc10;
        src50 <= 12'h8ab;
        src51 <= 12'hb0;
        src52 <= 12'hd61;
        src53 <= 12'h666;
        src54 <= 12'h5e0;
        src55 <= 12'hefa;
        src56 <= 12'hefc;
        src57 <= 12'h933;
        src58 <= 12'h41d;
        src59 <= 12'h9b8;
        src60 <= 12'hede;
        src61 <= 12'h47c;
        src62 <= 12'hcf0;
        src63 <= 12'h5ee;
        exp <= 18'h20596;
        #1
        src0 <= 12'h145;
        src1 <= 12'h35c;
        src2 <= 12'hbb5;
        src3 <= 12'h1ed;
        src4 <= 12'haeb;
        src5 <= 12'ha0d;
        src6 <= 12'h415;
        src7 <= 12'h6c4;
        src8 <= 12'hfd9;
        src9 <= 12'hc7a;
        src10 <= 12'ha1e;
        src11 <= 12'ha15;
        src12 <= 12'h53;
        src13 <= 12'hdb7;
        src14 <= 12'ha40;
        src15 <= 12'h32e;
        src16 <= 12'h37b;
        src17 <= 12'hbbb;
        src18 <= 12'h92c;
        src19 <= 12'hfde;
        src20 <= 12'h2e7;
        src21 <= 12'hd33;
        src22 <= 12'h339;
        src23 <= 12'h496;
        src24 <= 12'hfe2;
        src25 <= 12'heb7;
        src26 <= 12'h2f2;
        src27 <= 12'heef;
        src28 <= 12'h1bf;
        src29 <= 12'hc17;
        src30 <= 12'h2da;
        src31 <= 12'h4aa;
        src32 <= 12'h627;
        src33 <= 12'h11f;
        src34 <= 12'h53f;
        src35 <= 12'hef3;
        src36 <= 12'ha9e;
        src37 <= 12'hef;
        src38 <= 12'h57c;
        src39 <= 12'hf98;
        src40 <= 12'haf4;
        src41 <= 12'hcad;
        src42 <= 12'ha18;
        src43 <= 12'h6f;
        src44 <= 12'h5f4;
        src45 <= 12'h825;
        src46 <= 12'h274;
        src47 <= 12'h12b;
        src48 <= 12'hff0;
        src49 <= 12'h147;
        src50 <= 12'h5fd;
        src51 <= 12'h812;
        src52 <= 12'h9d6;
        src53 <= 12'h7d9;
        src54 <= 12'hdb1;
        src55 <= 12'ha5d;
        src56 <= 12'h8a3;
        src57 <= 12'h635;
        src58 <= 12'h8a8;
        src59 <= 12'h12;
        src60 <= 12'h761;
        src61 <= 12'hb2d;
        src62 <= 12'h7f6;
        src63 <= 12'heeb;
        exp <= 18'h1fe0c;
        #1
        src0 <= 12'h6f1;
        src1 <= 12'hbfc;
        src2 <= 12'hd16;
        src3 <= 12'hea1;
        src4 <= 12'h659;
        src5 <= 12'h1b8;
        src6 <= 12'h9a5;
        src7 <= 12'hc5b;
        src8 <= 12'ha4b;
        src9 <= 12'h63a;
        src10 <= 12'h119;
        src11 <= 12'ha6d;
        src12 <= 12'hea0;
        src13 <= 12'h508;
        src14 <= 12'h5d;
        src15 <= 12'h9b8;
        src16 <= 12'h26b;
        src17 <= 12'h6c9;
        src18 <= 12'h5b9;
        src19 <= 12'hb0;
        src20 <= 12'h8ac;
        src21 <= 12'h590;
        src22 <= 12'hb9d;
        src23 <= 12'h507;
        src24 <= 12'h1bb;
        src25 <= 12'hc66;
        src26 <= 12'h37e;
        src27 <= 12'hfc2;
        src28 <= 12'h305;
        src29 <= 12'hb2a;
        src30 <= 12'h65c;
        src31 <= 12'h772;
        src32 <= 12'hd1;
        src33 <= 12'h82;
        src34 <= 12'ha4b;
        src35 <= 12'h8f9;
        src36 <= 12'ha10;
        src37 <= 12'heed;
        src38 <= 12'habe;
        src39 <= 12'h343;
        src40 <= 12'h761;
        src41 <= 12'hba5;
        src42 <= 12'hfb3;
        src43 <= 12'h233;
        src44 <= 12'h8a1;
        src45 <= 12'hf51;
        src46 <= 12'h4be;
        src47 <= 12'h50d;
        src48 <= 12'heb0;
        src49 <= 12'h5fd;
        src50 <= 12'hb31;
        src51 <= 12'hcb0;
        src52 <= 12'heb0;
        src53 <= 12'h793;
        src54 <= 12'h204;
        src55 <= 12'hc9f;
        src56 <= 12'hf1d;
        src57 <= 12'h622;
        src58 <= 12'h7ee;
        src59 <= 12'h169;
        src60 <= 12'h70e;
        src61 <= 12'h152;
        src62 <= 12'hfee;
        src63 <= 12'h50d;
        exp <= 18'h201fb;
        #1
        src0 <= 12'h111;
        src1 <= 12'h12b;
        src2 <= 12'h2d2;
        src3 <= 12'h5cd;
        src4 <= 12'hcd1;
        src5 <= 12'h907;
        src6 <= 12'hfb;
        src7 <= 12'h99;
        src8 <= 12'hf13;
        src9 <= 12'h197;
        src10 <= 12'ha10;
        src11 <= 12'h740;
        src12 <= 12'hc24;
        src13 <= 12'h940;
        src14 <= 12'he35;
        src15 <= 12'h269;
        src16 <= 12'h9c8;
        src17 <= 12'h2e1;
        src18 <= 12'h4d3;
        src19 <= 12'h1a8;
        src20 <= 12'h7de;
        src21 <= 12'h81b;
        src22 <= 12'hf23;
        src23 <= 12'he8b;
        src24 <= 12'hd73;
        src25 <= 12'h243;
        src26 <= 12'h23a;
        src27 <= 12'h168;
        src28 <= 12'hf88;
        src29 <= 12'h2c2;
        src30 <= 12'hf4;
        src31 <= 12'heb7;
        src32 <= 12'h44;
        src33 <= 12'h3f2;
        src34 <= 12'ha04;
        src35 <= 12'hb91;
        src36 <= 12'h2fd;
        src37 <= 12'h67c;
        src38 <= 12'ha97;
        src39 <= 12'hdde;
        src40 <= 12'h3ae;
        src41 <= 12'hb93;
        src42 <= 12'hbfb;
        src43 <= 12'h5d;
        src44 <= 12'he02;
        src45 <= 12'h20f;
        src46 <= 12'hf57;
        src47 <= 12'h792;
        src48 <= 12'h2c2;
        src49 <= 12'h500;
        src50 <= 12'h3d6;
        src51 <= 12'hf2e;
        src52 <= 12'h982;
        src53 <= 12'h7a9;
        src54 <= 12'hfd5;
        src55 <= 12'h197;
        src56 <= 12'heb9;
        src57 <= 12'ha1f;
        src58 <= 12'h394;
        src59 <= 12'hbed;
        src60 <= 12'h99;
        src61 <= 12'hbef;
        src62 <= 12'hff4;
        src63 <= 12'h325;
        exp <= 18'h1e3fe;
        #1
        src0 <= 12'hf64;
        src1 <= 12'h52a;
        src2 <= 12'he24;
        src3 <= 12'h3ca;
        src4 <= 12'h14b;
        src5 <= 12'h294;
        src6 <= 12'hd46;
        src7 <= 12'he2d;
        src8 <= 12'ha23;
        src9 <= 12'hae3;
        src10 <= 12'heea;
        src11 <= 12'h8fd;
        src12 <= 12'hd91;
        src13 <= 12'hdf1;
        src14 <= 12'hdaf;
        src15 <= 12'hbd9;
        src16 <= 12'h279;
        src17 <= 12'h31;
        src18 <= 12'h1ce;
        src19 <= 12'he18;
        src20 <= 12'hc16;
        src21 <= 12'hfb1;
        src22 <= 12'h97d;
        src23 <= 12'h708;
        src24 <= 12'hc49;
        src25 <= 12'h811;
        src26 <= 12'ha92;
        src27 <= 12'h155;
        src28 <= 12'h25f;
        src29 <= 12'h6b8;
        src30 <= 12'hbe3;
        src31 <= 12'hee5;
        src32 <= 12'h8f0;
        src33 <= 12'hcee;
        src34 <= 12'h354;
        src35 <= 12'ha14;
        src36 <= 12'hb10;
        src37 <= 12'h96;
        src38 <= 12'h754;
        src39 <= 12'h9d3;
        src40 <= 12'h2bc;
        src41 <= 12'h289;
        src42 <= 12'h286;
        src43 <= 12'h3ab;
        src44 <= 12'h59;
        src45 <= 12'h72d;
        src46 <= 12'h68f;
        src47 <= 12'hc5e;
        src48 <= 12'hd7c;
        src49 <= 12'hca2;
        src50 <= 12'h743;
        src51 <= 12'hce;
        src52 <= 12'h496;
        src53 <= 12'hdff;
        src54 <= 12'h919;
        src55 <= 12'ha53;
        src56 <= 12'hbe0;
        src57 <= 12'hc1c;
        src58 <= 12'ha12;
        src59 <= 12'h5d8;
        src60 <= 12'h9c1;
        src61 <= 12'hed3;
        src62 <= 12'hc59;
        src63 <= 12'h96e;
        exp <= 18'h22f2e;
        #1
        src0 <= 12'h473;
        src1 <= 12'h304;
        src2 <= 12'hb2a;
        src3 <= 12'h965;
        src4 <= 12'hdfb;
        src5 <= 12'he4a;
        src6 <= 12'haa6;
        src7 <= 12'ha4d;
        src8 <= 12'h7ba;
        src9 <= 12'h681;
        src10 <= 12'h530;
        src11 <= 12'h452;
        src12 <= 12'h16e;
        src13 <= 12'hd8b;
        src14 <= 12'hd8b;
        src15 <= 12'ha5d;
        src16 <= 12'hc01;
        src17 <= 12'h120;
        src18 <= 12'h29d;
        src19 <= 12'h65b;
        src20 <= 12'hb1a;
        src21 <= 12'hd6b;
        src22 <= 12'h72c;
        src23 <= 12'h147;
        src24 <= 12'hc8a;
        src25 <= 12'hc9;
        src26 <= 12'h705;
        src27 <= 12'h320;
        src28 <= 12'h9ea;
        src29 <= 12'h49f;
        src30 <= 12'h5eb;
        src31 <= 12'h9be;
        src32 <= 12'h385;
        src33 <= 12'h596;
        src34 <= 12'h875;
        src35 <= 12'h388;
        src36 <= 12'h375;
        src37 <= 12'hb39;
        src38 <= 12'h3f4;
        src39 <= 12'h3aa;
        src40 <= 12'hc88;
        src41 <= 12'he26;
        src42 <= 12'h240;
        src43 <= 12'hb0e;
        src44 <= 12'hac0;
        src45 <= 12'h5bb;
        src46 <= 12'h6cf;
        src47 <= 12'hf50;
        src48 <= 12'h43b;
        src49 <= 12'h737;
        src50 <= 12'h804;
        src51 <= 12'hb07;
        src52 <= 12'h8ca;
        src53 <= 12'h1f0;
        src54 <= 12'h4e1;
        src55 <= 12'h479;
        src56 <= 12'h242;
        src57 <= 12'h966;
        src58 <= 12'h922;
        src59 <= 12'h436;
        src60 <= 12'hdcc;
        src61 <= 12'h7c7;
        src62 <= 12'h897;
        src63 <= 12'h3d0;
        exp <= 18'h1e01c;
        #1
        src0 <= 12'hbdf;
        src1 <= 12'h93b;
        src2 <= 12'h411;
        src3 <= 12'h743;
        src4 <= 12'h8fb;
        src5 <= 12'h824;
        src6 <= 12'ha8e;
        src7 <= 12'hdf4;
        src8 <= 12'ha99;
        src9 <= 12'h165;
        src10 <= 12'hc91;
        src11 <= 12'h490;
        src12 <= 12'he8;
        src13 <= 12'hddc;
        src14 <= 12'h8a8;
        src15 <= 12'h94b;
        src16 <= 12'hf74;
        src17 <= 12'h362;
        src18 <= 12'h594;
        src19 <= 12'hd84;
        src20 <= 12'h7e5;
        src21 <= 12'hc78;
        src22 <= 12'h714;
        src23 <= 12'h4f3;
        src24 <= 12'h8af;
        src25 <= 12'haaf;
        src26 <= 12'h22;
        src27 <= 12'hb8a;
        src28 <= 12'h309;
        src29 <= 12'hef0;
        src30 <= 12'h164;
        src31 <= 12'h7ec;
        src32 <= 12'hcd0;
        src33 <= 12'h255;
        src34 <= 12'h5cd;
        src35 <= 12'he44;
        src36 <= 12'hab5;
        src37 <= 12'hb83;
        src38 <= 12'h859;
        src39 <= 12'ha37;
        src40 <= 12'he66;
        src41 <= 12'hf5c;
        src42 <= 12'h6f8;
        src43 <= 12'hd87;
        src44 <= 12'h82;
        src45 <= 12'h608;
        src46 <= 12'hb39;
        src47 <= 12'h4f9;
        src48 <= 12'h56b;
        src49 <= 12'hcf6;
        src50 <= 12'h712;
        src51 <= 12'he93;
        src52 <= 12'heef;
        src53 <= 12'he70;
        src54 <= 12'hc67;
        src55 <= 12'h156;
        src56 <= 12'h5d1;
        src57 <= 12'h5fa;
        src58 <= 12'hd8e;
        src59 <= 12'hf16;
        src60 <= 12'h37;
        src61 <= 12'h116;
        src62 <= 12'h89f;
        src63 <= 12'h44c;
        exp <= 18'h2274e;
        #1
        src0 <= 12'h662;
        src1 <= 12'h85b;
        src2 <= 12'h79f;
        src3 <= 12'hd37;
        src4 <= 12'hc23;
        src5 <= 12'h470;
        src6 <= 12'h9c;
        src7 <= 12'h5e1;
        src8 <= 12'h6ee;
        src9 <= 12'h1f;
        src10 <= 12'h589;
        src11 <= 12'h79c;
        src12 <= 12'hed;
        src13 <= 12'h958;
        src14 <= 12'hee1;
        src15 <= 12'h17e;
        src16 <= 12'hdd8;
        src17 <= 12'h548;
        src18 <= 12'h707;
        src19 <= 12'hd01;
        src20 <= 12'h4d8;
        src21 <= 12'h16a;
        src22 <= 12'hba8;
        src23 <= 12'hb70;
        src24 <= 12'hd6c;
        src25 <= 12'hd41;
        src26 <= 12'hf71;
        src27 <= 12'h489;
        src28 <= 12'h2f9;
        src29 <= 12'hedf;
        src30 <= 12'h6f6;
        src31 <= 12'hc60;
        src32 <= 12'h851;
        src33 <= 12'he14;
        src34 <= 12'hbe5;
        src35 <= 12'h251;
        src36 <= 12'hb2a;
        src37 <= 12'hf39;
        src38 <= 12'hd12;
        src39 <= 12'he5a;
        src40 <= 12'h5c5;
        src41 <= 12'hb1e;
        src42 <= 12'h2c0;
        src43 <= 12'ha0f;
        src44 <= 12'hb0b;
        src45 <= 12'h155;
        src46 <= 12'ha6;
        src47 <= 12'h649;
        src48 <= 12'hd19;
        src49 <= 12'h910;
        src50 <= 12'he69;
        src51 <= 12'h947;
        src52 <= 12'h964;
        src53 <= 12'h7a4;
        src54 <= 12'h421;
        src55 <= 12'h1a3;
        src56 <= 12'h765;
        src57 <= 12'h812;
        src58 <= 12'h9de;
        src59 <= 12'h385;
        src60 <= 12'hac3;
        src61 <= 12'h62c;
        src62 <= 12'h346;
        src63 <= 12'hc8d;
        exp <= 18'h20f7c;
        #1
        src0 <= 12'h815;
        src1 <= 12'h3fa;
        src2 <= 12'hc6a;
        src3 <= 12'h67d;
        src4 <= 12'h246;
        src5 <= 12'ha8b;
        src6 <= 12'h25e;
        src7 <= 12'h587;
        src8 <= 12'h3c7;
        src9 <= 12'h569;
        src10 <= 12'h4b4;
        src11 <= 12'hd15;
        src12 <= 12'hff1;
        src13 <= 12'h193;
        src14 <= 12'hea4;
        src15 <= 12'hfd8;
        src16 <= 12'h47f;
        src17 <= 12'h4e;
        src18 <= 12'h2f4;
        src19 <= 12'hc28;
        src20 <= 12'h6e6;
        src21 <= 12'h17;
        src22 <= 12'h13e;
        src23 <= 12'h5a4;
        src24 <= 12'h338;
        src25 <= 12'h2d7;
        src26 <= 12'hf78;
        src27 <= 12'h8f6;
        src28 <= 12'h2d8;
        src29 <= 12'h5d6;
        src30 <= 12'h9d3;
        src31 <= 12'h420;
        src32 <= 12'hac5;
        src33 <= 12'h78e;
        src34 <= 12'hb26;
        src35 <= 12'hbda;
        src36 <= 12'h3c9;
        src37 <= 12'h43e;
        src38 <= 12'h55b;
        src39 <= 12'h5cd;
        src40 <= 12'h2c0;
        src41 <= 12'h23d;
        src42 <= 12'hb16;
        src43 <= 12'h3b2;
        src44 <= 12'hfa8;
        src45 <= 12'hd31;
        src46 <= 12'hce8;
        src47 <= 12'h9ba;
        src48 <= 12'h928;
        src49 <= 12'h14c;
        src50 <= 12'h970;
        src51 <= 12'h743;
        src52 <= 12'h213;
        src53 <= 12'h2de;
        src54 <= 12'h141;
        src55 <= 12'h54c;
        src56 <= 12'hd2f;
        src57 <= 12'hdb1;
        src58 <= 12'hd98;
        src59 <= 12'he1d;
        src60 <= 12'h2d9;
        src61 <= 12'h1be;
        src62 <= 12'h630;
        src63 <= 12'h8ad;
        exp <= 18'h1c9fb;
        #1
        src0 <= 12'h1ea;
        src1 <= 12'h8ed;
        src2 <= 12'ha40;
        src3 <= 12'h5bd;
        src4 <= 12'h643;
        src5 <= 12'h8ca;
        src6 <= 12'h871;
        src7 <= 12'h17f;
        src8 <= 12'h67e;
        src9 <= 12'hdc8;
        src10 <= 12'h2bd;
        src11 <= 12'h31e;
        src12 <= 12'ha02;
        src13 <= 12'hc84;
        src14 <= 12'h7c2;
        src15 <= 12'h377;
        src16 <= 12'h176;
        src17 <= 12'h16;
        src18 <= 12'h4c7;
        src19 <= 12'hd8a;
        src20 <= 12'hbdd;
        src21 <= 12'h58c;
        src22 <= 12'ha64;
        src23 <= 12'h4ae;
        src24 <= 12'heb6;
        src25 <= 12'hfc1;
        src26 <= 12'h818;
        src27 <= 12'h8d6;
        src28 <= 12'h4d4;
        src29 <= 12'h200;
        src30 <= 12'h750;
        src31 <= 12'h96a;
        src32 <= 12'hc85;
        src33 <= 12'h484;
        src34 <= 12'h5c4;
        src35 <= 12'h4ea;
        src36 <= 12'h6a3;
        src37 <= 12'h5ad;
        src38 <= 12'h1d1;
        src39 <= 12'ha09;
        src40 <= 12'hc5f;
        src41 <= 12'hbb0;
        src42 <= 12'h31a;
        src43 <= 12'h8bd;
        src44 <= 12'he82;
        src45 <= 12'h9c7;
        src46 <= 12'h2d1;
        src47 <= 12'h2a0;
        src48 <= 12'h26d;
        src49 <= 12'h7a4;
        src50 <= 12'hf78;
        src51 <= 12'hbdb;
        src52 <= 12'ha37;
        src53 <= 12'hb1a;
        src54 <= 12'h1e7;
        src55 <= 12'h70d;
        src56 <= 12'h4ca;
        src57 <= 12'h5a0;
        src58 <= 12'h1c2;
        src59 <= 12'h41;
        src60 <= 12'h524;
        src61 <= 12'hd3a;
        src62 <= 12'hd05;
        src63 <= 12'hdaa;
        exp <= 18'h1dda0;
        #1
        src0 <= 12'h2e0;
        src1 <= 12'hadf;
        src2 <= 12'h970;
        src3 <= 12'hf46;
        src4 <= 12'he7e;
        src5 <= 12'hf0d;
        src6 <= 12'haed;
        src7 <= 12'hdf0;
        src8 <= 12'h5b4;
        src9 <= 12'hb0b;
        src10 <= 12'h3f;
        src11 <= 12'hc38;
        src12 <= 12'hcf0;
        src13 <= 12'hfa0;
        src14 <= 12'h2a4;
        src15 <= 12'hd58;
        src16 <= 12'h284;
        src17 <= 12'ha7e;
        src18 <= 12'hbdc;
        src19 <= 12'h2c7;
        src20 <= 12'h27c;
        src21 <= 12'h12b;
        src22 <= 12'hdb9;
        src23 <= 12'h103;
        src24 <= 12'h409;
        src25 <= 12'ha10;
        src26 <= 12'h372;
        src27 <= 12'hcb3;
        src28 <= 12'h879;
        src29 <= 12'h5c1;
        src30 <= 12'h2a2;
        src31 <= 12'h784;
        src32 <= 12'h141;
        src33 <= 12'h5c3;
        src34 <= 12'hfc5;
        src35 <= 12'h7e7;
        src36 <= 12'h66a;
        src37 <= 12'hc32;
        src38 <= 12'hca8;
        src39 <= 12'he76;
        src40 <= 12'h481;
        src41 <= 12'h589;
        src42 <= 12'ha36;
        src43 <= 12'hce5;
        src44 <= 12'hf1e;
        src45 <= 12'h45e;
        src46 <= 12'h3cf;
        src47 <= 12'h475;
        src48 <= 12'hda2;
        src49 <= 12'h9c0;
        src50 <= 12'hce9;
        src51 <= 12'ha0c;
        src52 <= 12'hdd9;
        src53 <= 12'h82c;
        src54 <= 12'hd03;
        src55 <= 12'he30;
        src56 <= 12'h6d9;
        src57 <= 12'hb19;
        src58 <= 12'h970;
        src59 <= 12'h122;
        src60 <= 12'hcb7;
        src61 <= 12'h7cc;
        src62 <= 12'h4aa;
        src63 <= 12'h84;
        exp <= 18'h22a58;
        #1
        src0 <= 12'hfd;
        src1 <= 12'hc7b;
        src2 <= 12'h529;
        src3 <= 12'h4d1;
        src4 <= 12'hbb2;
        src5 <= 12'ha59;
        src6 <= 12'he84;
        src7 <= 12'h918;
        src8 <= 12'hb7a;
        src9 <= 12'h4a;
        src10 <= 12'h99e;
        src11 <= 12'h4b6;
        src12 <= 12'h56b;
        src13 <= 12'hd88;
        src14 <= 12'he04;
        src15 <= 12'h289;
        src16 <= 12'h4d1;
        src17 <= 12'hc72;
        src18 <= 12'hc71;
        src19 <= 12'h993;
        src20 <= 12'hf61;
        src21 <= 12'h5fa;
        src22 <= 12'h6ac;
        src23 <= 12'h6dc;
        src24 <= 12'hda6;
        src25 <= 12'h990;
        src26 <= 12'h253;
        src27 <= 12'h60;
        src28 <= 12'h527;
        src29 <= 12'h600;
        src30 <= 12'he1;
        src31 <= 12'h6ab;
        src32 <= 12'h46e;
        src33 <= 12'h9f5;
        src34 <= 12'h179;
        src35 <= 12'h590;
        src36 <= 12'h697;
        src37 <= 12'h124;
        src38 <= 12'hc8;
        src39 <= 12'h27d;
        src40 <= 12'h234;
        src41 <= 12'h949;
        src42 <= 12'h2e9;
        src43 <= 12'he9b;
        src44 <= 12'he59;
        src45 <= 12'hfe7;
        src46 <= 12'hc70;
        src47 <= 12'h68d;
        src48 <= 12'h6bd;
        src49 <= 12'hcf3;
        src50 <= 12'h845;
        src51 <= 12'h328;
        src52 <= 12'h5a;
        src53 <= 12'h36;
        src54 <= 12'h9ce;
        src55 <= 12'haf7;
        src56 <= 12'h2bb;
        src57 <= 12'h151;
        src58 <= 12'h757;
        src59 <= 12'h944;
        src60 <= 12'hd2e;
        src61 <= 12'h288;
        src62 <= 12'h827;
        src63 <= 12'h1b4;
        exp <= 18'h1cacb;
        #1
        src0 <= 12'haa6;
        src1 <= 12'hefa;
        src2 <= 12'h8e7;
        src3 <= 12'h525;
        src4 <= 12'hb6a;
        src5 <= 12'h363;
        src6 <= 12'h3e9;
        src7 <= 12'h1f3;
        src8 <= 12'ha7f;
        src9 <= 12'he7a;
        src10 <= 12'h16b;
        src11 <= 12'h564;
        src12 <= 12'hef5;
        src13 <= 12'h955;
        src14 <= 12'h62e;
        src15 <= 12'h28d;
        src16 <= 12'h8c0;
        src17 <= 12'h434;
        src18 <= 12'h79;
        src19 <= 12'h8db;
        src20 <= 12'hd43;
        src21 <= 12'h41d;
        src22 <= 12'ha61;
        src23 <= 12'hdcd;
        src24 <= 12'h99c;
        src25 <= 12'h294;
        src26 <= 12'h79b;
        src27 <= 12'hdb8;
        src28 <= 12'h9b0;
        src29 <= 12'h2b1;
        src30 <= 12'he57;
        src31 <= 12'h850;
        src32 <= 12'hcd6;
        src33 <= 12'h89e;
        src34 <= 12'hb0c;
        src35 <= 12'h1ec;
        src36 <= 12'heb0;
        src37 <= 12'hb23;
        src38 <= 12'hfbf;
        src39 <= 12'h293;
        src40 <= 12'hf16;
        src41 <= 12'haef;
        src42 <= 12'hf4b;
        src43 <= 12'h5ce;
        src44 <= 12'hfd9;
        src45 <= 12'h445;
        src46 <= 12'hf52;
        src47 <= 12'h8e9;
        src48 <= 12'h7a4;
        src49 <= 12'hb62;
        src50 <= 12'he1c;
        src51 <= 12'h223;
        src52 <= 12'hbcf;
        src53 <= 12'h191;
        src54 <= 12'h164;
        src55 <= 12'hb72;
        src56 <= 12'hbfd;
        src57 <= 12'hae2;
        src58 <= 12'hc57;
        src59 <= 12'hb50;
        src60 <= 12'h8d9;
        src61 <= 12'h2eb;
        src62 <= 12'h764;
        src63 <= 12'hfe8;
        exp <= 18'h23a9c;
        #1
        src0 <= 12'h5b1;
        src1 <= 12'h9f1;
        src2 <= 12'h879;
        src3 <= 12'h901;
        src4 <= 12'h2ad;
        src5 <= 12'h911;
        src6 <= 12'h52;
        src7 <= 12'h7f4;
        src8 <= 12'h52f;
        src9 <= 12'h230;
        src10 <= 12'hb4;
        src11 <= 12'h856;
        src12 <= 12'h4b2;
        src13 <= 12'ha76;
        src14 <= 12'h75;
        src15 <= 12'h8f9;
        src16 <= 12'h720;
        src17 <= 12'hfeb;
        src18 <= 12'h89;
        src19 <= 12'h6e3;
        src20 <= 12'he4e;
        src21 <= 12'h71e;
        src22 <= 12'hf87;
        src23 <= 12'h35a;
        src24 <= 12'h103;
        src25 <= 12'hc08;
        src26 <= 12'hf9e;
        src27 <= 12'h3e3;
        src28 <= 12'h3f2;
        src29 <= 12'h10f;
        src30 <= 12'h9ee;
        src31 <= 12'h8eb;
        src32 <= 12'h8f9;
        src33 <= 12'h4ba;
        src34 <= 12'h1f1;
        src35 <= 12'h691;
        src36 <= 12'h421;
        src37 <= 12'hc12;
        src38 <= 12'h3dc;
        src39 <= 12'hfcb;
        src40 <= 12'ha2c;
        src41 <= 12'h211;
        src42 <= 12'h677;
        src43 <= 12'h462;
        src44 <= 12'h1e6;
        src45 <= 12'h174;
        src46 <= 12'h8b1;
        src47 <= 12'h3e3;
        src48 <= 12'h281;
        src49 <= 12'hfe3;
        src50 <= 12'hd8e;
        src51 <= 12'h2e8;
        src52 <= 12'heb4;
        src53 <= 12'h50b;
        src54 <= 12'hca3;
        src55 <= 12'ha77;
        src56 <= 12'h74d;
        src57 <= 12'h59e;
        src58 <= 12'h14f;
        src59 <= 12'h10;
        src60 <= 12'hcc0;
        src61 <= 12'h6cd;
        src62 <= 12'h7b8;
        src63 <= 12'hd2f;
        exp <= 18'h1c2cd;
        #1
        src0 <= 12'hd79;
        src1 <= 12'h352;
        src2 <= 12'hacd;
        src3 <= 12'h16c;
        src4 <= 12'hf6f;
        src5 <= 12'h736;
        src6 <= 12'h49e;
        src7 <= 12'heff;
        src8 <= 12'h9d1;
        src9 <= 12'h7ef;
        src10 <= 12'hba5;
        src11 <= 12'hcf0;
        src12 <= 12'haba;
        src13 <= 12'h2da;
        src14 <= 12'h20b;
        src15 <= 12'h6e;
        src16 <= 12'h64e;
        src17 <= 12'hedc;
        src18 <= 12'ha5a;
        src19 <= 12'hce3;
        src20 <= 12'h58d;
        src21 <= 12'h851;
        src22 <= 12'h9a0;
        src23 <= 12'h854;
        src24 <= 12'h6b3;
        src25 <= 12'h798;
        src26 <= 12'he99;
        src27 <= 12'ha68;
        src28 <= 12'hce8;
        src29 <= 12'h2f3;
        src30 <= 12'h8ce;
        src31 <= 12'hd31;
        src32 <= 12'hd8e;
        src33 <= 12'haa0;
        src34 <= 12'h7d2;
        src35 <= 12'h470;
        src36 <= 12'h285;
        src37 <= 12'hbe7;
        src38 <= 12'hc7f;
        src39 <= 12'hd57;
        src40 <= 12'h317;
        src41 <= 12'hd51;
        src42 <= 12'h617;
        src43 <= 12'hc9c;
        src44 <= 12'hb75;
        src45 <= 12'hc80;
        src46 <= 12'h20f;
        src47 <= 12'h1a4;
        src48 <= 12'hfc2;
        src49 <= 12'hd5;
        src50 <= 12'h965;
        src51 <= 12'h143;
        src52 <= 12'hdb5;
        src53 <= 12'h8e3;
        src54 <= 12'he55;
        src55 <= 12'hf7;
        src56 <= 12'h5f5;
        src57 <= 12'he3c;
        src58 <= 12'h180;
        src59 <= 12'hd5a;
        src60 <= 12'h81f;
        src61 <= 12'h91e;
        src62 <= 12'h2b9;
        src63 <= 12'h98;
        exp <= 18'h21f38;
        #1
        src0 <= 12'h7ea;
        src1 <= 12'ha4e;
        src2 <= 12'hb03;
        src3 <= 12'h695;
        src4 <= 12'hf10;
        src5 <= 12'h21a;
        src6 <= 12'h6bb;
        src7 <= 12'h7da;
        src8 <= 12'hb0c;
        src9 <= 12'hea3;
        src10 <= 12'ha42;
        src11 <= 12'hbac;
        src12 <= 12'h340;
        src13 <= 12'hb75;
        src14 <= 12'h498;
        src15 <= 12'hc98;
        src16 <= 12'h78e;
        src17 <= 12'h34d;
        src18 <= 12'h6e1;
        src19 <= 12'h90;
        src20 <= 12'hf13;
        src21 <= 12'h4b6;
        src22 <= 12'hf22;
        src23 <= 12'h310;
        src24 <= 12'hbfa;
        src25 <= 12'he7e;
        src26 <= 12'hf43;
        src27 <= 12'hcd;
        src28 <= 12'hbdf;
        src29 <= 12'h99b;
        src30 <= 12'ha79;
        src31 <= 12'h8b2;
        src32 <= 12'hd81;
        src33 <= 12'h2f7;
        src34 <= 12'h9e4;
        src35 <= 12'h1e1;
        src36 <= 12'hcf;
        src37 <= 12'hc2;
        src38 <= 12'hc87;
        src39 <= 12'h272;
        src40 <= 12'h217;
        src41 <= 12'h510;
        src42 <= 12'hb5f;
        src43 <= 12'h237;
        src44 <= 12'h86e;
        src45 <= 12'h53;
        src46 <= 12'h77b;
        src47 <= 12'h65c;
        src48 <= 12'h3f9;
        src49 <= 12'ha47;
        src50 <= 12'h850;
        src51 <= 12'hcc0;
        src52 <= 12'ha6c;
        src53 <= 12'hdcb;
        src54 <= 12'hced;
        src55 <= 12'hc36;
        src56 <= 12'h650;
        src57 <= 12'h7fc;
        src58 <= 12'hee6;
        src59 <= 12'hc0d;
        src60 <= 12'h6e3;
        src61 <= 12'hb6e;
        src62 <= 12'h97d;
        src63 <= 12'ha1d;
        exp <= 18'h21a75;
        #1
        src0 <= 12'h3e;
        src1 <= 12'hdf5;
        src2 <= 12'he2c;
        src3 <= 12'hcce;
        src4 <= 12'h7d9;
        src5 <= 12'hcf3;
        src6 <= 12'hc1d;
        src7 <= 12'h780;
        src8 <= 12'h5fa;
        src9 <= 12'h928;
        src10 <= 12'h7c5;
        src11 <= 12'h81f;
        src12 <= 12'hd03;
        src13 <= 12'h3cb;
        src14 <= 12'h5ca;
        src15 <= 12'h34;
        src16 <= 12'h8c0;
        src17 <= 12'h458;
        src18 <= 12'h630;
        src19 <= 12'h2b4;
        src20 <= 12'h62e;
        src21 <= 12'h83e;
        src22 <= 12'ha30;
        src23 <= 12'h713;
        src24 <= 12'h50c;
        src25 <= 12'h93a;
        src26 <= 12'h63d;
        src27 <= 12'h78d;
        src28 <= 12'he41;
        src29 <= 12'hcf9;
        src30 <= 12'hd48;
        src31 <= 12'h27a;
        src32 <= 12'h505;
        src33 <= 12'hfdb;
        src34 <= 12'hea0;
        src35 <= 12'hb0a;
        src36 <= 12'hd3e;
        src37 <= 12'h9e9;
        src38 <= 12'h52c;
        src39 <= 12'he05;
        src40 <= 12'h96f;
        src41 <= 12'hfe8;
        src42 <= 12'h9a8;
        src43 <= 12'h806;
        src44 <= 12'ha1d;
        src45 <= 12'hea3;
        src46 <= 12'hd28;
        src47 <= 12'h706;
        src48 <= 12'h489;
        src49 <= 12'h4f3;
        src50 <= 12'h24e;
        src51 <= 12'h1e1;
        src52 <= 12'he43;
        src53 <= 12'had6;
        src54 <= 12'hf14;
        src55 <= 12'hc23;
        src56 <= 12'h3b4;
        src57 <= 12'h62d;
        src58 <= 12'h821;
        src59 <= 12'haed;
        src60 <= 12'h519;
        src61 <= 12'hbe;
        src62 <= 12'hf8d;
        src63 <= 12'h74b;
        exp <= 18'h2308d;
        #1
        src0 <= 12'h78b;
        src1 <= 12'h950;
        src2 <= 12'hcae;
        src3 <= 12'h649;
        src4 <= 12'hae6;
        src5 <= 12'hff6;
        src6 <= 12'h9ef;
        src7 <= 12'h580;
        src8 <= 12'hbf4;
        src9 <= 12'h59f;
        src10 <= 12'h767;
        src11 <= 12'h634;
        src12 <= 12'h466;
        src13 <= 12'h39d;
        src14 <= 12'h284;
        src15 <= 12'h657;
        src16 <= 12'h8bf;
        src17 <= 12'h157;
        src18 <= 12'h932;
        src19 <= 12'h76;
        src20 <= 12'h8af;
        src21 <= 12'he4b;
        src22 <= 12'hf6b;
        src23 <= 12'h481;
        src24 <= 12'h92f;
        src25 <= 12'hb4f;
        src26 <= 12'hf98;
        src27 <= 12'he6a;
        src28 <= 12'hc29;
        src29 <= 12'h5ba;
        src30 <= 12'hfb;
        src31 <= 12'hbfe;
        src32 <= 12'hed3;
        src33 <= 12'h2;
        src34 <= 12'h99d;
        src35 <= 12'h472;
        src36 <= 12'hd85;
        src37 <= 12'hbef;
        src38 <= 12'hfb6;
        src39 <= 12'hd6e;
        src40 <= 12'h481;
        src41 <= 12'h42b;
        src42 <= 12'ha1;
        src43 <= 12'hc42;
        src44 <= 12'hc84;
        src45 <= 12'ha98;
        src46 <= 12'h955;
        src47 <= 12'h8aa;
        src48 <= 12'h39d;
        src49 <= 12'h779;
        src50 <= 12'h8cd;
        src51 <= 12'hb06;
        src52 <= 12'hc66;
        src53 <= 12'hf30;
        src54 <= 12'hc9;
        src55 <= 12'h24f;
        src56 <= 12'h4a;
        src57 <= 12'hf57;
        src58 <= 12'he2e;
        src59 <= 12'ha29;
        src60 <= 12'h8ce;
        src61 <= 12'hb95;
        src62 <= 12'he22;
        src63 <= 12'hc6c;
        exp <= 18'h234cf;
        #1
        src0 <= 12'h4ec;
        src1 <= 12'hf94;
        src2 <= 12'h15a;
        src3 <= 12'he1e;
        src4 <= 12'hbb9;
        src5 <= 12'h521;
        src6 <= 12'h3cc;
        src7 <= 12'h8b;
        src8 <= 12'hf2a;
        src9 <= 12'hd05;
        src10 <= 12'h310;
        src11 <= 12'hec3;
        src12 <= 12'h759;
        src13 <= 12'hb9f;
        src14 <= 12'ha1f;
        src15 <= 12'hd99;
        src16 <= 12'h305;
        src17 <= 12'ha4e;
        src18 <= 12'hd9c;
        src19 <= 12'hfed;
        src20 <= 12'hfe9;
        src21 <= 12'h7e;
        src22 <= 12'hce8;
        src23 <= 12'h84d;
        src24 <= 12'h318;
        src25 <= 12'h589;
        src26 <= 12'h61d;
        src27 <= 12'h432;
        src28 <= 12'h3c1;
        src29 <= 12'h8d9;
        src30 <= 12'h839;
        src31 <= 12'h685;
        src32 <= 12'h8b6;
        src33 <= 12'hf7b;
        src34 <= 12'h330;
        src35 <= 12'h475;
        src36 <= 12'h860;
        src37 <= 12'h359;
        src38 <= 12'h1c;
        src39 <= 12'heb3;
        src40 <= 12'h83e;
        src41 <= 12'h244;
        src42 <= 12'hb1;
        src43 <= 12'h9aa;
        src44 <= 12'he83;
        src45 <= 12'h81f;
        src46 <= 12'h445;
        src47 <= 12'ha15;
        src48 <= 12'h266;
        src49 <= 12'h39e;
        src50 <= 12'hd2f;
        src51 <= 12'h91e;
        src52 <= 12'h852;
        src53 <= 12'hfc9;
        src54 <= 12'hb6c;
        src55 <= 12'h2f2;
        src56 <= 12'hc77;
        src57 <= 12'he1d;
        src58 <= 12'h986;
        src59 <= 12'h60c;
        src60 <= 12'h8db;
        src61 <= 12'hd99;
        src62 <= 12'hc1;
        src63 <= 12'h7a8;
        exp <= 18'h2109f;
        #1
        src0 <= 12'h425;
        src1 <= 12'h9f3;
        src2 <= 12'hf67;
        src3 <= 12'h996;
        src4 <= 12'h4e6;
        src5 <= 12'hdd7;
        src6 <= 12'hdad;
        src7 <= 12'hc6b;
        src8 <= 12'h40b;
        src9 <= 12'h8aa;
        src10 <= 12'hc86;
        src11 <= 12'h8e6;
        src12 <= 12'h5fe;
        src13 <= 12'hdd4;
        src14 <= 12'hf99;
        src15 <= 12'h34e;
        src16 <= 12'h8fd;
        src17 <= 12'h162;
        src18 <= 12'h69c;
        src19 <= 12'ha20;
        src20 <= 12'h39e;
        src21 <= 12'hfa9;
        src22 <= 12'hc40;
        src23 <= 12'hee7;
        src24 <= 12'hd97;
        src25 <= 12'h99f;
        src26 <= 12'h3b8;
        src27 <= 12'h2e8;
        src28 <= 12'hed3;
        src29 <= 12'hd36;
        src30 <= 12'h3c4;
        src31 <= 12'h26e;
        src32 <= 12'h3c2;
        src33 <= 12'h3b0;
        src34 <= 12'h352;
        src35 <= 12'hfa7;
        src36 <= 12'hd2a;
        src37 <= 12'hc9c;
        src38 <= 12'hc71;
        src39 <= 12'hc24;
        src40 <= 12'ha80;
        src41 <= 12'h9d3;
        src42 <= 12'h52;
        src43 <= 12'hdda;
        src44 <= 12'h398;
        src45 <= 12'h318;
        src46 <= 12'hd5e;
        src47 <= 12'h38c;
        src48 <= 12'h684;
        src49 <= 12'hdce;
        src50 <= 12'h35e;
        src51 <= 12'hfaf;
        src52 <= 12'h4ef;
        src53 <= 12'h7d2;
        src54 <= 12'h404;
        src55 <= 12'h22c;
        src56 <= 12'h734;
        src57 <= 12'h4f3;
        src58 <= 12'he75;
        src59 <= 12'hd91;
        src60 <= 12'h7cd;
        src61 <= 12'hd9a;
        src62 <= 12'h104;
        src63 <= 12'h2a;
        exp <= 18'h2264f;
        #1
        src0 <= 12'hb51;
        src1 <= 12'he56;
        src2 <= 12'h8cd;
        src3 <= 12'h640;
        src4 <= 12'h106;
        src5 <= 12'h29e;
        src6 <= 12'hcd5;
        src7 <= 12'h357;
        src8 <= 12'h923;
        src9 <= 12'h49;
        src10 <= 12'h30;
        src11 <= 12'h6c2;
        src12 <= 12'hd74;
        src13 <= 12'h3ff;
        src14 <= 12'h48;
        src15 <= 12'he0;
        src16 <= 12'h60d;
        src17 <= 12'h190;
        src18 <= 12'he7a;
        src19 <= 12'h2e7;
        src20 <= 12'h223;
        src21 <= 12'h78c;
        src22 <= 12'h924;
        src23 <= 12'h507;
        src24 <= 12'h7a1;
        src25 <= 12'ha06;
        src26 <= 12'h389;
        src27 <= 12'hdab;
        src28 <= 12'hfe4;
        src29 <= 12'hc6;
        src30 <= 12'h70a;
        src31 <= 12'hc99;
        src32 <= 12'hbf7;
        src33 <= 12'h273;
        src34 <= 12'h81f;
        src35 <= 12'ha9;
        src36 <= 12'h14;
        src37 <= 12'hed5;
        src38 <= 12'h724;
        src39 <= 12'haf3;
        src40 <= 12'h4e3;
        src41 <= 12'hf43;
        src42 <= 12'h7b3;
        src43 <= 12'h9d8;
        src44 <= 12'h65e;
        src45 <= 12'hebb;
        src46 <= 12'hdf7;
        src47 <= 12'h4d;
        src48 <= 12'hfcc;
        src49 <= 12'h8ad;
        src50 <= 12'h4af;
        src51 <= 12'hfcc;
        src52 <= 12'h813;
        src53 <= 12'h7ca;
        src54 <= 12'h2f6;
        src55 <= 12'h19e;
        src56 <= 12'hd45;
        src57 <= 12'h25c;
        src58 <= 12'h247;
        src59 <= 12'h41;
        src60 <= 12'h3e8;
        src61 <= 12'h215;
        src62 <= 12'hc62;
        src63 <= 12'h926;
        exp <= 18'h1c7d0;
        #1
        src0 <= 12'hcbc;
        src1 <= 12'hf56;
        src2 <= 12'h101;
        src3 <= 12'h6aa;
        src4 <= 12'h674;
        src5 <= 12'hb07;
        src6 <= 12'hb38;
        src7 <= 12'h49c;
        src8 <= 12'h78d;
        src9 <= 12'he9a;
        src10 <= 12'h26e;
        src11 <= 12'hd08;
        src12 <= 12'h10e;
        src13 <= 12'h167;
        src14 <= 12'h685;
        src15 <= 12'hff9;
        src16 <= 12'hc6f;
        src17 <= 12'h32a;
        src18 <= 12'hce4;
        src19 <= 12'h3d9;
        src20 <= 12'h757;
        src21 <= 12'h36f;
        src22 <= 12'h254;
        src23 <= 12'hf2d;
        src24 <= 12'had2;
        src25 <= 12'h7f5;
        src26 <= 12'h4b;
        src27 <= 12'hd9;
        src28 <= 12'h754;
        src29 <= 12'h84;
        src30 <= 12'h7e1;
        src31 <= 12'hb4f;
        src32 <= 12'hb00;
        src33 <= 12'ha6c;
        src34 <= 12'he44;
        src35 <= 12'h298;
        src36 <= 12'h2f8;
        src37 <= 12'h2f;
        src38 <= 12'h15;
        src39 <= 12'h430;
        src40 <= 12'h595;
        src41 <= 12'hee3;
        src42 <= 12'hadb;
        src43 <= 12'he4;
        src44 <= 12'hb5f;
        src45 <= 12'hfd4;
        src46 <= 12'he14;
        src47 <= 12'h9e8;
        src48 <= 12'hde0;
        src49 <= 12'h6f0;
        src50 <= 12'h30a;
        src51 <= 12'h5e5;
        src52 <= 12'h66;
        src53 <= 12'hb1a;
        src54 <= 12'h2e4;
        src55 <= 12'h629;
        src56 <= 12'h297;
        src57 <= 12'h4a8;
        src58 <= 12'heeb;
        src59 <= 12'hecd;
        src60 <= 12'he37;
        src61 <= 12'h7bf;
        src62 <= 12'h841;
        src63 <= 12'h768;
        exp <= 18'h1ed28;
        #1
        src0 <= 12'h42c;
        src1 <= 12'hd55;
        src2 <= 12'hfb8;
        src3 <= 12'h59e;
        src4 <= 12'hc2d;
        src5 <= 12'hcd4;
        src6 <= 12'h346;
        src7 <= 12'hee6;
        src8 <= 12'h49;
        src9 <= 12'h3c;
        src10 <= 12'h99e;
        src11 <= 12'h1c7;
        src12 <= 12'h188;
        src13 <= 12'h3e3;
        src14 <= 12'h41e;
        src15 <= 12'h946;
        src16 <= 12'h5b8;
        src17 <= 12'hcf9;
        src18 <= 12'h7ac;
        src19 <= 12'h5d8;
        src20 <= 12'h32c;
        src21 <= 12'hb90;
        src22 <= 12'h1ce;
        src23 <= 12'h509;
        src24 <= 12'he75;
        src25 <= 12'hd60;
        src26 <= 12'h14e;
        src27 <= 12'hae8;
        src28 <= 12'hca6;
        src29 <= 12'he9;
        src30 <= 12'h880;
        src31 <= 12'h83f;
        src32 <= 12'h53e;
        src33 <= 12'h424;
        src34 <= 12'hb69;
        src35 <= 12'hbc8;
        src36 <= 12'h4e5;
        src37 <= 12'h73;
        src38 <= 12'h5b6;
        src39 <= 12'hc50;
        src40 <= 12'h83d;
        src41 <= 12'h179;
        src42 <= 12'h46a;
        src43 <= 12'hb58;
        src44 <= 12'h2cb;
        src45 <= 12'h517;
        src46 <= 12'he0a;
        src47 <= 12'h56b;
        src48 <= 12'h28f;
        src49 <= 12'h7ad;
        src50 <= 12'hd0;
        src51 <= 12'h659;
        src52 <= 12'h9b7;
        src53 <= 12'h93e;
        src54 <= 12'hca;
        src55 <= 12'h6b5;
        src56 <= 12'he84;
        src57 <= 12'h2bd;
        src58 <= 12'h3b;
        src59 <= 12'h756;
        src60 <= 12'hfa5;
        src61 <= 12'hcd8;
        src62 <= 12'h580;
        src63 <= 12'h308;
        exp <= 18'h1c34e;
        #1
        src0 <= 12'ha88;
        src1 <= 12'h41;
        src2 <= 12'hd91;
        src3 <= 12'he92;
        src4 <= 12'h8c1;
        src5 <= 12'h7e5;
        src6 <= 12'h830;
        src7 <= 12'h40f;
        src8 <= 12'h4c6;
        src9 <= 12'h8f5;
        src10 <= 12'hcb1;
        src11 <= 12'hbbd;
        src12 <= 12'h337;
        src13 <= 12'hb11;
        src14 <= 12'h4fb;
        src15 <= 12'h298;
        src16 <= 12'h72e;
        src17 <= 12'h241;
        src18 <= 12'h275;
        src19 <= 12'h630;
        src20 <= 12'h9f2;
        src21 <= 12'hf9;
        src22 <= 12'h2eb;
        src23 <= 12'hb87;
        src24 <= 12'h142;
        src25 <= 12'ha93;
        src26 <= 12'h335;
        src27 <= 12'hf69;
        src28 <= 12'h478;
        src29 <= 12'hbb3;
        src30 <= 12'h7ef;
        src31 <= 12'hf43;
        src32 <= 12'hc62;
        src33 <= 12'h919;
        src34 <= 12'hc96;
        src35 <= 12'he04;
        src36 <= 12'hda3;
        src37 <= 12'h1e7;
        src38 <= 12'ha59;
        src39 <= 12'h93c;
        src40 <= 12'h1c9;
        src41 <= 12'h1af;
        src42 <= 12'h7eb;
        src43 <= 12'h734;
        src44 <= 12'h9ff;
        src45 <= 12'h6f9;
        src46 <= 12'he60;
        src47 <= 12'hdc7;
        src48 <= 12'h99d;
        src49 <= 12'h867;
        src50 <= 12'h3c9;
        src51 <= 12'h3f7;
        src52 <= 12'h5e7;
        src53 <= 12'h45b;
        src54 <= 12'hbc7;
        src55 <= 12'h63e;
        src56 <= 12'h801;
        src57 <= 12'h1d2;
        src58 <= 12'hdaf;
        src59 <= 12'h6a;
        src60 <= 12'h89a;
        src61 <= 12'h44c;
        src62 <= 12'ha3a;
        src63 <= 12'h92;
        exp <= 18'h1e9a9;
        #1
        src0 <= 12'hac7;
        src1 <= 12'h88d;
        src2 <= 12'hb3d;
        src3 <= 12'h8cc;
        src4 <= 12'hfca;
        src5 <= 12'hdb0;
        src6 <= 12'hd7c;
        src7 <= 12'h9db;
        src8 <= 12'hbc5;
        src9 <= 12'hd8b;
        src10 <= 12'h7e6;
        src11 <= 12'h442;
        src12 <= 12'h7b9;
        src13 <= 12'hdfe;
        src14 <= 12'h20a;
        src15 <= 12'h9ab;
        src16 <= 12'h592;
        src17 <= 12'h2d;
        src18 <= 12'h69d;
        src19 <= 12'hd3b;
        src20 <= 12'hda1;
        src21 <= 12'h5ab;
        src22 <= 12'h688;
        src23 <= 12'hdde;
        src24 <= 12'h53c;
        src25 <= 12'h6d2;
        src26 <= 12'h871;
        src27 <= 12'hfd1;
        src28 <= 12'h4f4;
        src29 <= 12'hf65;
        src30 <= 12'h636;
        src31 <= 12'h40f;
        src32 <= 12'hb65;
        src33 <= 12'h9a7;
        src34 <= 12'h5a6;
        src35 <= 12'hbf4;
        src36 <= 12'head;
        src37 <= 12'h571;
        src38 <= 12'h428;
        src39 <= 12'hfb3;
        src40 <= 12'h2f7;
        src41 <= 12'hc4f;
        src42 <= 12'h433;
        src43 <= 12'h3ce;
        src44 <= 12'h5b0;
        src45 <= 12'h542;
        src46 <= 12'heaf;
        src47 <= 12'h68;
        src48 <= 12'h4ea;
        src49 <= 12'ha21;
        src50 <= 12'h58d;
        src51 <= 12'h246;
        src52 <= 12'h995;
        src53 <= 12'hdd3;
        src54 <= 12'hf69;
        src55 <= 12'ha60;
        src56 <= 12'h702;
        src57 <= 12'h814;
        src58 <= 12'hd9d;
        src59 <= 12'h4e3;
        src60 <= 12'h3a;
        src61 <= 12'hb63;
        src62 <= 12'hdee;
        src63 <= 12'h42c;
        exp <= 18'h22e94;
        #1
        src0 <= 12'h71c;
        src1 <= 12'hd2c;
        src2 <= 12'hec0;
        src3 <= 12'h346;
        src4 <= 12'h5b4;
        src5 <= 12'hd26;
        src6 <= 12'h44e;
        src7 <= 12'h603;
        src8 <= 12'h20b;
        src9 <= 12'h4bd;
        src10 <= 12'hb3b;
        src11 <= 12'h17d;
        src12 <= 12'hf60;
        src13 <= 12'h987;
        src14 <= 12'hae2;
        src15 <= 12'h465;
        src16 <= 12'h919;
        src17 <= 12'hd59;
        src18 <= 12'h387;
        src19 <= 12'hc03;
        src20 <= 12'h3fe;
        src21 <= 12'h8b8;
        src22 <= 12'h698;
        src23 <= 12'h632;
        src24 <= 12'h824;
        src25 <= 12'h841;
        src26 <= 12'hc46;
        src27 <= 12'hb0c;
        src28 <= 12'h888;
        src29 <= 12'hb51;
        src30 <= 12'hd3c;
        src31 <= 12'h546;
        src32 <= 12'h42c;
        src33 <= 12'h6e7;
        src34 <= 12'he69;
        src35 <= 12'h3b2;
        src36 <= 12'hcf9;
        src37 <= 12'h271;
        src38 <= 12'hb36;
        src39 <= 12'h876;
        src40 <= 12'h87c;
        src41 <= 12'h34a;
        src42 <= 12'hed;
        src43 <= 12'h574;
        src44 <= 12'hcf5;
        src45 <= 12'h703;
        src46 <= 12'h19f;
        src47 <= 12'hf3a;
        src48 <= 12'h2b6;
        src49 <= 12'h41c;
        src50 <= 12'hee4;
        src51 <= 12'h32e;
        src52 <= 12'he70;
        src53 <= 12'h659;
        src54 <= 12'h56a;
        src55 <= 12'h54d;
        src56 <= 12'hd07;
        src57 <= 12'h326;
        src58 <= 12'h905;
        src59 <= 12'h39;
        src60 <= 12'h5ea;
        src61 <= 12'h66f;
        src62 <= 12'hb94;
        src63 <= 12'hfd2;
        exp <= 18'h1fd7f;
        #1
        src0 <= 12'h29e;
        src1 <= 12'hc39;
        src2 <= 12'h1d8;
        src3 <= 12'ha3;
        src4 <= 12'ha25;
        src5 <= 12'hda5;
        src6 <= 12'h388;
        src7 <= 12'h6e7;
        src8 <= 12'h3cd;
        src9 <= 12'ha0;
        src10 <= 12'h331;
        src11 <= 12'h176;
        src12 <= 12'h34f;
        src13 <= 12'h886;
        src14 <= 12'h2de;
        src15 <= 12'h549;
        src16 <= 12'ha07;
        src17 <= 12'h714;
        src18 <= 12'he40;
        src19 <= 12'h7e6;
        src20 <= 12'hcf7;
        src21 <= 12'h670;
        src22 <= 12'h238;
        src23 <= 12'h2d2;
        src24 <= 12'h1f6;
        src25 <= 12'h70d;
        src26 <= 12'h8c7;
        src27 <= 12'h707;
        src28 <= 12'h69e;
        src29 <= 12'h232;
        src30 <= 12'h821;
        src31 <= 12'haff;
        src32 <= 12'h85c;
        src33 <= 12'ha96;
        src34 <= 12'h8b2;
        src35 <= 12'h8c5;
        src36 <= 12'h3cc;
        src37 <= 12'h245;
        src38 <= 12'h576;
        src39 <= 12'h911;
        src40 <= 12'h954;
        src41 <= 12'hb6f;
        src42 <= 12'h4e0;
        src43 <= 12'h39f;
        src44 <= 12'h2dd;
        src45 <= 12'h9f0;
        src46 <= 12'ha14;
        src47 <= 12'h70e;
        src48 <= 12'hd41;
        src49 <= 12'hefd;
        src50 <= 12'h5dc;
        src51 <= 12'h869;
        src52 <= 12'hd31;
        src53 <= 12'h940;
        src54 <= 12'ha8b;
        src55 <= 12'hbaa;
        src56 <= 12'h137;
        src57 <= 12'ha33;
        src58 <= 12'h5c9;
        src59 <= 12'h22e;
        src60 <= 12'hdd9;
        src61 <= 12'h96;
        src62 <= 12'hb63;
        src63 <= 12'h6fc;
        exp <= 18'h1c498;
        #1
        src0 <= 12'h3f9;
        src1 <= 12'h47a;
        src2 <= 12'hdc9;
        src3 <= 12'h7a1;
        src4 <= 12'hff1;
        src5 <= 12'h7bc;
        src6 <= 12'h307;
        src7 <= 12'ha80;
        src8 <= 12'h4cd;
        src9 <= 12'hd72;
        src10 <= 12'hdab;
        src11 <= 12'hbc4;
        src12 <= 12'hb78;
        src13 <= 12'h220;
        src14 <= 12'h443;
        src15 <= 12'h5d7;
        src16 <= 12'h2bd;
        src17 <= 12'he;
        src18 <= 12'h40e;
        src19 <= 12'hd88;
        src20 <= 12'h7d3;
        src21 <= 12'hf89;
        src22 <= 12'h9cd;
        src23 <= 12'hc25;
        src24 <= 12'hc6a;
        src25 <= 12'h1ed;
        src26 <= 12'h140;
        src27 <= 12'h4a9;
        src28 <= 12'h5a7;
        src29 <= 12'h6df;
        src30 <= 12'h6df;
        src31 <= 12'ha5;
        src32 <= 12'h2fc;
        src33 <= 12'hfe;
        src34 <= 12'h600;
        src35 <= 12'h72f;
        src36 <= 12'h882;
        src37 <= 12'h490;
        src38 <= 12'hc16;
        src39 <= 12'hcc;
        src40 <= 12'h65e;
        src41 <= 12'h470;
        src42 <= 12'h6a9;
        src43 <= 12'h373;
        src44 <= 12'hbaa;
        src45 <= 12'he61;
        src46 <= 12'h1ea;
        src47 <= 12'h396;
        src48 <= 12'h58e;
        src49 <= 12'hb8a;
        src50 <= 12'hef2;
        src51 <= 12'h87e;
        src52 <= 12'h80c;
        src53 <= 12'h62e;
        src54 <= 12'ha1e;
        src55 <= 12'hb1f;
        src56 <= 12'ha49;
        src57 <= 12'h663;
        src58 <= 12'h545;
        src59 <= 12'hc7;
        src60 <= 12'he9d;
        src61 <= 12'h187;
        src62 <= 12'h5ad;
        src63 <= 12'hdec;
        exp <= 18'h1d670;
        #1
        src0 <= 12'h91c;
        src1 <= 12'h1c9;
        src2 <= 12'h1e0;
        src3 <= 12'hb8f;
        src4 <= 12'h502;
        src5 <= 12'hb57;
        src6 <= 12'h5c2;
        src7 <= 12'heb;
        src8 <= 12'h526;
        src9 <= 12'h6d;
        src10 <= 12'hd47;
        src11 <= 12'h261;
        src12 <= 12'h3bd;
        src13 <= 12'h854;
        src14 <= 12'h109;
        src15 <= 12'h31a;
        src16 <= 12'h623;
        src17 <= 12'haac;
        src18 <= 12'hb44;
        src19 <= 12'h48d;
        src20 <= 12'h155;
        src21 <= 12'hc4d;
        src22 <= 12'h9c2;
        src23 <= 12'hf77;
        src24 <= 12'hb45;
        src25 <= 12'h31d;
        src26 <= 12'hd5e;
        src27 <= 12'hedf;
        src28 <= 12'h959;
        src29 <= 12'he27;
        src30 <= 12'h523;
        src31 <= 12'h8ef;
        src32 <= 12'he29;
        src33 <= 12'hf35;
        src34 <= 12'h1b3;
        src35 <= 12'h592;
        src36 <= 12'h2e2;
        src37 <= 12'hf56;
        src38 <= 12'hbfc;
        src39 <= 12'h98a;
        src40 <= 12'ha56;
        src41 <= 12'he6a;
        src42 <= 12'ha67;
        src43 <= 12'h333;
        src44 <= 12'h21e;
        src45 <= 12'ha9b;
        src46 <= 12'hcf2;
        src47 <= 12'h23c;
        src48 <= 12'hd09;
        src49 <= 12'h379;
        src50 <= 12'hdf8;
        src51 <= 12'h2f;
        src52 <= 12'he3e;
        src53 <= 12'h873;
        src54 <= 12'h566;
        src55 <= 12'h60a;
        src56 <= 12'h8aa;
        src57 <= 12'hd0e;
        src58 <= 12'h63f;
        src59 <= 12'h303;
        src60 <= 12'h97a;
        src61 <= 12'h2d0;
        src62 <= 12'h356;
        src63 <= 12'h516;
        exp <= 18'h1ef91;
        #1
        src0 <= 12'hc45;
        src1 <= 12'h25a;
        src2 <= 12'hba8;
        src3 <= 12'hf6f;
        src4 <= 12'hab8;
        src5 <= 12'h15d;
        src6 <= 12'h693;
        src7 <= 12'h1e1;
        src8 <= 12'hd56;
        src9 <= 12'h139;
        src10 <= 12'hcb0;
        src11 <= 12'h3e5;
        src12 <= 12'he80;
        src13 <= 12'h634;
        src14 <= 12'h778;
        src15 <= 12'h43e;
        src16 <= 12'h7ba;
        src17 <= 12'h16b;
        src18 <= 12'h6f0;
        src19 <= 12'hb8c;
        src20 <= 12'hd8b;
        src21 <= 12'h8a4;
        src22 <= 12'h33a;
        src23 <= 12'h3e5;
        src24 <= 12'hb3f;
        src25 <= 12'he5e;
        src26 <= 12'h829;
        src27 <= 12'h9c5;
        src28 <= 12'hd7;
        src29 <= 12'h38;
        src30 <= 12'hda2;
        src31 <= 12'hc2c;
        src32 <= 12'h3bb;
        src33 <= 12'hecb;
        src34 <= 12'h98d;
        src35 <= 12'ha2;
        src36 <= 12'h8d4;
        src37 <= 12'h705;
        src38 <= 12'he66;
        src39 <= 12'h547;
        src40 <= 12'h9ca;
        src41 <= 12'hc66;
        src42 <= 12'hc16;
        src43 <= 12'hb8b;
        src44 <= 12'h898;
        src45 <= 12'h275;
        src46 <= 12'hfd5;
        src47 <= 12'hb65;
        src48 <= 12'h219;
        src49 <= 12'h413;
        src50 <= 12'h58d;
        src51 <= 12'h829;
        src52 <= 12'h37b;
        src53 <= 12'h36b;
        src54 <= 12'hb57;
        src55 <= 12'h8e9;
        src56 <= 12'h12;
        src57 <= 12'h668;
        src58 <= 12'h9e0;
        src59 <= 12'h356;
        src60 <= 12'ha2e;
        src61 <= 12'hcb2;
        src62 <= 12'hfa4;
        src63 <= 12'h303;
        exp <= 18'h1fdb6;
        #1
        src0 <= 12'h156;
        src1 <= 12'h958;
        src2 <= 12'hcd6;
        src3 <= 12'ha9c;
        src4 <= 12'h731;
        src5 <= 12'h37;
        src6 <= 12'h63;
        src7 <= 12'hcff;
        src8 <= 12'h337;
        src9 <= 12'h68f;
        src10 <= 12'h86e;
        src11 <= 12'ha4b;
        src12 <= 12'h430;
        src13 <= 12'h8a4;
        src14 <= 12'h397;
        src15 <= 12'hd8a;
        src16 <= 12'h669;
        src17 <= 12'hd45;
        src18 <= 12'h16;
        src19 <= 12'h26d;
        src20 <= 12'hef6;
        src21 <= 12'h67a;
        src22 <= 12'h60;
        src23 <= 12'haee;
        src24 <= 12'hb5;
        src25 <= 12'h385;
        src26 <= 12'h70c;
        src27 <= 12'h6b3;
        src28 <= 12'he7c;
        src29 <= 12'he11;
        src30 <= 12'haf2;
        src31 <= 12'he1e;
        src32 <= 12'haf4;
        src33 <= 12'h41f;
        src34 <= 12'hb2f;
        src35 <= 12'h312;
        src36 <= 12'heb6;
        src37 <= 12'hac9;
        src38 <= 12'h5d6;
        src39 <= 12'h9da;
        src40 <= 12'h8a4;
        src41 <= 12'h756;
        src42 <= 12'h3ec;
        src43 <= 12'h944;
        src44 <= 12'h58d;
        src45 <= 12'hc3b;
        src46 <= 12'h24c;
        src47 <= 12'hc;
        src48 <= 12'h64e;
        src49 <= 12'hc8;
        src50 <= 12'h9e;
        src51 <= 12'hb54;
        src52 <= 12'hd19;
        src53 <= 12'h153;
        src54 <= 12'hf82;
        src55 <= 12'h901;
        src56 <= 12'h3e5;
        src57 <= 12'h3f8;
        src58 <= 12'h850;
        src59 <= 12'hd98;
        src60 <= 12'h7e;
        src61 <= 12'h82d;
        src62 <= 12'h5d3;
        src63 <= 12'h591;
        exp <= 18'h1d37b;
        #1
        src0 <= 12'h9be;
        src1 <= 12'h1c1;
        src2 <= 12'h973;
        src3 <= 12'h316;
        src4 <= 12'h49c;
        src5 <= 12'h2a2;
        src6 <= 12'h65;
        src7 <= 12'h6bf;
        src8 <= 12'h91c;
        src9 <= 12'h956;
        src10 <= 12'hf09;
        src11 <= 12'h1f7;
        src12 <= 12'h35d;
        src13 <= 12'h8c6;
        src14 <= 12'h781;
        src15 <= 12'h939;
        src16 <= 12'hc4b;
        src17 <= 12'hf3;
        src18 <= 12'h22d;
        src19 <= 12'h37c;
        src20 <= 12'h926;
        src21 <= 12'h319;
        src22 <= 12'h4b8;
        src23 <= 12'h91f;
        src24 <= 12'h293;
        src25 <= 12'hba1;
        src26 <= 12'h321;
        src27 <= 12'hc91;
        src28 <= 12'h968;
        src29 <= 12'h9db;
        src30 <= 12'h6f6;
        src31 <= 12'hb7;
        src32 <= 12'h2d5;
        src33 <= 12'h130;
        src34 <= 12'hb51;
        src35 <= 12'hca9;
        src36 <= 12'h661;
        src37 <= 12'hdd1;
        src38 <= 12'h993;
        src39 <= 12'hc75;
        src40 <= 12'h2a9;
        src41 <= 12'hdc9;
        src42 <= 12'hdfb;
        src43 <= 12'h520;
        src44 <= 12'h9f7;
        src45 <= 12'ha04;
        src46 <= 12'h909;
        src47 <= 12'h44b;
        src48 <= 12'hd2f;
        src49 <= 12'hcaa;
        src50 <= 12'haee;
        src51 <= 12'he8;
        src52 <= 12'hae9;
        src53 <= 12'h8d0;
        src54 <= 12'h205;
        src55 <= 12'h399;
        src56 <= 12'hfe3;
        src57 <= 12'h6ec;
        src58 <= 12'h315;
        src59 <= 12'hbd0;
        src60 <= 12'hd87;
        src61 <= 12'h3b8;
        src62 <= 12'h730;
        src63 <= 12'h514;
        exp <= 18'h1d9de;
        #1
        src0 <= 12'h9f4;
        src1 <= 12'h66a;
        src2 <= 12'hec2;
        src3 <= 12'ha7b;
        src4 <= 12'h528;
        src5 <= 12'hd65;
        src6 <= 12'hae6;
        src7 <= 12'hbb;
        src8 <= 12'haa6;
        src9 <= 12'h686;
        src10 <= 12'h57d;
        src11 <= 12'h3b;
        src12 <= 12'h140;
        src13 <= 12'h1d;
        src14 <= 12'h1b2;
        src15 <= 12'h1ae;
        src16 <= 12'h909;
        src17 <= 12'h379;
        src18 <= 12'he06;
        src19 <= 12'h2a;
        src20 <= 12'he83;
        src21 <= 12'h24c;
        src22 <= 12'h2fb;
        src23 <= 12'hfce;
        src24 <= 12'h11b;
        src25 <= 12'h691;
        src26 <= 12'hf4a;
        src27 <= 12'h875;
        src28 <= 12'he68;
        src29 <= 12'hc8c;
        src30 <= 12'he9b;
        src31 <= 12'h1d3;
        src32 <= 12'h4f8;
        src33 <= 12'h6f9;
        src34 <= 12'hfc9;
        src35 <= 12'h903;
        src36 <= 12'he9b;
        src37 <= 12'h936;
        src38 <= 12'h4d;
        src39 <= 12'hbab;
        src40 <= 12'h901;
        src41 <= 12'he15;
        src42 <= 12'hb3e;
        src43 <= 12'h2cc;
        src44 <= 12'h9;
        src45 <= 12'he7b;
        src46 <= 12'h4e5;
        src47 <= 12'h78a;
        src48 <= 12'h91f;
        src49 <= 12'h294;
        src50 <= 12'h922;
        src51 <= 12'hf59;
        src52 <= 12'hacc;
        src53 <= 12'h297;
        src54 <= 12'ha6c;
        src55 <= 12'h9f6;
        src56 <= 12'h992;
        src57 <= 12'hf4e;
        src58 <= 12'h5f2;
        src59 <= 12'hca;
        src60 <= 12'h555;
        src61 <= 12'h1a3;
        src62 <= 12'hea5;
        src63 <= 12'hc10;
        exp <= 18'h1fc56;
        #1
        src0 <= 12'hd35;
        src1 <= 12'h88f;
        src2 <= 12'hfb7;
        src3 <= 12'h748;
        src4 <= 12'hd25;
        src5 <= 12'h374;
        src6 <= 12'ha70;
        src7 <= 12'h70e;
        src8 <= 12'hf46;
        src9 <= 12'h17e;
        src10 <= 12'h470;
        src11 <= 12'h7a2;
        src12 <= 12'hb5b;
        src13 <= 12'h11f;
        src14 <= 12'h4ed;
        src15 <= 12'h5c3;
        src16 <= 12'h903;
        src17 <= 12'h897;
        src18 <= 12'hf7b;
        src19 <= 12'h9e6;
        src20 <= 12'hc06;
        src21 <= 12'h744;
        src22 <= 12'h3d7;
        src23 <= 12'h4a5;
        src24 <= 12'hfba;
        src25 <= 12'hbf3;
        src26 <= 12'h261;
        src27 <= 12'h839;
        src28 <= 12'he26;
        src29 <= 12'hb36;
        src30 <= 12'ha54;
        src31 <= 12'hf37;
        src32 <= 12'h92c;
        src33 <= 12'h3bb;
        src34 <= 12'he9c;
        src35 <= 12'h673;
        src36 <= 12'hf5b;
        src37 <= 12'h974;
        src38 <= 12'h933;
        src39 <= 12'h4e0;
        src40 <= 12'hbbe;
        src41 <= 12'h8b5;
        src42 <= 12'h73a;
        src43 <= 12'hc07;
        src44 <= 12'h34c;
        src45 <= 12'hf3c;
        src46 <= 12'hb7a;
        src47 <= 12'h302;
        src48 <= 12'h9d3;
        src49 <= 12'h696;
        src50 <= 12'hcd3;
        src51 <= 12'h51e;
        src52 <= 12'hfb6;
        src53 <= 12'h7c7;
        src54 <= 12'hd4;
        src55 <= 12'hf13;
        src56 <= 12'hdca;
        src57 <= 12'hc11;
        src58 <= 12'hed1;
        src59 <= 12'h295;
        src60 <= 12'h444;
        src61 <= 12'h1f;
        src62 <= 12'h246;
        src63 <= 12'hb52;
        exp <= 18'h23b53;
        #1
        src0 <= 12'h692;
        src1 <= 12'hfb5;
        src2 <= 12'h960;
        src3 <= 12'h87;
        src4 <= 12'hed2;
        src5 <= 12'hea2;
        src6 <= 12'hf46;
        src7 <= 12'h211;
        src8 <= 12'haa0;
        src9 <= 12'hf7a;
        src10 <= 12'hbdc;
        src11 <= 12'h52b;
        src12 <= 12'h11a;
        src13 <= 12'h937;
        src14 <= 12'h57b;
        src15 <= 12'h80;
        src16 <= 12'h7fc;
        src17 <= 12'h69e;
        src18 <= 12'ha5a;
        src19 <= 12'h975;
        src20 <= 12'h7b5;
        src21 <= 12'h23b;
        src22 <= 12'hd91;
        src23 <= 12'ha7e;
        src24 <= 12'h276;
        src25 <= 12'hded;
        src26 <= 12'hb92;
        src27 <= 12'hf96;
        src28 <= 12'h10b;
        src29 <= 12'h655;
        src30 <= 12'hee1;
        src31 <= 12'h580;
        src32 <= 12'h3f4;
        src33 <= 12'h3b7;
        src34 <= 12'h359;
        src35 <= 12'h22a;
        src36 <= 12'h357;
        src37 <= 12'h43d;
        src38 <= 12'h974;
        src39 <= 12'hcf1;
        src40 <= 12'h5b;
        src41 <= 12'hd4;
        src42 <= 12'h858;
        src43 <= 12'hc96;
        src44 <= 12'h76b;
        src45 <= 12'h6e7;
        src46 <= 12'hdc4;
        src47 <= 12'hf6d;
        src48 <= 12'he0a;
        src49 <= 12'h7e1;
        src50 <= 12'h316;
        src51 <= 12'h3b5;
        src52 <= 12'h930;
        src53 <= 12'h19;
        src54 <= 12'ha1a;
        src55 <= 12'h33;
        src56 <= 12'h994;
        src57 <= 12'h3a6;
        src58 <= 12'h8d7;
        src59 <= 12'h53e;
        src60 <= 12'h193;
        src61 <= 12'h119;
        src62 <= 12'h855;
        src63 <= 12'hb93;
        exp <= 18'h1e510;
        #1
        src0 <= 12'hf74;
        src1 <= 12'hda1;
        src2 <= 12'he19;
        src3 <= 12'h30c;
        src4 <= 12'h17e;
        src5 <= 12'h594;
        src6 <= 12'hcfb;
        src7 <= 12'h9f1;
        src8 <= 12'h396;
        src9 <= 12'h321;
        src10 <= 12'h7d5;
        src11 <= 12'h682;
        src12 <= 12'h391;
        src13 <= 12'hf92;
        src14 <= 12'ha88;
        src15 <= 12'hcef;
        src16 <= 12'ha12;
        src17 <= 12'hbcb;
        src18 <= 12'h776;
        src19 <= 12'h935;
        src20 <= 12'hffa;
        src21 <= 12'h200;
        src22 <= 12'h282;
        src23 <= 12'h67f;
        src24 <= 12'h51e;
        src25 <= 12'h874;
        src26 <= 12'hbc2;
        src27 <= 12'h9eb;
        src28 <= 12'h4a2;
        src29 <= 12'hc49;
        src30 <= 12'hb9a;
        src31 <= 12'heaf;
        src32 <= 12'h90c;
        src33 <= 12'h524;
        src34 <= 12'h480;
        src35 <= 12'h864;
        src36 <= 12'h25;
        src37 <= 12'hbb6;
        src38 <= 12'h27f;
        src39 <= 12'hec4;
        src40 <= 12'h604;
        src41 <= 12'hb9e;
        src42 <= 12'h4eb;
        src43 <= 12'h6a8;
        src44 <= 12'h7d4;
        src45 <= 12'h81e;
        src46 <= 12'h6c6;
        src47 <= 12'hd7b;
        src48 <= 12'habd;
        src49 <= 12'hdba;
        src50 <= 12'h531;
        src51 <= 12'hade;
        src52 <= 12'hec2;
        src53 <= 12'h2df;
        src54 <= 12'hbcd;
        src55 <= 12'h54e;
        src56 <= 12'h61d;
        src57 <= 12'h803;
        src58 <= 12'h6ab;
        src59 <= 12'hbf1;
        src60 <= 12'h9e4;
        src61 <= 12'h2c6;
        src62 <= 12'hd41;
        src63 <= 12'h4d9;
        exp <= 18'h22032;
        #1
        src0 <= 12'h7d9;
        src1 <= 12'h60b;
        src2 <= 12'hc0d;
        src3 <= 12'h764;
        src4 <= 12'hce5;
        src5 <= 12'ha29;
        src6 <= 12'hdac;
        src7 <= 12'h478;
        src8 <= 12'h6d2;
        src9 <= 12'hbe2;
        src10 <= 12'h3c5;
        src11 <= 12'hd58;
        src12 <= 12'hb2b;
        src13 <= 12'hf4a;
        src14 <= 12'h456;
        src15 <= 12'hd91;
        src16 <= 12'h5f;
        src17 <= 12'hfb0;
        src18 <= 12'h2d3;
        src19 <= 12'hef0;
        src20 <= 12'h197;
        src21 <= 12'h8b1;
        src22 <= 12'h9de;
        src23 <= 12'h244;
        src24 <= 12'h7f7;
        src25 <= 12'he50;
        src26 <= 12'hc77;
        src27 <= 12'hb1;
        src28 <= 12'h8d9;
        src29 <= 12'hf09;
        src30 <= 12'h5f4;
        src31 <= 12'hc09;
        src32 <= 12'h5ae;
        src33 <= 12'ha21;
        src34 <= 12'h39c;
        src35 <= 12'he32;
        src36 <= 12'h298;
        src37 <= 12'h490;
        src38 <= 12'h517;
        src39 <= 12'h671;
        src40 <= 12'hd11;
        src41 <= 12'h369;
        src42 <= 12'h9e9;
        src43 <= 12'hfea;
        src44 <= 12'h16;
        src45 <= 12'h1b5;
        src46 <= 12'h984;
        src47 <= 12'he6e;
        src48 <= 12'h950;
        src49 <= 12'h4c5;
        src50 <= 12'h6c3;
        src51 <= 12'h853;
        src52 <= 12'h8d8;
        src53 <= 12'hf45;
        src54 <= 12'he8d;
        src55 <= 12'h260;
        src56 <= 12'h3e;
        src57 <= 12'h8ee;
        src58 <= 12'hb22;
        src59 <= 12'he39;
        src60 <= 12'h66c;
        src61 <= 12'h1a7;
        src62 <= 12'h43f;
        src63 <= 12'hce2;
        exp <= 18'h21a85;
        #1
        src0 <= 12'h993;
        src1 <= 12'h7d3;
        src2 <= 12'h914;
        src3 <= 12'habb;
        src4 <= 12'h14a;
        src5 <= 12'hf54;
        src6 <= 12'h4aa;
        src7 <= 12'hf64;
        src8 <= 12'hf9e;
        src9 <= 12'h354;
        src10 <= 12'ha96;
        src11 <= 12'h9b6;
        src12 <= 12'h6a1;
        src13 <= 12'h76e;
        src14 <= 12'h729;
        src15 <= 12'hb00;
        src16 <= 12'hdff;
        src17 <= 12'ha34;
        src18 <= 12'h7c7;
        src19 <= 12'h2a1;
        src20 <= 12'h538;
        src21 <= 12'hd23;
        src22 <= 12'h1bc;
        src23 <= 12'h86a;
        src24 <= 12'hff1;
        src25 <= 12'h3cc;
        src26 <= 12'h6af;
        src27 <= 12'had2;
        src28 <= 12'hac7;
        src29 <= 12'h564;
        src30 <= 12'h5fc;
        src31 <= 12'h69f;
        src32 <= 12'hf0f;
        src33 <= 12'h953;
        src34 <= 12'hf26;
        src35 <= 12'h9db;
        src36 <= 12'h851;
        src37 <= 12'hb1;
        src38 <= 12'h9b3;
        src39 <= 12'ha1;
        src40 <= 12'h527;
        src41 <= 12'h113;
        src42 <= 12'he6e;
        src43 <= 12'h70e;
        src44 <= 12'hcde;
        src45 <= 12'h5f3;
        src46 <= 12'h873;
        src47 <= 12'h7f3;
        src48 <= 12'h999;
        src49 <= 12'head;
        src50 <= 12'hb74;
        src51 <= 12'hb85;
        src52 <= 12'h37e;
        src53 <= 12'h7dc;
        src54 <= 12'hf9f;
        src55 <= 12'h7f2;
        src56 <= 12'h26a;
        src57 <= 12'h79c;
        src58 <= 12'hcf0;
        src59 <= 12'hbb5;
        src60 <= 12'hcc0;
        src61 <= 12'hd7b;
        src62 <= 12'hd89;
        src63 <= 12'h9fc;
        exp <= 18'h23cb2;
        #1
        src0 <= 12'h24f;
        src1 <= 12'hcbc;
        src2 <= 12'h7e7;
        src3 <= 12'h7db;
        src4 <= 12'hd95;
        src5 <= 12'hd5;
        src6 <= 12'h1e6;
        src7 <= 12'h4c9;
        src8 <= 12'hb36;
        src9 <= 12'h3e9;
        src10 <= 12'h8a3;
        src11 <= 12'hb44;
        src12 <= 12'hecf;
        src13 <= 12'h9e5;
        src14 <= 12'hfb8;
        src15 <= 12'h180;
        src16 <= 12'hf16;
        src17 <= 12'h465;
        src18 <= 12'hf84;
        src19 <= 12'h66;
        src20 <= 12'hfac;
        src21 <= 12'h362;
        src22 <= 12'h75f;
        src23 <= 12'h54c;
        src24 <= 12'hddd;
        src25 <= 12'heb2;
        src26 <= 12'h534;
        src27 <= 12'hc1d;
        src28 <= 12'h8b4;
        src29 <= 12'h79;
        src30 <= 12'h77b;
        src31 <= 12'h7f;
        src32 <= 12'h6b7;
        src33 <= 12'hdb0;
        src34 <= 12'h53e;
        src35 <= 12'h894;
        src36 <= 12'h2ce;
        src37 <= 12'hc21;
        src38 <= 12'h580;
        src39 <= 12'h9b8;
        src40 <= 12'hdc7;
        src41 <= 12'he76;
        src42 <= 12'hef8;
        src43 <= 12'h39e;
        src44 <= 12'he2f;
        src45 <= 12'h1be;
        src46 <= 12'h214;
        src47 <= 12'h162;
        src48 <= 12'hfc8;
        src49 <= 12'h4ac;
        src50 <= 12'hec8;
        src51 <= 12'h5cf;
        src52 <= 12'hecf;
        src53 <= 12'heeb;
        src54 <= 12'he2c;
        src55 <= 12'hdd2;
        src56 <= 12'h247;
        src57 <= 12'hf21;
        src58 <= 12'h54d;
        src59 <= 12'h1eb;
        src60 <= 12'ha45;
        src61 <= 12'h7bf;
        src62 <= 12'hdbf;
        src63 <= 12'h359;
        exp <= 18'h22412;
        #1
        src0 <= 12'h286;
        src1 <= 12'h835;
        src2 <= 12'hb10;
        src3 <= 12'h6c0;
        src4 <= 12'hc05;
        src5 <= 12'h27d;
        src6 <= 12'h4b0;
        src7 <= 12'h16c;
        src8 <= 12'h211;
        src9 <= 12'h5a5;
        src10 <= 12'hed7;
        src11 <= 12'h96;
        src12 <= 12'he0a;
        src13 <= 12'h94f;
        src14 <= 12'h8f5;
        src15 <= 12'he07;
        src16 <= 12'h9b4;
        src17 <= 12'he27;
        src18 <= 12'hfb3;
        src19 <= 12'h911;
        src20 <= 12'h569;
        src21 <= 12'hec0;
        src22 <= 12'h68c;
        src23 <= 12'h5ef;
        src24 <= 12'h379;
        src25 <= 12'h8fd;
        src26 <= 12'hb6c;
        src27 <= 12'hee7;
        src28 <= 12'h16b;
        src29 <= 12'h55d;
        src30 <= 12'h57;
        src31 <= 12'hae5;
        src32 <= 12'h192;
        src33 <= 12'h1ed;
        src34 <= 12'h7ab;
        src35 <= 12'ha09;
        src36 <= 12'h93a;
        src37 <= 12'hcad;
        src38 <= 12'h177;
        src39 <= 12'h242;
        src40 <= 12'h8fb;
        src41 <= 12'h713;
        src42 <= 12'h3bb;
        src43 <= 12'h5f1;
        src44 <= 12'h5f4;
        src45 <= 12'h687;
        src46 <= 12'h4cc;
        src47 <= 12'h4fc;
        src48 <= 12'hdcf;
        src49 <= 12'he10;
        src50 <= 12'hd16;
        src51 <= 12'hcde;
        src52 <= 12'h537;
        src53 <= 12'h38c;
        src54 <= 12'hc5f;
        src55 <= 12'h68b;
        src56 <= 12'h8aa;
        src57 <= 12'hb56;
        src58 <= 12'haf2;
        src59 <= 12'ha7;
        src60 <= 12'h3cc;
        src61 <= 12'hec4;
        src62 <= 12'h839;
        src63 <= 12'h885;
        exp <= 18'h1f3e8;
        #1
        src0 <= 12'he47;
        src1 <= 12'h4d4;
        src2 <= 12'he62;
        src3 <= 12'he34;
        src4 <= 12'h410;
        src5 <= 12'h27b;
        src6 <= 12'hf3b;
        src7 <= 12'hac7;
        src8 <= 12'hb33;
        src9 <= 12'h174;
        src10 <= 12'h909;
        src11 <= 12'he4e;
        src12 <= 12'hbc4;
        src13 <= 12'hd2d;
        src14 <= 12'h77c;
        src15 <= 12'h100;
        src16 <= 12'hcb8;
        src17 <= 12'h64d;
        src18 <= 12'h4c1;
        src19 <= 12'h358;
        src20 <= 12'h37c;
        src21 <= 12'h8eb;
        src22 <= 12'hcc6;
        src23 <= 12'h325;
        src24 <= 12'h302;
        src25 <= 12'h679;
        src26 <= 12'h230;
        src27 <= 12'h2cf;
        src28 <= 12'h5c5;
        src29 <= 12'h2c4;
        src30 <= 12'h41c;
        src31 <= 12'hca4;
        src32 <= 12'hcc8;
        src33 <= 12'h1be;
        src34 <= 12'h23d;
        src35 <= 12'h979;
        src36 <= 12'h569;
        src37 <= 12'h76e;
        src38 <= 12'hf3f;
        src39 <= 12'hfdc;
        src40 <= 12'heb5;
        src41 <= 12'ha32;
        src42 <= 12'hba7;
        src43 <= 12'hba6;
        src44 <= 12'h346;
        src45 <= 12'h850;
        src46 <= 12'h8fa;
        src47 <= 12'h4e0;
        src48 <= 12'he9b;
        src49 <= 12'he0d;
        src50 <= 12'h50f;
        src51 <= 12'h66e;
        src52 <= 12'h36b;
        src53 <= 12'h194;
        src54 <= 12'h2dc;
        src55 <= 12'h1b3;
        src56 <= 12'hf21;
        src57 <= 12'hd99;
        src58 <= 12'h7e3;
        src59 <= 12'h677;
        src60 <= 12'h1e0;
        src61 <= 12'h353;
        src62 <= 12'h6d4;
        src63 <= 12'hd86;
        exp <= 18'h1fb02;
        #1
        src0 <= 12'h697;
        src1 <= 12'hb1f;
        src2 <= 12'h240;
        src3 <= 12'h4cb;
        src4 <= 12'hf92;
        src5 <= 12'hd1f;
        src6 <= 12'hc61;
        src7 <= 12'h7bd;
        src8 <= 12'h21e;
        src9 <= 12'hfec;
        src10 <= 12'h8d0;
        src11 <= 12'h698;
        src12 <= 12'hf90;
        src13 <= 12'h19d;
        src14 <= 12'h7d5;
        src15 <= 12'h584;
        src16 <= 12'h6a7;
        src17 <= 12'h1a6;
        src18 <= 12'h70a;
        src19 <= 12'hf3c;
        src20 <= 12'hed4;
        src21 <= 12'hc9;
        src22 <= 12'h6c3;
        src23 <= 12'hff0;
        src24 <= 12'hbbf;
        src25 <= 12'hfda;
        src26 <= 12'hb1e;
        src27 <= 12'h405;
        src28 <= 12'hc2c;
        src29 <= 12'h354;
        src30 <= 12'h1f5;
        src31 <= 12'h3c8;
        src32 <= 12'h64a;
        src33 <= 12'h9bb;
        src34 <= 12'hdda;
        src35 <= 12'h9a5;
        src36 <= 12'ha09;
        src37 <= 12'h64e;
        src38 <= 12'h802;
        src39 <= 12'hdb2;
        src40 <= 12'h16d;
        src41 <= 12'h250;
        src42 <= 12'he53;
        src43 <= 12'ha4e;
        src44 <= 12'hc7;
        src45 <= 12'h356;
        src46 <= 12'he04;
        src47 <= 12'h93f;
        src48 <= 12'h75f;
        src49 <= 12'h4bf;
        src50 <= 12'h4f3;
        src51 <= 12'hc3d;
        src52 <= 12'h222;
        src53 <= 12'h70f;
        src54 <= 12'h1eb;
        src55 <= 12'haad;
        src56 <= 12'hbf3;
        src57 <= 12'h5ad;
        src58 <= 12'h408;
        src59 <= 12'h624;
        src60 <= 12'h12d;
        src61 <= 12'heb9;
        src62 <= 12'h10c;
        src63 <= 12'h995;
        exp <= 18'h1fd1b;
        #1
        src0 <= 12'h849;
        src1 <= 12'h27e;
        src2 <= 12'h97f;
        src3 <= 12'he2b;
        src4 <= 12'he5c;
        src5 <= 12'haa9;
        src6 <= 12'h8ad;
        src7 <= 12'ha6b;
        src8 <= 12'h2bc;
        src9 <= 12'h148;
        src10 <= 12'h557;
        src11 <= 12'h704;
        src12 <= 12'h5d7;
        src13 <= 12'h404;
        src14 <= 12'hf93;
        src15 <= 12'h5b6;
        src16 <= 12'h323;
        src17 <= 12'hb1b;
        src18 <= 12'h6fe;
        src19 <= 12'h2d4;
        src20 <= 12'hb8d;
        src21 <= 12'h88f;
        src22 <= 12'hd23;
        src23 <= 12'h77;
        src24 <= 12'hb99;
        src25 <= 12'heaf;
        src26 <= 12'h318;
        src27 <= 12'ha45;
        src28 <= 12'h9a2;
        src29 <= 12'h7e5;
        src30 <= 12'hf46;
        src31 <= 12'hc95;
        src32 <= 12'hd7d;
        src33 <= 12'h109;
        src34 <= 12'h2d;
        src35 <= 12'hc4a;
        src36 <= 12'h39b;
        src37 <= 12'had;
        src38 <= 12'h3c2;
        src39 <= 12'h338;
        src40 <= 12'h61f;
        src41 <= 12'ha98;
        src42 <= 12'haa8;
        src43 <= 12'hc6a;
        src44 <= 12'h159;
        src45 <= 12'h139;
        src46 <= 12'hf;
        src47 <= 12'ha55;
        src48 <= 12'h67e;
        src49 <= 12'h73e;
        src50 <= 12'h678;
        src51 <= 12'h65;
        src52 <= 12'h68a;
        src53 <= 12'h163;
        src54 <= 12'hc87;
        src55 <= 12'h4dd;
        src56 <= 12'ha7;
        src57 <= 12'h320;
        src58 <= 12'ha50;
        src59 <= 12'hbb;
        src60 <= 12'h30d;
        src61 <= 12'h479;
        src62 <= 12'h735;
        src63 <= 12'h2c5;
        exp <= 18'h1b618;
        #1
        src0 <= 12'h876;
        src1 <= 12'h209;
        src2 <= 12'h813;
        src3 <= 12'hb12;
        src4 <= 12'h323;
        src5 <= 12'hee4;
        src6 <= 12'h1e2;
        src7 <= 12'h28c;
        src8 <= 12'hbaa;
        src9 <= 12'h7c6;
        src10 <= 12'hf2a;
        src11 <= 12'h84b;
        src12 <= 12'hde0;
        src13 <= 12'hd83;
        src14 <= 12'h5dc;
        src15 <= 12'hc04;
        src16 <= 12'h715;
        src17 <= 12'heeb;
        src18 <= 12'hed0;
        src19 <= 12'hc45;
        src20 <= 12'he5a;
        src21 <= 12'hc33;
        src22 <= 12'h38d;
        src23 <= 12'hf13;
        src24 <= 12'hb14;
        src25 <= 12'h9de;
        src26 <= 12'h90a;
        src27 <= 12'hc38;
        src28 <= 12'h21a;
        src29 <= 12'hf01;
        src30 <= 12'h701;
        src31 <= 12'h4ca;
        src32 <= 12'h79;
        src33 <= 12'h863;
        src34 <= 12'hd7f;
        src35 <= 12'h5cb;
        src36 <= 12'hfe5;
        src37 <= 12'hdf9;
        src38 <= 12'he00;
        src39 <= 12'ha39;
        src40 <= 12'hea1;
        src41 <= 12'hb61;
        src42 <= 12'hbc8;
        src43 <= 12'hbab;
        src44 <= 12'hfc;
        src45 <= 12'h134;
        src46 <= 12'h623;
        src47 <= 12'hf01;
        src48 <= 12'h211;
        src49 <= 12'h47b;
        src50 <= 12'h8e2;
        src51 <= 12'hb5d;
        src52 <= 12'h9b4;
        src53 <= 12'ha08;
        src54 <= 12'hcc5;
        src55 <= 12'hbbf;
        src56 <= 12'ha8d;
        src57 <= 12'hcb9;
        src58 <= 12'h4fd;
        src59 <= 12'hb17;
        src60 <= 12'h6c1;
        src61 <= 12'hbce;
        src62 <= 12'h93;
        src63 <= 12'hf61;
        exp <= 18'h25d8b;
        #1
        src0 <= 12'hd74;
        src1 <= 12'h79e;
        src2 <= 12'h447;
        src3 <= 12'hf36;
        src4 <= 12'h9d8;
        src5 <= 12'ha52;
        src6 <= 12'h3c8;
        src7 <= 12'hb4b;
        src8 <= 12'hd8b;
        src9 <= 12'h33e;
        src10 <= 12'h3d9;
        src11 <= 12'hd22;
        src12 <= 12'h8e3;
        src13 <= 12'hb16;
        src14 <= 12'h7ff;
        src15 <= 12'ha9;
        src16 <= 12'hdea;
        src17 <= 12'h4ea;
        src18 <= 12'ha2a;
        src19 <= 12'h83b;
        src20 <= 12'hab5;
        src21 <= 12'h4e0;
        src22 <= 12'h294;
        src23 <= 12'h996;
        src24 <= 12'h797;
        src25 <= 12'he22;
        src26 <= 12'h8de;
        src27 <= 12'h28f;
        src28 <= 12'h10e;
        src29 <= 12'h60c;
        src30 <= 12'hfc;
        src31 <= 12'hedb;
        src32 <= 12'ha0c;
        src33 <= 12'h1ed;
        src34 <= 12'hd83;
        src35 <= 12'h94f;
        src36 <= 12'h1e4;
        src37 <= 12'h3d7;
        src38 <= 12'hc97;
        src39 <= 12'hb32;
        src40 <= 12'hb8c;
        src41 <= 12'hfb5;
        src42 <= 12'h79d;
        src43 <= 12'h3c5;
        src44 <= 12'h33c;
        src45 <= 12'h6bf;
        src46 <= 12'habc;
        src47 <= 12'hf92;
        src48 <= 12'h3e3;
        src49 <= 12'hef;
        src50 <= 12'hdf;
        src51 <= 12'h939;
        src52 <= 12'h122;
        src53 <= 12'hf3;
        src54 <= 12'hc46;
        src55 <= 12'hc87;
        src56 <= 12'h729;
        src57 <= 12'h535;
        src58 <= 12'h2ed;
        src59 <= 12'h170;
        src60 <= 12'had;
        src61 <= 12'hef4;
        src62 <= 12'hded;
        src63 <= 12'h6d7;
        exp <= 18'h1ed67;
        #1
        src0 <= 12'haca;
        src1 <= 12'hc84;
        src2 <= 12'hc15;
        src3 <= 12'h2c9;
        src4 <= 12'h8c9;
        src5 <= 12'h6e1;
        src6 <= 12'h8d3;
        src7 <= 12'h558;
        src8 <= 12'h31b;
        src9 <= 12'h3d9;
        src10 <= 12'h139;
        src11 <= 12'hddf;
        src12 <= 12'h6ac;
        src13 <= 12'h781;
        src14 <= 12'hc4b;
        src15 <= 12'h79f;
        src16 <= 12'ha19;
        src17 <= 12'haf2;
        src18 <= 12'h13f;
        src19 <= 12'h134;
        src20 <= 12'hb99;
        src21 <= 12'hd4c;
        src22 <= 12'hb2c;
        src23 <= 12'h572;
        src24 <= 12'haef;
        src25 <= 12'h135;
        src26 <= 12'h21b;
        src27 <= 12'h75a;
        src28 <= 12'h844;
        src29 <= 12'h701;
        src30 <= 12'h53a;
        src31 <= 12'h182;
        src32 <= 12'h11e;
        src33 <= 12'h8a9;
        src34 <= 12'hba9;
        src35 <= 12'h64c;
        src36 <= 12'hd41;
        src37 <= 12'h869;
        src38 <= 12'he69;
        src39 <= 12'h412;
        src40 <= 12'h9cf;
        src41 <= 12'hffe;
        src42 <= 12'hbe6;
        src43 <= 12'he2e;
        src44 <= 12'h5ec;
        src45 <= 12'h2ea;
        src46 <= 12'h80d;
        src47 <= 12'h8f0;
        src48 <= 12'hc61;
        src49 <= 12'h786;
        src50 <= 12'h401;
        src51 <= 12'h7a0;
        src52 <= 12'h6c0;
        src53 <= 12'he82;
        src54 <= 12'hbaa;
        src55 <= 12'h5e9;
        src56 <= 12'h8aa;
        src57 <= 12'hd9a;
        src58 <= 12'hf89;
        src59 <= 12'hbfe;
        src60 <= 12'h94e;
        src61 <= 12'ha2a;
        src62 <= 12'h1;
        src63 <= 12'he76;
        exp <= 18'h2146b;
        #1
        src0 <= 12'hb17;
        src1 <= 12'hed4;
        src2 <= 12'h28f;
        src3 <= 12'hedf;
        src4 <= 12'he27;
        src5 <= 12'h97f;
        src6 <= 12'h6f2;
        src7 <= 12'hdb4;
        src8 <= 12'hed2;
        src9 <= 12'hb77;
        src10 <= 12'ha34;
        src11 <= 12'h39e;
        src12 <= 12'hfe5;
        src13 <= 12'hcf6;
        src14 <= 12'h2d3;
        src15 <= 12'hc29;
        src16 <= 12'h3eb;
        src17 <= 12'h602;
        src18 <= 12'hf21;
        src19 <= 12'h117;
        src20 <= 12'hf59;
        src21 <= 12'ha47;
        src22 <= 12'hb6f;
        src23 <= 12'h8b0;
        src24 <= 12'h10b;
        src25 <= 12'h462;
        src26 <= 12'h799;
        src27 <= 12'h9d6;
        src28 <= 12'h9b;
        src29 <= 12'h99e;
        src30 <= 12'he73;
        src31 <= 12'hf26;
        src32 <= 12'ha2f;
        src33 <= 12'h62e;
        src34 <= 12'h12e;
        src35 <= 12'h486;
        src36 <= 12'h392;
        src37 <= 12'hfba;
        src38 <= 12'h161;
        src39 <= 12'h172;
        src40 <= 12'h7ef;
        src41 <= 12'h8e3;
        src42 <= 12'hbdd;
        src43 <= 12'h8a5;
        src44 <= 12'hdeb;
        src45 <= 12'hd97;
        src46 <= 12'h7ce;
        src47 <= 12'h329;
        src48 <= 12'hf3;
        src49 <= 12'h4f8;
        src50 <= 12'h6b;
        src51 <= 12'h5d4;
        src52 <= 12'hd6e;
        src53 <= 12'haa0;
        src54 <= 12'h1f0;
        src55 <= 12'hc6e;
        src56 <= 12'hf9f;
        src57 <= 12'h98b;
        src58 <= 12'hba0;
        src59 <= 12'hbf0;
        src60 <= 12'hfed;
        src61 <= 12'h3f;
        src62 <= 12'ha74;
        src63 <= 12'hb9d;
        exp <= 18'h233b3;
        #1
        src0 <= 12'h774;
        src1 <= 12'h61f;
        src2 <= 12'h3ad;
        src3 <= 12'h52e;
        src4 <= 12'h4de;
        src5 <= 12'h17e;
        src6 <= 12'h3c2;
        src7 <= 12'hf9e;
        src8 <= 12'h3a8;
        src9 <= 12'hdff;
        src10 <= 12'h824;
        src11 <= 12'hf83;
        src12 <= 12'hb18;
        src13 <= 12'ha3d;
        src14 <= 12'h11e;
        src15 <= 12'h76;
        src16 <= 12'ha54;
        src17 <= 12'he57;
        src18 <= 12'h598;
        src19 <= 12'hee9;
        src20 <= 12'h643;
        src21 <= 12'h86;
        src22 <= 12'h860;
        src23 <= 12'h2c;
        src24 <= 12'h9a1;
        src25 <= 12'hdb2;
        src26 <= 12'h52c;
        src27 <= 12'hccc;
        src28 <= 12'hc79;
        src29 <= 12'hbd9;
        src30 <= 12'h6b8;
        src31 <= 12'he3b;
        src32 <= 12'hd69;
        src33 <= 12'h85b;
        src34 <= 12'h9a8;
        src35 <= 12'hf23;
        src36 <= 12'hedf;
        src37 <= 12'h56e;
        src38 <= 12'h2fc;
        src39 <= 12'h7c2;
        src40 <= 12'h2ad;
        src41 <= 12'hfdf;
        src42 <= 12'h18d;
        src43 <= 12'hcdc;
        src44 <= 12'hda7;
        src45 <= 12'hb56;
        src46 <= 12'hda2;
        src47 <= 12'hc5e;
        src48 <= 12'h978;
        src49 <= 12'hec;
        src50 <= 12'hecf;
        src51 <= 12'h8bf;
        src52 <= 12'h870;
        src53 <= 12'ha4e;
        src54 <= 12'h309;
        src55 <= 12'hbe9;
        src56 <= 12'h30f;
        src57 <= 12'ha1c;
        src58 <= 12'h42f;
        src59 <= 12'he95;
        src60 <= 12'hdc8;
        src61 <= 12'he81;
        src62 <= 12'hca3;
        src63 <= 12'hc82;
        exp <= 18'h23dfd;
        #1
        src0 <= 12'h457;
        src1 <= 12'hb4e;
        src2 <= 12'h13d;
        src3 <= 12'h687;
        src4 <= 12'h4b;
        src5 <= 12'h464;
        src6 <= 12'h298;
        src7 <= 12'h9b3;
        src8 <= 12'hfda;
        src9 <= 12'h4a9;
        src10 <= 12'hf95;
        src11 <= 12'h32e;
        src12 <= 12'h1f7;
        src13 <= 12'hbd8;
        src14 <= 12'h1fc;
        src15 <= 12'hb65;
        src16 <= 12'h87b;
        src17 <= 12'h46;
        src18 <= 12'he96;
        src19 <= 12'h55e;
        src20 <= 12'h75f;
        src21 <= 12'ha95;
        src22 <= 12'h780;
        src23 <= 12'h1b5;
        src24 <= 12'h189;
        src25 <= 12'h77c;
        src26 <= 12'hc13;
        src27 <= 12'hc60;
        src28 <= 12'hbe7;
        src29 <= 12'h8aa;
        src30 <= 12'hb72;
        src31 <= 12'h1fb;
        src32 <= 12'h8d7;
        src33 <= 12'h690;
        src34 <= 12'h89f;
        src35 <= 12'ha73;
        src36 <= 12'h2d4;
        src37 <= 12'h8a3;
        src38 <= 12'h4ce;
        src39 <= 12'h7c8;
        src40 <= 12'hd3e;
        src41 <= 12'hc93;
        src42 <= 12'h3db;
        src43 <= 12'h7e1;
        src44 <= 12'h794;
        src45 <= 12'h2e1;
        src46 <= 12'hdc1;
        src47 <= 12'hd21;
        src48 <= 12'hfd7;
        src49 <= 12'h846;
        src50 <= 12'habf;
        src51 <= 12'he36;
        src52 <= 12'hbfa;
        src53 <= 12'hbd8;
        src54 <= 12'h972;
        src55 <= 12'hd65;
        src56 <= 12'h790;
        src57 <= 12'ha2f;
        src58 <= 12'ha31;
        src59 <= 12'h519;
        src60 <= 12'hbf6;
        src61 <= 12'h35;
        src62 <= 12'h32b;
        src63 <= 12'h33;
        exp <= 18'h1fbe4;
        #1
        src0 <= 12'h3c0;
        src1 <= 12'ha8e;
        src2 <= 12'hc07;
        src3 <= 12'hbae;
        src4 <= 12'hc44;
        src5 <= 12'h8ae;
        src6 <= 12'h161;
        src7 <= 12'h21b;
        src8 <= 12'hf6e;
        src9 <= 12'h364;
        src10 <= 12'he3c;
        src11 <= 12'h76;
        src12 <= 12'ha46;
        src13 <= 12'hf7c;
        src14 <= 12'hfa5;
        src15 <= 12'h484;
        src16 <= 12'h500;
        src17 <= 12'h5ed;
        src18 <= 12'hd11;
        src19 <= 12'h78f;
        src20 <= 12'h1c5;
        src21 <= 12'h41e;
        src22 <= 12'hf3;
        src23 <= 12'h9c3;
        src24 <= 12'h324;
        src25 <= 12'hd6f;
        src26 <= 12'ha7d;
        src27 <= 12'he5;
        src28 <= 12'h7a2;
        src29 <= 12'h81;
        src30 <= 12'h3c7;
        src31 <= 12'ha9d;
        src32 <= 12'he53;
        src33 <= 12'hac1;
        src34 <= 12'hd31;
        src35 <= 12'hea9;
        src36 <= 12'hae6;
        src37 <= 12'ha8b;
        src38 <= 12'h666;
        src39 <= 12'hc0a;
        src40 <= 12'h1b9;
        src41 <= 12'h351;
        src42 <= 12'h24d;
        src43 <= 12'haca;
        src44 <= 12'hb4c;
        src45 <= 12'hefd;
        src46 <= 12'ha0;
        src47 <= 12'hd64;
        src48 <= 12'h61c;
        src49 <= 12'h8f0;
        src50 <= 12'h9f0;
        src51 <= 12'hdf5;
        src52 <= 12'h81f;
        src53 <= 12'hf9b;
        src54 <= 12'h216;
        src55 <= 12'hd74;
        src56 <= 12'h893;
        src57 <= 12'hb6e;
        src58 <= 12'h977;
        src59 <= 12'h8c;
        src60 <= 12'h5a3;
        src61 <= 12'hd5e;
        src62 <= 12'h40c;
        src63 <= 12'hd03;
        exp <= 18'h21808;
        #1
        src0 <= 12'h2ce;
        src1 <= 12'h801;
        src2 <= 12'h4c6;
        src3 <= 12'h10c;
        src4 <= 12'he00;
        src5 <= 12'h923;
        src6 <= 12'hadf;
        src7 <= 12'hd17;
        src8 <= 12'h8e1;
        src9 <= 12'h4c6;
        src10 <= 12'hb43;
        src11 <= 12'h857;
        src12 <= 12'h72b;
        src13 <= 12'h3d6;
        src14 <= 12'h4f1;
        src15 <= 12'hda5;
        src16 <= 12'h519;
        src17 <= 12'h868;
        src18 <= 12'hfa5;
        src19 <= 12'h409;
        src20 <= 12'h556;
        src21 <= 12'h7f;
        src22 <= 12'he35;
        src23 <= 12'h1e8;
        src24 <= 12'h6c9;
        src25 <= 12'h856;
        src26 <= 12'h81c;
        src27 <= 12'h857;
        src28 <= 12'h34d;
        src29 <= 12'h18b;
        src30 <= 12'hebb;
        src31 <= 12'h45d;
        src32 <= 12'hd19;
        src33 <= 12'h8e3;
        src34 <= 12'h825;
        src35 <= 12'ha1a;
        src36 <= 12'h2e7;
        src37 <= 12'h115;
        src38 <= 12'hf55;
        src39 <= 12'h5ea;
        src40 <= 12'hd41;
        src41 <= 12'h911;
        src42 <= 12'h1f0;
        src43 <= 12'h48c;
        src44 <= 12'hb7;
        src45 <= 12'h811;
        src46 <= 12'h82c;
        src47 <= 12'h8d0;
        src48 <= 12'hb31;
        src49 <= 12'hf2d;
        src50 <= 12'h194;
        src51 <= 12'h81;
        src52 <= 12'hde0;
        src53 <= 12'h1f4;
        src54 <= 12'h7bd;
        src55 <= 12'hf59;
        src56 <= 12'hfb6;
        src57 <= 12'hb5;
        src58 <= 12'hca7;
        src59 <= 12'h162;
        src60 <= 12'h3ce;
        src61 <= 12'hdff;
        src62 <= 12'h825;
        src63 <= 12'h500;
        exp <= 18'h1e600;
        #1
        src0 <= 12'h850;
        src1 <= 12'h370;
        src2 <= 12'h7bf;
        src3 <= 12'h1e4;
        src4 <= 12'h785;
        src5 <= 12'hef9;
        src6 <= 12'h73d;
        src7 <= 12'hcfa;
        src8 <= 12'he38;
        src9 <= 12'h4e8;
        src10 <= 12'h55c;
        src11 <= 12'h412;
        src12 <= 12'h7e3;
        src13 <= 12'h31c;
        src14 <= 12'hbd3;
        src15 <= 12'h348;
        src16 <= 12'h4b4;
        src17 <= 12'h3b2;
        src18 <= 12'h19f;
        src19 <= 12'h437;
        src20 <= 12'hed6;
        src21 <= 12'hb51;
        src22 <= 12'h58;
        src23 <= 12'haf9;
        src24 <= 12'hf67;
        src25 <= 12'hadc;
        src26 <= 12'hb8e;
        src27 <= 12'h671;
        src28 <= 12'h7dc;
        src29 <= 12'h654;
        src30 <= 12'ha7d;
        src31 <= 12'hcc2;
        src32 <= 12'h3dc;
        src33 <= 12'h190;
        src34 <= 12'h511;
        src35 <= 12'hd6;
        src36 <= 12'he79;
        src37 <= 12'h167;
        src38 <= 12'h3c2;
        src39 <= 12'h371;
        src40 <= 12'h4f;
        src41 <= 12'hc72;
        src42 <= 12'h1b2;
        src43 <= 12'h9d5;
        src44 <= 12'hefd;
        src45 <= 12'h9e2;
        src46 <= 12'hb36;
        src47 <= 12'h31c;
        src48 <= 12'h9c4;
        src49 <= 12'he83;
        src50 <= 12'h8a7;
        src51 <= 12'hcd2;
        src52 <= 12'h48c;
        src53 <= 12'h60a;
        src54 <= 12'h295;
        src55 <= 12'head;
        src56 <= 12'h535;
        src57 <= 12'hb82;
        src58 <= 12'ha56;
        src59 <= 12'he3d;
        src60 <= 12'h880;
        src61 <= 12'hb60;
        src62 <= 12'hbb0;
        src63 <= 12'h1a7;
        exp <= 18'h1f21d;
        #1
        src0 <= 12'h462;
        src1 <= 12'h41;
        src2 <= 12'h268;
        src3 <= 12'h1c4;
        src4 <= 12'hc02;
        src5 <= 12'h7cf;
        src6 <= 12'h7a4;
        src7 <= 12'he28;
        src8 <= 12'h787;
        src9 <= 12'h687;
        src10 <= 12'hefd;
        src11 <= 12'hb87;
        src12 <= 12'he56;
        src13 <= 12'h740;
        src14 <= 12'hd12;
        src15 <= 12'h5ee;
        src16 <= 12'h800;
        src17 <= 12'hbc3;
        src18 <= 12'hc1b;
        src19 <= 12'h439;
        src20 <= 12'h5c3;
        src21 <= 12'hfda;
        src22 <= 12'h329;
        src23 <= 12'h174;
        src24 <= 12'h4b3;
        src25 <= 12'hfb8;
        src26 <= 12'h9f2;
        src27 <= 12'h760;
        src28 <= 12'h3ef;
        src29 <= 12'h8b1;
        src30 <= 12'he9f;
        src31 <= 12'h272;
        src32 <= 12'h169;
        src33 <= 12'hbde;
        src34 <= 12'h874;
        src35 <= 12'hcd0;
        src36 <= 12'h655;
        src37 <= 12'h82c;
        src38 <= 12'h561;
        src39 <= 12'h687;
        src40 <= 12'h218;
        src41 <= 12'he44;
        src42 <= 12'hfe1;
        src43 <= 12'h90c;
        src44 <= 12'h8a4;
        src45 <= 12'h99d;
        src46 <= 12'h8a6;
        src47 <= 12'h8a1;
        src48 <= 12'hfa8;
        src49 <= 12'h9f9;
        src50 <= 12'h751;
        src51 <= 12'hf5e;
        src52 <= 12'h66a;
        src53 <= 12'h3d4;
        src54 <= 12'he7;
        src55 <= 12'he19;
        src56 <= 12'h697;
        src57 <= 12'he37;
        src58 <= 12'h83;
        src59 <= 12'h362;
        src60 <= 12'he5;
        src61 <= 12'hade;
        src62 <= 12'hcf9;
        src63 <= 12'hd72;
        exp <= 18'h21787;
        #1
        src0 <= 12'h479;
        src1 <= 12'h95a;
        src2 <= 12'hefb;
        src3 <= 12'hf71;
        src4 <= 12'hf57;
        src5 <= 12'h7ea;
        src6 <= 12'hf77;
        src7 <= 12'h368;
        src8 <= 12'h7c9;
        src9 <= 12'hba7;
        src10 <= 12'h9bf;
        src11 <= 12'h61a;
        src12 <= 12'hbe;
        src13 <= 12'ha39;
        src14 <= 12'h42;
        src15 <= 12'h2db;
        src16 <= 12'h2aa;
        src17 <= 12'h587;
        src18 <= 12'h95c;
        src19 <= 12'h883;
        src20 <= 12'h958;
        src21 <= 12'h504;
        src22 <= 12'hf4f;
        src23 <= 12'h91;
        src24 <= 12'h58e;
        src25 <= 12'h979;
        src26 <= 12'hf2e;
        src27 <= 12'h27c;
        src28 <= 12'h5bf;
        src29 <= 12'hcf2;
        src30 <= 12'h48c;
        src31 <= 12'h136;
        src32 <= 12'hac9;
        src33 <= 12'h15b;
        src34 <= 12'h3e7;
        src35 <= 12'h83;
        src36 <= 12'hcd4;
        src37 <= 12'h907;
        src38 <= 12'h64f;
        src39 <= 12'h879;
        src40 <= 12'hab3;
        src41 <= 12'hc0;
        src42 <= 12'h632;
        src43 <= 12'h911;
        src44 <= 12'h785;
        src45 <= 12'h11c;
        src46 <= 12'h63e;
        src47 <= 12'hbd8;
        src48 <= 12'h971;
        src49 <= 12'h4ec;
        src50 <= 12'hb64;
        src51 <= 12'hea5;
        src52 <= 12'hc2d;
        src53 <= 12'h705;
        src54 <= 12'h722;
        src55 <= 12'h191;
        src56 <= 12'hdd9;
        src57 <= 12'hd87;
        src58 <= 12'h2d3;
        src59 <= 12'h69e;
        src60 <= 12'h421;
        src61 <= 12'haf2;
        src62 <= 12'h2e;
        src63 <= 12'h262;
        exp <= 18'h1de89;
        #1
        src0 <= 12'h6be;
        src1 <= 12'hed;
        src2 <= 12'h302;
        src3 <= 12'hff7;
        src4 <= 12'ha23;
        src5 <= 12'hc88;
        src6 <= 12'h62c;
        src7 <= 12'hd05;
        src8 <= 12'hb14;
        src9 <= 12'h318;
        src10 <= 12'h24c;
        src11 <= 12'h703;
        src12 <= 12'h57c;
        src13 <= 12'h99c;
        src14 <= 12'hc8f;
        src15 <= 12'hf7d;
        src16 <= 12'h73d;
        src17 <= 12'hc4f;
        src18 <= 12'h55d;
        src19 <= 12'haf4;
        src20 <= 12'hc3c;
        src21 <= 12'hcaf;
        src22 <= 12'h2cb;
        src23 <= 12'h6d5;
        src24 <= 12'hb5c;
        src25 <= 12'h2c1;
        src26 <= 12'hd37;
        src27 <= 12'he56;
        src28 <= 12'hf11;
        src29 <= 12'h9ca;
        src30 <= 12'he7c;
        src31 <= 12'ha58;
        src32 <= 12'hd96;
        src33 <= 12'h9d5;
        src34 <= 12'h476;
        src35 <= 12'h99f;
        src36 <= 12'h42d;
        src37 <= 12'h56e;
        src38 <= 12'h35a;
        src39 <= 12'h3a6;
        src40 <= 12'h590;
        src41 <= 12'h1cc;
        src42 <= 12'h221;
        src43 <= 12'h747;
        src44 <= 12'h21d;
        src45 <= 12'hc0e;
        src46 <= 12'h73;
        src47 <= 12'h2df;
        src48 <= 12'hd64;
        src49 <= 12'h2c3;
        src50 <= 12'habf;
        src51 <= 12'h2c1;
        src52 <= 12'h989;
        src53 <= 12'hd7a;
        src54 <= 12'h9e3;
        src55 <= 12'hd7c;
        src56 <= 12'hf38;
        src57 <= 12'h9ba;
        src58 <= 12'h4da;
        src59 <= 12'he4c;
        src60 <= 12'h52d;
        src61 <= 12'hadd;
        src62 <= 12'heb9;
        src63 <= 12'hccb;
        exp <= 18'h224eb;
        #1
        src0 <= 12'hc03;
        src1 <= 12'ha28;
        src2 <= 12'he3b;
        src3 <= 12'h2f6;
        src4 <= 12'h58a;
        src5 <= 12'hf29;
        src6 <= 12'hfce;
        src7 <= 12'ha4f;
        src8 <= 12'h542;
        src9 <= 12'h3fb;
        src10 <= 12'h4da;
        src11 <= 12'h5;
        src12 <= 12'h308;
        src13 <= 12'h5a4;
        src14 <= 12'h9c6;
        src15 <= 12'hf81;
        src16 <= 12'h269;
        src17 <= 12'hf05;
        src18 <= 12'h33c;
        src19 <= 12'hea4;
        src20 <= 12'h988;
        src21 <= 12'hc40;
        src22 <= 12'h401;
        src23 <= 12'h13b;
        src24 <= 12'ha09;
        src25 <= 12'h246;
        src26 <= 12'hc46;
        src27 <= 12'h6fc;
        src28 <= 12'hd7c;
        src29 <= 12'h5a0;
        src30 <= 12'ha44;
        src31 <= 12'h821;
        src32 <= 12'hea6;
        src33 <= 12'hb84;
        src34 <= 12'h507;
        src35 <= 12'hcb3;
        src36 <= 12'h93;
        src37 <= 12'hd52;
        src38 <= 12'h52;
        src39 <= 12'h9b4;
        src40 <= 12'h5f;
        src41 <= 12'hbe6;
        src42 <= 12'h111;
        src43 <= 12'hfc5;
        src44 <= 12'hfe0;
        src45 <= 12'h5ac;
        src46 <= 12'h14;
        src47 <= 12'ha34;
        src48 <= 12'hfe5;
        src49 <= 12'hf63;
        src50 <= 12'hdd6;
        src51 <= 12'hc45;
        src52 <= 12'he0b;
        src53 <= 12'h6c3;
        src54 <= 12'h7a2;
        src55 <= 12'h4b;
        src56 <= 12'h2a2;
        src57 <= 12'h9e;
        src58 <= 12'hfeb;
        src59 <= 12'hed5;
        src60 <= 12'h489;
        src61 <= 12'h435;
        src62 <= 12'haf7;
        src63 <= 12'hd45;
        exp <= 18'h22375;
        #1
        src0 <= 12'h947;
        src1 <= 12'haf7;
        src2 <= 12'hc2f;
        src3 <= 12'ha61;
        src4 <= 12'h37e;
        src5 <= 12'hfb;
        src6 <= 12'hd19;
        src7 <= 12'h15c;
        src8 <= 12'h79;
        src9 <= 12'h436;
        src10 <= 12'h4ca;
        src11 <= 12'h21b;
        src12 <= 12'hdf9;
        src13 <= 12'h601;
        src14 <= 12'hd5b;
        src15 <= 12'he42;
        src16 <= 12'h873;
        src17 <= 12'hebc;
        src18 <= 12'h7c4;
        src19 <= 12'h857;
        src20 <= 12'h5c6;
        src21 <= 12'hdb4;
        src22 <= 12'h934;
        src23 <= 12'h3a8;
        src24 <= 12'hd8c;
        src25 <= 12'h8e2;
        src26 <= 12'h205;
        src27 <= 12'h818;
        src28 <= 12'h99c;
        src29 <= 12'h9f8;
        src30 <= 12'h628;
        src31 <= 12'h3c0;
        src32 <= 12'h643;
        src33 <= 12'hc75;
        src34 <= 12'hf88;
        src35 <= 12'h6ec;
        src36 <= 12'h954;
        src37 <= 12'ha38;
        src38 <= 12'h432;
        src39 <= 12'h747;
        src40 <= 12'h385;
        src41 <= 12'h305;
        src42 <= 12'hc76;
        src43 <= 12'h258;
        src44 <= 12'h62b;
        src45 <= 12'hdef;
        src46 <= 12'he4d;
        src47 <= 12'hfd3;
        src48 <= 12'ha33;
        src49 <= 12'hdd4;
        src50 <= 12'hf6;
        src51 <= 12'h95b;
        src52 <= 12'h70f;
        src53 <= 12'h67b;
        src54 <= 12'hbbb;
        src55 <= 12'h555;
        src56 <= 12'h756;
        src57 <= 12'h11e;
        src58 <= 12'hc7e;
        src59 <= 12'hed8;
        src60 <= 12'h74b;
        src61 <= 12'h2fc;
        src62 <= 12'hc0;
        src63 <= 12'hbce;
        exp <= 18'h209e2;
        #1
        src0 <= 12'h1fe;
        src1 <= 12'h143;
        src2 <= 12'h80e;
        src3 <= 12'h786;
        src4 <= 12'h615;
        src5 <= 12'h29e;
        src6 <= 12'h36c;
        src7 <= 12'hc54;
        src8 <= 12'h124;
        src9 <= 12'h58b;
        src10 <= 12'h778;
        src11 <= 12'haa6;
        src12 <= 12'h1e4;
        src13 <= 12'h1f3;
        src14 <= 12'h37;
        src15 <= 12'h9d3;
        src16 <= 12'h3b6;
        src17 <= 12'h5;
        src18 <= 12'hdba;
        src19 <= 12'hcba;
        src20 <= 12'hfe6;
        src21 <= 12'h4ae;
        src22 <= 12'he;
        src23 <= 12'h8e3;
        src24 <= 12'h297;
        src25 <= 12'h1b1;
        src26 <= 12'he94;
        src27 <= 12'h55b;
        src28 <= 12'hb14;
        src29 <= 12'h74a;
        src30 <= 12'h4a0;
        src31 <= 12'hae6;
        src32 <= 12'h519;
        src33 <= 12'h89e;
        src34 <= 12'hfd2;
        src35 <= 12'h6c4;
        src36 <= 12'h326;
        src37 <= 12'h67;
        src38 <= 12'h32e;
        src39 <= 12'hfec;
        src40 <= 12'he00;
        src41 <= 12'he4e;
        src42 <= 12'hc61;
        src43 <= 12'h7e0;
        src44 <= 12'h9a8;
        src45 <= 12'ha8d;
        src46 <= 12'h486;
        src47 <= 12'hac8;
        src48 <= 12'hcc9;
        src49 <= 12'ha64;
        src50 <= 12'h801;
        src51 <= 12'hd;
        src52 <= 12'hc05;
        src53 <= 12'h3bb;
        src54 <= 12'h847;
        src55 <= 12'he6e;
        src56 <= 12'h60d;
        src57 <= 12'hdc0;
        src58 <= 12'h82;
        src59 <= 12'h945;
        src60 <= 12'hff5;
        src61 <= 12'hd3a;
        src62 <= 12'h97f;
        src63 <= 12'hcb5;
        exp <= 18'h1ed72;
        #1
        src0 <= 12'h299;
        src1 <= 12'hb3f;
        src2 <= 12'h1e3;
        src3 <= 12'hbee;
        src4 <= 12'hdf5;
        src5 <= 12'he83;
        src6 <= 12'h51d;
        src7 <= 12'hed6;
        src8 <= 12'he0f;
        src9 <= 12'hdba;
        src10 <= 12'h6b2;
        src11 <= 12'hc0a;
        src12 <= 12'h2f;
        src13 <= 12'hf5c;
        src14 <= 12'h20c;
        src15 <= 12'h2d7;
        src16 <= 12'h63a;
        src17 <= 12'hf40;
        src18 <= 12'hcc8;
        src19 <= 12'ha8a;
        src20 <= 12'h68;
        src21 <= 12'hbd9;
        src22 <= 12'h264;
        src23 <= 12'h5d6;
        src24 <= 12'h83a;
        src25 <= 12'hc3;
        src26 <= 12'h92d;
        src27 <= 12'h5d0;
        src28 <= 12'h6ae;
        src29 <= 12'hc9b;
        src30 <= 12'h7d2;
        src31 <= 12'he61;
        src32 <= 12'h586;
        src33 <= 12'h4ba;
        src34 <= 12'h6ff;
        src35 <= 12'h609;
        src36 <= 12'hd32;
        src37 <= 12'h7f3;
        src38 <= 12'h57b;
        src39 <= 12'hf5f;
        src40 <= 12'h53d;
        src41 <= 12'h7f1;
        src42 <= 12'h559;
        src43 <= 12'h97;
        src44 <= 12'h546;
        src45 <= 12'h1e7;
        src46 <= 12'hd41;
        src47 <= 12'h38f;
        src48 <= 12'h6c8;
        src49 <= 12'h33c;
        src50 <= 12'h3cd;
        src51 <= 12'h242;
        src52 <= 12'h32a;
        src53 <= 12'h1d5;
        src54 <= 12'he3;
        src55 <= 12'h419;
        src56 <= 12'h713;
        src57 <= 12'h533;
        src58 <= 12'h769;
        src59 <= 12'h8e0;
        src60 <= 12'h22;
        src61 <= 12'h89;
        src62 <= 12'hab6;
        src63 <= 12'heb7;
        exp <= 18'h1cedb;
        #1
        src0 <= 12'h705;
        src1 <= 12'h125;
        src2 <= 12'h10f;
        src3 <= 12'hcf3;
        src4 <= 12'hbb1;
        src5 <= 12'h69d;
        src6 <= 12'ha91;
        src7 <= 12'h83b;
        src8 <= 12'hb43;
        src9 <= 12'hc9a;
        src10 <= 12'h15d;
        src11 <= 12'h4b9;
        src12 <= 12'hb7c;
        src13 <= 12'h51c;
        src14 <= 12'h8ff;
        src15 <= 12'h602;
        src16 <= 12'hb5f;
        src17 <= 12'hde3;
        src18 <= 12'h61a;
        src19 <= 12'h74c;
        src20 <= 12'h6e9;
        src21 <= 12'h5ee;
        src22 <= 12'haa9;
        src23 <= 12'h56f;
        src24 <= 12'h541;
        src25 <= 12'hffc;
        src26 <= 12'h1f6;
        src27 <= 12'h573;
        src28 <= 12'h56c;
        src29 <= 12'h256;
        src30 <= 12'h52a;
        src31 <= 12'h3d3;
        src32 <= 12'h883;
        src33 <= 12'h4ba;
        src34 <= 12'hf40;
        src35 <= 12'h21a;
        src36 <= 12'h426;
        src37 <= 12'he3;
        src38 <= 12'h248;
        src39 <= 12'h1e2;
        src40 <= 12'h75a;
        src41 <= 12'h724;
        src42 <= 12'h8a3;
        src43 <= 12'hb93;
        src44 <= 12'h69a;
        src45 <= 12'hcbe;
        src46 <= 12'h546;
        src47 <= 12'h7ae;
        src48 <= 12'h9dd;
        src49 <= 12'h66b;
        src50 <= 12'he5e;
        src51 <= 12'hd6f;
        src52 <= 12'h263;
        src53 <= 12'h675;
        src54 <= 12'hc6b;
        src55 <= 12'hf73;
        src56 <= 12'h5e4;
        src57 <= 12'h997;
        src58 <= 12'h36e;
        src59 <= 12'h37e;
        src60 <= 12'h89b;
        src61 <= 12'h4ee;
        src62 <= 12'h730;
        src63 <= 12'h607;
        exp <= 18'h1d68a;
        #1
        src0 <= 12'h17;
        src1 <= 12'h484;
        src2 <= 12'h9f2;
        src3 <= 12'h30a;
        src4 <= 12'h4a3;
        src5 <= 12'h382;
        src6 <= 12'hd4b;
        src7 <= 12'hbde;
        src8 <= 12'hb7c;
        src9 <= 12'h9c9;
        src10 <= 12'ha3f;
        src11 <= 12'hf0a;
        src12 <= 12'h464;
        src13 <= 12'h2a0;
        src14 <= 12'ha26;
        src15 <= 12'he7;
        src16 <= 12'h91;
        src17 <= 12'hcbc;
        src18 <= 12'h521;
        src19 <= 12'h8c9;
        src20 <= 12'h181;
        src21 <= 12'h9b6;
        src22 <= 12'he55;
        src23 <= 12'ha5;
        src24 <= 12'h2c6;
        src25 <= 12'h2d2;
        src26 <= 12'h36d;
        src27 <= 12'h317;
        src28 <= 12'h7df;
        src29 <= 12'ha6e;
        src30 <= 12'hbe;
        src31 <= 12'h48e;
        src32 <= 12'h95;
        src33 <= 12'h4f7;
        src34 <= 12'hd24;
        src35 <= 12'h123;
        src36 <= 12'h11b;
        src37 <= 12'h8d0;
        src38 <= 12'h2e;
        src39 <= 12'hf88;
        src40 <= 12'h6e7;
        src41 <= 12'ha50;
        src42 <= 12'hbc5;
        src43 <= 12'h547;
        src44 <= 12'h351;
        src45 <= 12'h952;
        src46 <= 12'h21f;
        src47 <= 12'hedc;
        src48 <= 12'hd70;
        src49 <= 12'hc46;
        src50 <= 12'h4ac;
        src51 <= 12'hb6a;
        src52 <= 12'he6e;
        src53 <= 12'h251;
        src54 <= 12'h57b;
        src55 <= 12'ha09;
        src56 <= 12'h3be;
        src57 <= 12'hcbc;
        src58 <= 12'h1af;
        src59 <= 12'h638;
        src60 <= 12'hcb2;
        src61 <= 12'haf7;
        src62 <= 12'hc07;
        src63 <= 12'h402;
        exp <= 18'h1c418;
        #1
        src0 <= 12'h5e0;
        src1 <= 12'h830;
        src2 <= 12'h526;
        src3 <= 12'h7ba;
        src4 <= 12'hf8b;
        src5 <= 12'h517;
        src6 <= 12'haf3;
        src7 <= 12'h984;
        src8 <= 12'h573;
        src9 <= 12'he5f;
        src10 <= 12'hf8;
        src11 <= 12'heb0;
        src12 <= 12'hdfc;
        src13 <= 12'h2ba;
        src14 <= 12'hf71;
        src15 <= 12'hf6c;
        src16 <= 12'h42;
        src17 <= 12'hf3e;
        src18 <= 12'h46b;
        src19 <= 12'h94c;
        src20 <= 12'h498;
        src21 <= 12'h8c8;
        src22 <= 12'hf83;
        src23 <= 12'h7a2;
        src24 <= 12'h667;
        src25 <= 12'h4db;
        src26 <= 12'h2ee;
        src27 <= 12'hb0c;
        src28 <= 12'hd50;
        src29 <= 12'h78c;
        src30 <= 12'h8e;
        src31 <= 12'hc4a;
        src32 <= 12'h7de;
        src33 <= 12'h984;
        src34 <= 12'h4b6;
        src35 <= 12'hefe;
        src36 <= 12'h97f;
        src37 <= 12'hd61;
        src38 <= 12'h34f;
        src39 <= 12'hefc;
        src40 <= 12'ha14;
        src41 <= 12'hae;
        src42 <= 12'hdaa;
        src43 <= 12'h39e;
        src44 <= 12'hc09;
        src45 <= 12'h4eb;
        src46 <= 12'ha23;
        src47 <= 12'h753;
        src48 <= 12'h36e;
        src49 <= 12'hbbe;
        src50 <= 12'h2b9;
        src51 <= 12'h1eb;
        src52 <= 12'h91c;
        src53 <= 12'hcdc;
        src54 <= 12'hc7f;
        src55 <= 12'h8d1;
        src56 <= 12'h301;
        src57 <= 12'h5b5;
        src58 <= 12'hc41;
        src59 <= 12'hd1e;
        src60 <= 12'hcbf;
        src61 <= 12'h2ce;
        src62 <= 12'h201;
        src63 <= 12'h780;
        exp <= 18'h21ab2;
        #1
        src0 <= 12'h322;
        src1 <= 12'h57a;
        src2 <= 12'h70c;
        src3 <= 12'he28;
        src4 <= 12'h35;
        src5 <= 12'h70b;
        src6 <= 12'hae1;
        src7 <= 12'h9da;
        src8 <= 12'h11;
        src9 <= 12'hc5e;
        src10 <= 12'h43;
        src11 <= 12'h79a;
        src12 <= 12'hf6f;
        src13 <= 12'heda;
        src14 <= 12'hfee;
        src15 <= 12'haa1;
        src16 <= 12'he24;
        src17 <= 12'haf;
        src18 <= 12'h141;
        src19 <= 12'hb57;
        src20 <= 12'h489;
        src21 <= 12'h4a5;
        src22 <= 12'h31;
        src23 <= 12'hd86;
        src24 <= 12'hf5f;
        src25 <= 12'h7a6;
        src26 <= 12'h8f8;
        src27 <= 12'h6b;
        src28 <= 12'h11d;
        src29 <= 12'h38e;
        src30 <= 12'h8ec;
        src31 <= 12'h4ec;
        src32 <= 12'h136;
        src33 <= 12'h358;
        src34 <= 12'h107;
        src35 <= 12'ha5a;
        src36 <= 12'h9cb;
        src37 <= 12'h878;
        src38 <= 12'h96f;
        src39 <= 12'h60e;
        src40 <= 12'hade;
        src41 <= 12'h78;
        src42 <= 12'hbef;
        src43 <= 12'hf8c;
        src44 <= 12'h5a2;
        src45 <= 12'he26;
        src46 <= 12'habd;
        src47 <= 12'hdd4;
        src48 <= 12'h14f;
        src49 <= 12'h6ae;
        src50 <= 12'hea4;
        src51 <= 12'h41a;
        src52 <= 12'h5e2;
        src53 <= 12'h8f8;
        src54 <= 12'he8d;
        src55 <= 12'h107;
        src56 <= 12'hc30;
        src57 <= 12'h486;
        src58 <= 12'hc71;
        src59 <= 12'h8dc;
        src60 <= 12'he87;
        src61 <= 12'h455;
        src62 <= 12'hb2b;
        src63 <= 12'hfee;
        exp <= 18'h1fe24;
        #1
        src0 <= 12'hcba;
        src1 <= 12'h7be;
        src2 <= 12'h117;
        src3 <= 12'hc7e;
        src4 <= 12'hd68;
        src5 <= 12'had8;
        src6 <= 12'h949;
        src7 <= 12'h1d1;
        src8 <= 12'h971;
        src9 <= 12'h3e2;
        src10 <= 12'h58;
        src11 <= 12'h34c;
        src12 <= 12'h76c;
        src13 <= 12'ha4;
        src14 <= 12'h5b2;
        src15 <= 12'hc9b;
        src16 <= 12'h85f;
        src17 <= 12'hab8;
        src18 <= 12'h461;
        src19 <= 12'h84d;
        src20 <= 12'heb7;
        src21 <= 12'h5d5;
        src22 <= 12'h79d;
        src23 <= 12'hf53;
        src24 <= 12'hf68;
        src25 <= 12'h363;
        src26 <= 12'ha6f;
        src27 <= 12'h829;
        src28 <= 12'h56d;
        src29 <= 12'ha6a;
        src30 <= 12'h38f;
        src31 <= 12'h6d5;
        src32 <= 12'h26;
        src33 <= 12'hbeb;
        src34 <= 12'h8ca;
        src35 <= 12'h972;
        src36 <= 12'h31a;
        src37 <= 12'h239;
        src38 <= 12'hb79;
        src39 <= 12'h4a8;
        src40 <= 12'ha7b;
        src41 <= 12'h16e;
        src42 <= 12'h776;
        src43 <= 12'h344;
        src44 <= 12'heb3;
        src45 <= 12'h8e2;
        src46 <= 12'h3c;
        src47 <= 12'hfde;
        src48 <= 12'he18;
        src49 <= 12'haab;
        src50 <= 12'he0a;
        src51 <= 12'h8a3;
        src52 <= 12'h8fb;
        src53 <= 12'h3d5;
        src54 <= 12'h1d6;
        src55 <= 12'h328;
        src56 <= 12'h390;
        src57 <= 12'h97b;
        src58 <= 12'h9b1;
        src59 <= 12'h14a;
        src60 <= 12'h163;
        src61 <= 12'hd39;
        src62 <= 12'h9e5;
        src63 <= 12'h157;
        exp <= 18'h1e0c9;
        #1
        src0 <= 12'hb1c;
        src1 <= 12'h8c4;
        src2 <= 12'h744;
        src3 <= 12'hff0;
        src4 <= 12'h16a;
        src5 <= 12'h409;
        src6 <= 12'h976;
        src7 <= 12'h1d0;
        src8 <= 12'h6ef;
        src9 <= 12'hd1a;
        src10 <= 12'h6e5;
        src11 <= 12'hfc8;
        src12 <= 12'hdef;
        src13 <= 12'h5e;
        src14 <= 12'h26f;
        src15 <= 12'hd2c;
        src16 <= 12'h7b8;
        src17 <= 12'hc47;
        src18 <= 12'h32f;
        src19 <= 12'haf3;
        src20 <= 12'ha58;
        src21 <= 12'hed8;
        src22 <= 12'hb89;
        src23 <= 12'h3dd;
        src24 <= 12'h125;
        src25 <= 12'h9fb;
        src26 <= 12'h44a;
        src27 <= 12'h7e6;
        src28 <= 12'ha7;
        src29 <= 12'hc2;
        src30 <= 12'h3b9;
        src31 <= 12'h9c8;
        src32 <= 12'hf5b;
        src33 <= 12'hae;
        src34 <= 12'h7cb;
        src35 <= 12'h9a9;
        src36 <= 12'hb28;
        src37 <= 12'hf2c;
        src38 <= 12'h80a;
        src39 <= 12'h54f;
        src40 <= 12'hc30;
        src41 <= 12'h9ab;
        src42 <= 12'h70a;
        src43 <= 12'hc65;
        src44 <= 12'h2c0;
        src45 <= 12'h410;
        src46 <= 12'h906;
        src47 <= 12'h561;
        src48 <= 12'h2ce;
        src49 <= 12'hc85;
        src50 <= 12'hc22;
        src51 <= 12'he6e;
        src52 <= 12'h600;
        src53 <= 12'he3d;
        src54 <= 12'hf9e;
        src55 <= 12'hb62;
        src56 <= 12'h6fc;
        src57 <= 12'hd67;
        src58 <= 12'heb8;
        src59 <= 12'had;
        src60 <= 12'ha32;
        src61 <= 12'h8c2;
        src62 <= 12'hc34;
        src63 <= 12'ha37;
        exp <= 18'h2234e;
        #1
        src0 <= 12'h97f;
        src1 <= 12'h5b8;
        src2 <= 12'h1b0;
        src3 <= 12'h746;
        src4 <= 12'h355;
        src5 <= 12'h197;
        src6 <= 12'h2ee;
        src7 <= 12'h52b;
        src8 <= 12'hfb3;
        src9 <= 12'hc41;
        src10 <= 12'he90;
        src11 <= 12'hff1;
        src12 <= 12'he26;
        src13 <= 12'h15e;
        src14 <= 12'hf0;
        src15 <= 12'h523;
        src16 <= 12'h857;
        src17 <= 12'hb3;
        src18 <= 12'ha2;
        src19 <= 12'h396;
        src20 <= 12'hab6;
        src21 <= 12'h787;
        src22 <= 12'h6e4;
        src23 <= 12'ha20;
        src24 <= 12'hf17;
        src25 <= 12'h268;
        src26 <= 12'hb80;
        src27 <= 12'h56a;
        src28 <= 12'hfbc;
        src29 <= 12'h9db;
        src30 <= 12'hdd8;
        src31 <= 12'h8d0;
        src32 <= 12'hc9e;
        src33 <= 12'he63;
        src34 <= 12'h95;
        src35 <= 12'h476;
        src36 <= 12'h1c8;
        src37 <= 12'hcaa;
        src38 <= 12'h635;
        src39 <= 12'h2f9;
        src40 <= 12'h19b;
        src41 <= 12'h8da;
        src42 <= 12'h3d3;
        src43 <= 12'h67e;
        src44 <= 12'h7b0;
        src45 <= 12'h6c5;
        src46 <= 12'h5a7;
        src47 <= 12'h9d4;
        src48 <= 12'h1df;
        src49 <= 12'h4f4;
        src50 <= 12'he66;
        src51 <= 12'hf15;
        src52 <= 12'he17;
        src53 <= 12'h781;
        src54 <= 12'h33e;
        src55 <= 12'hb70;
        src56 <= 12'haea;
        src57 <= 12'h983;
        src58 <= 12'h7a6;
        src59 <= 12'hd3e;
        src60 <= 12'h4cb;
        src61 <= 12'h266;
        src62 <= 12'h92b;
        src63 <= 12'h603;
        exp <= 18'h1eb0f;
        #1
        src0 <= 12'hbbc;
        src1 <= 12'h984;
        src2 <= 12'h73f;
        src3 <= 12'h10e;
        src4 <= 12'h28d;
        src5 <= 12'h918;
        src6 <= 12'hb44;
        src7 <= 12'hff4;
        src8 <= 12'h81f;
        src9 <= 12'he7e;
        src10 <= 12'h82e;
        src11 <= 12'h190;
        src12 <= 12'h9f2;
        src13 <= 12'h6e;
        src14 <= 12'h834;
        src15 <= 12'h9bc;
        src16 <= 12'h5b0;
        src17 <= 12'h25c;
        src18 <= 12'h7e5;
        src19 <= 12'hb53;
        src20 <= 12'ha10;
        src21 <= 12'ha22;
        src22 <= 12'hfd;
        src23 <= 12'h683;
        src24 <= 12'he16;
        src25 <= 12'hc3f;
        src26 <= 12'h50;
        src27 <= 12'h689;
        src28 <= 12'h7a0;
        src29 <= 12'h23e;
        src30 <= 12'h5e1;
        src31 <= 12'hcab;
        src32 <= 12'hb42;
        src33 <= 12'h97;
        src34 <= 12'h142;
        src35 <= 12'h53a;
        src36 <= 12'h7c9;
        src37 <= 12'hde1;
        src38 <= 12'h451;
        src39 <= 12'h6fe;
        src40 <= 12'h6f5;
        src41 <= 12'hece;
        src42 <= 12'h3b2;
        src43 <= 12'h4e7;
        src44 <= 12'hcb8;
        src45 <= 12'hd4f;
        src46 <= 12'hf7d;
        src47 <= 12'hd6f;
        src48 <= 12'hdc0;
        src49 <= 12'hcf5;
        src50 <= 12'h465;
        src51 <= 12'h4f;
        src52 <= 12'ha2f;
        src53 <= 12'h65b;
        src54 <= 12'h93d;
        src55 <= 12'h85b;
        src56 <= 12'h1c7;
        src57 <= 12'h6fd;
        src58 <= 12'h98f;
        src59 <= 12'he0c;
        src60 <= 12'h3c8;
        src61 <= 12'hc81;
        src62 <= 12'h419;
        src63 <= 12'h780;
        exp <= 18'h1fc0c;
        #1
        src0 <= 12'h35;
        src1 <= 12'h58e;
        src2 <= 12'hf34;
        src3 <= 12'h948;
        src4 <= 12'hb16;
        src5 <= 12'h9b7;
        src6 <= 12'h93d;
        src7 <= 12'h329;
        src8 <= 12'h54f;
        src9 <= 12'had3;
        src10 <= 12'h818;
        src11 <= 12'h6ee;
        src12 <= 12'he72;
        src13 <= 12'h6ce;
        src14 <= 12'hdb0;
        src15 <= 12'hf6;
        src16 <= 12'hd3;
        src17 <= 12'h892;
        src18 <= 12'h40;
        src19 <= 12'h2b5;
        src20 <= 12'h674;
        src21 <= 12'hfcc;
        src22 <= 12'hee9;
        src23 <= 12'he46;
        src24 <= 12'h200;
        src25 <= 12'hb62;
        src26 <= 12'hab5;
        src27 <= 12'h988;
        src28 <= 12'hff4;
        src29 <= 12'h789;
        src30 <= 12'ha14;
        src31 <= 12'h7a1;
        src32 <= 12'h808;
        src33 <= 12'h6f3;
        src34 <= 12'h97d;
        src35 <= 12'hf76;
        src36 <= 12'h316;
        src37 <= 12'h815;
        src38 <= 12'h815;
        src39 <= 12'h34;
        src40 <= 12'hfbe;
        src41 <= 12'h9ee;
        src42 <= 12'he15;
        src43 <= 12'h51;
        src44 <= 12'h6b5;
        src45 <= 12'h5b6;
        src46 <= 12'h6b2;
        src47 <= 12'h39;
        src48 <= 12'heb7;
        src49 <= 12'hf5c;
        src50 <= 12'hb24;
        src51 <= 12'hf4d;
        src52 <= 12'hfe6;
        src53 <= 12'h64;
        src54 <= 12'he04;
        src55 <= 12'hc74;
        src56 <= 12'hc50;
        src57 <= 12'hde2;
        src58 <= 12'h62a;
        src59 <= 12'h3d;
        src60 <= 12'h13a;
        src61 <= 12'h7c2;
        src62 <= 12'he79;
        src63 <= 12'h2b6;
        exp <= 18'h221ee;
        #1
        src0 <= 12'he2e;
        src1 <= 12'h24;
        src2 <= 12'h8a5;
        src3 <= 12'hc63;
        src4 <= 12'h444;
        src5 <= 12'h6c3;
        src6 <= 12'h9a5;
        src7 <= 12'h722;
        src8 <= 12'h19c;
        src9 <= 12'h6b7;
        src10 <= 12'hb41;
        src11 <= 12'heac;
        src12 <= 12'h1d1;
        src13 <= 12'h3d1;
        src14 <= 12'h70d;
        src15 <= 12'h96f;
        src16 <= 12'hf20;
        src17 <= 12'h13e;
        src18 <= 12'he34;
        src19 <= 12'h908;
        src20 <= 12'hbcc;
        src21 <= 12'hf16;
        src22 <= 12'hba0;
        src23 <= 12'h16e;
        src24 <= 12'h10c;
        src25 <= 12'h46c;
        src26 <= 12'h459;
        src27 <= 12'ha2;
        src28 <= 12'h30f;
        src29 <= 12'h6a5;
        src30 <= 12'hf3f;
        src31 <= 12'h8de;
        src32 <= 12'h89b;
        src33 <= 12'h425;
        src34 <= 12'h8a3;
        src35 <= 12'hb9a;
        src36 <= 12'hd74;
        src37 <= 12'h69d;
        src38 <= 12'h489;
        src39 <= 12'h752;
        src40 <= 12'h82d;
        src41 <= 12'he25;
        src42 <= 12'h492;
        src43 <= 12'he5a;
        src44 <= 12'hb5e;
        src45 <= 12'ha59;
        src46 <= 12'hef5;
        src47 <= 12'hd26;
        src48 <= 12'h914;
        src49 <= 12'hc6f;
        src50 <= 12'h57c;
        src51 <= 12'hb2b;
        src52 <= 12'hb0e;
        src53 <= 12'h461;
        src54 <= 12'hd03;
        src55 <= 12'h32b;
        src56 <= 12'h965;
        src57 <= 12'h77c;
        src58 <= 12'hd82;
        src59 <= 12'hece;
        src60 <= 12'h8c5;
        src61 <= 12'hc1e;
        src62 <= 12'h666;
        src63 <= 12'h53;
        exp <= 18'h21de1;
        #1
        src0 <= 12'h8f9;
        src1 <= 12'h2a6;
        src2 <= 12'h42b;
        src3 <= 12'h825;
        src4 <= 12'h4a7;
        src5 <= 12'h8e;
        src6 <= 12'he09;
        src7 <= 12'hfc2;
        src8 <= 12'h6de;
        src9 <= 12'ha6d;
        src10 <= 12'h396;
        src11 <= 12'h725;
        src12 <= 12'h678;
        src13 <= 12'h27e;
        src14 <= 12'h7b7;
        src15 <= 12'h474;
        src16 <= 12'h1e2;
        src17 <= 12'h581;
        src18 <= 12'hb94;
        src19 <= 12'hc90;
        src20 <= 12'h94f;
        src21 <= 12'hdba;
        src22 <= 12'hcbc;
        src23 <= 12'h44;
        src24 <= 12'hc56;
        src25 <= 12'hd0;
        src26 <= 12'h898;
        src27 <= 12'h329;
        src28 <= 12'hd5f;
        src29 <= 12'h5d7;
        src30 <= 12'h7a8;
        src31 <= 12'h504;
        src32 <= 12'h61f;
        src33 <= 12'h622;
        src34 <= 12'h440;
        src35 <= 12'h4c7;
        src36 <= 12'hee0;
        src37 <= 12'h41c;
        src38 <= 12'ha91;
        src39 <= 12'hf48;
        src40 <= 12'hfcb;
        src41 <= 12'hd1b;
        src42 <= 12'ha63;
        src43 <= 12'hcc1;
        src44 <= 12'h481;
        src45 <= 12'h15b;
        src46 <= 12'hcb1;
        src47 <= 12'hfc;
        src48 <= 12'h4d7;
        src49 <= 12'h944;
        src50 <= 12'h9ca;
        src51 <= 12'h559;
        src52 <= 12'hc3b;
        src53 <= 12'h249;
        src54 <= 12'hcab;
        src55 <= 12'h2dd;
        src56 <= 12'hf42;
        src57 <= 12'hbc5;
        src58 <= 12'hf3c;
        src59 <= 12'hd1a;
        src60 <= 12'h6f5;
        src61 <= 12'he7c;
        src62 <= 12'h8c1;
        src63 <= 12'h351;
        exp <= 18'h20649;
        #1
        src0 <= 12'h5dc;
        src1 <= 12'h28d;
        src2 <= 12'h8a7;
        src3 <= 12'h482;
        src4 <= 12'h157;
        src5 <= 12'h72c;
        src6 <= 12'h998;
        src7 <= 12'h77a;
        src8 <= 12'haa;
        src9 <= 12'hafe;
        src10 <= 12'h955;
        src11 <= 12'h8b8;
        src12 <= 12'h909;
        src13 <= 12'hcea;
        src14 <= 12'hed9;
        src15 <= 12'h798;
        src16 <= 12'hc67;
        src17 <= 12'he6a;
        src18 <= 12'h55d;
        src19 <= 12'h153;
        src20 <= 12'h26b;
        src21 <= 12'hbed;
        src22 <= 12'hd53;
        src23 <= 12'haed;
        src24 <= 12'h44d;
        src25 <= 12'hac3;
        src26 <= 12'h64d;
        src27 <= 12'h3bc;
        src28 <= 12'h392;
        src29 <= 12'h340;
        src30 <= 12'h5;
        src31 <= 12'h167;
        src32 <= 12'h98c;
        src33 <= 12'h316;
        src34 <= 12'hc2b;
        src35 <= 12'h8cb;
        src36 <= 12'h37a;
        src37 <= 12'hbda;
        src38 <= 12'h970;
        src39 <= 12'h5bf;
        src40 <= 12'hb1f;
        src41 <= 12'h1d8;
        src42 <= 12'he28;
        src43 <= 12'hed;
        src44 <= 12'h789;
        src45 <= 12'hb5;
        src46 <= 12'ha38;
        src47 <= 12'h1a7;
        src48 <= 12'hb41;
        src49 <= 12'h101;
        src50 <= 12'h998;
        src51 <= 12'hce4;
        src52 <= 12'hed5;
        src53 <= 12'hebe;
        src54 <= 12'h2fe;
        src55 <= 12'h66f;
        src56 <= 12'hea8;
        src57 <= 12'hcc1;
        src58 <= 12'h723;
        src59 <= 12'h9aa;
        src60 <= 12'he1;
        src61 <= 12'hb11;
        src62 <= 12'ha87;
        src63 <= 12'h6e7;
        exp <= 18'h1e648;
        #1
        src0 <= 12'he31;
        src1 <= 12'h74f;
        src2 <= 12'h3b8;
        src3 <= 12'hb3;
        src4 <= 12'hc1f;
        src5 <= 12'h8fc;
        src6 <= 12'ha49;
        src7 <= 12'h3ca;
        src8 <= 12'he0d;
        src9 <= 12'h6db;
        src10 <= 12'h42;
        src11 <= 12'h81f;
        src12 <= 12'h32f;
        src13 <= 12'h762;
        src14 <= 12'h2fa;
        src15 <= 12'hda0;
        src16 <= 12'h3f7;
        src17 <= 12'h8c2;
        src18 <= 12'h285;
        src19 <= 12'h904;
        src20 <= 12'hb19;
        src21 <= 12'h892;
        src22 <= 12'hd41;
        src23 <= 12'hd40;
        src24 <= 12'h626;
        src25 <= 12'hbeb;
        src26 <= 12'h64f;
        src27 <= 12'hf38;
        src28 <= 12'h6a9;
        src29 <= 12'hdc0;
        src30 <= 12'h511;
        src31 <= 12'h610;
        src32 <= 12'hec0;
        src33 <= 12'h8bd;
        src34 <= 12'h91d;
        src35 <= 12'hed2;
        src36 <= 12'h4a6;
        src37 <= 12'he44;
        src38 <= 12'hd9e;
        src39 <= 12'h681;
        src40 <= 12'ha16;
        src41 <= 12'hef4;
        src42 <= 12'h6ef;
        src43 <= 12'h768;
        src44 <= 12'h745;
        src45 <= 12'hbc0;
        src46 <= 12'h38;
        src47 <= 12'h786;
        src48 <= 12'hb6f;
        src49 <= 12'ha22;
        src50 <= 12'h80f;
        src51 <= 12'h284;
        src52 <= 12'h481;
        src53 <= 12'h932;
        src54 <= 12'hc3b;
        src55 <= 12'h8d4;
        src56 <= 12'h6bf;
        src57 <= 12'hf49;
        src58 <= 12'h1e9;
        src59 <= 12'h62;
        src60 <= 12'hf24;
        src61 <= 12'he1c;
        src62 <= 12'h3b5;
        src63 <= 12'hcd;
        exp <= 18'h218b1;
        #1
        src0 <= 12'h855;
        src1 <= 12'h73c;
        src2 <= 12'h852;
        src3 <= 12'h5a7;
        src4 <= 12'hb1;
        src5 <= 12'h71f;
        src6 <= 12'h5e6;
        src7 <= 12'h23b;
        src8 <= 12'hb59;
        src9 <= 12'ha41;
        src10 <= 12'hd46;
        src11 <= 12'hbe2;
        src12 <= 12'hbe3;
        src13 <= 12'hbce;
        src14 <= 12'h766;
        src15 <= 12'h1f1;
        src16 <= 12'h713;
        src17 <= 12'h802;
        src18 <= 12'hf06;
        src19 <= 12'h97f;
        src20 <= 12'h750;
        src21 <= 12'h2cc;
        src22 <= 12'hcef;
        src23 <= 12'hd4b;
        src24 <= 12'h996;
        src25 <= 12'h614;
        src26 <= 12'hdde;
        src27 <= 12'h122;
        src28 <= 12'hc50;
        src29 <= 12'hd56;
        src30 <= 12'h33f;
        src31 <= 12'ha;
        src32 <= 12'h66a;
        src33 <= 12'h4eb;
        src34 <= 12'h65f;
        src35 <= 12'hc76;
        src36 <= 12'hf9f;
        src37 <= 12'h519;
        src38 <= 12'h3f9;
        src39 <= 12'hbc4;
        src40 <= 12'h4e3;
        src41 <= 12'h351;
        src42 <= 12'h76e;
        src43 <= 12'h35b;
        src44 <= 12'h950;
        src45 <= 12'h44f;
        src46 <= 12'h52f;
        src47 <= 12'h77d;
        src48 <= 12'h252;
        src49 <= 12'h3d4;
        src50 <= 12'h2d6;
        src51 <= 12'haf3;
        src52 <= 12'h12e;
        src53 <= 12'h5b4;
        src54 <= 12'h5ed;
        src55 <= 12'he52;
        src56 <= 12'hc05;
        src57 <= 12'h2be;
        src58 <= 12'hd53;
        src59 <= 12'h789;
        src60 <= 12'hf2a;
        src61 <= 12'h583;
        src62 <= 12'h2a6;
        src63 <= 12'h1e8;
        exp <= 18'h1e09f;
        #1
        src0 <= 12'h368;
        src1 <= 12'h8e5;
        src2 <= 12'h19d;
        src3 <= 12'h6a7;
        src4 <= 12'h68d;
        src5 <= 12'h5ec;
        src6 <= 12'hd73;
        src7 <= 12'hf21;
        src8 <= 12'h9a2;
        src9 <= 12'he20;
        src10 <= 12'h434;
        src11 <= 12'hb5b;
        src12 <= 12'h64a;
        src13 <= 12'h9d5;
        src14 <= 12'h612;
        src15 <= 12'hb85;
        src16 <= 12'hed7;
        src17 <= 12'h350;
        src18 <= 12'hb90;
        src19 <= 12'hc2c;
        src20 <= 12'h16d;
        src21 <= 12'hdb8;
        src22 <= 12'h90f;
        src23 <= 12'h58f;
        src24 <= 12'h610;
        src25 <= 12'h9a4;
        src26 <= 12'h75b;
        src27 <= 12'h521;
        src28 <= 12'h465;
        src29 <= 12'h2e8;
        src30 <= 12'he7b;
        src31 <= 12'hee7;
        src32 <= 12'h177;
        src33 <= 12'h471;
        src34 <= 12'h56f;
        src35 <= 12'h3a7;
        src36 <= 12'hec1;
        src37 <= 12'h22;
        src38 <= 12'haa4;
        src39 <= 12'hd51;
        src40 <= 12'h2fa;
        src41 <= 12'h4a9;
        src42 <= 12'h1f6;
        src43 <= 12'he63;
        src44 <= 12'h19f;
        src45 <= 12'h417;
        src46 <= 12'hb26;
        src47 <= 12'hbea;
        src48 <= 12'hbfc;
        src49 <= 12'h12b;
        src50 <= 12'h63f;
        src51 <= 12'h707;
        src52 <= 12'h76c;
        src53 <= 12'hc19;
        src54 <= 12'h2a3;
        src55 <= 12'h84a;
        src56 <= 12'h287;
        src57 <= 12'h9f7;
        src58 <= 12'h2e1;
        src59 <= 12'ha3;
        src60 <= 12'h63e;
        src61 <= 12'h14b;
        src62 <= 12'hc86;
        src63 <= 12'h3ac;
        exp <= 18'h1da5e;
        #1
        src0 <= 12'hd35;
        src1 <= 12'he7d;
        src2 <= 12'h3b6;
        src3 <= 12'h22b;
        src4 <= 12'h8e7;
        src5 <= 12'h2d4;
        src6 <= 12'h678;
        src7 <= 12'h9d7;
        src8 <= 12'hb3f;
        src9 <= 12'h92;
        src10 <= 12'h8c7;
        src11 <= 12'hd59;
        src12 <= 12'h41b;
        src13 <= 12'hf9d;
        src14 <= 12'h7fc;
        src15 <= 12'hd55;
        src16 <= 12'hea;
        src17 <= 12'h9e4;
        src18 <= 12'h1e5;
        src19 <= 12'h55;
        src20 <= 12'ha10;
        src21 <= 12'hf5d;
        src22 <= 12'hde0;
        src23 <= 12'hb4;
        src24 <= 12'he2c;
        src25 <= 12'hbe2;
        src26 <= 12'hdc6;
        src27 <= 12'h9e4;
        src28 <= 12'ha41;
        src29 <= 12'h1;
        src30 <= 12'h6df;
        src31 <= 12'h264;
        src32 <= 12'h48c;
        src33 <= 12'hd3;
        src34 <= 12'h243;
        src35 <= 12'ha22;
        src36 <= 12'h82;
        src37 <= 12'hb28;
        src38 <= 12'hdec;
        src39 <= 12'hc99;
        src40 <= 12'hba6;
        src41 <= 12'h56d;
        src42 <= 12'h9a9;
        src43 <= 12'hd22;
        src44 <= 12'h40;
        src45 <= 12'he36;
        src46 <= 12'h5ca;
        src47 <= 12'hbff;
        src48 <= 12'h134;
        src49 <= 12'h659;
        src50 <= 12'hb93;
        src51 <= 12'h47a;
        src52 <= 12'h855;
        src53 <= 12'h85e;
        src54 <= 12'hc;
        src55 <= 12'had7;
        src56 <= 12'hd0;
        src57 <= 12'hb70;
        src58 <= 12'h198;
        src59 <= 12'hba0;
        src60 <= 12'h748;
        src61 <= 12'h5d0;
        src62 <= 12'ha09;
        src63 <= 12'h1f9;
        exp <= 18'h1e8af;
        #1
        src0 <= 12'hc4e;
        src1 <= 12'hb8e;
        src2 <= 12'h1c5;
        src3 <= 12'ha2a;
        src4 <= 12'hffb;
        src5 <= 12'heae;
        src6 <= 12'hd0c;
        src7 <= 12'h332;
        src8 <= 12'he5f;
        src9 <= 12'h7ac;
        src10 <= 12'hffb;
        src11 <= 12'h6e4;
        src12 <= 12'h54f;
        src13 <= 12'hfe3;
        src14 <= 12'h6ef;
        src15 <= 12'h9d7;
        src16 <= 12'h117;
        src17 <= 12'h985;
        src18 <= 12'hc16;
        src19 <= 12'hdc1;
        src20 <= 12'ha58;
        src21 <= 12'hed4;
        src22 <= 12'hf98;
        src23 <= 12'h3d4;
        src24 <= 12'hfda;
        src25 <= 12'hebb;
        src26 <= 12'h596;
        src27 <= 12'hc9c;
        src28 <= 12'h2a2;
        src29 <= 12'h418;
        src30 <= 12'h46f;
        src31 <= 12'h982;
        src32 <= 12'hbd3;
        src33 <= 12'h63e;
        src34 <= 12'h7ba;
        src35 <= 12'hcd7;
        src36 <= 12'h73b;
        src37 <= 12'h386;
        src38 <= 12'he40;
        src39 <= 12'h525;
        src40 <= 12'h431;
        src41 <= 12'h939;
        src42 <= 12'h566;
        src43 <= 12'hd0b;
        src44 <= 12'h78;
        src45 <= 12'h7b1;
        src46 <= 12'hcd3;
        src47 <= 12'h269;
        src48 <= 12'hec7;
        src49 <= 12'h1a4;
        src50 <= 12'hf1d;
        src51 <= 12'h927;
        src52 <= 12'h812;
        src53 <= 12'hc24;
        src54 <= 12'hbb4;
        src55 <= 12'h428;
        src56 <= 12'hf9a;
        src57 <= 12'h99e;
        src58 <= 12'h2dc;
        src59 <= 12'h530;
        src60 <= 12'h3de;
        src61 <= 12'hacf;
        src62 <= 12'h570;
        src63 <= 12'h611;
        exp <= 18'h2404c;
        #1
        src0 <= 12'h141;
        src1 <= 12'h21;
        src2 <= 12'h44c;
        src3 <= 12'h62a;
        src4 <= 12'hefb;
        src5 <= 12'h816;
        src6 <= 12'h829;
        src7 <= 12'h173;
        src8 <= 12'h45;
        src9 <= 12'ha1b;
        src10 <= 12'h376;
        src11 <= 12'h241;
        src12 <= 12'h8ec;
        src13 <= 12'hf45;
        src14 <= 12'h3fa;
        src15 <= 12'h778;
        src16 <= 12'h435;
        src17 <= 12'h7c6;
        src18 <= 12'h838;
        src19 <= 12'hc89;
        src20 <= 12'h4ee;
        src21 <= 12'hb76;
        src22 <= 12'h843;
        src23 <= 12'h40c;
        src24 <= 12'h3a2;
        src25 <= 12'hadf;
        src26 <= 12'h2a2;
        src27 <= 12'hba0;
        src28 <= 12'h879;
        src29 <= 12'he7f;
        src30 <= 12'h253;
        src31 <= 12'hc3c;
        src32 <= 12'h112;
        src33 <= 12'h3f4;
        src34 <= 12'h99b;
        src35 <= 12'h972;
        src36 <= 12'hc3b;
        src37 <= 12'h5ec;
        src38 <= 12'h13a;
        src39 <= 12'h5c2;
        src40 <= 12'hee6;
        src41 <= 12'h331;
        src42 <= 12'h43b;
        src43 <= 12'h2a4;
        src44 <= 12'hd82;
        src45 <= 12'haf;
        src46 <= 12'h3d4;
        src47 <= 12'h778;
        src48 <= 12'h26;
        src49 <= 12'hc31;
        src50 <= 12'h73d;
        src51 <= 12'h431;
        src52 <= 12'h717;
        src53 <= 12'h42c;
        src54 <= 12'heb;
        src55 <= 12'h3b9;
        src56 <= 12'he4;
        src57 <= 12'h4f5;
        src58 <= 12'hda3;
        src59 <= 12'h165;
        src60 <= 12'h34d;
        src61 <= 12'hcee;
        src62 <= 12'h2b0;
        src63 <= 12'ha5e;
        exp <= 18'h19d77;
        #1
        src0 <= 12'h997;
        src1 <= 12'h4b7;
        src2 <= 12'hf49;
        src3 <= 12'hb35;
        src4 <= 12'h67b;
        src5 <= 12'h3c1;
        src6 <= 12'h88b;
        src7 <= 12'h9be;
        src8 <= 12'hb69;
        src9 <= 12'h1bd;
        src10 <= 12'h483;
        src11 <= 12'hc49;
        src12 <= 12'hdf0;
        src13 <= 12'hdba;
        src14 <= 12'h1a3;
        src15 <= 12'h327;
        src16 <= 12'h99;
        src17 <= 12'h2c9;
        src18 <= 12'h269;
        src19 <= 12'ha16;
        src20 <= 12'h47f;
        src21 <= 12'h87c;
        src22 <= 12'h522;
        src23 <= 12'haa8;
        src24 <= 12'ha23;
        src25 <= 12'h2d1;
        src26 <= 12'h312;
        src27 <= 12'hb0e;
        src28 <= 12'h6c;
        src29 <= 12'hd4f;
        src30 <= 12'h541;
        src31 <= 12'hdf5;
        src32 <= 12'h8d3;
        src33 <= 12'he40;
        src34 <= 12'h891;
        src35 <= 12'h9a4;
        src36 <= 12'hb46;
        src37 <= 12'h317;
        src38 <= 12'he35;
        src39 <= 12'h229;
        src40 <= 12'ha91;
        src41 <= 12'hbf6;
        src42 <= 12'hc3b;
        src43 <= 12'hc48;
        src44 <= 12'hf2d;
        src45 <= 12'h786;
        src46 <= 12'hb9e;
        src47 <= 12'ha30;
        src48 <= 12'hc7d;
        src49 <= 12'ha9d;
        src50 <= 12'h5e8;
        src51 <= 12'h5e4;
        src52 <= 12'h11e;
        src53 <= 12'hff4;
        src54 <= 12'h570;
        src55 <= 12'heac;
        src56 <= 12'hed0;
        src57 <= 12'hfdf;
        src58 <= 12'h4c4;
        src59 <= 12'h968;
        src60 <= 12'h240;
        src61 <= 12'h881;
        src62 <= 12'h7c8;
        src63 <= 12'h9d1;
        exp <= 18'h22139;
        #1
        src0 <= 12'h9d9;
        src1 <= 12'h785;
        src2 <= 12'h165;
        src3 <= 12'h4e7;
        src4 <= 12'h8a3;
        src5 <= 12'h15;
        src6 <= 12'h4ec;
        src7 <= 12'h491;
        src8 <= 12'h7b7;
        src9 <= 12'h817;
        src10 <= 12'hab9;
        src11 <= 12'h8ed;
        src12 <= 12'haae;
        src13 <= 12'ha03;
        src14 <= 12'h9c1;
        src15 <= 12'hdc2;
        src16 <= 12'h671;
        src17 <= 12'hed7;
        src18 <= 12'hb04;
        src19 <= 12'hc45;
        src20 <= 12'h75c;
        src21 <= 12'he32;
        src22 <= 12'h420;
        src23 <= 12'h32c;
        src24 <= 12'ha75;
        src25 <= 12'h2a7;
        src26 <= 12'h562;
        src27 <= 12'h9af;
        src28 <= 12'h7fe;
        src29 <= 12'h8d;
        src30 <= 12'h448;
        src31 <= 12'he88;
        src32 <= 12'h7b4;
        src33 <= 12'h28c;
        src34 <= 12'h1fb;
        src35 <= 12'h4e6;
        src36 <= 12'hf51;
        src37 <= 12'hdae;
        src38 <= 12'h1f5;
        src39 <= 12'h33e;
        src40 <= 12'h334;
        src41 <= 12'hf50;
        src42 <= 12'h938;
        src43 <= 12'h245;
        src44 <= 12'h6eb;
        src45 <= 12'h78a;
        src46 <= 12'h84;
        src47 <= 12'h7f7;
        src48 <= 12'hed2;
        src49 <= 12'ha04;
        src50 <= 12'he0f;
        src51 <= 12'hf2c;
        src52 <= 12'hd92;
        src53 <= 12'h3c9;
        src54 <= 12'hb60;
        src55 <= 12'h638;
        src56 <= 12'h252;
        src57 <= 12'h813;
        src58 <= 12'he1c;
        src59 <= 12'h977;
        src60 <= 12'hd16;
        src61 <= 12'hcec;
        src62 <= 12'hd9b;
        src63 <= 12'h1fa;
        exp <= 18'h20751;
        #1
        src0 <= 12'hc6c;
        src1 <= 12'h34e;
        src2 <= 12'he22;
        src3 <= 12'he77;
        src4 <= 12'hf33;
        src5 <= 12'he09;
        src6 <= 12'h90;
        src7 <= 12'h50f;
        src8 <= 12'h2ed;
        src9 <= 12'h9cc;
        src10 <= 12'h92e;
        src11 <= 12'h9dd;
        src12 <= 12'hf2a;
        src13 <= 12'h3d1;
        src14 <= 12'h395;
        src15 <= 12'hc6e;
        src16 <= 12'h802;
        src17 <= 12'hcb;
        src18 <= 12'h343;
        src19 <= 12'hbc;
        src20 <= 12'h99a;
        src21 <= 12'h908;
        src22 <= 12'h4e3;
        src23 <= 12'hd64;
        src24 <= 12'h3f5;
        src25 <= 12'h888;
        src26 <= 12'h6de;
        src27 <= 12'ha32;
        src28 <= 12'h882;
        src29 <= 12'h25f;
        src30 <= 12'hc4d;
        src31 <= 12'he63;
        src32 <= 12'hd21;
        src33 <= 12'hf7d;
        src34 <= 12'hcad;
        src35 <= 12'h48;
        src36 <= 12'h143;
        src37 <= 12'h20c;
        src38 <= 12'h7c5;
        src39 <= 12'h7bf;
        src40 <= 12'h170;
        src41 <= 12'hc3f;
        src42 <= 12'h651;
        src43 <= 12'he84;
        src44 <= 12'hde3;
        src45 <= 12'h342;
        src46 <= 12'h201;
        src47 <= 12'h502;
        src48 <= 12'h3b8;
        src49 <= 12'hf13;
        src50 <= 12'h5e1;
        src51 <= 12'hdf5;
        src52 <= 12'h81f;
        src53 <= 12'ha99;
        src54 <= 12'h9cf;
        src55 <= 12'hede;
        src56 <= 12'h741;
        src57 <= 12'h424;
        src58 <= 12'he05;
        src59 <= 12'hf3c;
        src60 <= 12'h805;
        src61 <= 12'hee;
        src62 <= 12'ha51;
        src63 <= 12'h5d1;
        exp <= 18'h21196;
        #1
        src0 <= 12'h21a;
        src1 <= 12'hf26;
        src2 <= 12'h20f;
        src3 <= 12'h71b;
        src4 <= 12'h612;
        src5 <= 12'h5f1;
        src6 <= 12'h208;
        src7 <= 12'he92;
        src8 <= 12'h4f3;
        src9 <= 12'hefc;
        src10 <= 12'h887;
        src11 <= 12'ha6c;
        src12 <= 12'h665;
        src13 <= 12'hf91;
        src14 <= 12'h4a2;
        src15 <= 12'hbe;
        src16 <= 12'h600;
        src17 <= 12'h7a3;
        src18 <= 12'h452;
        src19 <= 12'h43c;
        src20 <= 12'hedb;
        src21 <= 12'hb66;
        src22 <= 12'hf45;
        src23 <= 12'h1ef;
        src24 <= 12'hca3;
        src25 <= 12'hf53;
        src26 <= 12'h610;
        src27 <= 12'h9b1;
        src28 <= 12'h9f1;
        src29 <= 12'hf28;
        src30 <= 12'h46e;
        src31 <= 12'he57;
        src32 <= 12'h6d1;
        src33 <= 12'h577;
        src34 <= 12'h7f8;
        src35 <= 12'h23e;
        src36 <= 12'heba;
        src37 <= 12'ha3a;
        src38 <= 12'hbc3;
        src39 <= 12'h894;
        src40 <= 12'hbee;
        src41 <= 12'hfca;
        src42 <= 12'h4a8;
        src43 <= 12'h9c5;
        src44 <= 12'hbbc;
        src45 <= 12'hdd6;
        src46 <= 12'hc8d;
        src47 <= 12'h5a5;
        src48 <= 12'hf11;
        src49 <= 12'he2;
        src50 <= 12'h882;
        src51 <= 12'h169;
        src52 <= 12'he08;
        src53 <= 12'hdd6;
        src54 <= 12'hd80;
        src55 <= 12'h2f5;
        src56 <= 12'h10d;
        src57 <= 12'h5a0;
        src58 <= 12'h232;
        src59 <= 12'hcc4;
        src60 <= 12'h90d;
        src61 <= 12'hbb9;
        src62 <= 12'h118;
        src63 <= 12'h238;
        exp <= 18'h22016;
        #1
        src0 <= 12'hc;
        src1 <= 12'hb42;
        src2 <= 12'h581;
        src3 <= 12'h2f4;
        src4 <= 12'ha93;
        src5 <= 12'h705;
        src6 <= 12'heb5;
        src7 <= 12'hd98;
        src8 <= 12'hb79;
        src9 <= 12'h4e4;
        src10 <= 12'h6a4;
        src11 <= 12'h406;
        src12 <= 12'h7c8;
        src13 <= 12'h72d;
        src14 <= 12'h816;
        src15 <= 12'hdcb;
        src16 <= 12'h852;
        src17 <= 12'h1cf;
        src18 <= 12'h4b0;
        src19 <= 12'h351;
        src20 <= 12'h3aa;
        src21 <= 12'hf82;
        src22 <= 12'hcfe;
        src23 <= 12'h814;
        src24 <= 12'hee3;
        src25 <= 12'hf49;
        src26 <= 12'hace;
        src27 <= 12'hc20;
        src28 <= 12'hbdf;
        src29 <= 12'he5;
        src30 <= 12'h6c0;
        src31 <= 12'h16f;
        src32 <= 12'h780;
        src33 <= 12'hfbc;
        src34 <= 12'hd69;
        src35 <= 12'hd01;
        src36 <= 12'h590;
        src37 <= 12'h1b7;
        src38 <= 12'hf7a;
        src39 <= 12'h5bf;
        src40 <= 12'h3c5;
        src41 <= 12'hddd;
        src42 <= 12'hf04;
        src43 <= 12'hded;
        src44 <= 12'hb64;
        src45 <= 12'hec2;
        src46 <= 12'h85a;
        src47 <= 12'hdc9;
        src48 <= 12'h8d8;
        src49 <= 12'h7af;
        src50 <= 12'h626;
        src51 <= 12'h36d;
        src52 <= 12'hfeb;
        src53 <= 12'h158;
        src54 <= 12'h3b4;
        src55 <= 12'h4ce;
        src56 <= 12'hfba;
        src57 <= 12'h316;
        src58 <= 12'ha66;
        src59 <= 12'ha4f;
        src60 <= 12'h496;
        src61 <= 12'he23;
        src62 <= 12'h98b;
        src63 <= 12'hfd1;
        exp <= 18'h23a6d;
        #1
        src0 <= 12'hb44;
        src1 <= 12'h78e;
        src2 <= 12'hde3;
        src3 <= 12'ha5c;
        src4 <= 12'ha1b;
        src5 <= 12'h48b;
        src6 <= 12'h3d6;
        src7 <= 12'h854;
        src8 <= 12'hb6e;
        src9 <= 12'haba;
        src10 <= 12'h972;
        src11 <= 12'h5fa;
        src12 <= 12'hb5c;
        src13 <= 12'ha1f;
        src14 <= 12'hf2a;
        src15 <= 12'ha53;
        src16 <= 12'hbfc;
        src17 <= 12'h55e;
        src18 <= 12'h7f3;
        src19 <= 12'hf;
        src20 <= 12'h609;
        src21 <= 12'h5b8;
        src22 <= 12'heee;
        src23 <= 12'h7fe;
        src24 <= 12'h6c3;
        src25 <= 12'h1f3;
        src26 <= 12'hf01;
        src27 <= 12'h33a;
        src28 <= 12'h36e;
        src29 <= 12'hed4;
        src30 <= 12'h7d0;
        src31 <= 12'h71a;
        src32 <= 12'h547;
        src33 <= 12'he21;
        src34 <= 12'hc98;
        src35 <= 12'h4b4;
        src36 <= 12'h519;
        src37 <= 12'hb88;
        src38 <= 12'h2c5;
        src39 <= 12'hf16;
        src40 <= 12'h5ec;
        src41 <= 12'hd1e;
        src42 <= 12'h8d;
        src43 <= 12'h118;
        src44 <= 12'hbcd;
        src45 <= 12'he10;
        src46 <= 12'h3a0;
        src47 <= 12'h7c6;
        src48 <= 12'h287;
        src49 <= 12'hea1;
        src50 <= 12'h139;
        src51 <= 12'h1c1;
        src52 <= 12'h54b;
        src53 <= 12'ha7b;
        src54 <= 12'h424;
        src55 <= 12'h3f9;
        src56 <= 12'h21c;
        src57 <= 12'h34f;
        src58 <= 12'hbb;
        src59 <= 12'h9c3;
        src60 <= 12'hbe3;
        src61 <= 12'h1d6;
        src62 <= 12'hb2b;
        src63 <= 12'h3d0;
        exp <= 18'h1ec57;
        #1
        src0 <= 12'hdcb;
        src1 <= 12'h72;
        src2 <= 12'hc5e;
        src3 <= 12'h5bc;
        src4 <= 12'hdf8;
        src5 <= 12'h46;
        src6 <= 12'hc0b;
        src7 <= 12'h5ea;
        src8 <= 12'hbb5;
        src9 <= 12'hf60;
        src10 <= 12'h721;
        src11 <= 12'hf08;
        src12 <= 12'h63;
        src13 <= 12'hd8c;
        src14 <= 12'h641;
        src15 <= 12'h580;
        src16 <= 12'h48d;
        src17 <= 12'hff8;
        src18 <= 12'he29;
        src19 <= 12'hd3d;
        src20 <= 12'h5f7;
        src21 <= 12'h870;
        src22 <= 12'hcdd;
        src23 <= 12'hba3;
        src24 <= 12'hb13;
        src25 <= 12'hd90;
        src26 <= 12'h841;
        src27 <= 12'ha36;
        src28 <= 12'hf2d;
        src29 <= 12'hdb;
        src30 <= 12'hda1;
        src31 <= 12'h33f;
        src32 <= 12'h861;
        src33 <= 12'h1d7;
        src34 <= 12'h8df;
        src35 <= 12'ha98;
        src36 <= 12'h9dd;
        src37 <= 12'h16b;
        src38 <= 12'he67;
        src39 <= 12'hb38;
        src40 <= 12'hf65;
        src41 <= 12'h393;
        src42 <= 12'h378;
        src43 <= 12'hc3e;
        src44 <= 12'h421;
        src45 <= 12'hf08;
        src46 <= 12'ha32;
        src47 <= 12'h354;
        src48 <= 12'hfe0;
        src49 <= 12'h1cc;
        src50 <= 12'h995;
        src51 <= 12'h1a0;
        src52 <= 12'h721;
        src53 <= 12'h66b;
        src54 <= 12'h6a5;
        src55 <= 12'h529;
        src56 <= 12'h7f4;
        src57 <= 12'h462;
        src58 <= 12'had7;
        src59 <= 12'heae;
        src60 <= 12'h69b;
        src61 <= 12'h6b1;
        src62 <= 12'h797;
        src63 <= 12'h847;
        exp <= 18'h22d7f;
        #1
        src0 <= 12'h2b;
        src1 <= 12'he76;
        src2 <= 12'h9be;
        src3 <= 12'he0b;
        src4 <= 12'hd54;
        src5 <= 12'ha07;
        src6 <= 12'hbfd;
        src7 <= 12'h326;
        src8 <= 12'h33d;
        src9 <= 12'hef6;
        src10 <= 12'h2ce;
        src11 <= 12'h145;
        src12 <= 12'hc5f;
        src13 <= 12'hadb;
        src14 <= 12'h929;
        src15 <= 12'h987;
        src16 <= 12'h3aa;
        src17 <= 12'h3fa;
        src18 <= 12'hbaa;
        src19 <= 12'h452;
        src20 <= 12'h9e4;
        src21 <= 12'haaf;
        src22 <= 12'h78d;
        src23 <= 12'h2bb;
        src24 <= 12'hf2a;
        src25 <= 12'h67a;
        src26 <= 12'hc49;
        src27 <= 12'he9c;
        src28 <= 12'hba6;
        src29 <= 12'h6fc;
        src30 <= 12'h5a5;
        src31 <= 12'hc2d;
        src32 <= 12'h217;
        src33 <= 12'h6a8;
        src34 <= 12'h5ef;
        src35 <= 12'hb1f;
        src36 <= 12'hf22;
        src37 <= 12'h787;
        src38 <= 12'hd42;
        src39 <= 12'h1af;
        src40 <= 12'h5b0;
        src41 <= 12'h45b;
        src42 <= 12'haeb;
        src43 <= 12'hbcb;
        src44 <= 12'h7d1;
        src45 <= 12'hd9b;
        src46 <= 12'h44b;
        src47 <= 12'hdf0;
        src48 <= 12'hd1b;
        src49 <= 12'h5c5;
        src50 <= 12'h627;
        src51 <= 12'h218;
        src52 <= 12'h911;
        src53 <= 12'hb36;
        src54 <= 12'h529;
        src55 <= 12'hdb5;
        src56 <= 12'h38b;
        src57 <= 12'h4e9;
        src58 <= 12'ha8b;
        src59 <= 12'h559;
        src60 <= 12'h804;
        src61 <= 12'h6fd;
        src62 <= 12'h825;
        src63 <= 12'hf12;
        exp <= 18'h22133;
        #1
        $finish;
    end
endmodule

