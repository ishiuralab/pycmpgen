module gpc1_1(input src0, output dst0);
    assign dst0 = src0;
endmodule // gpc1_1
