module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [19:0] src21;
    reg [18:0] src22;
    reg [17:0] src23;
    reg [16:0] src24;
    reg [15:0] src25;
    reg [14:0] src26;
    reg [13:0] src27;
    reg [12:0] src28;
    reg [11:0] src29;
    reg [10:0] src30;
    reg [9:0] src31;
    reg [8:0] src32;
    reg [7:0] src33;
    reg [6:0] src34;
    reg [5:0] src35;
    reg [4:0] src36;
    reg [3:0] src37;
    reg [2:0] src38;
    reg [1:0] src39;
    reg [0:0] src40;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [41:0] srcsum;
    wire [41:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3])<<37) + ((src38[0] + src38[1] + src38[2])<<38) + ((src39[0] + src39[1])<<39) + ((src40[0])<<40);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc0f8501ca933627f45463a97baba1bba1f3befed7bbe09949de68ecf046703bdaac39aec75a043bab2e35211afc41f8a1b75626af63e71;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf31aad891c336b0253ed89c46d2c3b6bcb7aa37839735954ea38f319bf2fcbd07722ebcc6d4a6d06b70b1651047179a5ef43a501acf558;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4f968f129416b88299bdcacbe1b3bed6ee7be8d337f50cb2ea4b8f9f366b03808340c7c4485bfb2a020bbfb2badf85875df7e3e687bc9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fa09e99fa1dd723c38319819deb36a2be0baee13613df1b2c78ec0f3b52361300b46409b16adb8e0ff0edc6f15e0a932d1f4cf021eda17;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1242e162ae97857ce36e9012815f989a1d9370644e7434e9dd1b8c28435b652abdee60699691dc5dc8056c8272b6a78972f1d63bb9bac56;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13223d08e5f66493bb84c7d0cb65c57e2e1a1e828bfe01fa8e98e0d41c1228a2b0f3d9c0b316aca5f34c22f129a1a643ee178fbaea3c96;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13d907c5173baf14ff35602f42f191d95c18d35d1dfa8e6b9b9047216d4a6e3d478ced242e90e8abb6649f32a95815263dd035ed1d4857b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7a350e491320f87ed7d2236ad27fbed0db0eb651a701a75e07dec41c6e358685cf6ba54b4abcb87e588a138e8932e93e655b5e6926df03;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h953f5a6ef40f61b13e88918dbfbdc7e740ea19a46d378c6a3bfb8597835aa2fe1de580295e2a2cb3414292607a3c4e9cc379de96b590a7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb9339730501f5413c71beed507def6514758afea7f7d5ae4aefcad37950e70feda476f61db8810576c46b6895e309dac6f44fa92a02060;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h122ca36aba42651c74f31a21892ea49b572cbd22bfdc310bb28c5b98e8413f4e1be7c8236ce3f84c948deda96e943ed7eaa0e8d962869c9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a56e30f3f1a6480d37d7a4ef4cc19a515151c336d0de495e2a5b27db72e145d6716927ebfd4ac1a0034a9f44717305303c93aedca016a9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9917a19aad69f1dad57ead6272b1fa11d7787fe41c54c033887b2687b80eafb96dead6f07a4e19b769293551c3760ab6912a016aa6f5d9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12e8dd5559da22af0651e04a3a02367d8693909834c7dca7dab1c8995a213d9172763f1aec06c8e5a5d9f50f82d1589984a2e376bd1c7ce;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfaae4540dc4d986928b47947097761bdde1c693a5da02604bf6c3c151984bd62fbd2fdd2f49bd568d1f58ba18877a337f88103e1c416dc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b308b32a3bfb8fe451a82434aa30ce9c0484581bf1be9f073dbe89cc077a24a2876c655b5588ee97fb07e6b309352449b153fd8a6c5e5b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cccc5e880891f775e4d89c718e467bef2697b4250a3dc1d07dd8de5f408a48d333e022617d4091bed65a9cc3b4b77220d21dfad80e94e5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h179118a1201dedab23e9d0736550a8c20729cc609a4ac5a1022531eb39711e65e4716d223a8447cd635c32fb21feab827fa979f9698eb7b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5fa7648d20b01c44d0430085140155395c0b4cee26fc0b9b922a51469c03503fd4bd17aabde13c7e9e02e3d262e2ebde96c7581cadf38d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3f81933078bd664cb989a6d27b1e2c1560d4af31f5fa72c9c191af9e73a57f7f23a66b879abfb6664f0be93f63d602a2b95e417a5c0af9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h519b9ee6bb1f4aeee6d998eacd5212ad9e0f507c583a095b44594c61fc70d7fcf9340c190235ce59ef9a78893b4a9dda58c0941182cede;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12d081422914ef88da16ef2569f1e554b0f14f3d727246bf4f5eb1a8e71e211e282f23945e7647420609cee267ad1cb2f2c782df184b743;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e141d6474723ca1567cabccf95f8079b419a10f208b9749219ddada53caf45cab6368982963b0fe656d86ea4b44da372e759be3e7dfdc6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11bc8cf2d3a1279ff72619d37b75cac004c87ac0814972b4d1c3a67f74761ae12e4e52266bdbba5a9936b8fe18783387341dc42651a08f6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ac83656878292e5a21aacdc2ee891883aee1eb218878c8d6b246cc6b34569582443727d200c9ea6e897447b2cd1dee21c2753d69ee178b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16e70448edc76cbd9320174de5f18b938b241e7ee258b0cd82af2d6724046f200c473c1055c98a99a51914fb1408f862c6d816ecd7b872a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13755aa2ba03c70e9ef98e9c9ef61968044aaa6c42f0d30bb33cf9e18253f083c0c408ba8c071479109150d7eb8ef15f44b84bc99495c49;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha679348a54ca7028eaa0c2ca251abdd6eddf6366c36eda11142a193eb38a2b8518327c8cff1ea55da4c6d7e339d3656077b30261c0492;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf385b0dc422b6eafd4db104dde66589c8d714dc8c6fd64c5cdc0d2f8e6e2b844c74d27ec97881afce57580c8aa3c8a3b422133a4580c1d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1101bd008339983baa04088fc5787b58d195c9fee10859cf65080a25e1a4424d587cbbf68e6c6e86a0cc3ea55c748d27de99729ae94bfd8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16e0ec384f6a643a77d1554112d18e4761db64dd57cf89c418e2dea994a1725dc92fd07e2fb046cf992c1c365077fbdefe0de77e2319c09;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7d969c5038d2f654d348cd61ee7ced26d287aeda9386d433502f6f022d7bc7632aa589338c732f8c27ee9eb848b13429ac6daa857681bf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h101d9e3e306206e55fae6ccdf46eaedbcae2e011488d700ba1c1fa38c0de350f692c3979b30769cc3e91d78484077d551323fa3ff5ad73f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c967e0ba302a066c0a6c098837a931f1fc0d24948fbe38ddbed04f88dd3eb74e3dff9df56eba2ab5539ed9638da7e1306bbe2f92c9c1b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb899adb2030aeeb41f3a8cbde3e23c0dcdcc4a904cca9eedf562a169aff256d646c499873f3e3d8d76600dad8b3fb0f99a77de1b648ad0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h94c6e3b15e52151c55ccbac472904b74b9f84a6242ab3606685588d09cc5b773ed2d35099f9f22b515ef1a70b614b418f4d238f6e4d21a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d3737976ba5c21df43f9d161b53afd03b6055bc457c550c48ccdb5aa6d9a7dac1baa9d393699048342a07733a31452c5b3083c4dd17d8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h127ca0914a383af276bed7dd041d2866a76baf6684831b845bb2629c1501bca95bf4ddf77e2679fa68f25f35f59e7b4b27de59ea18a5bd9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd78dd8c62dac0ee588ec6269cc69048ae06b3b31fb0ccfd989f441f757a38dd4acfe80bcecd03c105c2800ace753ec14e0e42c09bdd8fd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a62236e55836388fb14797450bb8247c186ac342cde62d8ff15b6c4f700908f1caa2773e3f1b85f6474e9d1cba1fb62e1c3e93a0078b21;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h140bbb2a6d2a70680cb9ff63b67977d4144c1f4f6d1dbc9484d73c9c5070ed50c28e383cb83e16f1e5a363afb8bedd6ea78c3c3b126dc24;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heeb5930e38c69e928612676f355b0f37ed7f2bca4f5059e7a8ced41a82547b86affe98911bf97fa9bb2908c1d819f403181d262e428420;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb0b7b71caeffda696749279bf7f7589074d425f714669aa158957704f0b15ab0b4d9f713266013b5cb64267f684148e3ec221f3551f268;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h27b35e23a985a986476920d271f2b761a3599f30ac5adc0c9d0efdab3dbd4e7473017867ad1ba8974d77becd11b2826305e89321df8e6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfc5289cc7d972350b629ead71c21214d74afe9e1c0ab09506f4fa0e7b30512de0323b3421e35d1bb6ad571c2dc3611de4fc7f552e6dd61;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8f09d77876e9640ee7755b2f0e84ea97690888c35a6b4eed894c1faa5cdfd3baaec42da70043708cb63d1b24c02f8cd01ac351c3616ab6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h132c891298c1b53871c0d2253db35fa41f1f6a3e97a03cb61607c8250e57fc39c518f7ab02b9bb6f26f899a2757eeb37e132e4ece74b80a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2fe9408aca95258f958c1bcdbe10561fcf56fc90599b2aaf09db7eb974447d504730d16cb0efef03bb6cc5469df231511282b8c6ba5b8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1929d2814e205f5bc4e0bc3e76e2f67802ab56b53e278c8f431db6475e05396824f0822159f624829c36497fdd794446d6577ec940555f3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h172fe6cb7e57f389845ad2bde332ddda5849da1b9de8c6350d5b873da4c951aee15a3ccc037ea7bebb28ddd47844a2e671641dcba499a22;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h124f6b9cac907a68bf7c505f0e2f728a8820c662cc6b41c29669be4bb11729b9434ae7844055b7d78ae4f8cde1a6d418ac975029bcc1b10;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13f73cf3ccebc03902663565f99b9a4a28b9a9e7f7b7c032dc4b44d0666a679b6648f07bee780c50e3beee537babcab894bc2bdb54804a2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15204d2e6fb6de5af7b3b9314e4fba54781f64f3fd588bf9bd4a247bafb8393fe060a60b13a64c49c2ef22205c32dd81494e5a8b7f3a68c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ed1be6e7f468446baab0277d180c4649bd1d9bb9810ba4a315d89e8c4ab5d632b54b94130c5527e6cb7a28cf7a88db63cf0ac6aa37a8be;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h819a23e2704ec7c92ddb1a9e4368dfbdaaf5854716205661fe9f1e905736aee26897c7d9817bf4a70a13a1354f31591ca3673a1a0e868c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14dfbfa6ec27b338f4e07ebc20ca4a4e2e596ca8a902e6c4a19ab34330571c76ef145663d3b130ba64e0a19d3f7789ab78e6fa22ce3fdf4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1afe16a1528e597f6dae825b970dcdb45e24bbbd40693a5b72a08a96e8c8da5235624c564c7b67e6b1ec38eeb96e2b0e89afb7ee91dc768;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd927e9b59bee1775e0f86df4abfc63c4d8498726e22c54d3a85757cd2a535b9bea6baf748824aa824ba6d6dce6118c7ca288ce0e2fd545;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h615664eaf3414e2b8240f3573df0788e01ed35f12bff8b947b838a2768865fa05009107db281653917697cc538d7d06741769156a2d303;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14273b17c833f4f4ddd7e5be82b49b40c7ab9053f488f22357b4a572bbac2738ddbe1a5832921fdd88f5317045d67ab456f69eb92a44e93;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h117cab0238c3775a56562519a3df7a62767f978780186ea676707bcb647489fc6b8b9716f40fe24092dccdc1d56a4ec8c878c58386148d4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d6f23a70983414675c140ea55369a8d187cb9b935ff0c625b9cc3e5ef32d02e54d04bea0c33984d5e9e81739bf1b968576eb3e4162d227;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc4ea911dfbb312299df3259b75317633c7673d0ad576eb71f4ceea62833a35ffa16e21bc372baee294c0b243a5f8e244b9cf69f1b6ea16;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h902518577e43f0021ac744a0f7770d31c1d85c702ba2133ba3db6435111c5994fb89e9d09ec565fdb4a2e6ee0f4d6a2db6879b623534ca;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha5a057162be4424fd13fd5d8073eadb26792d39b5d554ddf640106adb3eb0bc21cb2192e66e04138b6b779a77ca78c4a042b534d752bfd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hba5cc0c9d43ac0e0f2b5d7733c0ea4045ac59d726e8d69c22d9d3c8ac6bed696015d02d4a9f978f3deb24335cd269fae031592969bbd34;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14e233379b053808d00625dec6745be96610b159ae6714d759a7dfe204dcef6ed10634a7c200be25115a2755d6d145c0fd60efa25a22810;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eff6ad9b76452ebca376ef452f916648c1c16642fd042541964a1cdcdcb634331665b3907a4b21e6ecef3fac05722c7e4e679358d49880;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h132a35673c4c326c273b28ae006b689976c37f021b2bb624a23356d7184c09f0241130a2c5259a188af271f717a8350586bb67b2e4db78e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17dcf0e84bed0af414a5af473f5d1c18913b8dd775ba2acae0b23a38f0b7713e7077a1cf274da5c36dc9fddef07e4a718646fefb92e84e0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1da680300460124bdf5818a98a08350ffc7d0fc3f3b00c60bceecbc7fb9b08393bdce19fd88d24d0d0d477c41344f610c447cab2e4e9e80;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha8ed9df8a32ab378fe44f6b9416cda2cd60588e0153239ab711d7224f05cf5c73d701d8511384d65b9434b7076ddcdb0d842914ace2f91;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dec24fb8d8d0a6ebdfcbcddf989f8e6a865dde31d1961414c3c278ca682c749e81315e91d4f35b2866e59a0b4e532fd90c82f4de0a29ec;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5c7713c4efcc742446bd1f2ee409f1e4149949124ce9a0fce56e031a8977d20cdc9c432ba685612a2cc4376cbc573d7802b2729bbd102;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19482a54f602ab3be813c2e577b470f064f1a32d71f9debe9963dc13d7b77491348b6547625b717513f1e56e10877f9fd9cb11384bd3359;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1deba09e4a8e6bcec9ca37a63a89766a1ad2f7fc4c6c765a84f1e239e734fed4f905461d34f83dcf0141dff122da406e9f65af637d0e676;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b683f8704c0a649f6c1d586e3c1a043c2c20049858b9c057ac4730bca06a52d7469cf18c424ab3b5067c66d9815ddc134d063b71e25924;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5262303bc7649a9a2b3b992610446aece1fe34694aca7b293f31a13a9105ff3fd4b42a9cc20c23a7d69a3b0158108e732e5cd1ba4a1c4c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h29695c60357644f662a69fddc96e774773d48a9a2050cab57c5d18173a286e65664dc2b915389644d4fa2838806a7c7a271598bc7cb41;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10bd0a1d0277e4d56344c20b0f7f87b3bcd9bbe9e1ebd3ff43287e5bce5b6fd0346984365dce709522f34801fca4f8f6e78e0b31d31778e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a6ffe2e1a36d1f0cdeea7918eedd9767045e451378268c9e3967f741279e639a4092a4bab8514cc2e2984c34488db55f698a8791ab597a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11945ac0cffc9f0a947afc6915e7bd1a0e630a888f8f160da3339e1ba8b68a7683d8a7f835529d856d98b7786d3467d814f5ec054e443d5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f29be622e933fb4e4983ac7e44e7af2178ee1717cef2641cbe4165ad73aa4c19005dcbbb9ba15b4476bc7079f9fd38ae4b69e6c0e4bd33;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13482fe7c0102885e83be9b6e86517fd77e0dc1825eda4c887c02cd1eb3d7dcdeea851d48298778131e1281437c0c5adad873a583b4f0a7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h115d1510cd3d18a2d8b3eb0580b984914335a3d6a0e21c83956678fe31963cc76300c7b60edff5730431cd187129b1ac4fa1a5d7923e52e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h141d8cf9b2193701b9ac4da4c9cbd2cd6df06883da0a401990af8731584e8bc20e5407628194c5113857fb1a9afe87bf9f53102fa9cf414;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h180b465703a97de0f34eb72114ac79b04a0a2f16b7ded963f24693d62ae04b777c8b52ecf488bd7d10b7c53c3f7c29e0284d516aef40e6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb5e6d659a3820d0b0640d0df23562cf3bb93d0e5b11ce1c1259fbb758e98513dfb482205e2e777417701aa56dac84b07cc968227dc70e2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h54b57b9ed6d7af413f110d64a4594bedb64454528d858db5623c4a3329e02414804ecc793b33a1993ecd0a461a84ecfb17d9cfa83ce2c9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf6aea8aae415458ad1031b0c4fa3b0a27b2a61f27b17f37184191ad1170d43be7d45fba8ee198e86490d1f9c48bbf601feeb324e430e5f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h137888c2783f5da7a71524f503f3c21690f5fab85b1f753aacfe59a1bd910065cb1f12231b836fcd5bdd63ba366059716618da2199e34cf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18bf9a1fea2dff7910710a3399dd6122364ae9fa49a0b58700059b185efb7f2221666569ff4475b59b5a43d6c9ba0834034ce71401e955e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hce619980b5a4419e3352416a0b7012bdb23acaed5fb5f06044c7790479b5fa8dc0e2aae799005ffefc3c6492cc6c6b8f02243c6b1a9b6c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18651216297554c926639b37184f692b48390b44e43cc6619d8470ef357b5edf302bd7d6eb56a27a86fce973fa2ca455f0ba487a1ce9034;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7950703d2da05a4768acf6d1bd33170379c385a27929c2b666ab92a2928c9115b3543584bd15b7b119507e1c974a524747ff0f277b2c0e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h103337cfc2a58cfa71e131d2f71feb8de9001493a20cfc0e131f00aa126e35b039a109288156ceebb11fc4f2892c674dc480892b66cf740;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ddcfc999db586f361f706d14b5906df096c4235197611ae69e42598de0bfcf37a4f559e1a215d90548c72885a6dc195a2b9022f39ded58;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h77a40fa0ede13a32c7c79d21636194e4f4422d8e8e9265ffcbe2ddbf89d26c35e5431e0225d1dd8250887c82e97121d144991cbdf6dc68;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1765d518cd9427f2077d42e19653423281566fd8bbe1f1077bfeda452c017bff5f7184555bfbd8f8bf5c3ba391e5fa874fe2a17a653489d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf02306fd037646d0168b013482a51bf83d57a608f560c9758c1537f4ea386b40bf0c6adaa042af3bbed84e8aba0cffaf2ec107579752a7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a340dc48af5018e90729e7399cf6b653a20b7ff677ecec7f48092c317c74c2a2dd55c10cf0cf82016696db438b69e53db38fc4858a585d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2b2cfc95d823aa747e94f849085f7b53e76d4d92647fd2569c443325713addc8c78d9a3422810e596d791894700c4da8cc748a7e4c1291;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c6916535cb184de9e6d68440f19599ca9f2af2942d8e0d0464a650f0ba4bbccbb6a61e5fb9fff64160139d9e0c6c9009868fd7ca746bc4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h135b0d6ae2cc06cc9a75d1936d6451f42f6d4168acd33b5f5694eb3b30e41ecd144cb96724ea1af99bd2d4a66a0216e3b8279bd182ea9c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h33b9c42434bb55b953c8851d5737e421b09b1f5638dbe9a395fb5e4a31c720b9e2a294069004a4b81677e53e92a04245fd6445b254f2df;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbe742a5f1ed157bd17fc3c269bb105c47400a4d265bb61b042a0ec4e5b72ee5a4883bcb6c84d1f510c765855f0a58528397324f1a4ff14;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c21e38adddf807cc9e0d0b2858e4e8386c32596721c77e5b3a5fc18949f2540a97635a9fdc99216c3219b3221fbfc7b43ce819efcfa229;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8c5a8783c7872a63aa964c145fe956556618aec5fa257bdde0fdc385baf6765a2f9b2b7442cffac759d3e3519203c281dd527c58d12329;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6396fc48c4ee5f5e1cdaf556d25e83c0e40cbac1e7c99beb80ce43166ce95a8a89335a6012566b4a196e1bfb445092860288f1fd881f61;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h263a2f5df0f32e47cad050030983fc28a7f61c5f03e2adf8720378defb8df2061fc3e2f9e80a27525aea3ca30e4d5326b8de1d4c93d86f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15bef604ac90575fde9e3ede054ac0adb2e9b6e4c1f41b0f958a83f22deeb02e72c3f81054acd32af4981b630149ebd2b8cb3a60b987582;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h165d8adc7e26c0c5b77e9bf58862a486c6811f9e1c6929836bed8203196735615df1f70e2ae925fe5f8f7da5ea5b20ac86c4a6125dae06f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haec908af0ad7baebe97239925130acc49079cd54dfbb642eee274f18a05538ad406bdb7003b57c95a661937009dd24c7174f8b8ba0100b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he27ae1cffa4242196054bf05a4fc46b0d828b06198eb597a04eb06e2ba76b0af435917bb9a9761215e33fa649992bc19d3e975e69bd465;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h133db4d0549558c7edb51816b11d23c49d1d253c217ffed62e7debecec83c011bd9d367596b75e156dc3f0461bed2a2ef73d326813c4bb7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha9307f985e40d0521c0c47ba808cc5ebc142c32167eca7a65a0260fb36d352132c7e95e75d3b8cbc9005a66a5ed3bd9d3e928a81a61c13;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haf36cfdf7d4870319d3892cd4b752c600a4403800c4ef95aed97d1d804244307b186ec66391c3dd838d2690ac30756b85df1d814a2559c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4bdeb3b94806bcf49ac111c605454638bb27ca4a22a8c7dad085c76337ebd5aa860f6ff264d3c1b847aeb7fd5a401967a4badb5e70420a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h33c9cfc1b6eca2b3dd6578f9947bd55014277926f2d29f90582a96f8fac5832f85ac515d8c6929ed5f812b344d8884dc29cd8d59b1236d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h860169fa3c28c4b1f5866de3cdebb5dfc61fdbe8cb7ba89eec529b4145f3b9c2b411ddb6138357894a8a8aa15634a68b5ec6628c098165;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h101f360a1203791d021f41dac6e1711c4f6e96f6c56ab9b62cecbeaed7aa8b9c3d02d9732e6270dba3d2e1ff1caf309fd6ef54ac96a732a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb7bb2ea5fd798cde87dc590199c11560b5fbfe10d7e9749a5185981cc1932a8be81010993dea1dba5af914e71f06c163c275a04c0bcc8a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10d366c5c1cace36c1e26b2a04bbe85267964e83f5739742d8941c4878f0bc901fd4b01f591c5f502f2bd8bfe9efd1b25a563677a414bff;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c318b7e72a61776b06a00bb701a647841f3d659eb029136fc828a2bdc827ab5f19ba0041f2ea020eb6517202827229a722f6414420586d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10648c4491677a6d274b055ffc623c44117d13fe552fe2c883167bb66d1c2b667e87ea2a44528ad74b485b397e62edbdca775c64f90d2e9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e8edde8598fbd91febfac1adcc93f728f5a8429c20b63473f23c762681701124ec1ded4370beb2615ef8d62b8693a9e37b42126ae4ecec;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h961d80122b15604bab9ab28a1b4208d295192240470d619b3eb018466061eb8b94c567b27c0651638fdc36fccfabc8ed3259c273a27a00;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb9476ed26003168599d1e07cef48653dc217701ed4d61fa16b178cc817b2160a91a34f00a63f8bde129399ebf06bb07e4672a11efae4e7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f46e37de635d4c7a057232edef9482065c43f01a7755175055e8b8fd4708954e66e8352a32850734e7f1854fb283ab7b87aa3bcff48e71;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10712c7fc46bbc5ae5abf417dc35d3bc2821dffa65e3a5821fbd0f90870aff3d776bc7911def0dd52bcd51ac74fdb6800cbe3b8d42c464d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfc5e600c404afc339fa3266ef0ec40305bb67fbbdd3f49cf6d802c0b3b7165f8c2eed7de1109010c899c0db9c59439e2794297b797c685;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcf171d6033f7fa48ea2ead37e848f5ff78d497ff18e24a75ea536fe93c832fe1102b1df55d0513315336c953c1905e44c00f592bdd70ac;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e6336c03701f96cea030d42b2738dd8a0cf201c657278df942a6554e2814a321d3ae249ebf6af6ad5642f2330013478cf37e9f9d60a9c2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha085445ca0bcd5d148a762656a0ab626cf6e363d1d3bfb66a47311dff328d3e2e7b934440db4b2a6b0b758ded618d1cd843ae4529edcfc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc0bd3098b05f00fe115b9e7c7bc0b7ce00538b807effdd4a963b4dd9bd50a206c6d9993f21202d19a86a31cdd2684eecbe8e1b055a887;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2215276f1d676c8ccb1993e4784e3c5dc24552f014a8193fbf03fb45bf3aa17bbb289aa08d64536d20bd7f0af7e357081089baa83bd655;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bbca9db134ede5d20b0d686e65b1f7cee0e17c212ac519b9a159119527f0c5679df6718827bdfa882ede3c1fd1858bcf70761e3c09a0d6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf9f761399365b5f091830d02564a044f5ab28b6ac277a17f3633dc4e0b9a1fc06f17016ec61fddad8627ee6f8b287656336765fbaecb5a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h103566c78a1cd627343620a9e9d40302a63866acad6142ca937ff851e6143e932807fe4b1f40e748e33e4ecb432f1c8fe4d33eb420e716c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h121b4e6a9f4797f8727f9c87ba8185521b0f43644ae095c28d4977feb5227eab9497c04131496dd5373f19513c4d2cf9d3edeb429cfb1d4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdd2fb5a59a453963aabe789403d325ebf536cdc1840d955c79e90f98f3e5fe98052810dbf3c5093bbfc77a5c03dc21c01024b3e529774a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h67af65554186ec7f9dfef554d6f6f1de1e57357e192ef49093ef71b8810e63ba36f83532b93f534795d13fa0c5e3820b2fec288d9cf6d9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h31c5f790be64b74edf8a4f711106ae9664a43b18920407ba6e162dcf2686dcd0dff295362771f7d441f82f732bf45a8c0ae0dd911895de;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h132f485bbc99219098b2856960328f3d469a81dc87942fe22f442c685f8f8ff5344eeaa325b8b1e6f90d35d61448b25b4a48f1b6423fda2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf30297f209368b40ce4d1d771d13db186473282b5bb94d3d161710d8c835dd1aac9fc7f7a5bc32167044c486bc6e1aa49441b2501a2e00;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h142713a978523df08cc0f9df4902d9a44f2a1a5cbf3ef2bb3d5756b7c6afa02288e57317c1ca0d80ccf1ab44b3b8d76ad9cc37ac451c309;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13a1f6482141e927cc1d4770632bd8b675810b6562ade791d82f1e624c69c23aa10ff10f9db077b322d0335213b519f1f12f7b6ba7aa52b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cf79e44cbcb71eeb88d0ed54beb7d893c609aa580b69053a6cac252bf5528c54bfa920b81ca598ba24633d98a21132dd230ef717269408;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7b68482a949c657d49d456746c510001116776e71fb7329e7933aa4db694bf0af30a162adcda5730b5173e3e3c48cffbf48f9395bb0251;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9b2048ad9f5c062cec6fde1a7e99bf8ed91f2b0ab67b4bde75c3fece61968a85caed17af8391c6be7379493255d1e64fec52ff6dcfa4ca;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dc5c52a7f918b4db8d2b7e907b294d1414b3f5e2e3bc67d9e85892dc7b23c51315bc57892ca4447f3c022368e83896afbcee404870579a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15da800e5db404f4abd4259f4252825f35f705f6b724d3bed682f07fd0d32eb3122b1fb43e1bcf7c4690b3ebb0a3a3f876dbe26bf6e0fd1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h75697f16bdf014c5c22654ccfcf40ab856647e264df6cfe43fc49310b38b52a1f8fcca3b928076817329b03eef9adb0b113a89e0b3b67e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h110648d06717742629e45ddfbc8f196d7a989d87216578d370ab699947dea4ef7dc56a4b6bff1850db26897b423f00ea7c9b77ce065240;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12e617b2a39b72d30502771770dbb4316839c29e7ba47354c0c6371064d973da7ca8e481071f2e5629222c1a0a02f96648538a0b0754b95;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h55ec6fdaca8f1d6a0dcb798ac49240f779a545e4f34f891e4cd1bd77b6cbd334c9cdafe7c98d51584f7804f3f8dc8ea5cfd132a28a5f7a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hadce4e6c1967733449818fe05c7558ffeede5fd712e7b5695b2d42553fd73101fb8458f90d1ee0a77ed29c73a304f7895e175a34db4b1a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h139c0ecdf1e386b40936b64ed6ec42433ad6452b20cef81878c79cb15ab12a478c23f0e1497d833ec62c183902cfb4b62a856c203d6a6cf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f4dd553ff9b8855981a819e467fc6a0e2e227aaea546173eba8109983d079c9a2be7620e479ea4408eac6ccffe34c0cdbf6db0bfd15138;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10bb32e8c7707bed80281968dfa9f0777695ac6e169bbcb25c93cf8d102a158f0924964a21c22890e849ae39ce1f91ecbe205f02502a96d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2d69e6f38186477e7909091e075870bdd20213719df85da9705a971d144af2a57e9b550cf7532502a7ce5ffc6f53296d591b4fee6b2196;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7102898d7f8de395ccbdc8a11ad63d4cd587e2251bb501ff83045feedf02beee8b7ad2667349236e8bf87c7666f2fa95b01d03c92b00ec;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c1218f0e5245323e189b34c26c4546048f90abd2033a09add0ee3b8c8b11375f439038be421fda5704ca0708de848cefcdda18da31b5c5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1511a9e55b99380d4afc12d3945a2fbf5fa34e6cf2285b77cc895081473be9c58eb7bed9f1b46b22eaf48d1493afc0b952d50a4be864c36;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19ae2d0cdb9f5349ef2ed9b4d5c6369d2bb423f232b49c1f943e2c5c8c70568769f01575a6efd2e944a8fa239b12f065fbe784c5fdaa573;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1863dc34d4b106cedfb8566f50d33e455ce735be3ee08599f9481ae1fca68e77b07bf40db6bb943b72682933f476bd1cf9c7aa29d4d238a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc1afa63aedfed02a1c3950c41dc391374d28abb21c7e492a5d687d4e1450fae780877b735d63f2564684126639a525853fc067e2ad9ad1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he9d4bc3d65348ac1003706599bb48baa1d716902a4c7afbcd0e9ded25682183ecd538bb0f6183c483b6b4931a1ff9f04b98d769f581296;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h56f56865d5377d15e66fbc12e52e61485e945eca2d89218f322c7e30ea9434b76fa5f1582dbdaa72e7313e34879988c83fe85a7188c399;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b6ce5dae64508bf6b39153a4a3822350366277a29a0546511ebf1e499110b10f34420e3e0ccf79e06ed04a560c0b4534272958427e932;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5fae3198fa71fb2c04c805314ebf3cb31dac3728a05a8b0724f270eaf838a713eec8f00146cadc48575504ad937c39500dff75c4796844;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f50d264ece9f7e1332f1abd5195edaa5116c14df4276bf6f1bf84d2179169b188d0a1032ef4074fa5423a577daefaae0833cf3bb9d1175;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3ceb847ecf335d8c2992f90e7bf8685ad8bbe540b365ef12f798245a9dfb56bb45ac3642bd63be595b26b91a71549290ce8fe75a591ba5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9d0bdebf9fba3b23e733ff857f02a1c7fa65ee677896d57c24f374a0c0723db0c0c6af1416f65e8aefd6f473da3819959f58164ce0c519;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd9df98d2d202f1b315c67406b015acbd7a197c92d5c36507b19d7c45312f64665441736f1ec358e2ca414970c94e89ef2315e039774155;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16f33bfc4f709615e28f526895da378bc31eab9ebdb10ef277bb5f18f1c760a51a553ac8ed5e17285c83ecded619b26b2420deb70482484;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6a960f38d18c34dc5654f492245310655110afb63cb3028907ab42ea49d74e6ff1f4cc84fd3b2b74e1058a706227be58d143172a4d13aa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5733d016960be96682e85484009d446e36bfbc3fbce86bacb402c09de2413849660ce3dc6a37b92b3f1db38878ba5b4c9c6724b4438057;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e43951cbb092727e0a0e6aeca211045326c9d2b45ba38fa959aa4a906d29628a145203491a3effd32910edd7807423fe70fd985c68d208;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13ef7c810ebcf7b51d698fc277e821f040a00ffcdf3df8aaa4900a2d31942213c69d02919514929ec7cf65995d2f2e3879f5a8350b7781c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h66ae060d0fa1031933b83b4d70d3443479c3b1f4833b6fefd22da881fc5728b0741de5f24a00d770195b565db84c1818eeacb9e335117e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h425a586e544812a881c0ff3e58fd46e60983220ae5c4e860d260093db12cd076d71bc451587c24d193fa88f600edb731aae7ae508395b4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdf2b376378634119de9734e205cbf65013447331e33b781c4a84a2771a88ab2af536d08267365850b08c128d01f9b23e9ff419cb814435;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8c42f9b2cef720662bfd522da8a99e819d28f4afab8c51467772bb90fed795e2df82d9c01ed799894a986d143cf6f5b65b9cdffd72e6a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a487eb83b5471f9f9191f4f6ef8ebd7136cb9b11f9da49840bc026e2364fe47b0036fca08ef3399a4623792aeaa22d70541c1d84a126d4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dfaec01e6cc16cfe32a8467d00c7a89813fa30f8c85a212d267bde2515cea5a68e98b1b2978692517f0a5a98c0dd5dd43e568b7772bafc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h918c5ea5609b57004a43730cce9453527d639712d896fafe4241294af425f547d50544577100622e2e514f3fb0fd85b1bfbbb5ab61c8a3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e21a7e86d640b3345f2680efc044f96e311184a69d3c4dda6bda18a519d7f37c19102208d69a12130f742d16e5fd7c7bedceb6a3df5871;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h158224bb371351af934e19dfff912e1b525210cfcb6bdcd1b5dfdd16a7dbb3c10e58e13ce1f3bf2f40205983f831fd28f507a5a0613a36;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c15ec6572d58507d60124dabbb7c96f8c15400d7d910927507729ddc2f2d792828bc64887d7981080c27c7b22562d2ca5429d58fbc3911;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e98820b0e63b7fcf2fd68c9926be5606e7a0772961d42bca899b8f2fdba2767a25d048abcc8a9b80c517dae1e69c18b5bfbd208b27858d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11fd480103edc2cdd1566b910d379a9f9cea00dfafc3cd36f200bc38a76a9dbc36264e008e51005f4e7bf569c0d8583f3ea90f6af917857;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d8878a2bdb79d7a1c52f390ddc5d72bd0a36bb788b66463928d1b6a2108e9157786e3b17189be7ecafa7e3183104d80d115ce4e44ef750;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1179a737a2c1cb11e004916ba42efcf8b37978ecac4db23dc47ed20c61f821f276c9b845427eda89e79c61bcc8c905d9c09a1c3fb6d2f48;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8e1a507dda7c98d91e1f2aefaea318e9e032401aa232ca8b545531dc20caebdde7713f2436bbc6d09a44bb3ddc51118517982d101c1ac2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h119b71e2491cadf64db4a305fed538322c996780e13429b8e05cd6d53b8bdfaed2c1a7a303f2bf3429497f236a21dee6c3a3268851e9391;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h366b529bc0e72ecaeb6d666a23ce0642820fa768f3b465e9baf44b554abf8e0c970bc2cfdcfe6f29425b4c0bcfebcb735847d8b45089cb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f0d0a3f66fd3e56df9774cc5aca4555545c7c65c8619a56e0adfdda7f4feb2473341b17c28d12c6b00745f48bc9d493ab7a34a89188476;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd75f53fb8322ed9ddf79c957267a1007f03bd640153f78257e935a80b3db9f9750bb4ddab41181a88a40191ceb80b5ef5e1abafb5ed05;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha8e34eb32e75f5eb0e6a6c006ebf55a2518b40536989db9c04e4967169d10383e7b618da04ef026d0a6059e96a06ed66408a4feb1cf1db;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h23c68bbc14bb207688fd6197611775ee391de645a96c89d3c7a17f59fe74052671e07abd6d0d87a48e0152e7e546aaf996e9d82366a728;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h177642c2cd4d276364cc9313cb3b0ed759fcba654fc24872e39722bab467143c612d3cf1c647b7d72f08a67e1e04e55f48529247d94e952;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h388ed10d89fdb3618accb48f3fb62831f3b1624ebd3bb1443e8fb0875a8dc0f77cb4c3b70a8752fa35251ecccb0adc55b5e1a4b703c0c0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbb4462e1417f686aecb062300e284304f61504df0a6600adbd78a00e6351a40cd239be6403ac00800d29fd35432989399e2a2a1610c557;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h467e191c4ca38cfc8219732a2bb13ffe17344384bfeb99917bdc53088bfaf24832be2170115ddc8272a2ed0ce879e6810b807e718ffa02;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12dd1a434c75cc808843417eb56a1ae1dcf155fc6db90fdf76981b01c0e54f6a4582380f9515ad4d1ca7761175c0a17eb4260416a92e139;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12209658a86cdde20b6fa92bd9ace779790e5057dc116d74e3e2e7be57003d973f622357d408439a2ec506185df3edd5305829803abf4af;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fa3fff05ba54dcfa397bceda12c807e8a8d6d3f2b638bfa97ec6758b077d3511dc3889a4df7a9c69f815c9e4410485acc4064356e769cc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h181d2131c13abe5f7b2100ce09c7b40e36f432901abd54087a74c59271e45663d6b6dc737e841553ba9b0e781564bc60e671f1d2bd09f71;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4cabba64b2b95cc040beadee3dd4e9426a505899c4ad4354e1201755de3906b9d1543f8b7d163352cb08edbb12de899c1638ed3468fdea;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3955307f1181fe2733fbfe62b1e19005aabcf83b974247deaa6cddfef94cd6053fc4c93584163cb2f60bd61117329350c7f75496e43fe4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h53d25065c767bb8cc065ca0445e7544db9036398952420d86f29dbb40692ebaa1d374e2b831f2dc339e7117eeb8c27ab6a9fcfc0237121;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdc6d9c785516254abebbb6eb0612055cb794aeb7fb92ff1b8d7d3afcc5c64eaf6215313a72f5d92e11861d9dd0668b7911555ad709936a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h294afabc5f26e028d41be4c690d970016fbe8c918ff7937157e116799223f39e9550a247e71298adc21614ae2e876fb69e04571d1d1208;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eb050b912434bd1d7eaf1efec35cdd6c12cdd9a1014bec114bb3248dafb2e01b6b144fb004dae0c165a2de1f8a57f46fb85106206a637d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a45bd17331f915cf63cbe8c15fbb9a44d6e02e2fc31a594b455f7aa87bd791e63f29b5a92c99a82a7d31be646c3f6636821431b05b070a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h173ea20633fd65fc9e7ab16f3e3c6aeec4c0e97b96d3e0b84edf032ba10be2450361edc1bfc9d0edeaefce2b96d2dc8c0cb30d44516127a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h166144b15a072c90603881c854fa4b8bc82251ad37c1fc7be951f671062016263d8b7a8dcf842661a9b379add25766060fb4b3cf346c447;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h34c6124fa12fc5c5d29b1f9f53763095f505332dd5a21eeb3817626c3b6003c0771180ce6b2a9f8c1208ff7cc00609c95aeecc87211ed6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ea43442e9c84b391d825688a63fd8663bfb366b5be546b6a52b1a64c72e73d367a61e3fb9e413df5961e2d4fd6868d01016530d652af38;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfbb3599e0e21b8c0e21c4fd58645662c38faa615576ceda8e1c1f3ba30bfadc4ad2d71b8d87d6125ff4d4cf0fbf6156d19f4e538fabe1c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'had581b103bac73ed6eb10117b65330c4a102cd2ea42effedd506d97cdb56f76b947ab96977ce6707a6ab43bc3b449c9720e329d058bf39;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1adb23f414c4d5cbed51fe392035fb1bef3b94b534a750747399c186951c59881c0b016cb964bd548557c560cddd462ee151809164c0695;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdee008c3d289dad4e8b7457b195a25bf189b7adc676650af6fb47adb2aacf95589f701b47d52feea7b85c360b98fffb6d8ffefa0ed9826;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c71b2ddd9b2eb240307199d00e93f1d3fd37974f8eb25f9294eef03985568e349ba63f0596eeb7aa04231eed2727a59b2f5e2088951f98;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1732e4907e62cc21b6788e5d0981f4a49242057aa0671b208865b43bcb83a281d1eb3117766c73bd4041def5caee0ca4fc68d8b6746507d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha075986ce610bcad5aa253946e137461babb535f84219e173348b04df8cfe0eabbd1706616e0bd8838761860ef2df7045eeeacb8440458;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h548e17f2bf3e051572e3a558e3cc00f80d22e6ac6ce7610579f9dee4ef3e62c89f53cac9a680178ca66987ff3c9e044385dbc9d3427b5d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2ae8ba8e60a21619cccad84f842da7b865138eb757a5893a42a59000c13d5e7733dba5febba90bbda6cde9abacba5799fd89dcb6cb276e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14396401ec6c9ead4c5f792ce14d0f55dee5498b671ca0e81a61d2189e3e614efc1f7dc227645e125d4874955b19ac5c1d31c8694ff3825;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb6f0efa5c283dac8fee86c1eb6566fcdcaabdc0e936f4e3bfff8dbfd56ccd3efbfadb7c6f4fd45a1b4ca3c31ccea9fe8ac55c70b1b3ac;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8b3af6266bee6f51b1538ce58d311bcdd16c4b1cbbdd949766a4ca6224bd15ff7a0d7c734cf0791efc154c74c1cddec5c98615596aab2f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c438c6c2efb3731160ad4059b1823cc9838c333255165cf8e6a4d040acd0c381b226591d01d9a4cfc78c44915ba65a3a0f0f5255cc3a0c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h91b240ae41a9997617d6f856169e7d3d82d6c1991661cb384e4a7d5758209f42af5abe8b309eb0d6cc8eddfc2ceab0b7da49f7dd400701;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha907d854196bd7225a6d9c18d9926a5e8f19ddd91e18f9c74a7a9053294f6ddde4adebc0596e1d4743d1197d7f02b4ae9d221e93959faf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb093aedcc83d0033018c595b6ab8e72c2e965ccac8ed529cb2634dc1d7561d263321c8a2da27a0c9f507733839789cf853fef7250d09cf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h20e55866f60406a45ac8b93b88470659fb636cdc95be2349fa6b934375b5c24d7b402793b783cc3d6f8ef191b88a453c309102034a1d8e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5369b9296474fbb4c12193ce34763eeedbdceaca2ca3263c172f21a1c3b2d7bb0b8ed79817ef180d186d83d36fbcbadddf1d5d85c804d4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15598acb3dd33e4456f423b6755a362ca35b327cc608d4bd43921fc5849179ee9670e4b8e6e078a99adf9582c388c1e3e77b83e1c066673;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1673076f23b1a389daa3ab7ca8df5027ca29e48ea266685ad783794d14af37de75fe907dc3926e44ab9f13d1a54dac424852de6fffa2326;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha66b27a67874f9199d54dec4caa3a3b75d4281cd9a987c364ef90b29bee2dc009fe1a225ae85b0f0e197f8e9970ca0e68e4ad7febac871;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dbfecaecfa10eb18549e506dd6adb19e32182b2b35182c61be1fc353a3cdb524594f6c5bc5f380524d459f4dafaa9c01a60f0b02dc173d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4564a6a308b4207532552876a3948cc1e27bc7e2d1440104b251db441e73fd36da9bdda71ed22d6fc78a62f230ec2b85d9662be4e0d8ab;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h140b233bee8f13d5c7ebb3c716fc4bd6014a56c57548e72161be777e86b3a19ef0931cc59e16cee8fcac262042a7a022da80e1e0c64f101;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h71bd160c323467ba81ffe6abb325314e9e0ef4aa9ff1dfe24ce89315db93775e257095269f86647db659d384b855031ff9ac586971de2b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d45ea89e482818263261627428cb7d74c101a0c11d42cd504f27a43eb786c27bd856bd223cbbd722c57a3d5decdc89cddf6d97de4cbfa9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h92a89cdbf16320645364b59aefd8aff8a6750c3f8b59dec5cf861eb1e09303f3d1b398e584c9fa1854c0a3f4c86fc392baf327b1acecc2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b82d7fb1e63752ac57d90972641e7dd0975f1a6d4dd583d9b013bd9a60eee21222053cb9daa50dca387e44394ac9520810ebef290f9d0d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd06c3934402fab821936ccd0e1a818007b5cf705c72b5b470edae596f199884dd48a75c4df65a225ba67d269ac9d00baa1e3f439b0d9ab;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h90b21e5a2d1929a90a3a8a90dc974ed9a02cbaac7c5cb240bbf51318d3d741cf085fa26fbf88621759baeaae63f3dde8292f13a11a881c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7f323957b0fa14e059f5cfcf7eb07bd3ffe22f17d6e5216e73fb0fbab9cb603e95eab764fd1b6ed61a65bbeafee8a5b20d5ea3ae0affde;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd0c2e6a82d3728aebb7baa7240e3dc24662b4abd0ec77fdcb84118326712ba292d852c9db003e1634b007e6c8de9e6dc803b511b18d6f5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfd382a5da7398f7367881a135cd6c394917df06bfa268da4f4b5b758623f096bbdf75f985090fcdda6cef83da2f86742101dfffc7f87f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16827ad1f0fa79df896492de98893e372eb2b1924434e5bb294b555ba768a86bd71734d08be7bb6aae93298338a203bf4addbe74eb8a4bd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8e09bc206530119b693ab8c0097607284320cc168b37990d20aa2a180cc50a2378de9cdabcb1ae9c95342fcae81babe724e3f6c9b48407;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h57c13636e01ef64aa72cec6884203a9b8fa32850cc4a8124c60bca62129c12a2215e893f135a07d66c2f5c5e7b2dd5cc60a594171d59ae;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hed18365118411c3330b27444f4be59b45f4b439b62a6a657b8932c0813cdb99741f40c22add9be6c87146c277f75a0580e74b62da42723;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h157fc88d885eca74f136029edc7fd178a404c1ec4bf85b301680a894a8f6f8a63642b8a1016096321a9251db383d6ba00afee45b5d379bf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5186bbb21239c7ffe2c7c90879841e974a6cbd0d1c6f6df36bc52f5f31217a11834cc1d63e16daa220c3222e05a76a955cfcca21cf2617;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ccb6b60a6b384a54826b3dd0643278661dbb7d97aaab0d4d500d18b6922fe142c5c5b580a34086572955d3b1e69800cbfb90df049c6afb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7e1d293de303fc696499605c698549dd9fac6910db3c8a29f3ce81ee3711fc5fa628f3db26dde808ac450b710a124594b6f9389a063942;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16a854a2150988e8870e00a13115990ebd133564f79ab181a700872644596a6e95828aa9054ed38b54701a1143cabcb66ca832da745665d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h841e1c5b039359951b5d2b47c3a4cc31667f951e3a7bf3116ceaeb936a5ef9bbd59ab019108d10dad4c8cfb2d75591837e117079b91d9f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h140bb555d0a0e85a1ff7cbd30384667f57923ba4bc3b080435376cce7aef2b288354862f5d941500ee417378c43afdccbd2f20167544256;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a22693c973e441dc3b6fa66e1607b38e05a861fba9f4c5e878ad5f56682942ccda0880c48d8e84c6e05ceec56b0ad0d51db04fbd250bdb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdc5ac368cf538546d1b0aca97fe48f954cef751226ca7f5c3f9c8615d84ae6ed09e8996af1b8d50f59f228d038cdeeb058cb69e66f20df;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha153ae7ff6fe233ef17183bd3b46d5a9d50674eda95f0fe9d04c9dd78b3dd97c61899f3674a4b7e4e7dc0045f60bd42f1e99c1f1c55f35;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h51eeb3569ca6c8b6277231949e762018024a2891458726c1701b38d5e7ce07145c0c597be34ea3a0ae64768643e8f1168c7ab2cc2ec7a6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h73af0dbda1026f3fb9823a29ec1e91672b8b7fd9b8b8649796b1eab443e0009446878d0ef07d2b7dfc41ac3cd98a4ccfead2e1130cb79a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c2f76e0d8bcedd0dc36c0b5ce5899624359b0c5883981d3e6f155fac1e2613fc4b1104debf63c75c8ba20bb8e1267629b5f12502020dc9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13be712b370bff7236478a94f28eb93c7af17ed37f2d3ae3ae300f8399589e95b5a2a99b283b05b533ecc428a3a34d3b57cb5867c234884;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1749b21860f23d28f47387f780fd869893c0887f928a900bfd17a642aa6379429e78f2463590e4da117dee37a967021001e623fec4b2e63;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8b1b3f248380fe7ae5b8f429047cbadd603c27c01b914f4e52aba5288c9b432f25071de144ee3aad0c9bec57e41fcc182fc011e3ae8664;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13acd29e6a1ba33a208540dcc5e17b3c3cff73c115e2bc9a4aa9d4102d5d4977e9a0fee83067a01cc36c0b917c578501b859a1acb6ebe1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h124710aaee350ceb1e4f0cc2728e5db2aeadd73d58d03c18078a350c51884e2dd53274e1c79f75613db7882fe90e893e2bbf19fe30ea492;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c567e2af68e4834708a51ea1fbb0d9db355752b3a76cc2dd6ebe310532bf6df13f907ac9ecbd35a23cbf6f9bb43c01003ffad20968b5bc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8866c5a9e104d3f9ab2ce2ff107201d612d77bdb734f50df33d3efc16b41630a11fbab46cbe7ce96a21437146b02e269f81a476bdc8650;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9c8805b0c92c02ca5beba00b6137d9a35247d57ce9b69e4695f4bd2bb9f4119940fa25b72dfee496aa70e6ab1d708e585a4ace6f08b260;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h899c57fb6b661786ddb37b7aec41fe77dafc062617cc9a11e2d86d186da24c0fc05bb3d7f7423f39459e614393195946909317e0e93bb7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h131e07942f45502b3d45772e44e04206c2d9530a4e8c8dafe0bb83a2abc39fcd0656d8a6bf4acb193002c311134ebdd1bf11e2d1bc768a7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h134d8f6b730f2c8eb003728ca8494e5294b1d8230a1da94219a38ba6645875ba8b337913c504e4c521a3b6456b4000c3843ee1833f52961;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7a2760a1e2ad43972a9953fb1ced66d7d28257f5d97ae8e832660f4102d5b0794fa4c4f8973c9dfce5d5953de6b0e3ea405542a8cfd6e0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h191b44c82fd4a4c4e456193fbf93b0924d1173e3256b0f52b7ff70c99205065abf30e9fd18504f2bd2c92cbd775abea9acecb7a4d1e9f7d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f793a8bf7a57f78eb29eb3c5ed6e5ab464e430045a320457fac40b233e59c25085fa3b29efd291bfe2d98ccf3f1c9b470898874899c57e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h157bf95db038a58924bf90ed55911a29fd426fc33bda65f9d8eac49b21daeea70cadea3e1b25f36f5e66e5a9f2de80bd197c69883df2d32;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16bbc2f4653cb0bb9be9b412bf4929ad0889dd636f555de7eb9b36c432e9ffba54e69010b402d1fb4931f72eb93516aedf9c7f35f4a2e63;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15e4fccf1ed9c9199e8a0a1f661ffdf62e911f427d5273779b6609ef4e80fbebfddd7dbe32acee538881a37653fe8fe6630aa75d4f36445;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a51c77f3ac680bae453dd3a1ed8d2c83c43af12ba41cbda88944c55dc3facef2def184da36fbf9ab534d72e932efeb4ee760c67cb35e76;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14f8d682c17deda26e358480288ce1704cb0b75125efd8398065bae78f47cc3e4f650493c05512297989b29b99935fff5c32a87248f0b34;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10f488c6d24a9a7366b3cb360e34a685aaa6c9406e9b478a7bba4cc41a30f6cc0e7286df3dad53c6109aa2f2a10bfc0490d093e986ba216;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hee58600d9c8c004848e2b69be4b568afab0d5965ba8e64fe6e1bdea01dcbcff0cf173a2354c02eb19fdeb37524971c0f04000908596274;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h44e3bf7ac600abbea22d0f1964ad0172c685c37fd562bb01f1d94b042b160b4a6f9d551bc806dbfb9b61414d6de6459e0a39693f86f07f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bcfa5f451394c67f974e67f4b15fdf6319b815e0ee5d667a7b57c5a8a1a69fc34591ba185feb5c88512d6348bf787877485e5b43c834a4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17456b06a5a5c82e07cc8973c9f6d03e229fbba6ba9c0388fe8053a84ec5f460937f9efbb265a242a3d5ad0d4f1aaf8984d83666e14a3fe;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14d3f1093d62182e0d9d0df7a610174e5bb4ef3324d684195afa92d26ef19632021d60f2c772e1434ceab4d9002ffcbdfaf745d3d30ba7c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f8f9407fa16e2b5564ae16a4f6e6d948920f46dea1cca3846665fd12e89653303676fb0b68f03bec8e9566ab37b981e01b9a98e3acf72;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc852bfc2f02da2673721629f125aa29c962a38c4c6bed3c18ce6f1ee4c82edd0dc26667f4c32e46d73b5711b8ab4370b50c45d3ae557ae;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7bd5a7c47c5a03534df45e93196da33bd76ba0d368ad57a468ea655cb1064e71f928d5ce66fff3da339a72ef636461d4fd2c632129d64;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11e153f81e433c734582bfa084b527794972988c291fcab5ad2f2be4361c61f8da8ff6d90bfefc667b41ec5c931fa850d5024e43add9b6a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h108401eaf4a047b20330820b29e4a379a762dd0240a2ac03e59986bf00f1f7333bf167a2d7b08d85665bb88e9d9e1998142dc5e3a14404a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h58c373d4a744993451a8de5e3e935aadd68a8fe13b7858b9bbb440fc4aa43299c63357264c06033a4d19d5156e4f6950e04bfa7f99cde6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hed5c9790757ead0670eea9044651efd21d43791ddbc2ae89ecb08f783b71d84e51e14aadca74f748d0ac708d98823b709981953d13a5df;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16293c4868e01bd24afc74247b54a885cbe4066daeffc115035803f49ee45739d904135e81f5cccae12e0de4a90e2529c65fce22fbaedaf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11e2edcedd8fde3248940594ebfe0b49d5f43663dc64147df16eb336ad6328fe6da9fbba8fcdafeabb961793375a012d764f4b10a43a91c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1aea21f644ea5bdbdf68abb52ea4a876a7eaffc307d6acd4a4e39134120178f1989ff324532e3a46de2e6929abe2438011ca1ff9d2818b0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h67b490c92bc11f12857299ab9e2127d29d85943b330434fd0fa09f1a0ff97405db79dcc0e06cbee77eeb0bdb458a0af65ba37a586a7832;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha459d8dd8447d6d2d1fa04dd48a122e5eccb3882f78110cb1605b8cce9715fe8b578224406e385e437b78df3f7a2e2fc6c24ea97d96fe2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h170b6f423f6ec0e487f4d1d17651260892040ef147c78cfaf011acdfc31fe8cfeb351a189376dd5f3bc7c5a982a8cc7d36bedca240cefa4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19510d23c0b9883dbba6dc77d0e7c02c3a505b0d6bd53ac186aa7aa2dd1b12f14c9087b733805cbb8911ab6d58f56aee1a9577b70fe18e4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h73519cc5462e04733076bb4459c9a9c9ff996d11295bb88694092cc9cba0d53441bf3a51c5e095bb19ae6ef2ac4b6b4352d0270441cb73;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9c2ebe86e9ee51e0169ede5d2e095fcc10ec68621f7330d7e762322055e9eae1390a5cf12e8374d292d68e51b5dd3548168c926d59ea8e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15ff4166dc25cd1ba7fa86b5773d95ae24ec28cb4b9053a7d98a6876982d2fbb79ce4474e561e3d10bb634455f8de63d7b98222e57c0969;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'had276564f625e80058a8c21af0eb5c6aa686c6d4d8b6310c7a52bdedd041017412b7b10c43ae3bd66c188f0f97fd81ede1a65eaf140fa4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15e5fc2cbf69ea8b888d25e2d24dc2f88c05481e45f4d070063137d6fef2a21e601b04ad1145a8c5ca167da3fde2b703557b2626dbb8cb1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1039fdce1a1607799b7cceeb6b34f1f3706332d0ba4901d45d8d46898ec858849a4829b0571106b4e0f66dc6edab4943c0f871e9c5fbbb3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1833711c1f5c64f10a5778914820899ed992703e60bfcc4b0bcd86e169966ab3505ae71a8819445c2a68c259104755318882572604f2803;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h24b7a34daeded3f7acf9d723a2f6ec4ab3dbc48dae8598ecde31a4fb57689f12506547659ddf6df39369ecebadbe9792a0849bfdeebc07;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3ee485d5bf43577a1b20d1a56cff374dc41254752fb9543c24998e91b3483811d1c6e91ad60841a40c1185f3e4f1243a61d168e16bc407;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h83cb3eb6a31dadfad4b4066e72641db0c5fa0acdefe9a7cea2b16844993001e1e905d27ae8143f705bfaa9a0675ae0b52d942151aa6eb2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a73b6f7410c5387774f7410ba9e4942a4397efabf98498e6d3241f9f4b9ca379249b719b0d3abfc2a254e3c06d8842936421e90e087bd1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14a4510ba6d2fef0632d7fdba4dc8230301dc79a407e34b8ba58c9029c36e85abf2581e38bca52e91874546be9e4fa8e35a40c824dee2cf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1688977a68250ef4ed04e57399c8745c811e6609fe70f3d9a79d4e030d66642e324acdbe1589f2f97ce67d3cb054466b9936a6a0757025f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1186acf6beffddb361006ac8e097ef248d1afa8da4058c516c1ae73ae934fa644b6343bca2f2fd91f29c73f37e9e0119e2dacd14a8f2da5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbd26ac0163f25ba8fad64836938698818a73767e31d82e3fa11a1b27c2facdc7583bb06ce6a2231326e6366cd3e88e215719d02bde827b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h92c6cd4ed351e9578643ed87385a5f01471c781589fda62cc17fa9a67da2ca64e8f655d950bd37f490f5b7371bf9f792c0ea4310549aec;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he0bc6c81454e725dfa6f517a80dfa3ca6096324e105d49bbacf10194c5a32b5a8e523e5375e8f93f96eb076962c6654ebb687e14cad4f7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfd6e8f8fd6977cd02006c61072ddb323e55a389255acd3db7f93a8f81d51bf77cb2acdbea257e65ac2ddc821ee4a695bc1ca5975e13d23;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8be7808aa3ad8f42045cfedbe048c536a3683de08c665658d2022477eefb7ee870b735bf78c1113541f03c8fe2eb1084fc6b6e42ae741e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc36702b45611334980f9220cf731ebf3a9684330f00995ae7b7253872048ac5b4b82ac6d3f73a3ce16ba388dc7eb23d6ab0b59a8849af9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1382ac3addc74762549d2b75a139342a151ebef3bee5ffb879e5ee404013a016c67c6574a86baf2a989b9705cc82849b09366eed9246cf6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11fd6fb79cfd8fdd53404aaf9fad3666c4a15ee900da8c98a0417c9a6852943a7b219d2fcc177d77134d1f2d9c04ca66da297bb0010f63d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h191b1e39b538275748100aa69915af9b960b8150c0bc65fa86e4981f67258512cb1608adfebf944eb437f4c764efbb62c370090477e1f90;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f3fe2db6f1e07cdfc60f0c540e64b3bbc52d206094134026acb42042f11b4587e3cf5b1f3ed15c83066c846f3a30332dcb50e6c3929225;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heb2df92c3ec9e7e141e77d5eb28ed8588ee4ba6657d7dfe9236b1d3b3a22eec531653d2bfe9b5cc5be2dc9a52aaa5b81e4426c9b327848;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h105ac6fb986149332fe207e9641a5bc6a6563651be1ec4c109fe865df8fe5d8a29793abef17b8a5ae8c105a16dac7cfd738bd29afa476af;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e3f982eb0d256b6bc431a794a14152ecf51ac18d8155b833ab71b8573e18433017a4b8009e08b2c69a948f909fa389b8994a06bd8b553;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h51c4f96b4878883b61486a554343ca98334b3d135df8530f17d61389e49f97f7d6e8e6bafc45ac5f4299fc4c71a8466c4b077703d25eee;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a8f2f33ff9a43330fc5849159c7542ee6d5f0b0b904535d193a455aee0c81e30a0c4e3f4b6a244472cad5dfc6bbcc2f8faaaa63b6fad7f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2251fbb61059fe4e1be7788ba5a00bf657bd487b76309b61516705b8ae71d77d5fec4e533cb8d457b55e4db68a03dbfd839acab88dc128;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcf6bf22fdae58870b95d13f872e164def2a2d83b4e8c169b3fd02f1ab5916bc83ece23b379dc5a69f561f7a860d8554202266e21bd7ff6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfa12eecc7a5c007d3d0ec46959683abeb5d4c3684eff0cb95db188c04d9979b7af4e94d165fab2d9f48ceced36a9397bf58dcb38c9cd11;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2bcfa0ff9336c3c2474872fc5cdcae6287723e468ca09a0dafe4285c5476cc3317e03c85dc45f4b38389e4254606662a6948191eeb8bac;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h34eefd3c7c60647cd9c933589fd4ac0a3e2121f0b455e465079125c0a3c083cf8ecf2c898e33b7339faaa4c8c66735ca7e11990909214e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d75c6adaa7043f9bd7c2a3e8d9ba7ec41c09505f4abfc053b3dc58ad55633190b10dd621d18e320aed1ebd79d7fc5ecd6f601ef4188d22;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h113aede47042cdfe29d526a709870515a21905697a2d5d9f8c815348a3bb8e9619d2f2b1e5f408afc2bd2a6ed0cc6ffba0cc1c5969d57d9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd372b251f4c9ac707c6451e47e177dec0577e5d3e1ad968816b046443b044aaf272e8c2631b6735abd4cab199519ddaf8efa41b90fa2e7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc93589c1232eb30dd00dc9e5dbff067613e0abce1c9feec5c9dcfaf8ebbb6bbe6f9ced8a543ac97ce99fbbc1306d03ebdf961eaceaab9d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1527baa0c21ce935cca4537a46efc53fdd5c5a1125ef9406a9ad354ebb8fde045b06d85b097a824327b884e520541cb0a2ed96dc2225508;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h78ef835ad74d56d63bf3f0e6d8f32785107da92d6183f8d018cb21810d8f8f38dbf98e6809dc13fdfc8da3a5c5864e9696ed63e2503daf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a57823913d685e27310abf5b570191e1e07d397c6618a77d3849793dd39503448c77003f58133e3788d6bae33237013ddfb66f7bd8814d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19ab5751a1297868f63f44633344c38bfb8c70ac7f81926ab3671544b4a9d4c16b285d66b9fa5ca6609b0834ad1cadfdd338df1677fa72f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c7d4d06a84420b43681e127db14f8ab3dbbb59d7766837a8f0d86fbdbd71b5ea64c1ce723324751069e0013b1f13f993d23fa90435a2af;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9b34c44acb281368763f793ba01a8b6140a09dd4954a2fdf1008a7b37abc6f0fd13a9f6fa737cb59c0946d4e45696db9be8af37ca24da8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hef4a303501ff6d09cc28031adebf254a58a7c996eb15044565e75734668324d20f189612420ee2d02c8a5146df657313ea8bec38c06533;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hde808c72a4e65b778f1618a13cc28dc528eed25f8f7f10db793f221b5311369eee7f28259a4663d631a15b70409dc1567ffd812ed24fad;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h81145c488d2e9309ad61c8939ec1af84403735dc10bfd14b81bc6327abc161ef140771527c8fb0f9c275d69332ac250640988edaa31dd6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14b3da3782b9eb4eeccac85d61c0d6eb38bd97ca3f0ca83eafa1f010496655568b6ff0f4060dbd1593492c853d67b491c127431b971b491;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h66f237b9bb85bb0b50ff541f1a7b8c07fc7ee0d945a26125a5b80667b798686877b9ad60760594fe0c45f08db9055f04132a92a0830b08;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6db8fadb36b0e1efb22bc5f1ffd8bb119d618a7f51dce5ad311ba1529d9e4848b8960e5e361742078de52db8bbe0960b46c7cfc551c409;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h80d3a96bfd8977476efd531f5ed7ddcc430fdf5d4ec7443b7aefa97668f498dcdbe243bcf3d857e0f1041a6f9c0da21addb6b762c2b187;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c256549501efab80f925899f9a91db5c75cc7f156d94b11afa0efc4d1ecd43dd342afe52ecaf8bb453c2a67bd4ef850fa71c93758d43e5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he2e81d5c492f8924ade56bd5917493075dd61faedbb655a609143ea440d37c5a8411e6a31a779c4454af756e40c0109c6635a6564d847;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1de0eda2df6e7549c8bdcbe5a09bc87c59a50bf08019f1e771e214719350762678a6675d4d1b84f1cf536e18967fc3f5d004f9a4f665793;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2a8efe6db0d77ed58500de267069712793964ba362caa9a324e820eb6343ecf9e3960fccf969c7cf801b33ea104cd49d4e5e0e43eb4827;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fa4e8a3de92a7739ec2aa0e6f7d265e018bf30958f6178b5da8ae6f365a4738855d43a32b3a60bfcba018973e2722c4682266de29b1c77;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he2e6f6a75d53b1eafdfc4cd4e76baa9efd3b89093c551a9cab778a568596221d93010d3d89777cc5b703fcc42cee0be677724bba39467c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he0824ad3349cda59d9a5abde3162251d11c3e01b457ca58045977b85d3a32520368026a40b1b0260c5de294805f2db3e881fe4dab8ed8d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e0fa6b57f86fcc20ee4f228a0e4b2180fc16bc635acceae65417f6d73a16bd677a47886903828d52d369001c8ca83fb902c61889cb71d6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15175c8a9be7c7d3383500cd3404ae2672dba33289b116dd9056e76875796ad236f509f400e2aab032ac6ff93a1dc2f419f08dc882ab011;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h560bd0fc5d26f195d756627c4ab7369593efb4d64c2bcafee3b4258b8b28275689d54958394cfe9503537150f375ce8dd29b39dca46048;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1da1b010ee44cff7452cc7a95dd49732b21caa55d9cea69a2f12bd100fdcd23467f7bd61f465078afba39c73558da5e5ed5042dce7c51bc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h81dd241ac8816d0f1924fa82c49c335e8bc81a53b50c095b5a9bd798e6a41ac58c2acbadace6a9f3a3dcd63b31fd8a30a325d5f45d651c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb3a6a3dfb73bb32fc5db5a9f3076da28932bd48e49fe41adecfa9606e031ee7d050ef87fb2f08835c3f1546e4adfecc8540ddb4a43abe2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14daf2c460b3d67b785d629b2c372bd9dadd53d85f98b02034cda2244162be66096b9f6b7f976dc37803ebc1e9efdb42f5653327a2a8f11;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ea01782d88b3d01772a6ed6223f188eabb8c2184f2413dacc4eab76e825df04adc797c10623aed7bbdd73e98fab464ab38530307d11b85;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he9e706f86dbd9073ec646e0587cd015416f2f0ca0500e4a36ca282964116507509be2a200e7ed6f43bdf908f7893626fa08bfcfc5043d2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1925dab67ffcbf263c54feb5db7dad68d0204f8713b46a4161e867ca3437d8910f050a4a1caa7b69b54dedf9bd1dead93f5f239e84eda86;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ad5e009d7d3955861cb3791101f5887f81fd72c5ba9eb7f9e6a0f8e069b503050576052eeacac69de05dfab731cf5998dead63d7a2c7da;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hff17632e379997a1f30ea4108b4b8b10efda62450e9d5ba073a77d5b85ea5d2bd940696831fba6735dac68c89c8262e871f9fb1aaec008;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hae7633de30c74dca661964c378f84125508c06d89a775e8a8aa474cdc4d18ed1c12991206b0f0a18cc8aec12a5de284bfff57ad323b96c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcdc7ff071cec94a9a6cb67f12480afc6c728eabb252df55c9322d1caf4ff71b610b64dfc5110601cd386419d159c3cacc07e2931d0f535;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf295ad9a88ec7895ef0a3cfcb260fbb70c8d87bba2de3449df19b29a25511c7e57848f67a05561eae9709d971c23bf8552f5f2d41ff38c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h156627ef6b1e873e423742bf16dcfb8506665468f416225b0b4fdc2af79567e597ffd2cf2c2d5e992e358febafc311e774e646776226aec;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1258f0c72c53ab44244769f012b0fcaeb1c39ebc7ac4fd166d11cd9c27904cc9c77958c721fe933be089a4110aecb86d3d9efdb458f771;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15d5daeca03ff13a7ff08318c499586d65503d211926d02643af569421eaccea2dca844484b15438b2fda7cb726e66884905dec2e1716a7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1475d897127345cbc306c73eac7fa6197cc7ae3526498376a8f3f8d2dc41d9f77f0aa00514d89786b505138f5eae56119cd9e739a13c51a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf145633dd1b732760ba659385cc2485ac5e70ebd5f7cc2b074f8d1d481196203654df37a0eee47952b47d1c9b5626c42bd5b30a8663619;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h53661973c7d9a43ad1abf2ec8ed6816eb5792c2ae9e991715dd800dd4f072ef3c0e4bc27e68529aca7f23a7f9c2bab998f875e303c76f1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13cdbf2cba35ab811929abd0f4d3d007b1a7773a9f2a6a870922b3aa1fff864e55bf8edd224f77e5572dca2c6a9accd1df3266c5b4e3a21;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17065656a1a9d8c2cb93313cd7e9ebcbbdf4c4ba3031f63c10b3d51762c5c1d01e94553b6fa2bdbe26f27f713bf8dfb1ae1f14b8bea2c60;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha5ff137406216087a57426744d39dcb82756501c3bc4929201fbb23b2ddf7163588b53744e5258c93f681969d52958fede7f03d8d10968;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h834d0848d7894ca34dc4243749759d1bb78aa79b36854a7df970cbb7520ce4193292f05384f59b501d9721bbdc2e100078948272d20db3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a8f19f7928cacac2386a515c54d6a3b933b6211a78d1103c63796dba65c5625f09575a64fca261085ca9bf043fea8bdb303c3493f8559c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1592c882d93531e6b9e1f479b4557be6aa55c29919fa1b6d631ba24615aaa2a92cb1cd5e2959789d47d7c98f6cb684a1ae709c5c6aa1a19;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ca68a4042d32ce88e9379422461ffaf51d3a0d64fdb760cb73aaa64b0cc0afe01f44af897890aea49e6130cc6ecec94b0f54f3959551b2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7d614956df4d9dfe74d4d9dd04f58540b9e79487604cf111aa486884a1d82dce82cd2a35c531ca696c1b772efe568885a43925cf36635c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ea9c3986ea4146f838d21880c16f469be8f8b17a13895b4ef1cffcb8a5ad923e62d9193c511e301cc71d8f27043f2a928d5ecc92749d7b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1673eafea1ef40f232a0d118ed447048d08c0766db901376ab92e13e5a2f4e0797ed37fd3ab9aeedf63cf753672676582b67524ac9da6ea;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19244fcd65a8eaf901aee4ca087b866ae686a9914a1648f09cf5596462cb16008d1177ef73fdba477d3795a3c8bb9484e61b156b0c429ea;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb0d25bd32112a92638e409d35e971b64fe5f23b62b6344b2a31ae4d2d2aa71b43e9cda94e1be0ed0c36d9971a9d1af931f7440c3a85b3b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h140a8153ebc93eba2de1a2802a63a72ebcc88c19451503f6e25acda6ed6827c874c8a5d694146e91bb5a4afb8bff49d016014d851a18b05;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13c2b7fced3514062f9c1bfc2df27396c6b62bae250f986691f3de7d657dcdc153231696ef1b9407adb6bedf797ac2ca9f336c25f883c05;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc976507509d2764225bb721b7688f36ff3dcdea53e5c22314179d628016f9bbd510a7529ea38de349e475d9f2d5ad55d0551b6902852f0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h79e6b55449b9b52e1c044f3ae962b40980bf7829d4d5eae78dd6210fceaaf9bca4ed395884c09530210e5b104b5100ba1ba049c0059445;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hca3a7d9aae3b98f1f9887c4365e89f3978e925314e9d8ab8b7aaf4435623d7b989c9e548da83d29df58dc4d4bd6f29bc90ab78d4eb2ff3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d00ed2d12cc2899cc3c4786e3685795c589e0a9dde3cfbe2914f8ffb2821d7f69ee49fcdd8a73649d5cb60fcc8b3f5139e5f0c5533525a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he5d7dc51d8298e73f434baed2a60c35dc5e8dc6508c209a244542909b0ec754815a234b454cce93c8bd450199c207a21ccb34754d32dea;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5cedb38d2c7f6c9240cd90ed4c398da79bed263dfa91b66ff0494578d627378ebb48561caa9a9c7f4654d445c4e71ac3d7ac0a3fb6397d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14d031c31b207067cc7e9e9839b8a9b696ee11def30f313e025505705af626ffaf6a6ec5cfe9783ab20a7b2cb651da4be11db1cad6ac4c5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17868db0b1815bbe762ee23b0e7c899eef213536c29693d5cecd7df69c4744956bee8e679c739f1a8b21b60f5184100cfe4e7034e146b1b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17c833e232cb9746168199a92293ec5c27bfeeb33b8036d1a45d10828322aa469ad4063eb7e36ef1792cafa7a6e201c9824e678c190a553;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f221231d4d978b485d4eb6f639461031b12ffcbab68d143b8da31e430c2b4e4d2d1cb6d0a94c5b8561828b4820823a2af4078df4327394;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1548bdd9adfce15714ab71f18f3dbe99fe94f010b1fdd3a381f4d24f00e566efecb2c7c866297958e5c69daf9fdc0eef4c06ebbd4684fbf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdaf71d7dec906c01f690e93a099739cb790a3b7ce975b5527079307c5f53e95b84c32ed7f57955908d5c60ad538025fae29c6ea7d11f02;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f02343affbbeebec5223b98e3af8756813c6a0fbfa2b632da61522748683797aab872c677d7e839f703f5db3908394649bb2762af68d2e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9ab53237c7a954a70cf77edec3ea0a8760a85737010bef128473564520f9d8f6fb0377a4da569e924561741d0b455c658d4e27ec37d662;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcb64fa841b9cac585bd8398da01db4a93feb764d528751388062f25c88a8a38728f3a2f1c7213cd3415c77709b79c0700d87ea8467560a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he1e7b50438376cfdaffc2b8bcd7b94a34027782a6e4f5339e4eded745a028f797174574cbf6c3d5d5c3fe08817a7640ea26a76b7395cf3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2acdad7568473c91be5efaa27cbfc94841dcefd60743d7d485d95a4fad7c4c9c19eb066acaccf9f42e846b0f9cc35aa0d034cb6f224d65;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16ec59dd82230988f71ebcaa367802a3302546c5cf797c428632fdcabd750a0b1329d2653e3fa3a43ef7ba33dc9a9054d2d3b02325ea552;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14ce918c0d4c26707b7093f1bb91add0cf17f83afcfcb3c71e29b31745b730290d80e022953b0f32bb17653b67ed6173e98ce608c54c0fb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a2bbcb2387650a844b479298632b4d51a8ba2ce5b2460ab7b8db30c71de4c100b4d08e4e50e4b030aec52f1923b2ee63650171233f4318;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cf6797cd973fd97868867544374fe5f7da44b4d610380273cb0bd41cf0117537b64e0a6c8f397a65e6437b7e330e675570569ab2144e24;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c621d72a3ef29912d4d31a3d3c2d0d630b05606084c25b48e50e18a349dcba49ea7d5bcc40de2d1326a6be791c4b2b308cce993975ac63;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf39334c36c9da258a419b916317ccbdaf81b4829981b708fa72b2039e3b913b4bc56be7e145c63e87af46a43ab425f3ed1e291fbeb5269;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h352ae2ab9622c16fda26a4ae5ff707f8994bb11cba23ad8ab0d4eedccfbd58364327cd985c2a9998453bdb85ba516a49e9ad6539eec071;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e6db8a850681fcd648a0e40366099dbf2f762fac9e2978ffd9142aeaba13a4c0337c31e9ae0b07e4e4621aaa4702e3623256c905d19750;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c678b0be6e1c3370271aeff5fd6273332c2f95b31b117214d4004e0f96c9c6d4d4ea5dfb4c4278ffae5e59a0850b292712903c6cc3a7b3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf57c8b6e6f1110a6b302705936bacc5ff3e1e7b184a677f1eba50f3f79901add98822ba8ec62056fd6eb0e179d3d5583bab02b01b8018;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9e1cd13d470703f4a45b860f6502608b073c8b499fddb1e080ae0037be7d482a62407e184792bdf6d6b68ae2aa8cb9fe524608b7a6b77f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd0a00aaac1af937d4541e43ebd53cbfbc6bec988015610c4753369bb75c5a6c00626231aeeb82d798d57a27c1fbdff21dbf724e557605a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h46b77c8f954021ccff3e7a8c0823c5fee655928a1e973b1fb18d0f99678784fca57ebf9001f7a369ee77859f9797d1f5b6f5016dd74845;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha2611a8aee2a8c2adf0b2327f9235d6ae2ac90fd5adf1268b3d88bee770ee5383103202583c6931bb72bc1126b90390635daa1bcdbdd94;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fed5ab0864d788751876167915d7a3df037ba30733c611cf13443003cc45a14311be1dc8c57904ee908f784f031e6e04612975495c82ea;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16440dc0f9a4c0bdd064da09bd79af962d3d2f10867e0222288e0b6bed701d064cf5eba562602a6067d874a49429704a4948cb91b887969;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he97c91a8ae0728f51aa97582aa677336651020346d54422a67bc23330df39026febe1d3f3dc7f3669c830b8ad06ad659719810a99c0c10;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h146e08a1d3ccc44c300ff8a766c87f01803a3430ee8fe0bc836941de3bbf2089f8b4359d2c355af19bae0b1ff0c0c74391b61d0b88aeb0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h544385431a160c7cdff2406795a079f50025fa71d64cafab42b32c78e90e664b7211c9a664fa74b37416d75db5e483215e615e3b28d0df;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a9f655baff95e692aa19abde2087cc53a7c1074dc8908609e65d4efcd809f67bc7ad9b9e0ac6fe617584c8755729e509e3a5f015f81b93;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb3d9fb9f4fcbdf6c21d7b38d592285f900df1f468063c8aac9e9bb504ac227b766de52ac8ed6315e87da805d6efcdb4d7c8fa3c6982302;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heecaf029857850937c45f07a81f29505456801773f98736062c3cc8ba23964107e00f22b9386500c4201eb0ccde302bd55bbfdca1facef;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12134849bf1d4de34bc75f94abe6e524f8d8ea9099d3d6065f5d2459ca6f722125777169f19ea3867def977d61962590c46dcf61670100b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h146857ecae82ca5d0cf26201d4271fcf2c34bfa2a29799f32ee07992e62a54709bdbb0644082faf829ee1dd0abe72683a8781c704f6a27c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h99ccd9ea5f1f5f2ac8bed71fe21bb593d0ce64d97079f6bb9326ef661041532f279ddd7e6e6f04e2efa71e654ebc621ffd9dea3409d66a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9a39f5e488b81342d25ae9db38b7daa003bf1c80d31d1bd4d78f67f0a380cb970506682289eecf3ad3f35ac655772ccbc0694589b3e9fb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7b0c04ae0b7fb42d151734d0a649f50104c499cb60fc425bf7469bde527e3a57209581285624b246a88a1ad42a330230038cb30d853732;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1750f88ffbf54f7f0998d8c4f767ee9dfa0d34a6399d542794d804811506bf8a5669a550f79f0ad8bdb6f05d613b95360018559a74d549e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h127618be4799bf33c3795b11ad8fe7dbb571640a4fd358026bbbcea3083eb2a13ac311cd9e2a32030866722ce8e549c8d80b0f736305904;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a1452e046613d9ce410b44229d3629444a47ed8e14d384767bf01d0a2f0a44e65fc0581d404e5ad68d6f675d0394a91a1be3a4740956c8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb26edcc27cc43ad94c7976dc0938619ca85e4d0231b8f1e51eee4588e4a7fcf2844cdef71b7471a10d963399b90c002da7437b93fda8f3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16acfe562928372dfa6081ef7a965020b30b946b983a238f640fc612b58b7106f529c023c33098661c7370b054ea735167db0e5da8bdeae;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hde7ccf78e47cb2b7c034d5fcf3946d68554ce8263c20bb279e706331337298b509d0cc64d364c96da26c8416234db83df48b9d2d3fa3a8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e5d2a96a1928f80390fe1e1e6de99c31cc14f4d6c9f4afd3fd615a9c7d001af3b50be7d5d4559c43e0c07164378df2da7b781bd87d5d79;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc28fd36239af7ee9d138c1801029b00124054c2229eee3d73b7af651317925c33a239756647a760d058a35be748579e68ba66b2049bce9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11a0f3c881df0baf592ee6d0335ea8c8f2085317d9ce7113262b268ed045633f91dc4dd84d9444fd71b9c0470c0eea6260b3cd87452bfda;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h729be0ac590b9b571b770e33f7aaaaf8e9b2d8830b1b708447207f69ccdb8937f086c7c63509f6d85b47632b24306ef33c0845bbd9a26f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb8161897c3962d46a5e52ac1cfab1b06c4b49510aa008350c4992aa27bf1379078aed8e7e119d0c28b16c64af0626305c823e6f17e759;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hadb9fa62e85710b36423ba91b2f00dec7f7c3924449be9683af9f5b823c76999fe4d9c052b69d1de06896ce8b80e7a1dd3ab9d3e8ba411;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb5e10147dbb4dc251fc46ba2e4f900f64d3aa576f5214dd89e5069d43c0918c7631d91ec020c64cfc652a266a734fbad35bd3e4449d938;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1399f517921e383c979d49277c635a34e9a746148600de9d99d37933f7b393ba8d2b8ba85a6f0bcf7f5104e03672260a43f88ad0d45f3e3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcde9a67b2dd5b1627715aee661be54587ba72f1d88f66f425e7d057060f2d819591605d0dad7f989b9d0a74a1b9d912172ca9445c76051;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h142514444132b0dcc5473156841630d095a2adef585646ffb93589f9baa5efa6db8004e6fca78f953af89844623e8cc6ddbbda89582cf5b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3f63f7cf37253d69a7ff41a19923a287d4cb70a88fa64687572f958f97ce3bd1dc76097fece3d36ec7ee7029c6836ef77e2884c4c06363;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b8e36c75d303a61d4c7aacf59513cc3f59181731f4990548bc5f35af2c0f34aa0f4ada4b5ea168239e91925f852a707c7fb77b58f98740;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc517044e12a5e96527471980c3f45e2592707cfb622e8522509d4afcf2808793a7346581ea8578e0fc65fb54a42ab5e41386b140dc4414;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9830d3a473e02069a0ce5e8b62c204d9273486643d084532ab5b33cd7083622b1bd81256862e1bd741efacf86fd3f6661998de6208e59c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ca57724d7750ba70a47762b388c5f89b0a9cd3519d296f45fc5c26577f2601431a371eb5582c93f586b4f87a9949c58c2909241166bc1f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd1c8d456a7756473a582e4cf6133f77c77092ce70a1a26f8be093f7a779338f6c59663dcf990ea4aeb1800d5607d07edee4962983efe47;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bd2ff2cf57eecd252c01aadf34d8f2e3729981d862dd3089f35036b639ff74f81f7db24574f954cbc95b144b0a863396cd557de6b5fa5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha5dbfae2a181fc615a8cd84b756e24b6f386c6d07d3e1aa0adcd477ee41c1313ee5ea1b5d7f8559312d64249318fd91319e9ca794c9702;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7cd103c3df7a9917f3d49aa01dd44e7645146ad36c2bf8022025882a041593971b203cdbd409e3a9072f4b541df171073874566f695e7c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h110f108f2c29b779f279b4f498cc8da758170a993b7d31e5361ebd2a4dd9cbc791a1498fb1c267e7aabe25ac5b29cc3d06182303cd28d2d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4f6fca598608443fcc78b305a6bea1728f2bcb90fe59be535581500625b62f5c5a6665d677f70fe26cba3b69c8463544042c5ea965d998;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d0e3a8230eed2e8ce545653948d37e0abd8f0c219f7584ca9e7289b873b28510d884677fee71a93bc523382b4542ce34aad3c57b32a55a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e408ab03696d9089df56edfd9eae08590a3e32cd78990e15c2215b9a988236b08aaabdf9b6d42edb6357af1c66cebd2acdaa4ee1fe543b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd6e5faa6e5e314b8dc52696e7c6bad8505fdb024cefdfd5b69c77fc7ad7a280faac88f0a00ef290e9ecb5287c3b276643a64e5f8570f5b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15269bf88f966d540e533e81093641ca444b0b6251cdbd2264b53aa0b3042cd616311c7928fb6584fb6fca44fcf96ae4d8c84a800635cbf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13cac99bc723861a767daead3622f8a38fc833ba9735595490dab61706a95b4cc92015cc4f433613224dd74bf4398b79fc47c63e26f91db;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b888a26c57a085b439b44a6c41f51bb614b16ed8c3bc34a6970947e3f6d2b68708feac5e49f6cfad4650e981ff4548dbd2878af87df981;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13c0706f624726866ce71c832364a3a940c40ba890347b3b99dd59302065f5483ad101ebb8eff963add0af4204ee8b91aca2d9a352b0be;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2f6e1828dbf575f0d0165009085a4046372864cabbe0bc11e87b040f4d7f3c16d648bbb3ad0e7fa341add954f6848139ba4dddb7268807;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h184a2c49a2d6b110c634fbda0f2a1bcd70160443772d3d32d166a60617aa8075f9bbe5bf9cff5fb9ce1c817c0928e7ef931bca98bd3ead3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15178320990977a4df7f209c1d04baa208fef714a37016c3e087a88ff49b85d991adfd0007787332182b564d53e6f5b721aac6eb2cd83e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h121d9553273359151fd41245eabfb626f504f51c6fbf7138c61954995055c5cb9777e9ee6c59268db4696672be6a7390162ee73d57d6de9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d7138ba6a681782ea7598d867d8cae9dc5a814b3d1fadd25324d886a610782d8fda5f4e7fc2950b498e587b5d9f541695d7bac0cf09bd2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f579f6b005dc2bbbe867ceefe11961df95cb4b2a7421006cf1800164348f45e692b522ed243b1c5af5c50d976640a3ca26f49c04386b2c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb464eb8508682585aaf8520f4b2ebbe6c8d48995d43eee4be5b270096d14f6db9ccdc858da4b780e8485aef0b02b133e05dd0b723d8a5a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a670429c6cd941040866931b15116567864c13e095ab3f39f0998d8728e205c6fa609af19c442b8e53d59424e37130e8e7f120cc3e042a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11bea1373b85af644e26644f348318d855e54cec32689d5aa412409f09525d0a8635552f8fe9440159d8ccb6569f42bee228a1dddd9be6f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc8cb62bb859de68e64210971f4f35da78efb2ec98fc5ff1286fc435036a6292b3800f6f21f479ebb0ee76fc126e16bf5c6d065ade0bcfd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h47a5d7531e715f9d736af47d793b3a6ece2dc6a6c91294165d535ce69541977b4a35aa0a9a66820eea5966d27541c78b0efeb8ce318f65;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h194adf1a299df3dd348585e5408c4e3eecedb621f390bfd7e08b12ce70523475387d4b46f453698ad7a09de1d3b56681e025093fc2ac93b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haebc5eb77c1a847490185af2a247c8294d191d9be8f5c7073f51ebd4054d6fea22d3510504f933005cf865212f2955339a7a17514c7936;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbc3c41246dc701988398c989ce8f87a295b9c8a96d0389110e9a629510700be8b3030347d1502891bbd49ef91fdfc0bfcfdb4a6ca6a9c9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc5e972d46852118cd4138477b4a659224dd329b522b69d682699dabd8a0e5d64d6af363887fc39e8f2879f6ae2639a4245f4de707c1734;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b3389cc07b05738dcfad9c5dc4cff46c4bfb03b542c3559b02e5d80c4518f24d291b94818df7f6f7c47efca936d8066edcba2d235f38c7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4d2577b98d84402d85a4e11c70f796e1e2badae53e479236b7727c3a3af5041643fea82eaffa7712b0533eda0fac1d118b954dde259e0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1468c0d42904f3dae12a834ddbb2c544a35f40748bb23c57999fe8e8f61294bea3f41b9dcf94dfdbe05bb2ccd0d478491383e5cbfe3214b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17d6029a7354345d51680f53f7c9620c615f35149a4e6ffacfd43e4d1d3acd23fd0cfd26a6d60e9d88d585dd48b33a225c8bdeba7ec978e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h77a8d7c780381244eccea4293bd1a0474bde3fb3ed8055ed4eaf91f4eb90a16f4c0fb087adb9e865e1175498168f26a373c7fde2ed79b9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdc2964871af46954688cf303c52ba525ee077bffed95dec9fe9967a55b830630601454331709e0072d3b124edaf0205efc4940f9775006;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13b4552e62efab33bc2f1b3ad8e05a64867483951d980c313108fdb26eb6b2256f1ba8466284dc56ef7101010627fc4022a9c8cfbad856e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2a7768c73aadaaea5267a8c6159b172b6e670558e494297a276d5de5bcf648cad42cf60e9b63bfb9c50570140ed76dd517aa56aee13c00;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14ec6f4fd6e49541aee0a429ffb616c093826ec169291075974cbb46955bf1a2e7e41c48e1cf6bd799e1ecda2ffcf54f6922abbf5c5cbe1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7d308a98db9bf47ee33600479aa1ebd46b4757d5a886e0fd0f5135f0ac20842339b6e64b937826ce9c2ae979e080d3f313db41997d511e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha5675762919c5a0eb7f5f6f46dfe287cf4d2cfd8e106628ad7ef2d7b2ef85a5cd4afa554bb1973a3b0125747a0477e571d9e4a2b853ac7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ce566201b750ab603a76a5cbbbc46f4ab65821a3cc9f45efc4cb59a80846bf1432c1252775c3b43025729b160076405a196b3d61ac0c4d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h88adebb140dce4a0266cb20251a91f56df6f40b1c91ed33865b6b674ea5aa64784320a9fb800fe627c3facc69ebe3e8995bf52549917f5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16af3bec37bf63be823168dcd479519b4cadd0db836c6d7e7ae6edb8a45a9bf466ced889441b42fd090a722efd3294036e4231145e74dd3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd83e0436c771ab9dce2f98e820c539e314285ddf38e6acfb0a7bc62548aa3f9edb5b7d20b86123f6913e7c5ca15d44cefff459abc474a0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3a87ba3ef46627341358c0c173e34fde96492cba8c2acb3f2b59f76ed2b47509fb6748d77281eda414b8d62f2856206e5445cc24c226b5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b40ea97abe7f67dc11138a5be82a0f7808d7451943019b4f72652506c9565fad6bae902ad7c900768038699db6bd840efa00dff1679771;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1918e6a2975d935160b27297bbe7ef4ea65dca5a52766373ef6529f2012c2d18dc6cb592cdb4a0e6c7faa244549f2fc5c135546fbdaeaa3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc8cbf11be12c8f8ef8da35b0d3fdb3526062d83b1f646ff5a21c9e7dc1d62ee348cc7b53f52b8a9b406cd53b8d565436c2624038e93242;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2d9865bb57872a9645a8c717c692df1fa4d60e7a7fb85c7048bb428d4278cd4f2d4803824326ac54bcae5c6604a80d7665c6aee972fa62;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14543eef2002d818cafa18f58d38d12884609642482120f2a4f0bed4ba0effc0495c19d7c7c38906b18df96d119b24a45bb2c5234668360;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1441dc9df89c9ec67dc2796ca440dd5a27947a7f4c0945693996a15ac717d2ea428ce7244cccc6d819d7820166cf3a0924512151bb5a47e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7a260f1bee26d62ecaf1bcfcaca9784464e83d61a4e39f3febfdaa15cf5cea059ae503738a800f5669d4b55dc99a37f019674cefaaea15;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h66b01781e694c23f6956ce4b42e7c916eb85da863c88cdbf302b6f724bc90e900dc74653a1f046cdbce61e205247c52eae6a887d9d09e8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3d3bcaeb55a7bae2a73ced96bf4f6d86bd6c7b3951f6fc2140aed0b7a911b823320ecd00b653f6bee99d141df59c7f195e333d738aaaa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2ed5c24812456b039918eb1a08d6ca0ea2fc9542da91dff2a264f6c09188ad68283b516cbcb1722e00ea3e15632e96022a52deb060b0be;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1833d017a06330c7306b4fac02793484a43a4c9593a6f18adb8a57ae01ee6d1f761cdc4869057da637cdf2650e6a81f84b54318b508af80;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6cc6e1dbf3617d8bf38ccc4100c2b55b1b26201f2479df94f177f0389c199c8ff92819f7c2d21165d601902c84a50538f082ce1d14c7cf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h118cdcd67aca432e7a71fafc3e851e764e2517d648f2ba7c6012d6f60216486db74a3478116b887e97f9e58b650833b03cc59db67fa446f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h90ee7b8fae8bde7985888289e66deb17d84eb782c2794259efe0a5fbb702d9f6f1571098e346497b963d5be89d3b90880045ac0f87742b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bef4ae698cee45a0926a009aac36ce583c32b12d971f8c9eb67d4180d1d8dc4068b03ea535472bf8ff7e9d6566d6cc11d6d4b33c9f5852;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1920f5da02a1a24035debaa1293e52d66347c3ea15d845768c5354dd7a86c3f7ec91bf3d8c021a1a2aff939a3d932341c3292a272a37085;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h94e199e23c4b02d93eb78166c74f7246838f509e63cf3a4c6e40cfa9491802cbf6182e7441cfd0dc9a2beecefc0dbe3c0863da01f8059;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h29da471eacfcbef8c5715c1ba1c1abaddb770ed8cbcacca6da30fa2845d36f2a9ff01a829b9025518308ea7c3632042699c62f942b8959;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h134eb1c5601a0122161a2027f3c86966cfc2868678127e410b8ec3751067a85a6f5f62d56492833f70293b38b35e88819450b3fc93a9111;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1db0000d21d8d2966d5746a6cbaf692548ba6018353e2eafa5850ca36483e48dcc49e92f993c8894cdebb84e2a3a02b0bfabf777d3efcda;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf49086a60352c94383cdbe085f1205cfa5b69f73d30ece415b5be8d70f39bba567a32c487eedd6b841e8aa112feb5dc52e4864d7c7be5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4f6cfa6a053e2e39aa2d50646852143b2a9dce767d4de430a573982575f135a3902801312c2052b5f1c8baca86726d8bd6e8203f4019d2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19cd45dd8dae842c68aea17456fff5814dbfa82daa7798d50ac243506d99a444e6177a7ce659446e4a80f47cc7c007e625f4f22c51753ff;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h130de857f1dd19c5c4a85661f4506f80d587f7d6a92a80a2b0c8bd068d1fcf34db42c1171eedec44fb489220396bd68658c0dfb26c1f09e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1573ffb8ddc3f9c6a981f8d8c3d56f552542d8c20e66deb84d7c91dd33f4001aeb25c60b01c1c7290b003605227e71df93f79891e35e595;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9ad3218cd7630adb25ab2cc06dcde594ec93991cbd3116599dc31d86e1be42771db3c73737af5d76eede317b5669fca7883bec5f9d691;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1653da504273e06f05cb6f663ef0af781c72f4e165053d0241994ac121477e63385d29176a3b8e8af21ebbdee987419318bf2bed9c82536;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cf2e6870bb171a916264b48f2580244dabf69319b269eb0f0cec215ae67e0686f15c1d0e37d1f0635b6928a82e6ea267760958da6c6899;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h135fd9bd3fd54d2ac1b3e82b1922702fa57dc1759a01dcfc9b288577766e83b04dc2a741646ba4fbc2385e490e42e387720156b633deb88;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18ca9ff0aea0c2a976137bb0f66ec2d8b49d69ba380d76c91e43dbb000d26c672d1a196f353ca42996a4dd7d0418d6a8a5cee4fcd61041;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5c685debbd556c52a3fa21bc3e4ef1dc1c2ec1c9b0c08bd65875efcfa323449378e57b8be3cb14ebef3a42905ea5a99497f6b658e46328;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a0fd26139f770e570af96933d5d9cb7ff9ff4944d0721702bf232663e37c84d9d5ffdd86f44939539ef75ef3b4b2c2eef1756765b809b0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2b63d05a04cd2e867e91e287ac44eff4b97fc73a9a657273dea532d772fbcd1720df571e64b748c5e5e0b14e847b89826e0cc7b2d3d2de;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h60be98b39fa1a5ae7685e259d3c09471285b3c30a32c4fbe7676e061db0b22838fa5791c6d5e16177e5e65172bc78c9ff352efd982ead8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcd5669539a373e4bc5fa26e1e37720340ef0f7c3bdfe0037cc83aab6263983d9172089d8df54fa2b9e2b639400548a112ac690cbdbead1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h22cc2d3d2be53aa6a37c6f9181d80d85f825cda37b1edc98c17d1f729c88193e4fe5ff6be89bbe104f9b7ac70ebdc8c9ac2f63a84e1933;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10c0850089179ceabf270c570af539fc3f64414b0aa6cfc1acbd5659689d870839117de61ae20fc62b4a294d5bba0d34a44bfaa72a4823e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3f9a919b2b76286f7b8ab841bef354516f8911058bdc3f319c2cefabec70f01881c658717da60c8671d58e49d14d706ebf6a3057e94d8c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9e3dd739cfcc6889048f6628ebda408e6a8d4fd4c678c5844a129d4339658b62d80fb630b3b5569c07b8f117110e445979a073ad76f467;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h121e2f989ea6b8340c9a6c4c3ba26da2d27f1eddabc4119bacb782b2aa28cbedc242e763df9c17a709e653c9851c24808c9d645ab37544f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc5b5e770cc75d102bb108d5ad712eb6286262bf8e055cf7bbef9cf1fe29d3b1cd9da49427bdfed6e09fe36561d22326d5c5168aa39e40b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h20b4d5b2d1d71abb88aa39f1c9f258897d1f2ae41d94092ce6ae33a965d97472f7afc85ef706a1b4c8a28677559458f4d409319d1ce5ef;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h129b47eb3cb8be335d4dea389677899866ef51d8ee9b0c5f67ad2c68e7668c471b371b9d05fcde799e27e0092c0d9bb193948a77867f08d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h132c782452284a7b9c5045a65576a56ba01ae761ddd7b9f7ba3fbaef2a6050766d4e784b1e9c4a13e843e09fb00094bf5fff783ed81ad6d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h118a4fb0c4447e151594f422589aab3f56c6bbab4df4d934d667a53f812599ea8cd8bb513f0f91bfa53ad34872bec797bb4ee602d1a6f48;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19bc27ee9922c00cbe49f8a636ce39a1c1a966645d2a913cb9d2848475c22eb3430f889fac16f80272d2967e8d72b0931eec64fa16ec1c9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1414d72e7405cdbfd30b8c9979231db14abcabff5cd2326e8df013f41040fac46f23f96bd2787a415d00de09e95a6d8318c564718828e9d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d5ebae9161b37ffd31e53fdd72f463992336d65456b85b82e6e03729151c5adec79ac1a0cb0b659bf2f4e262d31942ea75350dcd1879a4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h63079c3336b61b42b6e8f02d36448d9edb809e741128507576caafa4b7356e2fea4926f25c5ee2532d8b081543265e1c2bf6c88cf98220;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d57b1ecd0ab478aa8f1af6c1a87deb660ae34a31050ddd5f80ca85ccefcd5e94274030e60eb69590ccacba279a3004309a61a75c12d631;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he8462e42cdfcb6562423d342e7d5af17e31bec57746371f3cd52913aeee7bc7da19a000b8ccbba5d403b131fc7495059d8fa77fc1f90f1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c9bca40ef4f3b4a2c7414f4e32f1a721e058b78a7fd6ab8373b4054f621dca3a50773c54e01fbf1d034f1b4b7812809cdc5fe84fb6d514;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h107cf619b76672c8439cd1e2a27e8b903ef63c2a10abb1d99ca8f4056c2dc05e69595453c4b16f930ba93a3a5f2cf61195293f0d78a1f2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h79dc7f0567ad6c4ccb3c50fe6d877b427e76055d81d2b0498fabcf48dc779d753e61549afa98334ef838308432adb3359d7d64792746d2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e49a47119f40a33c3f2a6d4b98c880ba2a9810002ba8c0340b27c1303559d9bfe0fd7708c4928dbc8d323c2b1e9f85e9bdce756a07da09;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f1cb44783a5f45365c380138bdc281b6669450e8ec6f64a2eafad6ceb90617a8a165b10568b05c909be0411a1405e8510c6204bceba417;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h161ed442aaf9f4cf14448a24f616a36531067adabe1cf65ba97b129d13e694d2a207002ccc9e105687308595e0088b4d329f2a64c9d6fcd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13c4f8d967fff47cfdcfaf96721c942cbf9a6cf39d8672fe1988cab97d1c55b921d04c6e651633a27074c68fdefadcdb189a0256c883c2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h66d95bfb7c82263f353f124a71e4f8eb1f5210051be32305d08f2a76be3cb143d2d4b0c8c76faf616460ea0a8f6602012e2a74e001d503;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h109a86294d16966fa93f042d4cd7bac0e1688c3f686437e915b3bbec88062bcd708f567cdbaa0f7ef0902caa22deb53313eea586c6d15a8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h177d25f44b2f04036b745ce4b98037f66aae607ed7267d79891f14ef0f9e482477bd703f59f0cf070ee40e0e7cc5e393dbe8929778ea2e8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h102d95c3a5bd2c23e95406dcf6189805cc40667d46faceeaac230b6df472d7fa254cf393f641dd02a6e89c39549a704a22f06ee639bd7fd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfc6b2a80dd025ee50619871bfe4a8f82c012b34115d31553e6329c4b2acd7302dbc89bbc0352b9e35c70a856fbe944792a35c47e294353;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h160922b3b6fc93e19ec48b3f78a4f6c85bf46dcb3e9298ed3bd3b92712c5faff42185718e637b0d76b14b68db0f73b6795b2b304b961fa8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h123e296dab5385d3860004ade0290f71b183c399a48e61b133fb23f51370331e5f6952687d49e43051dd171525093313685e7ca0b385525;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ad34276046816ae8f64d0b4f6fc64c29932839b7a793815217b7c27a1dcbf6179a629e84c15591757a40320328054f7bb49e2ae84931d8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8e6b3e1022de0beee1f29c1e741788606099438010952b65e2c719a68b33003818371f5ddef4afb6b06d018e64173a77d82ec59be5dd34;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d74f04219890cd72fd64621b02f3e33120c7df343893b99bfadc857b43c60dff59172a3086d6262c1b3fc58b3f2f2faf564b86fa3830f9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12478cacc98522a962e6b2dca76680773ac14699364e80fe79687856be6ca15a7ec333344c39e2ceb3c66a20a7b84c85d7708494daf18da;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7f30dc367ef9f98e43f730e9d17eb36e921d89365557fb374707f70fe47bd0d730c8838031f6516d10bae5a27c5090dc2fd8cf36159e79;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11562400ee2fc2aaf93ec09f28689bc082999b335d0ec17d6c12d9477763f2e1d663dc439d5bab6373b6abf73f138c13a27f76c8523b90c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b9548068cd30e7b58485451ff271e5633e12b6f81cb1b16d82cc69be1e952a442a4c8b63eaa0810c0f8a95e4036b3faf47b28417c1ca77;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12f7a7f72935e01fb804cd8dad55f200a542bb999a095ffe59d07b682500f22eabbd4669631f132552a913aa01b7f80b3de4019f2af22bd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h42d3d57c046727006e1d10e0fdc341acc40062806b69386832dece0a0d7fb4b7eb9ca6cb4086a27720f6e503a0f6f8256c936f92a05d49;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hebfa023065217bdb419d6152ecd66fb3d3d2f94ae7e18151619edb556dd2393323b04e7b79baa78314553004607a0c4385488def2a5ebf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h199050bc6b97f34b47bc5517725533e74443b00ecbe7c30c11ddded14b101602490a0a53f9ec1a95389d4d3f7ff522ca9d0cd0ee8b2202;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ab2be71a94e8e3ad9971068480069f3011de7bf11cbc90c58ee314ea2505a70e9823464f650a24facab120713b8561d3ddbfda954afdd5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h97c8b28afeb7733b7e92426737926d7b046fafa39a057781651ba1613faa3603366c2a6dc334755d836031d0b7ae2540b8c15b97c1afc5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13dc1741a26c0211ebbcaf597e9fde3bafa33b9f031ac4d14b3a52aa54446eed1e0dd233cbb3252def832bcba9eb2239401b55713248669;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h88257b615a5dd5b5ea405b845c91cd435bc18f862bcba14b94bcee73c79527c2132d60e946c1fffa80e6d12c427eb1535011590f943d14;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11bee0a88922d4e1665c3bdba8fe532718f47682d81e6dc92dbc40663c1a02722f824c0eefd46b9718dfeb33ca0af4cb1dc30828e5c69f7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he913537995cfddaabfca6cbce37d3a7cea350ade1548c4b5b20d0cc2dba1cafe3e7378908c49150880e89d081c90fdf3bc92e47268fb4f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d9f46350fdeaf4af5eb71a0d4e9b0c47119d328a8a7cae5f489bf5708cfaa1dd49e0411b1ce0d94edc13e77de192a910d1a4c9cfc05162;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h37ae96c514732610b339a64eda42a4da315e1a49edb669f35c9e9b2008016961bab6d6ac54b784ab104b8bcfd9fe4c10c605f1133fc0e9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b2839d3029b788ea3dedc94bec932f512853147a9e43276900943efe718cd8987a1970f3b7aa747e779f6003ad183c2fd971e283415d1a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6b0a072d2a9b271b7141d557c4433163504659e66c498100e641323e4abd1ae9e5471f2484cb11eb4d0403a1332ea2b2591a19e57cfb07;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14c6999e3d64ce19e07b950ef4ad93c22da8d8801d0184bc207bf3dc4f968bb6a1b2e3fbaaf69cea4f9ad3d435468602535bce79562017a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfa14cf5dcd0d2c9735704f6b66116108fb58adc43baac055a13304f5184b83682f1dfb6505570b9345e4ebd1f7e7112bfa73e3e42b98dc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hac6038f7a10bd5eac24e7e9701d8fcd8222516df3e8a56ae946b5ec52e5ea20a935141349a0f3397e25bf7ecd26326c7962620dffd6f34;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4dcfdf114a22137c076af758877e3cce8f46f32a5d02a81a6d680d476b78b0e51c8fbac0d3475acb7b152df6ba2401a88647a84955690e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4eb9351cced1115006e9a8304b6abef10fa682209356f294c7185c3d471f46bd9f2b7177548a8531f914d91c6cb92fd5a2d90535ef26a2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13830dfd9d69fbf9ef31a224cc704995cc70806a19baccb3fb004f9eda32c838506799a06e4be65dd21da744e4bf39aab3aa6a3b4c28deb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14f24c4df3e3cdffe0b9df3f91a640c61cbc8c54d8c307d87372bb3816a9afb9f3a81c22627a0736684ec03f0187e82b233e4147be4b3d4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1960cd13a5c49565c5f3845715d07ae70b85dd8a9b7da02b3947f218b5729057faa540d945f07f53d43a1aa9ad29ea229c95ef47720ff;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11c76b77881dd080796c898dd67315f3058aa019ef35c283cace473e641efe7223b0a7035f882a07b520308bb324e1ebe4b708db9d6ba7d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d402bb1c94044e8fb1150a1d7a07e67e55574fe654de1774f5cce33914e5ddd89969b23b7b3c1e9d04a70b03521437869f35eb6763ae57;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b4bcea6be25de90553de2af1125024126c1a227145fa429aadaead204ab4d71ddc4e37c760bb2cb08f6ab1f8662c4528b8ecb4941fc433;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h58ed76777892741fb82c5abab75a9a160d74a4c7f247b220934259a57cffca951c8f025bc71b01367828dacedffc1b07a7e9febb1a84f0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h139b71bb0858c2fe420175333c513a4bb4225b24a17e2e2c2d7c75612ea742c7c6897e7a0f415409bb44e0d5ea0858e43b6b16de51c7804;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h77a017e9bd575c976cba1376a170bded418c9ecb81a03998276728d5dcba032d86c40f86e7aa90016d1b7706419963d057f794fe290c0b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f1a3049bf432753ebe7401f8ed250f35da53af95c76e908dd8a19a957573c4f6896ae222d20f40f4b0f11a5dafc23043311b3b7cb69541;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4c916f787a81e1bdd2694fe88fc43d9013f92b4aa138b5dd3d0e80e0b74bded3da6f609f7667456929c559181b356c535bd5d46d6d5fcd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf4bcfdc033d8910e85c85998e526c4ceb633f2a0a4f3c251faa38f3656841453be0372f80d80f157b0a4a81c54135f0de8cbc80c4bbfaa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bb8501cea6d38937acb9737185ff4e476f8b4e3ac0b444f8a5aadb07f903d87c67b37388e0836202f82df6621a0a59d2375f4a834cff13;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c48e81e2718fbe433a97f4cc7b3d883b8ba24d3bb228afe21f33a95e49e7792c26ddd1694c862dc236548416dccf88a56ca4b3c5ee77f0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2f1dec6af4b554e52ab3d0fdfa908108eb861cb2433ccafb6eac7e9d8b600db7b902f50aebeaab2b9196cd0bca440804fca9b3073fde3c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11df4eaca1c4e847f416885d35b93eee7c8e42f3cff27aa8d17582c197eecd4e850001a611231e2e35e4c18969bb83a1b69ec752b0a7c61;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17a3da8e7b483c50e6d25cc90d79d5e15ac448d6ac09c4b8f17674151e01667eedee3b97bff37605466c7e117af7d156b0ce9a180011d77;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h995621bec5a714eb0cd36b5aa17c6f1fdf8a2849813c3c29864f4dc3d0d0b7ea959da5239df88b794d309c41d6c433c15f2ba041b283d9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h549fbf094339e4e76828c881d81fd4317876d1977aa7ac1fb08afa9fe925517e68f018a17a5ab3ce394b51ec82feea1a7406b9cf46aa7b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hff797c645fa5129cc62456749c5878ab974324e5e2114edb9c3b19cfcc37e14c1be8e2f2d7f4d3f5016816dc40d11cd3caeb758166ab95;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h32e46f0687f61600334a25120343831c0063c424d0182883167f60e2404504ddccc62f810b668b1691813fad9835bba3342cfcf12c0732;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc1a9aa22c76e6a82eb6a1f0f0d374a024e801093e1a20512e96b726e43a5a69f607f240eefecdb969886aa81ff84443a351a59764257cf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e31005cbd9e53dbfbbb9cd82b71e6a97ad2f4cd6492beffa8681af048306beada64fe6665b46983ee62652ace7890659e46b4b84def41d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d63201c2ad1054afef8f5a0bfba0ad43de1278f27e016839788960c643d897cca68dd57c10e7991cc6e0dcdb14a1919212f7fb8ee4eea1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h185efbea432d93c0918ac755b1cc80954c02199406425533552033cf746445d6effc602c161f66e13e71a66bf6f768ba982367c9c5ee445;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9876ab9c651a24066e6b67aa0c5529eb169ec33517adce871db1063bd4b8452dce79be54e4f28fdbae55cb361db7eb020a8d27a4cacb07;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e8121b5fda133e00dff2d3faebe7e8512ccc8a1242a56f2d5d6ea636d9e7fcafe9f199a3f5a75d7974a1f0ebed9aa550e1c82ec0b7847c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h535cf5eb6fca4d259ede4bbc1550c14a88ed1a77433feee01f94db5f68a74081e6c32732d69bdc4e1d2076ad4efef0f16f9c272a7c8925;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12ed728f8df29a7c07f0f4e177bdcd02e9a8bec4c5af73f931e1bbcd0f123b883db50f70796216dbcf66312d0fe56e455f9c5ae9f371900;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e650b72617bad64f1db0a0a2324a523591fc16f6404c36efe1ea64120a5a17f3e7c750bae1c98c6d1ce77db6bd0452945df0b7eaff6afd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1313096e5d73c68029dd3b0cd910220b83d8d458669033e800e163663f697e6b4c920419cc3982833ccc3e13e7c4e0c8d0067185cbf3ab;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha465968a896d804bbabc3a2a31d4959a3a95b238890d679673a99f36ff4fce6afa203d470ed7ffd7a61d1406fab9738f815d2cffee83ee;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb5a965ac78772f3e121d806651fad89ccb96ecdbb92720a7d8e9b5cc511e27e1945bada3aca9e836ef6ac2ad89f8f66f93b44b7ab0887d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he68e53cf8b0ae66808bec500ef1bb390115381d804318473377cb0a0eac27560e5dd4bb010ae12a9d588d92cee9b57088c9bc273834594;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h412a62e27099bf9196b2fbc94d04da75f8f31ec5deb1e5c753c33e30759071db07c6b7041c06fda76ef52c2d157385d845d2a5b2390c9b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h399843d4f4d3a1bbf1fec96211277d7765b30478f1dbe1cb92f28305004130498b0c8f94c4d4f22a31072cf89f1018122d8103ac5380ee;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd5f1a1c16f8a1e54638a05885947e35e5aa445c05006f78faa160ed1667012ebd4de1a48d9db427c4b3ebaeb2b2b211dfb4fe877e484bb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h83815b89f8b610368e65885c18f25b8828026dae57fbf35dedbac7ca7d69f8266c513f3bf91ea94ca55f358a495361c2bd44b79a4436b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h95a36807667697b2dfe1f33619a18d713bf012e71ffc36b23f7841835ae12fbdd7c7886d149c93e1b496c1a68c4a7dc74e7479a8a34353;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h70c90c98f6ce97244705e82fdf50ec08fd1ef9427e8d7737c26ca34fbc1ac1e22459292650ee1b072b126163275766134d405281357d98;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dc40954650a97d8fec7d7488aa557c9f0a91f1c1fd27ff6fb628cea4c9a32d1a6b5ea1b6967b164814b3d503153f8ddca75197d7e8121;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e20a7e5cefc90f9ebc077eda86da47708a5a10caf59ee4d7f6a66c0cbc33f1364f9b4cf0310aa5c5fbf76a8ee081d357253f9e7f7dbaf3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c9c4983fc5af814edecc04ab3d960e3996d75824cc07636b82c7b1b90c3f88f17552bfcae7bb7a267f16d3d98f4f269d29f8bc966667b5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b686034829574092a0c73e00c5503979f8a6cc8a2d1b47e352cce0158e7b34743a4729ddd7c9240c96f638feb003d97f5c123a88eeea72;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h177bdd40bd12e61e773703a94c303773732be3279c7d95d061a7da623dfb188a1dd18e48f92b8ce9112012a786ad149847baa57dae1cec8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h683b5fa35169b3f414f6188e2498925ced24c3b136cc5f245fbdb74ce99070ef825ec32643643282785c3c628b2543efa5250f39edb1b5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8c38ed1a226bfbaf874fa187a64fce450c8b7c246f2638a58071e6ccd5a064c77a4c1500a384db97b6c011ff7345ed551dba7faddaddc3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h93156e11862ad81f9492d17161b61f38cc62fab2d628f72c9c7bb1895e8ff627267b65690a98c35ba199a8d485a349a40fcb9d18404ef6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb0d7480952306bdf31f09d1d4b1d9a8507a51a15e75bcb9ce1477f868e027ba43b4af79b47e90455741c9838c249767196a50c0a0c18a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13d62a2aaaaa3cb4821deb5141f5cdcdbed4593448adff6a95f268fedb50a00688dbe9eb456dbc131e704d952b87cde5abae28f4af195a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h140db65456fb468bf1f7815a3b900add27007edb5d9f937060851d0e099d954f30f5597c66eaeaec210e10e5a981961fb81004c47bcdb2d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a31115584719e7d9fd682577ed9712700ca1a4e68c651c59bb34e49adec8657bb5b90c3493a11d4b63b9d28919ad4b00eb60dbf6fceda1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h149ef2377939ba1827a3815010a04055dcb3bbd0bba18a1ab3274949beef9e57cb080b56a510a23617f7fa9789892c1765c1b36e25c1a1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h189606ff28a69af85317ba40a711d9cd90eb0162bae37fefd55a7cd9412fb7389c885b78c2c22e236e69492a7938a04241c156c4cec1c29;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b2069deb08348ae05b13ffa4c60e1f4bef6e5f93e257793edda01f185271fb4f1dc5ff7d75cab6f66cf4964f993395008c5a45af381282;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f292d626146a06febca60add5ebc05c87392e5cdf0adeb133e9172d82ae8531bb09d4085b2c9a97c21018a69772f3f0bf132469ba07777;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e1328fbe70bd729201082b4a09fad1074c6bb41fd20afc9b116071fff6b540a53ea5aba4754470ecfcc6def2aba79909566fc032a8eba6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h94e6e29a77609aa77c5a43e00d09175e7ae85cf74b58a6b5a9dc71930ba7aa77c6b8b6d6b6b8194364c424192bffba3d537231363548ba;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7317daaec9027c37f72e3d29ffb9903250e6aa25b5692ff0baafe58f700eda569a12406362a4df8d6808babf09c2bfdd1c1d710eb95c35;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4e297e62fca5c492f9d174d009ee5d15df05f8ff2bd9b48dfded4c8baaeb0363745332223e277927536b0a5b2592b5bcff011644c77a70;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16e88449d51e6fc59701372c16fc46c63a4d1ce0a2a4c940bc2ec458b17d4552689924308cde458fb266e60475802de989c86836fc3b181;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h649784551c4975f7357bbb7004bb417dd156f748aaa06d612b346490f0a40d329e870a8446c7154ec80fa042178d2ec4d6889495e1e54;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h644edd200bea148f047f9ab4a23724f5e7d5a4d7f45f116cdc0d68434ecaeab8dfdf32ddf6b65e2673350134616ca33d6135ce39f75f11;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15537f1175698685bdf0801538f1d93a87222c714781b583bbc731ed64ed2ca06e3a5f9c5ae55ab6f9689afc0791267300324175f4d7a7e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3f362ab94b81462fe87b633303a2b26b5dbaed7a84ce39839d81e60f6d9696d0dde6619d06bc2553dd50f6ed6d9d9e82af984044b2e997;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ab2008db6d390c0a3ddde3088465ee58b4dc96f7f83edfce6ec4b796c453b0b27f79e5cb772638f810d8796a7f410c42d10ce898b45cd1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hda840ea51fad5c7920a0b36573502041d079632dad425857850ab51f0ce174d11f9648fa0a130007ee6b4cb7b009b0a9beafa7d5bb46bf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h518a6c6aac0660bd15704ae81543fea2e558871acbb02213881944db5b1257506c3dbaa51ab8158df531793c2eac25b8e763e4ef340bcf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a66f1457ba6d9f148bc7ad2b0a677382ad75e5d3b1be3b859eab0d627a6e44ddac72a9e429cfea43ad373e4fece675b576c3ae13c1afb7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16b19fef56f6b3afb8d2d865b16ad4df2ba5f201530c0b832d029be0971cae0b8a8be8b2bdad7567e861db9f0aa7c46c2150a860ed6c334;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4204c2ecd8eac31219a5c691249dd0c04e20c47877d65f32ca245e7224f3d5b366ae22fda21fda326701f3c031bf0545b96f0741ca7c46;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h40d4f3258722eb2c7321d89ace12b76dda28fdfa87918e1e922406f9e79589f0262495c85380df923c78d50d5d73446214406326241614;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he18f6500a1749f1605c57d6b1a8292e37267d01010c8a513df17c02527137002b265b1c020498eab1909c90fe6ef5fcd1de3dab9bf6f93;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1506e931d4d73e14ef97429c49cf8592ffb94e625da9c82748a4b3be0721641a41682797621c9ca551c32e81e90d0eaac000b183287b515;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h63f2b4878b152a696fedf7f53984deb42a344ca9000c1805494788323ac1d405b91bacd59cc4b371ac9fff521e2c11ebaebeb1b5218882;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12a33bb4ebe85c2a072f52a3872f7aebb459a2d22db1525a6e7318179ca04fe2ead36d5dc30922fa14bf3934163da4a8a270f227eae31cb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1967e6f6ad934da5f3fcd80f3c86921537a5c73878e97240dcb3b30fff02beb96914036bcc3e469e7b46de37f70533e06219ac17f2319b4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ff14285aca1e82bd9f391f9a556ab6a2ba58f9bb6ac8bf3b422eaa752bec4c31255d1359b0a0b0f1c7f13ab1aa1c193446fe97714a5af9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfc5c18bb20947875dd02022676444fee50ad3f2de70c3265dcdc3abad9ef8bd925d03198989d2ba3962bf63fe84e0b911f11637508047f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h156e3f782ac41f2215b107b8e515643c5fe0405c9145853838f45f8106560fe74714ae20ad61f1c3abc855f4ca8033dc28c2b8438c76ab7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8dcb57606d1c3cc11e152255204197e1fee72a81b59aee90bd10cf75324791902abc6d4975148ed2a3559628bca3c73d9c3cdb2ac9c0e6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h133598194d4c838c2f380987ec137e463456fa6be09fb33f70367fea2b938346c8590754bc15d988792a5b867f9bf77a8bc8a9c1f4c066b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11802dabd389c5e594e1c3500ba692d6b6077e0c32c55ed7906b08d7350c77b98bc1ac89e22ef9e822705819f2940405d2724e567e6da88;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e3fa64b610b9ba2102f901059dab3433e17b7dc7bac9d17008fb1e07c9c828347bef4634f49d44117920d27aa727c5e7deee991daa6e76;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h138771a506da052da1be808c6954efc9c36a62c7fc43e278e48cb5b000384d102b65c62c276c40b70b618c20d56dee9b5b6a4d23c46b137;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h125932026b3a0d2949d6916d7ff91e87524f5bd931d3d3439906abdb2af3e5756f94746b33a657a030ecdd15a5339cd7d539eb8e1ef9883;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h152cae93bbca70bafaec52754ed59ddeafe63ef03e630ba176f2e800ac1e11d2b6a8c075219a1c9adf89768eeced783e8d80448baef17dc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h142e25535a0bc6130b8b9a808740d97394409f29db1242267b103bbd6ff2eed571f53bd479031f7944fe96e0dc7f7f7f63c1f30f8cb5c92;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ec511c293f0581d82278d18b2500ca0481f217d6742f29d08157b5e2ad8a58348a83d51a46d9c81d17e23a5122ddde88bd2a66a17cc662;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a185eec20c8068fefe144b0efc933ef6147059028717bd9d3637d42baa612eeef53e768397f7899f597ff78022ba88a0e3fa56acc2bebe;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd0da2bed207d09fac06b819015da76f06c2da313cfe6a816a933b5b01ff90a32b15cd8f76d2ee1e06d202b46aa3f34f62e6a385663d628;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfed94c615d49ef960f6fa016fd7b96c94ac690028bf3a01eb8f654555377c708acc9878a1f355cd5374186c91005824f8349237363d05f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18d9f826e96174c6d1f114eb86c6399547632805a1519a4607127e0545b67f4671ef242a6d91666318e4081740d9904eae03cd9c3ed0a86;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he879e51969a00e6d9e05b42425f99ce2a0ff3c3707b805393fd08b89f252f54fa971ec1aace43203e092ff341fc0f5b760f34e294d45c3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12862901d8afcec5aebaed38c2f7a70f461d7fa36f55384905afad9ae5a1c7ea30dae9aa03808596c5c339fc82e19078445def2fc1fa5d1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12952ce36d4b1e0205c4998f93dc20609dd7fef847780686efc241c10161d603cbff143f6c2148a841a44dcd983852da65ca1ed9d85026a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3b31aa078ada63e9bcc43f7c97e0fd722d0d638f2e4800118072488849559129e44dcea9069b09719098b0ba1c52486cce8f657c7501ce;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1379d7ca3fd4d14f81f844d51b5477c745b088b7bacc237a2eeaf71ffb30416c42da8aff397744d1f64bc2782ac30fb9449cd3a5be040d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c2f4054ab2b04ca2f8036415b6a5f434fdcf0a0dfbd527590ca0f1e38f07e0dee2cadac0fc174eed13aa4279767d0a2bb703156c838bb1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h629054b78a49a9068ea118c225fb89d553ccad2ed5fa56eb3ed9df87fb651f0d6fbc600a8f250f1fa1fe3a761d4ba811773d271ef8b25d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14a4e123601d8457e12f5af42ad5eaec4c74ec637abb1b2220aad66a8a007d3a1d85f9bb1ca1fee38664ef654f15d5849275cc0db3114c4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1143f818238375eef0aa5e97a04adccbeb7efba6339404aef9dd90756f0dac1bd8a00922cbe07b69f86786c5c71608f03e7a7f9e7b0d68b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f997384b2fb7dd0c47196ebf598ece0f3a9cc62d417e142d88e6c182809896f3e042befda52d3e84d5009cf40fe013f2d63ba334411a9a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18282bde6b175a2b64ad26ae428f707067f07c1438a9b96a0e7e3e2d54e5995c5d6b43113a9e6b8a5f856cf5a3c904ee33cf8b160c19991;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb75b7f420a05ec1576045bd4ac396b57916361a3146f5c00f3ff5d3f388a603ef55b756dbe6017bf2f9e5a38ad6f9903f499a588bdc3d9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19975a6d57addbf49612513bf1c612d92eeeadcb85bb54e504aebe2115ac5d18b33f7b37ebf642ae61df2a89b8ff803281bc84bef306e9e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h984881c21acb80b3d018f4f3325153c3fa91eabc67b4f82fc6ec2a7501051ed62c9a4611a92aef370771f74fecf2afcd4fa3c92b940621;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a512e91de2cd4956b36d21dc96f923a3e78f073f44962b9dfa7006bfe37a48b6be16b76dd47faac626c42859f082e05f1da92d788a8456;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h687e5f6ad9ad639fc53bc8296d137a7be26c976c262708d3f0ea50e4a4e173707aaa4ec99d199ed346ef30d5b3bb272029cd63a7ac5bc9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12d35842b712695914fcaca47102cb8537bda539a22c864d84eb7376926122cc6d0c286174f73b6a3adfc8db991715382dd2ee136e8f714;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdf1697b70885275a96b927681cc4a12a2e34c0b7daaf165527790e70b80356a2614aa56f8db69f4ae18a25422801d2b08d89f9f31a0099;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4bbbd755187f0b8e4a807fc6cb3066982d707c586781b30be439f02c9c2ed2f82a512f7e8053942d87e10e8fa87ea702ed2f2ff0c6e2fe;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11530e06277bee58515081259ffa0bda6825cbe353b877de4193cc4abd6f47446ad93dbb8c21f3737d6277abe35a15e50b054fd0d2c6232;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19fe5117d9eab470c1f6b3f296a2eb48d3c8045f7edaa68a33a5db3f5a6eff0c7a3bb68c6b08d7061b79f8dd26b1ff9fd0d00561f4b4171;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9f9e2fc8374ebf421e6dd0e1f60bde21aad0ef0893b17c1b40a27dda7e8971ee4cc02bda24937f0e110df5f26c58413c1edecf3316cf54;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e3562b4a926e358db574abaed1e1f947508a8ae0c35f6e654013e9ba180273d8318616f90567fda16a94e289e34d7cbed65b26c3b6b53a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h179196cbab9c26423cdde606463e7cf7bb1a58cf27f56ae9f59231b071a696f593645fc69ee5e77cd1941af79057ec81c827180aabcc0cc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18e21416408e4f09d8d91920538134e9cc152fa0a98a9294f4242b9f6dcc40e09d2efed2d2dda6f656d0637fb9b2f4592a14f8119a26662;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6930105dc84548e5992a0998e86f2ce522137fafd03d10b20afbce1e26e853b9b0fb0ee837dd840dfeeada36a10bd91cf7172fab3de45a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha31773d38e9858423fddfd0740e95baeac1b69c750eecdba6f0e0e773718c5ef94609c1a42b3b6ff523b96cf707657ed5c70bce3e8fc29;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h22c12608e2c7267084a42d09acff7fa67eac983cde458a551b7ee25f180a82278f7f287da3531379b6d355df1fa5002db6ff338541a18b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1663a0285d45d68126f84d1454f50995fc98f4ab86b6b710fff048b18fa1af74c19cf05bfdb50143a7a3d0eddb8e0493a67bffb6610ff6f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf97a97f2037f2bf6cd060d0276204cf43ac9158516687a22077b2def5fdbf8134f631e7dac2fd9c17964e9292a34cef575cde8cb7fb935;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcd44e5a7154cd32792fb9ffa5e30ce9bbb639040dc95b5b2c23932b5d030b0d9e4685f0b78ab4fdf040c602621e7ace11a5a2cc3a73a13;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h886b0edb939b3306159914bfe22938165b711ec954008c4bc4084e634751d703698cd0e640eb5258e90add57cab690bd1be28c6f236ffb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6a4248869387a72e551f0bc337540eb0fe5b67e63c37eb278f972bce60ecd3fbb83a6b0a55ef0fbfb1458ce4c380970dd8f1ceaa36f419;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h70a95e87fa864565972fda38895cf0239a76525d119e3501b87e1f1eee664d03619ab8078a79bfeb12479be01579fb4308ee1f0263590a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdabba0eb13a279d88da3236f8d1aa1c56584479755d91ead1b9782900188d33d6fdf4e6d38ff864b8cd0765709fe0e036b482a3a49b154;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15f402b801ba265f1ab17cf0413d277043422180dfb9513b03313e7ffc5d5efda8d0d5b49b806ac412ea23e4767bdf98461702238a752a0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11e8e8f863cbafcf1152e93b2d078477eea782e12dd7f292acc6fdc9d4826513c99f30a44b656c8b5a0c597041599bab4badccdfb1e9a80;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ed1d89684262f8f04dfb0a8550d593777dc34d95306be4007bfe627878688e8bdfb6223d15aaeb9d0fa97d28373c852e47a1f22c2c56c1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcbf1b50226c0ec98c30ad959cbc851a12130beec7a53f30c960c7110ff996cd617782ca0442ba8f467200426a87971ca4600fab57e71ce;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ed35ccd15da08aafea38e8284a382a8bc11a78aff61421fc80e1bac224598e2360968b5f7cd7588185d07ee7f747d2c29bc0492cecd50d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19ce95332ba96fb88c54413c440830be4e52b26d3f5570ee5fe0cb334e0c725894a2ea0f3a4c48351689dbdeb954973f9a77d0d3d08d1ec;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1de2f1b5c52f7d5e249a584b78d685e9f28b7bc0e70a0cc5823b74ee098b4d4f658ac7f2e038a6fabd2f6d048693957d97503c5d754894;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ca3160d02ef5e709ff31d4dce3bb9775dab56788d5722a81cbf2c5b5842763329fca7966ab5398bca959365cefba30f1ad4a4cb0f667a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h193283d56d35703f6ddc494efdea03e25799b6b87333535b66847aec7c0292ab1e25eda118cf130b7e27869864f974ea9d293d2be64b874;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19a207e9aa4b8a7bfa72e1d116f46bfef5db82666a63c1cb60d971704891cc6a276c9778a9f0d30410436b195bb73907ea08105d325be7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb9eddc7a1ddfc680b50ec6b4c4deee927261f5275db7682455dab498033efc58f96e5eb07a07a2eb496bc5a1cf59d248140a2dfd20c964;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbee5850243da63d45d041d7f840931734595165e2f12abb5c9b9f577bee0b77b141d7851907fb91e6405a087a39436aad88dd51eee6368;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf1a05649e26a261553d2c31e7c944ad9eeaeb6e8543504c76e362b76964cd18821238c29a605a162ea32e79bc3bb40115c794ccb5b4d1c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h46c890356ee814d8ae3d6ce32400da33c15741fb956a7cbea96693df101c998ab8326f273ba2c7c6707fea54bc390f581ba8cd9e597a3a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fc19d0216c2dab0ac080d36fa05cf6b9ceda2cd672193d41568003a322ff011aefbb2a10ef42b3e147369a897277c1bee80bc6b75db585;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha1d714c856a1b883815f6ef6b004ac014d9b4c14499b694864a45897a363c3855f95e52689c3815c4e70ca91f503972fd4d19c78a99364;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16d1f710d65f15b065f958541194145b9389a0ea776fcd09ec872c1486471648174253798199acbd59fd4dc715d8a6170aefca7434f9c66;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19b6c4e1108e37fe29105fbfd35ac9d2fe2133571c73f336d35bffe6218aa63ee6c6a437fd28ef415caae72882249d34383ef3086555f00;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14976456595a13c393f6c18e203040ba09e4ee0c94bcc946ec9152c931ab9f0e8c60be9e5e4e8b242909bb175e9e2386903304d6421c089;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb34ae3b9b5f7168cb051ee12a1ab6256881be68593e58ab3f4bac60c5642915f9d6e7ba701b1b2eff761a3a4d02b78b4cea6b034074660;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bb92214a615ac0d613cb393e01741fed02faa63b5bb40e380c79ba8993634e806d958e443ebfde00df393566a6316f9f8d6376d895b52;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h57989de7ff7ad5922b1ff4c2575f794f0fa4ceb2648c5f660bcb95d8d43d900d6c3da56c11632c608876b8f736620d63713ad807abb28;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13850beccd6fc260b7c94c4c2c2a2660d40f968770e5bf940a2124c51cb5edf695dbc10c454adb9af7008ffb2efebdab36e1b94a2d3f15b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h104cd57b43ecbf12af903a6fdcaeed3dd172a4ca739f2fbcce44ce3ef5a369fd54db35f006756dd0398deccac83f47bd039dfbb835abdca;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f2adc976d3a0103c25f16276338b8ca811362c8378311d1b8801d53594b64e544121c1f4c133e609b0f0cc3a872e18b0dc795f4aa55283;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ac99857453e8296629920b0a723f6d216933cf68d9d5775d30c2c0f5bd38ea95b1bedcc00780d95e87edbfb757117548f2ad8a3e7996ac;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a733b4c5ec4c9717cbbfd4b779e368c58afeb0b9b3ad0b00d2e4101c924f109bd7f4aff6efd380f5390d387a694a8b3070a93b051e1c9c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h73218d586c0c1b595f6eeb83ea98c9ce6c4f4638a182ae57d8db0eee0d110a3ad32e91374ce5f184a2a7e89afac4cdabd2ed767a62a1de;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h85912cb713c7716e295cce4d34c40c06e8530314c3618a2b4e6e9cbd5c8a4b0e487f88b5ad3d16abe48f64cadf75dd1ae2d2fd0188c895;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eb71e08472980897686bd52929d65bf96502a90e6f91d75fbbc9c660ca2a35a399f8a3199ae6c0fa08cc232c7c4f33433800d7c9489533;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h174435d8e083454a954ee3bf76f297ce64034e40f7bc5b05442e6130bfa9efa11b85e858454b8c10292d1945b374e6992d16234e9af2de1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h164c710989461f3f8d822dee72d7668f3d0e59914bb5c6ca27343a81f071fb60391a112dd4d627f82cd60762d4f8b1d6026c4f63e8d5c65;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he7ae376d9dfd322276075f2a9153f9a596b92b0835f85ff28c0c280b6f267c9770d718edd5863004ddad8422e21b3e5d37d27f0a5484c9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8f9eddf29e39a082130e131bb25b279a488d472cae8d41613954c2d57b4714d1dbbe5e97aabb33366e061682c20b16b8f72a2d9a8ed6fd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8c3a31599e9c4d8038b805eb4b8ca97d958cf9a906e30efaae325e3c50ef68c2ea14fda6c30dc602aba644aeade50c8809f5dc9219b49f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc96e3a0481ae839355396ce57cff4b19f7c4860249a36cbadb4370ed596927193de956e0ab3574943c8c3d0c5951ac7550d0ad09707764;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8232e1a5399bf948b257e432e303630039f2d5155c59d6532e9459daa74189a542a6eb9627deff3459c2d6479a98bea2184414523e081f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h57087a38b4e1e38b87ca2912a51455c612da4386ae86b6fa94811fa05cab8539a34ae8ea1da782eed9153f2a1e65e2dc09ce01fb08024e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf827bf1127c8180893467d4019ac154ed56f36c939c0bcc71c781c0103f29ac3bc421003929436ed9c60d979f05d1225737543507880ac;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h157a92b5fe8a4cf857deba9bcfeacf24bb861adea99d1675f316a0b26fd30aa9af6483b8c5fe18705e72eff4f37fc69654fe74f554674fb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h190b89942f7a3bcb0c517add6a8d3a0dcb90b86b0930d3511e603399c1866d5d830a34ee75a0337bc516c19c4ae6a2db190ef921a1ac47b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h269eb24bbf7dc8cd0718f8c17b159fe3fcf642a4346bbf67185c08c6ad5b696ccbabfa61140f67f8db62705d3e5a724eeb61b739726281;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h90f495358eaa420e4101e74fd5049f42b530da6929ffa9fddc5b27d709d19e941f535bf9c054997c10f5955d5314e4628a3bd4a1767eb3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f8dac18dc839977dd9329a5e2b212e19d597ccc8c561d37a0f61b1eb2ce39ca904ef1bfdf0b4c4453d9075f42a88c8454edb09cc0d9250;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1de1d022fb9f1f035dccafd1b325c529538d987cbb3577cb46a9607d9f703d67f180542ffed3dfc5617130c898b28c7934ffb93fb7e214a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h742bdb84422fc140f4a0016408045c90f743e581424ad237c4a4a112e5c3e208e3fb969ab430ce62b22bda4946603d6eab7f84ec30f7c7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16cda43b97f8a19ba2d61240123778500ea9990de8370f1ce8bd9499e30a4699b9db404677b38213bebea1ec41a447d603e45109fd8c707;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d1ecb73ccddfe1417f0ab13932f0efc32f7aa0fd4a3e2a7e650a4338ca0b8febf7d13e2d68a03daf8ffc73e0922a43c1ad3907ab39afa0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2799f77713c09fc339fb19cf3757d06c8d8ae0f68da84ea9c83eb905bf4f4acb90cc94996a7249a7d84d4778a559ae4135562eeb8b65fa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1276c201ed8f4647caaa5cb1e0b4f017bd89401c26cc3d645f7769fd261186fe47d4404f14116df632266f0f873bdb06688a6f68803fee4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h157ec06cb63e491f753ea47c9cdcf169c8d74f6752d7221d4ef9cb9d7209990f9efc1cca8eff83d137a2ee8ad4f3b38e33e1185840db940;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7897356f7858cefccc25752a83b8f3429b3c0225be5f6801a646f759f8e8ab32c2634f8d85fc448c188a1e11a033fbb154364acf2d4c45;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9211047610a7a7b38e424780388c4c4456fc35c8fddf87c2b77979db0d594f25cf564ca7a6bf65cb1530a71b58abf83c3c6bcc62b2dcc1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18c62adee715ffff811090e80006a677e1f2cb09e15ef988aeafc2c62ed2f346c33037cc66b3a2506d8e9844c50aa9c7e98c0906b943649;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10dc7026fc4e48f06e96320edbc296146b8b97d274f5b8bc2b79fc308b148e175b446d2d47f73e97ae4b396045118b717f47c587442310b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dd8578646be89fbc168dd42dfbb0cbab3b96a85da1498904683ed87017a921899cdae719ca2b3e66f245af0626ef66562d70b808745ccf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h73772f8dae4de1384abaf8f38d6f99bfef9516f8d579ef97187cef337c94ba3d1a5798bc1387de0e36013c6c186e7cb9ad24705ac0d47a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he393ebde216d830ad4ed1da92006191b673ac61fe157f61295f9b84abbf694d5248ce4e71de029ba87d81e4aafe42d834a4719a30c1c2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d61ec1d0855b7873a4d5cbe7e6fa61021f809c7f3411e4344275262225a3146cf8da7b0fc6c153690661531145597ecc6ab508edc1dfd4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h508c88b32393a047b3418ddf49bc1c4eb868a6f47c685cdcbe4bdfb5903371061aaec9f13a4a942b7c92ac65b3740ca20bebac6a34036d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b8b21c28b080a87726d9ae61898ec1ba6f5711f4d889c927cf6e4aef962e3e820a0a84f8f2d015669b25a97495ff230d09ec2d6cdd135b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12d7212f6e289ce0968535d7913c6a3846dea344a3c14809eac81b067c04ec44892d5e136aec3429b621a1cf9e8198de465261794c6b4e5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ab4c06b78db6c69eee9bb14247781ed51a4eefeeb00957604346f4262bc6a535b44b282bdffed7d679fce0a156b2fa2fa216411a3684c0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e92880adbf4036b4ecba2b9628a9ee01a1d47788a48398043c1facf7ca1cb6adbbc27a0b3c9abcce33edd8c2118e4bc0c0cc2d6e88dc96;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12e0f75294bac1569a641b8fb41c1d49c042b6f878e1051db5267a6c272f68355efcf4e704b7493c21dabba6c7a576207058e56309554d5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fc26a95f7234cf47122fe5d26ce127f5e3405805b876f5d00dfd6a731e693fa9d7ddaa7d3fbb5841959f27c30fc5612829da0e33f228c4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h164e309e828e85095dfa8c8c2a5d71d4c5c398b11fcdba71ce035c99392fa81daddcccfe672c7ecbb7aeba179885f637d5db6f8c45dce77;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h75ab0e6ca0b7715393ba0ecbe1c9cac9dcc0b1cded4d9e50de9c1f1895988f241cf585b3abb9a6dae8cf292d443c11e3f1d8b868c33c19;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e91a92235409242e92b0ede53377b95be841b90e562ece413f996fef3095d338de1fda265941dc5bb0388501961635e1675481adb90fcb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1300b4d56e30f2660fb0647d7d0589d8e96e7a5cb4abe5851c963ea066fdd6095ec120c02f64601baf9123e6fe2d6d4aaf4860ad3be114e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h61201b6efa3e9ea2ee19dfe801c3648d09748796aa9d4767597c999477b502a4746f5bfe794389b5e20dedcc9b083ea5b5620d91bef3cc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h131484dcae1ee119c4f87476d1748ef3fdf2b00b71be813bc534becbcab82c72571b01d2b9296b9fc70dab4e6214375d1d2523961010925;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f9fc61624ec388386f3b2d15a4fd9fa86aa388c3470626c2be7fae1b1b357d2be3943bffc979db7cae7375692dd24126fa06a9a545fffe;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h138ccb35e01b39503a75daf0fcd3df5084e98c2c167ce1f090711eefc773c0ed5527441504d0bfdc6fd188708e1640ea8a84995a5f7751c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1202272c6ca653f0ce9c25b667bda19758cd831c198b76caadae7000fbb95576ff738cbe16c736ceeb439b70d501cf20e98ec78bef4a815;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h132d0d070ed4953d5a1befd784f480ebcad3cb0d3a09c1aca461289f079d0875ddc60b72b3dccd2d84b219592f5e728fec720cd70fd4cc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e82e08f2ff55b9484ae64cd7a07ad9269c23371a07285db2895a264b88d44d62bd5ef5a54eece8fb5efed6590fa0f8244abfae2296d2e2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16c2fe5cadf1802097859efd6d2545d2a8731a42580eef8315cdaf419bc26050073879d05d4fd9283e93e73f0c6109074780ec080059d76;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18e7a03125f44c2f58baf36abf53a6c5ef7a6b5a5b81a22b23eeafa77994be33f99bedd29e678fb77d2713c80e23cd7e8adcf01b3ec482b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha837eedfa545b90ae3a5b050cac285eb6ea0395b6084cf96e6caf9d49bf52efdb381e242ba82550a884bb23ac7d262881e28471245d9f8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he6ad92c5c53af468c4e57a6b71a0132e28206b4eb95ef8dcb2859b62f81048580e0f247fadc1462721d6ec8808c38887f0169e65de48d9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h123e34208073d821699dc6b7a63bdacb8a17d55908835f6a0e8f6213a67657587c1d22ba176f8b382b9cfc3f4a92f28338f4bbabf37a481;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16254890b3ae241b183f836c7c2320ec41f263fa017341f7a2bce1c5300d46eaca1d1c3ed89654115dc6db28780fb2f2d423aed49f29ef3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18b07649e1ff2ae8783e1fa91787eb3921443376d18f0ac2c16c211c9d3ff41d46186b75d2c9d6065b145e20bfb6ba048246485e1509a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c639ed1ba27a01209a6327d90c1b78dcfd00ab3b12629b9fb0af25af8fdeafef4f119fc3329824bc8a7e066d585fa51874e488df0f9d2d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h999f0dea7885aa1f4571f45181aa2e2a037fa573d02eccc7f240187dc0a6b4961cf9cd7ba7086fbf83ad847ae6cfe4bb7175f907969b44;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h177d4a21ad6fc7aa9c447f40aca6bd6fe87ef48729c1551aab14b7d58b726b8b36a5286b5b67b8a7b65c2805bda22b965892a0562bbee88;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13ba95c67f5e8b1d902429c864f024d29e645da7df12c10f517ac18f40ee78fa5dc3f1fa2462fb62eab41f37a5cdfba4b87a53a483e22df;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ccd110562248413fa0baa693ad7294c5fbb5e1e45f14443d8f38b70cf9d551f15b048f3382b68ea83b8d792386bec3f7fd3d500fd5b041;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2c365ab749001d85cc5ed605d52aeda5e09fb1677570a9dbfdc4b3b17ff9e531d8313a5978d3fa893624b84c6d47ab8114ff51240e49b6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3697fdbae7104bad26d21f988b344bda52055c13544ab069c154a552afd5896b513ab2d035d9ae5976cd8872d365a0f71c6d2f3b57acf2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h675cdba200009bdd75040b92dfb8c40abf2e5b43e40a209f9c3c5c85ff4cdc72f5ec5c117defe76da42ea7827580954569bbcf91267a72;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h532b02b169f90b66f5200d92b3a4f4b2568924111723acc3388cc0da742b269fbe7e7c8b03c642f3e906fac6128a6ef55067b5167d7f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4eca4847bb3a82d8a83a5e4f20e82a9781c68437b299f6509e68c38fca4ef84ce10e846dfa492dd6f24b418bf798e4336f5e8943d2113e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h140cc7bcc8ae3a6bb257e31440d7c2aa53a442ddf416f13b804411bec98f15c2b45b67addf3e692bb4b85bf5264d5dbcfc703d71a2a4077;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4671d47efdd0df3a0b1c985ec5ff297ecfbf7ed8b809047f76fec2a11cf7a1146fcc301922c8d179b054adbcad2d85d1f54017d5794811;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15593899676539fae9e46fcf1b9aa27a41583f5d470696570dbb2acf03be4bdda8d93b3ec7969a4b7cace2e9cd70782a17c3a11bcbbf04a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11703442d59c76f388c6701e8136116fe75db79b47306ceaffae8c37173ede685500e5d6c01adda7c3b6e63501a77a3afe3def9c8ad931b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11412a46e9426c932a0753ced15a7fdf6136789f3def7411efeb820ae243cf22962d36073b2edd0ebc0211217c50cef6b77e87062eb063b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1422a9f85c9f2df89979b5ab6c2bef75e0dc49374fca87c93eefcb67ad46d928154c88974971db22e9026edf58b5613b9f990ad8ff8e058;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5f407b3479b2e765563a2a40b1fa88cdfef3b1465baac60aae277252e2ee7b799255cb35d6af84242dd811354a68c42e669a73ecc01a9e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcb4f940d1418c5cf016ad5b3c603c5acae4a2c91e69ad2dae1a47352bd1f1cd375b45df3cc41303d20802933dbee7461889f5a42e102b0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h84f495d5f90367261dfdc57ef403c7cb901b98ba9e5b889b2fbecb132e1e4a0c70a0128ca4b691a4532265f0f4bd1b4f671f91c0bd794f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha3c0b4f5599bb87c3392a9b03cbd5732ba629001b88e0a06aadb5b8d478212217c52d46d3bc71cdaf11a2f76d755f46da55f7e81ccbd4f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d55b78b01d44bde425d5c84ed04add1fe9c0a789147f4d6286ff12adcf5cb3ea03775c4f1e290ac8e353f4d82b5f78a93750de9ffd2358;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1919dd32d09ed8b271d708d689fddcdc338901fa684cdd56af916ff302da3d855b28eda66608d544d9c82f57fe53253926c1e8c1ecf83e3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1607952548089147e8ccfab5a8a0bd1861c22ce76a3933ab78477c329297c4b532e69ca47dd30061e67b8105103d857e7bae707eb100483;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14b5b5569a60f6be3ee3e7812d9e9098889b7ab927678f5a1782f4e93a65d3c54bc974146ded587f3658d34d20bd4f50488bd1332d5eb04;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bc8acb56fe072ce2373308666f91ec9a5b2b5a7bb03e42d7987bfb123717a4561e8c37982614f505ebb456dff380a979ddc0b8fd35eaf6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e09ffd5cefadc01591915e9b820ffc94dee6611e6db0bd3986ebc425792e59175b5fc424e38063c18230a3169fed4519675a93f9cd9f40;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha6849b55e2a933c28d25119f9b5a4526ef2d26d71591bb629b40423e38d35029d808758e5ff9b95748a586ebaa01607704329580fe04df;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e70b636cc0113bbb59df3d21d029e56dede2e1f767479c953194f13d415396185326409f42d15e53f06860843a32b217bb6eeb62395374;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h71a642348bc2ee9dc759ed2a1393767ae56476e9ea6d4f592da2d98de155484b1e4379b061a67c471e898aa11281443704336f8a10dcf3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he89140d92a9325654e03d28ec77715d4d827c2e4c380ba7ef36d6fd8711ae5abe871d5ef8ceeb4a77cbbfc394bf7e9145affe364a0440d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18cb59a4155899cfdb6a4eb26d04c0bb928a481654513e3cc68ec6980cf09824078e567c4160aa300f1da4ff451f7b62fbe914ec223bce5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b8b16ab23008dd4ed60770ce8303829ae541703223cdf4852b4ce5682a8d300faab15d3592342e3b274a3fe94a3cd20097688f431c4d79;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d07734d8849a42bbe68fa3aa58e772079f6ac5ec90561ed83e428a2b52df1e2a7721cb26d4410c75977e2d7e13ed98c160ae32d490d944;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a8983a47b9011386c56cfab256e1fe00e2e5b5743ea7824ccbfe1b0c8c068b68a188328cad94b154349458ddc836074e630d72b917859b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17778ff867eb45e55fb1e3119e458b594381bdd614ea8bc5cac5521b5d5831588687a1ba2e9bba42219d0df2909763a3e28df92967c3bfa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1709b08c8c59b9e64885001d3e4e3a67fddb31c7be6651cc03b30dfd83111729f4351eada2d7cfda48b139b831942b415a623da126f03c0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1714e7062d1fb7ed809b4ba1f83427d1ddce17f40ee6f76d03c3254d79ba692ddd3cc6424513a3e8b92cbd1a6e57d4a102f4ba345d74c26;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7eaa8662836637537f55aac99c3c238383ce3eda9d46597ea4a551b691520719bff70452aa47d536c07289d1ad594a6d507cbd3529837f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he3bb1e84a84653044f16b92ffd6505b000e178fc2b69fe91e91103548a3432a265d9a65d800daa4b9cc0529bf395ecb67b760e3b356355;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e78a383118ce6e990cde0bee05a0b9e25fd9d7b6432cadd418e1d47ae6c2886045e3bdadcde6347060b3685399206ef0b7bcdbd8a8725c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd9fbaa2df6c076de92c26e7374a52536439e9e61dfe284e3256640132c54366e708d41ea88eb259ae88d118baf1eccf0aa986b33609569;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f8e35857d7fb1d844cf3ad2a77d8eb44a2aee094acbf3c83dca2c096dbc843b6349a89035b997eb80b357dd2138b76f9de3b06126e1bd9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h71ecbc198d35f644b583eeec0a487c6287665b7f93dae85d0f55b2e362168e8f0910f32b08af52dde7c1122d92c170b2e131526dce7c76;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h156386ed2e1372106657873f621aabb95c7e764cf7c95deeeae783429a030bee2515db97dad947561f4a9b4260de28352ce3467ff964af9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f10d76789ac0b568d2c4faed0e46b9f6f0421d1f88507fea06f5d2aef23e1eb11ef20e8b731b28c7f26c9acf1412685d3f2f71915179b6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11983bde2637f833aff2bb2660ffdedeae4686a081334afa58a1c5f5bcfe9816ab2dca15ca685e2d5c499678adf8e1ec74ff387495415f6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc1380c7a137721313f843fd1131824edb5c049657af9403cfe6cb021c9a06c3772f81689a83465364cc81facf39cbe5ef0ca02bf68475c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6b37b0e0bc5e3599e9989201c0f04b986f0ec4f59b609af50019b1f15b2e38130def7c5651b09d21e34796e376711c11dc2bc6932274a2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfb1e86c647f2ca4d694c4418b22e5d7fe72173c2bf9346276b593bbe45bcf127ee21420f9aac84530f6e2b8968923c281f9f4c80e7ea96;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h39949bc689d67238b9e7ec6ab0567140ac91024cfcb47a48522037d8766f7fa40670e6c1763116490f6377a6bf601895e3d094a32bcdce;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19f86f9cf4bb6eb8750edd3313263d09a4137a639169b20d42f8b1f8be69db8dccf93c9fc35a825469d09ab9f33214a781767e0419bd737;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb35f770177a6f70ae6c65f32139f9815e7b4659bdf471153325c078b288981006e8c8060a7268c4a09bacadc32f9d206b5810a7362cca9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h164652dc89c670c242d5d0d82b206b83f4c86d7663f165295034936c3fd9d09cce38acdbaa856cfc8de9d640ffa8f4db10afc1e75b27f77;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h94f6ab8e56c1582b455de7ed653e1976e48985c3e4ab73a16b0559f25a9830311ead461e4ef18f08a5cc2a21011dec6c3f2ea37a15bb35;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3ba856a29fd3fd5a0b450d19a323f4504227938374ad7c1b34285f54d8252989ba93c66c88c4c741edb675f7034a3087a76fadd865833d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h169c76c955c79f9e92da9fb20b8c38cf5b3e70d92e191f890c676cd49578a01dde8b6a179763496825b7920df652841acab2b6b8dad3df4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c81a2dbc76da39d1e6ebc6790264cbdeaf04f116b2a94cb760da8e846caa416a6f16b5f455d3bbe5c072ae3143ff1392b680bfc749e0b9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ab05420412af9841a46fb2cd571ed2b9f17cd5e117262b99f5cbe440a4d11711cd44997c7cff2840bc5b41a9e28deee71306f52874216b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbc27199aaac117584ff52c284c9d3e71dafd3720766a85b06cbb8621e9a776d81c44f13bda89bddd6304a4e83c2b08a0a5a6f5ada3ba4a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h830d82015945fb7f8213e97aceea15bdf3b37d136e3cf43cd4db4223099fae9093be06341f58a159116b433503dd7431b24252cf3d2dad;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h98e095dad85efb244eea48523edb8b2b317f29fab7cbdb154915e19c2eea57a3c7209f8a8dc9894b409661a43cb8676bef227c93a1c2b1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fbc8cc24db75a7d9423db26c8ab34a5bd9c0471132ea6b0ff39d36e53e7805360aadadd335650e25da13bc784497281506a93e3ed39134;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd5d87ce7ad0d7f145fcd1d16f156a39be1b955342e4837c110f7f93e4d24be65717df89927855b9fb874e72fa03be7d87c19fabebea0d4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb4c572be86dbae1a6f06ac3545f1fa4ec55225efd638a516ae3306adba9741fda44ac5fb3e69e98fc8f0bf9e4ddee7b63aa1c39c0f308;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1137a2147bae4e151969bba2eca264f14a24ebbb115b8569b80ce5a1f0b1f688e9949f532315b5003a8cc90a2cce1165d29935641d08c4c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f103cae9194883d0a8dae03e76f3730a0fe6d4f17618c1c654e080cf20518c3e846657b6616adf394e818cc6bdc33e90177456c45b5142;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h91385f36a5eead4f72b21dd4e410835f8c5013e1ae5cac86eeecc9e96596fd56300d33c054f14b606d4d773e026a44883be459573f06cf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h38ea5820ddc9e7b379adc7de7f63f7da002ccf53894528e2bced260ea8d346eb748d58820ec398da281ab19c0deb93a0e25286f54bb572;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9339f9fffd792904a87b66026e6d1a57777ce261e0b22ab74fde600bebee72c2e83c0448a885b588ed5866ddac793ad4d2710ffd74615a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h139177d7a8bf5b4ae66060921e7ac98a636445b0b5f60ee22ee6791f57810247ce0426f6b5e25bd2ea1b4ad773c781a0b5c58cd9fb2fc8f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bd4bf61cf73c4eb53534373edcd2e9367f1452c8393ac2b5648f5149abf59d588e654f88269b30780c71cbd6b4bddb15c46ca1b8509859;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heaa5f07e072138b61fe13f8cbff8d49102d1f5daea87c5d4e00798b112c504b17ef9ad8252efde2e4f1238836a27a89e3c7821da73187e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he8a41c1d26eecfa57dbcb4af8575b369a4d7e9d2dd69a7e8ccb60ca66cf0898a1a1c5a98d78ab0f52e6229313144d417f49aabc2fa8ce;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1adbfab2225282c88ad88cf19b7df39084b7df6d71a0993e297975145ce455c14b09f394203f6978caef99fe283bbd6a0cc2eda4b7443d2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1872e0ec52e709950ddd744e7388a2b33b84f3dd464872c9a67cd2e883c249e4b8b4039e0c458622347ce1dbfa217dbe0efd848a2dc9fba;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b8d13ca29e5e08eeb220db70c642c4c9b8ba791c18127ccdf684396921834078da5735e43932819ff208447a11d11e336bc2ffe8612325;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcc28305a7513e0b7c90a6e9b5ffac84dbbed25022bd1a6b349b9f4cf3a4e52728e457be8d54e23e5ed61b991c73ab6a520750046241463;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8c4326f212ab1ac2b287ec445a690a52bb0d4660d1f22e85d5767d93cbd3a9d26e03deba500fd90de707d7ec8f6d16caab18ddd486750c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hed60751689ed272fb7a4cd594113c38bd084e585d050e4572a42d100b6990babad78274daa246f1b044b3c97b056ad43039dff98f9cb17;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e3f7767d01f6d82dad7dc81fe0e9c7caace60c756af5c91f8c20b1863d2c2ac438007c8bc511c57b15c431094b70800fda42c721690ce4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h173b1f3c452f877b19534750a272e19b3f957b84f7d8de9d22fd6bf21bd5e176b57792edd50b5786ab39fc2017ff295def4ae81027f3481;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1061370528382fa53cf17a1c37417f3b3e2426e9e31026940ea39768696cc96d4acecedc41266c978e3e516bcdacd299de37fda477c0cf4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1908c1d9c2eb7d0b917547a7b7799fae5b1e54770274e571938526d4f68eed9683f595d745aecfae04b9b94e40e406090479853a98f278b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h66749c448c4228971d81e8c9ac069fc408d2893912a34933872e4ad4c87c289d6a21f7a22554a580cbb5e96a299b612a5292af6bc3c91e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e7c699479804465ab36b8a52c538a451179df985c6f5f1405209be12219f30f513cc018c38cb6fcacf785d961f8546edd59a3945da85fe;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5c62a761d84aa380c1093dd3c949787cb19f25bdf21d5bceb17db3e18f4a584037dee553e34ddde31fcee69b9d91cfe838eb9a1aed4c1c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h133d2ff137e02aad8fde396e57b77df798e6607908d9d8df37c29661a2e731481cc3931ced65a0fb2c40dd7ceeb74615e90efa48327b917;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1134985c19906808d0704b21d66d09b0217d9318151920cd7a7ae6980ac00be8438e535efeb3e0a8f3eb55d58bfca99b0f253e39e6d7ec7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h64912cf7fe17d71cbb13aac6a8eb01b791584744fa8e100d9dd597416b9af57ca45125bd3e4a41d67a46f3c6ca47ef037f580feda1e48c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a46e9a71db0c05b81d894f26e8a1cb8b4b09da1f59226c5d586657234975e55a4eca49945417189426f6dec55abde2d85cc99da4535fcb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd31455339f8ad6e5e57646a646a00c69731a0acdf04870f024a40764e4ddcc6aa42f8d52564b6c39846884acd0812605486d2c05eea3ff;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17264ed0659692baa6c6dbe45f7bfbb3b5ee66e8d385afa006e2c9ca68d25eabcef8a45526abdeba13ca8fb0618bdd69ee3d884ce1bcb66;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6bd199ee0a57d57cfcc7fbeee7fe5e728091645a25777e0ee949f039f3036fb7496df6ebdd71392bdf39d4eeec5f223f67da248842134f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19cbc82be14bb120a8a7690370de8916ba20039881fae1210e7d1aa153b5594330742041cd7cdcd2413ae76de79e34ca88bec436d9e5b1d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h314b4409b9a356feefc748325b06f8bfe3cef7587ae48495e854770740bccbac4116414233339ac5d791d4312be4531d1a11abbf46cc99;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h133c95e352a56ac3564b8bf8852ecc10514504a3c0a6a951688e37541abe065748c2b09c5056962fa5fdc9f217e251a231a1a644ff1d783;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4efe185d9cac573c1b289419ae4f67ff279c8b41502fc10620ed71dd2c2e9a315194e091335a12bcecbf11d73a49f592894595e4f8631c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb6043fd02ec24d52e8ea210b1fa9bc808d321607343102b8e552f2afa696e1c70ed375263a0889a7f81cae6d60aa0fe7b9b7ed69e0e8b7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13b2756f9efdbf5df5e55a24831181ce05fa93fd598bb3fec263980c40dbb212034b291da2e9110af98b442f0e7d17c6fdbdfe39c7a1a9a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eafaf69556bc3ffe08497da083351eb98c6ec37181578e1f20468bef08b0b172ac6eae8eea6bab0c4bd00617ed768b821067b979286c74;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha211f5b342ea62005d00e34274e5ccf8690fe921e747d4c77519fd0a465272597fa6bc5e37cf84bcf4791c9c9078dc010f82caff5ef8b4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ed853ded0282a39bdabeae05e339ddc54012e8da54e0a9a1c6a45b0c3e782a2e9dd129c19c56f15992c716c68c69095954d4ff6547b288;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha2398c514070c00db3773175d5448e896b87e16b5e00162668d6f9aef54fa4f8d4a08b3a29f83c66c5031ca6b74aa8dcc421b7f71f2b21;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf179a2a307eea18e1ed183af273c2fb3e83c66bf97ae0ce84ea0355e4a392a23fcc103038b28df65fa654d40578c9cdcb6b44d9a29cab1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e764cb3cfee39955ad26b68bcfce8fff2c158baab778b050e1519f158bcd17f43b1b3306215b8db2de09ddc1561ec6a6dea2da000f29fe;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1aa9854403c8ec48a5c0507d2d76ad460eebcfc85a14b2306feac3387d68963d6c19e89727a372a77cffe854a82b82f7624d54c2c20ed23;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h432b48704fa99a382d441341d4e1752fcdc4f12c6db7bfa3979e0058c4bbfdff172557be73b6b514600ba39a8423e696c49c7c1b8df69e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h211a5dcdeaddd65379392c124367d48212e852e4373c7a921f6cf94172f40708430145064313c6f5145075980c43e5b19809a3da4397f7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15dfdb7aed1d778acb9ed89b57ea76c6fd8f347021b028b9c91ed21780c17f86de7f44af349dc2268add7f1c23425cc5ff1d665c8b31e6b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1762d847673b6c5e2270bc14ca7f839c2d362ecfbd64e28d9a81952047cd5e208044d79669aa08257f948a220b231156104acd3447d7725;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1659582333c04554d6aeede3aad40346d401353e4dc24f6c119f0d9f75f401d26d75934a52ecd1d2a95e30b227c5d4ba85f2744e133f1c8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdea548811d0a58ff651d5e05aee223f558e75cd72f6179476a9c8ad5597d17c4ca4f23f8b756a0e8869c1b99b53c4d44a7b205d251f2fd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11cf39efcbea5effa493cddbaaf758ad4bce97c4addee1c4fda298747bd03d2c4e240b0048baf253f9f806a336ac32f7e26ab5b6ab2b8d7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hea5cb956c279770b858226c6715aeb8b9fef1af845951a767758cf74233a42594c33c42c81c2928296ff34b03a1e704f0090f41a6a55a8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1937f2cac6d5f3d6db5c6b50a86db9c712f4475a60f300648a99f5d9543f5d6a79c049ffa3c3dc9f2327b0bb8057e56eb6811810730466d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f714d476239089654c105d2e1b96d27b53197e04d135635015e30f39887724634cfba6045825e5f192277bcef275aa2f640e1995d3a94;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1af42d52b548939fe3e53627970bebeadb9393227e2b3dda78e4f9eb6d052174e690c7b96dba3334c299103bc4eecdc84845ca049644e89;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5a0c6ed2e9470846e35109da6e74e4f37f26d3339226859ec6d1d092ed6748b57cb484f965672d9a6b4a505e6ade1f90945c5cf619371f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13924cd9406fecbb48de9f406cfb56a82b1d93a3ca2a7917fa41b237b6c6a3598cddbdbb962b8cac5aee79eb25cce03f3c1fe48383c2087;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c1926b934eb4aa64b707a35783eb2e0d148d0f44311f5a8709baddd4a8d13bb96b1b54054fd8d443608d8b664f1ede6780bb1e692787a4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cb330b845c54efb25a346e86a61b238190d0e2fcc7d5e9732f0faa4c0a8f6114a8bad673c0696b4e8be338246280fd6d890cd8e3f0d506;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bc7da7a306a8d027fb62acb24ffda888fafabd758cecccd61a1d7620f1a68bcca80b4118b53cab5413e8fbfc8b3d6114b4c386d5de0c2e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16a29944692a4176996a663d6a8562a526c617a6a0cf85e35906e5dcdc5620e32637368ed1bb3b74ac1f8358bcc7a8273601d7a67d15292;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d295d4365d20159cf4c03cae7b7bbe53f6fc9594333a3ff20abdbcf725e0684ba60ebd1c8749c2914c2ec683ae2fca3ec6a7e064f241cc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1aec629709f696859f28fb9db5364f00e80674b22d90c94ab3f4f8e053da4e0eb8e10a2010d392fed949f74e51b7abce022fe4e2be47279;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h793d1ffbce174f0d6459271bb4e2a16fc7ec974834b1403fe07d603690c153b1e09edd89e2482abb35f7623cd6674f1f871f4c3904524;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e154fab59802d5733accbb9c74c5be9f7b429e2010ed416d26486017f3a9e663b6001083d700a0fd4ba0d9244cdb443edc3f0cb93f0c37;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2980ea733a4dc386c2f4e705191ae8eba5be28f90bb302e2bc85d9149960ea01260f0bdf4d4e7af7348fcdf06e994b29c93782d960d3a1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c1ec9f944980c69eb4d516f896fc9e12523c4774ae652767af46ef8c1fc3a4941df1812809045e6702f4d3255a20330c754bc71a6285aa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h42735783e028f6c93d48d3056b84f388cec1252f86bf6167a87977aa2ea52104d8f5eada02ae1f7da0c1dd56bc5e062783fe0e74f35759;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c0ca35fd894298e12e4372787575467461913f0a73377e4906c3df9dd3b2855af1bf240aaa3c66a34aa0d7c117e8aa592d55c4c3202dbd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1db446caf62fbb9970a7f1e009b0f3f150a648856f4e20aba61e930086186cac80fe09e5f7261b67caf16742236ec55f19c3993f188b5bf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h95203dea43732e781ad974d5a3092c7379c722525ada20e4360e1beff1e1b4dc04bde0568f5667bd070f0528504394a1232d41fb014d92;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17bbf404bb86db12e0220886e5e6ac03cdcb0ee3098d694c097e8f0eb8d5415a5fae19b5077ed6b78c3535bfa63075e17040271b4bba6d9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19be887c8e536866def87c0da6266d5fdb75020cb36428a2854c972cede505721f374ac0806c549752a3ce6b282a37c58aa5bcdfc84540c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h969f27fd9a3e12176c06d143d11783f1ddf8718d3a15e104bc02ac47da76e29c8d6ed5f74bfc88c39549dde91ef0290a0df9f77f6d08ef;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ac95ca0464e607bdc955b5667b777588d26f286effd87d7ee847df7568bc3f1297d02bbd9c13886c765a440d65b931ee3967b359ed669d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ea99348514efb91bbd1aa35eae10ade1a1c4a08815aab38e6683f4eb06829162e7a68c86f1f8df71c400da5c2c631836f675abcbd5fc36;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9a25c61914b03fe587d99d21d2fbd19608443edee04eec5d71ae175212c77990934a2af8b3402e972c300c52e9b2b5fdca19e407b1b614;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdfba3cb62ebb7f56ede1d44ff50a0ca85ff49464cf780e2e20b5425a20087c36f09fa0800fee7cfdd32d3d897ca842b41049cab2d1a8b6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h191e2a13f2dbb4a40429291bd3f876db6f447d490cba7d466bd634918c569c842a068acc5f451e2b75dbf360228cf477a5c1c0f6c71c9c5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c6f53ff84c02e3935b3b58c7168498caf50517891f93cb8b2ad2c643bdf9345c0edc38cd080fcb6bf0a02ed4e79efde1e988fa6727aa04;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3d65ccb49075794e9bb52b20d50d2b4792ffad9f744f9e09ddb4dc2384d9be8a7a7477f7726a485723bbb44eedb29ff4adb4c1b0d25723;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d166a61c479aa6bc7077feef05b9db97f55806b50bd98a1162d13375c44bc40df3573c2d997a3590386f5db306d54df2dd057892209a83;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12585f700915e61d76c9eba76b5470627ef71fbe8a6f5b7bc1d1537f3e972f8fcb3878480707c1ba5e0b09143ab704938395a4e277d80ff;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2b02d6f3f31dab976bd4dee67a45b8c03475f87c8e99224e18747ec2447f64066937ccdbd4aa1459035edf57cc4802a05920657d0db9c6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h77ba25f7f084376e60d22a4b7922385390b8d718c4887f85255c4ce96997cd1fad3ff6671460d2a80f17854e72a9cacd30691c55d2004;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h141868827b4325011362bba1d559fd17dee74d17a76ae3fbf035d8ab0b894dc2d1f2f25df2733a00c9b3aef09a81a59b1c83c1210e88f12;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'had8d629eb7450d1a422afdcafa9f49d9ab06fa27f10f1b86b836403302575d924920dfebb7de105d243f938e84007cdc372277f873958d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bb16942032e00d00577767d2071767efc987ea4ded5ccea2cfb3d9100a8a1e3b712c7402ea6ec45afc8d6a21b3cf31b5e858f774fcb128;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h191b68ec2e1f9cb7655f7c3163e80e2f1b617ac5d0a8c0782a30746740922d7e4900ac227d2d53f0acbb280ca26073969dd2cf2be45e0a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9f4e4f9b945e218a4e0fd90c7a444173464dd7d099a8234665642bd205d0c3d1634e9890acdba9512e5b9c22a0575f3bfdc91bb9023431;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h196e31f416969a95afe4bc7e9678117bb70345945e1e4a7614eafca4bbf74b51f5ea3745b1c07632d782f94a2b09a548a80b159edba11ee;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ee1121e3a462b6b7517804db6c6027a793ace872db8fd84e9376fc292d487aa50fd6c7d004ef68662b534fd7ae8d3ce4fe9bacf6dd40d0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfbd5ce1ee3bbe3393acdadbe6fdf73ebab1b162bbe6d3b284241588c4674f76acafa77d5453e08e8dee8565d2e86c7ddc95afb151a7dc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf2c6248e441c538fe9fb466bf6a41c1650af1b2464c14739ae3c91f4309524896ebdd72d4052ffdcee859adab56395a558956229b5790a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1041e6d75814ede36987019daf24c48111844bd71234ec45b59c19d1050d3f284fac0bf10804b70ad2db477d2bf3d08ad599348a1b552ad;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e0ab19e8be2190b636cd936941659758adec09bc32bb9b0ab8c268b6644684db99da2880dfbaa75d492d1b41592528630e6fc52810ec1d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14c5894ce5f64663b40fb0f546675f5eecba94155d34864bd7c3dbcb0becdd1fb2bfae7d6d8f272eaa57004453855d503b73574881c5781;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16d2e682b132cbfe050443878684061bcd26f655ad233dca4ff5a1a716aac3c731f8e5ea7304b2e4efa37f2fcbedc43467d4fdaa4a515d1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1331949d9bcefdb4b5d13f19f26fa00ca64083195293a010eadb65128666124323e5c52b62b2dbc9aa4223bfb01ea8c72de8c480f9fa9a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h167b5cfcd4913a866935b2364b5420d589ee6f45ea2f8147f4f6ba2350147706a20d0654cca159a64478a91276f0d877d6a931b93ffca5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4482b43e83fa95c640a8ce9886e37a0828cf5ae9b9dc6223cbcc6f032cae9b32e80ef77c9c4c8f64bffd2551e9270b9ff51f7a36c6b6de;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h458f9acba79278d58919e16e3b47d69b5ca69dd5b7043fc6cbfcf4169db66b080c32494a7aff45064336523a1b564a815dff61558778c8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12c9816f57574b222d91121f77f14b7bde6397b6d4f321c5b52e3e97613a0859c9cdfdb48bcc3956c12c4ece5110d29ed51a9f0f97b5e5b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11f8fdb09bb8a0234ea0048da330b389c306d20d27d397bc28cfb45c009ef2b91302b0adf12c19f6523282c1e9dd099ce43c7ce28ca82bc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h71b9253b152df0ac3f134ba9aea603a25d0db672e2cbf29edb1a5316800634b42872df0076a6c4b840b8fb3a13a8c45a28e533b54a0d60;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h524d02e0900d801e4c8902c8fe7d1a8535592dd51f1542f6f1a42e1c27866e434df97f766ed40d8fe0dc9bb925607bee24efd0c530a2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h350f02a2fa57ae148c87954f7efac60f186b71b88c28291917554449ba125fba2017e4184bcc1e8847173175f9f4b6eaebd5384a7d63b3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14bd2d2a80f22de6fe0c81cb8488924d06035f192168a089d3b3f1b214e33986b5e767df2eea00590298bf7b0b84dd4c397fcff3828f9a0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h114737d89354263e9495f2860cf1cb82bf56bed566ec6ea52c717ee91fe2b18d05a504098750a90e41445d3c3a5d7abda9c2f7f87b80602;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1af6914a36e847cbb2cbf76f9dcf1b2e10d1ff3b8370ff30de0396a3469a87fa6b44a0341bb956a5ca8d993913f331de4ea3a04c3667c9c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f7296cee5d82539e7ca6049430cb73def864d391f29884222de4ee1230a765ba9259fa8e1356f808d115537c40991f3801f8b6d5ecdb1c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13529d0409fa3b874073f1606dc3a3dcc5ae3f44a37a02c633965cc9b544b45be7d2703832a07e78ba3a4124e4506eaed1fcc3d6edfc6b8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h22b4b2cfde9c4f3d25bd5035542152d8d11fb848ab82ffe0bac7c8c7077062c212e12ca3ac4af03b10204eb9555a060e55bcd35e95f5e8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d80376dc8d0858cf2174213fb654154fc5596be68e732c16fa4e6cf17cf5e1a7a0785be270183b7b0f64db217fd07bd5ee6556016841ed;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h51a6b370c2b0d5d47bd37273cadef806d1080f2cfadbea82e02a8ab982b0abd4d326d640af04d2bc404e6dfe83a33a83337ce039d85801;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13f2a374dcaaa3b324177cd0e8efb572b96063dd238a79e47286d5741d5414bc3b4ae77c32db2b56cd5f741e27c99ea8a3deaf26a1acf9e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4367d6c0739ab44b8bf70e7ca6ba2046b881bb8756bb0dac5a02ea342ee62dbc4a929a338bd1102a10469280f071603ad69e973d4627b2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c4492e5454717877fbec39c5060e895b6cdf0caad0836255188534e390b2895f4261a17f83b6a158fbd37694617eb79992ade710c15970;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h172f7c42a7133a5f672f1ac2c30af31d14e9c4630a5f28d0b621f2df5935ae69174875edb174baa20e4f1988500b2bdadc5c80ad7a7e1fe;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h337dad9dfd8f17181793609c2c3ffc4cba067e1cf0712eecdc8b7359eb15c79ad63c85160f40982c9e110d61f96a21a04aa77eb11f9f64;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10a4152ed87300aff67a83b2b879cde77f257d073fdcf84083e07fe316338aa10dd9ad75f853fbf2077f004fcd2263d824b492f13986e9e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4f4f8daabfaef456a276e6994b254e42c60f20ed10b93b554c22e6425f91c629ad6dde739929febec9f860a21314299dae44642bbc20d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5d7475e5013eb4dac9c6064d927e59a488c83f99335ba9af52c408b83af5da4645d8a39842d06b012194cc4f5501f50a79f0297de13604;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10471cabcf419b77b65c0b0328b9da4b6f59d4edde27d159def6f532c2d5c9c3b9e14676964a5949ae0022af3f5e821a236f241a0e4d2f6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c96574f6db13436dc4b06fc500bffcb46e29d038f24bcdb9522c580ff734b7ccbee8eef206c3ea20f71b911f0e392231f217b9a7d8abbd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d216d09be326dd4c3adc59fdd5c7fb610904456948b1cd06974d39805687ae3a0ce375a9ef580da6bff97f1aaec08ad1736f41c71bc552;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e0661ae217e61f33823fb0a790dd350df7a1f9eebf0b601a63ca7115c928b1df3650243b629191ebea2462873b64b774d9b40862e117bf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bbef27a15c1d60cd34aa1078c0cf7bdea0be229de1c275b2006efa2f14295cde849114f8ebe887fb58b69585d3552b78c3258b3689bb28;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1785f706263f8129a90ce783562e0115b56030e9a9a97b079a3351c1543bc185637ff38809e18558015e7a12bc9cb172690cee6f3f91c3f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5239795a2164e1c8081723874872113c08e1d8e13de9778dd386cf04c4a210c1550be6e67293409e0b85836d0bdfe6b6bd0f862dacfaed;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hab0b8c126bf2418d898cbb70454cb44420c7f5b4a67f9534293f94220fdb4973516cbf917bae0e23a7e113295f0308b5499ee81ae3ca7d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c1177ea6b4e6fafecdccd47dd6428eca589ce8841ccd02bbc51786605d634aa1e56d105276b6ca575e521931a3203419809a860b3310b6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1097737b8d6c30f5149a977c61029c3f7d52bce0387e7c83bba43b0bfa081aa418c9c4d570ccc6172f26c574f495d49d703281db840dd9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf2ccd960b6443aeee41e30f3fa4941b2f280cc6bc532677d17dcd77e74d538df51df84b38276d9660207064ce41e9250fd0efe9bcbb961;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8cb8d697c5319d97040dc80bf771b51879ccdd94b41d6dd8d60811ef6091e7e4d91bae2a383678838451dca45496017997ad222e1a7ef0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hca89d759e41fc04bc6319bb7bf2b190b2303fa7dc4f8bde414fa666f378868a37fccc8debd5b4fe8cd626d92076ef8345a04a8d923c2c1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15a67689b16cd9a8b19f15fa3eaa3c5617c2d56cbf94ee9555295743b27af18510710fbb96810f3656b66530971b4ce57a640e56132d0f7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b829a5914ab1a7850da8fa19a985627e1daf52e5af94d64911551a03d9d6053e74de2817c458db56deb0b59af34fadd1194ba7db3cfda9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h51a0213a55e58b8e51fa87675e59296e612245bc8accc600b4ab5619b6b4e52d6fe9ba09a80eff3f2d0ddddcdd2de6523b62235a3a216e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h42d9b960ab36448a557521fd961da0f32ff6f59eebbde315138aa71c651cf2537cf92b3dbf684e6ca8a18aa8d6494960cdb62e4a452cf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1894802375a1dbde6f7f7e029f5e3d9e1eb8cda671bcbdb50c71b45ffc346b21970c24e353fa8da34fdd247d7e73a8a97a39f05db59d30;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15a2de6908455be026bf32d732a3919bdfe622f18eab2b9360f05d6e3e1ad69d5d43ce754b5649ad0f0eae148fc9171073699dee8cc018a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c4df943cec615db2254516162137748b61cb7ced25a9cd32204b8c590eb4c15d4df0226c2d67227945303d3a810c80a8e22d95fcae0a79;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb96223a12314b08d58ed63d7a86746f54205b92a6e786d03b3a71161c876240ca897f02855e85184dde3f959cb127714043f5c6817be10;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h82f8be52b02e17e16b33e8473f336b3323b139dad0353dab227c6143dfcca97c93294995956bf81cf905fc2a98ef95497f4c4319f5a7ca;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2dfdd7462b392fe891c98d5afba0ce9eb9349c75114d7a0506764795c59a1462c93d1bdf231c862256efe3d90caaec8a120609abbfd152;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfa524b5504f2c2c30d0625dbd23e190e9f76f63a49706ce9116a158f09d7e9547681ba48fe7422b05402bdcd77c15c46dceec12a7b2d18;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17237f9d4ca41e6d2c00f6de025e70951c65fd8245eeeb2d1ac147a37b88510420d613ffa5d3514248f74a945873dda4d28ce1918698207;
        #1
        $finish();
    end
endmodule
