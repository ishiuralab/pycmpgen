module testbench();
    reg [24:0] src0;
    reg [24:0] src1;
    reg [24:0] src2;
    reg [24:0] src3;
    reg [24:0] src4;
    reg [24:0] src5;
    reg [24:0] src6;
    reg [24:0] src7;
    reg [24:0] src8;
    reg [24:0] src9;
    reg [24:0] src10;
    reg [24:0] src11;
    reg [24:0] src12;
    reg [24:0] src13;
    reg [24:0] src14;
    reg [24:0] src15;
    reg [24:0] src16;
    reg [24:0] src17;
    reg [24:0] src18;
    reg [24:0] src19;
    reg [24:0] src20;
    reg [24:0] src21;
    reg [24:0] src22;
    reg [24:0] src23;
    reg [24:0] src24;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [29:0] srcsum;
    wire [29:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h81596d6fa2fc7f9ba5bbb7027901e4cbe0e2f55b6477ec788e14c8ac164bf9ec882f635b4ad7333998775ebaffe914001076e67a177b3ab6323524ae612a3cf604994f159dadc30bff63a2869c3d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd88863328d14de56576686b45f96346378521db1d02699c231c57c770bb491d4fe2492d386042ee2e82fca48378d03bd97dd75c10d6f1071e1fc7a872886210085a0f3fa3d76e5422590bc2dd86f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14c19fc91a5e56c8d8911286a1660734bdbed2df92696a9fe01add9b3ddd37eec5321d248596cc64c1cc13a0c567b30dff6ac488f7fcc37554276082d4cfaa4d89ef40b850ccff43102a445964212;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h60d235ad429c4f8652f7fd2e0bb8faff13adca35006b83f6d37d9a973c668c3745936c2a1c8ddbf8dda6d71e15b1538615273fd524382edba060a66968945b51b5c23db43a2d3047a59e5caac61e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h113eab30e18b0b12191752bb273edfe3b6715bf53b275d305fa72a26438c70310b3a9e2ebaedab38e47aafbec4a9632e5f1592361cabff2f326dcb646ac3b5edeb30c2ed75a7476a18398671a90e5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcd567115d2b83b6589ca7dd2d4e8c06892ec2d9e2c7a4c5d453d19488d3eb33295bed7486ffe563baf9503bb76532a796ee8930eeb5c9e5a8665b7373f5f88bc9424c69738bfb65b90c604defe8e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc496de770cb87447a206ee0fe60e53fee5b8268b402765baa427288dcc11a08e8382d2300e22e4b62a45f98d414f0b08509e8d6a5697a8c0b3753ebce813650f7337301d1fd4f8af52cb335eaea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c5ad9c6209f30b025a0b521939f1ddf6500a3c0ed4c3b4cf7e45d2f65c3226c21bd3d62c71d240cae0e7c8b5adb3e0ffb73f646b01f7ab638b732b785ed6272afa17cf3c57e2c4ec702af3cc9521;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8513b903bd5527c995bbe43ff93fe704b7cc155570123371f3655afc114b5c95cbdcc5f55422b2534edab4925e299aa6069b5b6042c8e4039da3be5e7fd757837a819eb491977025dc8b94f27294;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he28d5caf61258b01c05b4877bec023878bde269f2973bc09a6e8f3203c2044d5bc5d4fe85a6464f74a9356e5165de6e544132920837b7d7826f25c9f8a77abb6bf91a676c294ce114e5420085c04;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc9c44fd6aedbd3ec5967b703c2e11729d2c3676e242d34116c68aba9d2c7104767e2b148e9e125607579e8c6733909e8a2c0d6f0d5af7d42cca9c8c1896051038e0fd459c7091c8fcf47937357b8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11b1731c94d66756e09a2789e2efd0f9ce85798eeea3bae11641673fa49a202eae1ca1f243881f102b61292e0e87f3580ceeea90f5a5deea533913a657d4e07acbf6d5b97991b09e6b58cf8b8eadd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd7715c9dec711be3a8e2cd9421d240f4ac2c17c314a69abd88cd98645bcbb3dbae588fa9ee21d45d459aa9b128b42811569f0f967ed147e1eaf91d3634e5774665816728645f8b5c99ae38f0081c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hed2750e0f7459f824d1e318095907c5f0e37f9f1f301e35d00557bf729efd6cce588349de689eb1218417b1b95823ead8051a6141b464c0e9f2d7c0ab010fa05285770f7c30f28eb4b669d5bb196;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f254ae17a906d2bfaa7ea0bbc02cef358dbe3f76b5c6d88a9f1fb73807577be48e4d1c63c8be9e7fd03b5cae1e224aa6ea7d43768c4ca422725c0eae5f1175e51ba32693dcd2d87160b90cdfc026;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9e67030b011b9a841cfad4f8611e30ca0a57cde7c66019d4328cd4e38797bf4158de559682ed33251ec5b19a44301fed65e2014329582dd16945331a6700130d1ef9dd1c380a60c5d5326344989f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd998d80bd12d8282f46d0b368fb2b81f92cae66d34572d648c625bcb5bbe8269779aebb4d93e6a8c015ce38e188a05cec4cf84e9da9490518598694336b5712b08538691782aaa98c8d49b383424;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he2c5789707d7486b16b35ea18d3462622d4d9b8d70fc2bdae17bfc0367626b51f65776cc258aab2433432edaafb527f590041b33fcb24ccb17c06b6a077a6889f931a0fd33bf1d78d2a70dfd315d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ea63233b269cd6f8e19414a3b6454d90505cd8a40df0a7dd40a431da1993307ff2ac714ed127a6c7d59cd86ac4325bae71cfbefcf6c68a905ed7f181a422ff3e391584ae374ed342f089c25c4659;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bfb9c19cee7baa8caecea1d931f752e48f23cfd37c5ba8f2a77ab996c71fea1c2e1f2316315af0221e39f3de01f232bdbfc6dde32aa7159bd88c106082adde2c7a18b1e3b0267b1ab6238963ab5a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbde075063d25e972ebef33ef922dd102a66cbcf43b109388dc248abf6898607a1528b229584ca00f787475b1ef6bd5a17696545a06e6ef471a74775efa01b7aae7203440a98bee741c386a51acf6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fd25e8d0243ccd00cdd18bb2bbccf810aee60a8ecd700a69939ca45ddf023e88fd3c61cbe9ee021974ddcfa4bc3d3098da4b2637a722a0bd46694525653c3be9c2d145647e7d88163b3aad97409e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha9fa904a732cc2a7e33535a9bf9f8328da9c8a8b69f4ab55792b38cb8d58d733a7f9e1c118a559771bd5b46637dc21fea51a98e444143a66e03f9961afd31750e6781e6e8c5375e491ddd8668064;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h45ccb28c783b7557c71f09d837b9d99f8b6b9f2a198749bc97a42eca2e421dc36bcca2e21b4c267ee3662cbeb60a84ac0c882040a35faca60936dfe2aa2546ec763258676d903d9da9dcdc26282;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h198a66dd85e622749ac8088115220d538d7dc60309ff2a51c422cd14296e7bbba35f6214ff51f6c52f63c4b4aa1cf1a9418259f65dc73c5c5162a9af19776239472a7be539b6bd0964ecef7544674;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h64fbf640c27026b8d5bab14559633b84f6b1aef3e3bd1b52747379272500d6b9726524a18bec8e26749b854f5f7ca1c3b22bee2b187f1d7ed68d8ef5af59570da7a58b55755dc337031f69ba0b62;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16e05b70baeb58b65693d3584cf9c6b82202e8580b3fbafbef4efe4d500a20a7e99ab68d94f55db7ff849b7b97c87bba77072638dd583eadb0eadca8a205a48dea4fab6577ad157498ca2cb9e7df6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3d9c487d6a7c63d382ecaac37e5d03592165f6555b8cb45c14de34782939580826a9b7d21a95632c73d3e8644b8c3993ffe64c217f89dd210c5e3a73501e6f5a9b2750bacadabe60e7f1d172eed1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1458906febba48c59cd617eea39c8d26b2b5efc609c0a22fe0d2f25d9d4aeaa94312d4d9300eb74159882bf435ddfa2bb9c64d66347b19b099f944c051f64d426c58cb657898cf053d21d4148d7ee;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1db3bb7cbeaf10c61cdbafbe528d8e74d64d976516d617e65707dac9dda1f057645aa77eed96c9085a2f67e7d50770ff795e18b496697edd0eb63ca7a88c7ec9d572711c4a34ab09e4d4d39298331;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1241ed856aa31d674147f86b0127a6c13d03f2ff931a1f8b2058aa5b4fb92c9710708858e32a653d9f21b18110486f18b6aaca39486b60b62c1450280315fbbacc633a89ce1dd082830df5a1c6e54;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d5a47f995a73cc987858814324ce44bd77641dd421858b0a2238a0e0cc7a4b08c78c683c1c905f47f7e7ef34a1d3e21aca8f676ddc086e61321e1f3e7e10e32ab26db9b7ac054f7c26bcfe4f1e42;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb42f7f7941cd6e6cff5fba48bac929b0dea47c957c8f3c24b611508e41115adeedf0521b73eec107da468bfc4c78bb6206b6bda4c63939ccf1183ea8790b7819189bf35926133a309e658b52cf38;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5e2ecb826bbbdce0d6c57f4e927701e29ccfe513c08995a2a524b548335cb066466f871d3ba3ab217475b81c08ec12fd5729bbd1ae3832fa067b5f9b68651d055434d061b2a5ac9dd3e597de9425;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h185f62c32bde3e8033a83b6e6417c0a99407a1b4acd5a1cd087e65697b1e740a1f749559a2ffb34ee459f9b504e851e3feb37b92aa9321e8a20989c47fbff2c0e5046af39e402d0fb2f456343f294;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h538760ed3103f541825b36efb1e2c66e87d1985cf787950e0c70abbf016bc5c859d371faa591176aebcb614a5bb883f9e59f32be71a8ce5ad29de18e1e5924b1a32161c567d5c914adc8f869b713;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd1b6312d1220715dc1cd2f9b54321e5ba605effd5e22bf2a38f09fe94464a194b9294eca70543bf0e3cfbadff557dc029444b358bd6fd2e83efecb5991cdd79ec77ae5e7a7ba0a78a6c7b6716b95;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ddcc0e01651b68e632fe0b355b4efbac14c0cb9f47f1c0fddd28638c3d0b1890e6364d7067b4921ffd7ecd58b52e6eb6bd461d0c9a0377d65ff5cf7055491a417e9ba6bd51865546d05fd68bebc6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc67e58d4aee7cfdfa98d1270f18ae7ef251ee6fb382ef575c3348a360914462ccc09b76cddeeb5786a831d7a30c4777235e5bca4bcfc5d24b7af1046316151767c60dc1672f9bbbfbaf8b00acded;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1850228650d5a470998bd2c9df6039c5eb4e422cfdbd8ab574fc377de0a8dc14bec783de07d58754fdcb95a3710113df879c1c49ebb00ff8fa1d99e01f48574109d9b9447d65577186dd65d99a040;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h163fc994e0c33c97e0b6de3ae2bb56f8cb5d3d10f2cce9833f86a81af6a1c05b57364202f524812f0f7f98e08d79b9dbc90d63c1c980f548ac8f50ce0682761979ac677683f5bb1fbf0931fcc10d4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd70968f372dc1a0fd9f9503f886032d0cd897663d22b8add035db6cefb32ae3ca6ea7f595653908a731c9660ef6c16b9010d737da951277fe9fab6ce04578db8e3970bf32fe29819d6f9a9585b4a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4ba6f0640e3a8362b3c37de90631162e564ba63cfe0dfcb2f43d92e94b7603a78f82f9f88f48d0109dd9102a4f31eb0b794cd3bab2e3a2974ffadb644f495a9defc3e147d638f928fac60dd92de5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1959b6dbcce2c33ff90723ca535477a5011029042d0627aec33df79ccccf5b516175d3e625f2ea3be4f1d747b0909d49b382ae11da33cc3ce95ce9be767eeef973bb1ae4f50bb199570e4753abebc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h87133343aafda1c4843232feaa4599c23ecc6fe2dc9e2c54970cabd75b3d15171923d4c9cdaeb489978eabbc51e42a7f244c67d9b263f588d2c22d7f4976df1f265120181ad88f33410aae475b25;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he87c00560ab143379890de00259d89d4957a4d86bf80880502aee608d551c8f01c4eede25d41b8da88af0e0875c258bcc8c1a27a8e8af8e713600ca059cf7cd11eef72f30901c494bb34b6573f8d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h55dc63baff9419bba794de60264151c80704049fd6ffcb66e3caa442e2b4acb8aaa717115e6e2bc987ea40cede954b3a07c61b9cfd7c3d83a23f861631621a61169dbafc8b9d23f1cf2919aab81d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h63a5a51ed822a0e09580a88a9736877fcf4e86ea0919628059049ac391d44a0d224e77cc0b0a2b7d24da150e2f99366c0c419966cf0e0c937f0353770e872a572a3a113faf2eaffb11d5a6fdd141;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9997d3f0a1c76ffd9ec5b52be3b537330278c455052558b7e51af7eaed258f90154594a47b1137a47cde8388b3e39c621293f9be91bd56b4d993a5c6b9d6294acddcf5b259c36afc7d7d373a38f1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13f8e3ee1377d42b25d22d60ce0c36f433f2bf9056df8e2a8fa45b47ca6bf11fc0bab01512a46fa1412ec6307c0956518fefade07ba91ba6e604539a0badeae461fd9b3ede25b976aa5aee016cc6d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfd818d3b5018dd415946280d75201fe923a76e8832c36a7cb2b325ab021a9f1936295444f9f501ce5a74392d20429e5df5211a672db5f018c02b0bb76ff6b65310244adcf9f7c6f2b8e42f5999a7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbefeeeaec3c91d98b9a328dac1d78f3e32abd0c4a48e9ba8009be395390e247cd12dc241232fab7b25af1aaddb65a367867daf1d06206d8358fc62f2d9e4be5146f8560c959259bc02599316e71a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1adbd009d58509c1d59f7b3c7e53e4947ecd5b3e913870a7e17ac91e03cd51d5683572a4202d19e1ae40d565a3831e1c583bf6ebf7fca73783daee8131d37d46daed3c73bdf467601478f932abbdf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5a6bb19177d20c61bc5b4f3683a2af9dffa1a9c813590cb0b858b86572cb12ccc2e249d31c6b86d108c52b9d38639395d7d773aa1b83421273c23e9ea61499d8085dbd52f26845431c7f09b39b47;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7e94e1996b22e87b6027b10ff8f66f2f7271266e6cfe18b4386ee4696e36bf30c0fd7911d95f0a660d9b6d4e5bb24b8f76275f51a7462962b4977e7ab8b7f9ae0f49fef3fb6bff3b7df9279da4c5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9f18e60d0bc5ae44caf4ff5aa9a24cdee957ef428a18795e1539c245a781d20ac0744801bf82a3b96558d685275e9f84379e4d8a767e7573ac8da5fa02247b4942477ca42ebbc6c8c1e7160adfb7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc38e81a3f51ef3c76093900db296a58bde63fab951d32024a7c782141c0f6d6e9752dab351794dfc54eb4a49670016214950fd01cd8115d24c152c1dd50cfa0ef6a9baaf3efbebd8f98b72bf1473;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cf395ffee27805a799c5d1636ea4bf0ef24b884938cac33d7fe312e304713ba495a151c7499955c38dfe0fc1b9056d47578ef6b87e5f6a429e3d7836050caa48f81af3b6f72bda69aae4b690e289;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ed27d32b0f8eabe6db2ab3569820df18b53f680a2a258616d63d756ec2bdb149ca554b91308f28073c65301f2cd5f6cdda94b1b46cb8a595ed499fcce5230c0056cea3e427f133d5d93e4ba08521;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h291aedb15d05ad3bd936d1d547b3be194bc110391fb11d15b55077e2cc813d7e59be18928e3e209f4fe271e255bd20ea7bc0a1f472399a0f9d681d1fc8494b8784208928eaff35809965ba35cb59;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3fe799e220bb9862b068474fe1bb18051887ba8120d8075f6941ffa027b209092c50b9a327e4c60a9cf1a1f885ac1becf17517c6c3748225d7097710439457474ea5a5b200891bb3b69832b41bc1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1890b99f709b7c0d5cbf2effffe2d0ee9b6cd546d8b67fd5666c551bbdd51c2ae326787236c4a569fcb18dfd7f3a796d75aecf6cd256e99db6bb27f79f0aef6e5e69d204645f1f0bd031b6c661859;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1854a51e75b3583ecfa3235b5d1a5560e886aea753d8833d9f99b87891c2f56b58f89f87f6b321991a9b9f40dc4e5ffa5e17bde2cd7cb96d047220d9ed2f92b5650f8d4a49dc09f34265a6f8ef0dd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h105e430a833b258680fa9b2416e6ad2da18e338856334cccf91bf1e2e7b06d982734d2c0fb4f7291ce47c4e684140da3fbe33f3a4a0f4b8bef429fc6d2065a23759b9916060bd08de8354521b1e3a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aaaafa77f6b470e74ac679466389eca1cf633cc67a004f77005432f3bde077aa560668f36c78ba3778b690a5dba9f027eaeced87cdaac0591181f0a047b73f0581271dde180f2071ff887ce21fa6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11b6b08034b905f1c965581ba3feb97130703bc5dd1de91e9125aeb403e1a88d7643cde24e9d7647698717514510dc0dcd98072c202e4cd478493f5f1ac97a411ed4382327829f0c6c80af6af7243;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha9d3ad908b7b53d72a2c23f5137b18196596ae7af333c910209da6d9735ba408520d8692184f7af53f59b0025f2d50a7470a51287f6e0507d6f58f8bf01c5c1de28a1ac4efd3a14f7677a2dc3d69;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h157b7398c6869944638bebc3f2a7c17dfb006912ecc08be6decc1fc5cca371bb10f1a9ece2bcb776a3fd12d46cd8a9d45e28f086b287e21e9042eae38ea570bdc63705889485acc6c3c9c7776c735;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6a6f0ac440c88ac93c6d9399a4da1bb7c8d49d13e20eeb5f889323212d5f581e2ae0b3af20ed335058f4094e4d63a903faaa16913e00ad661fe13968ac22c2f0d8cd8b273fface7102957746c67c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1acea283b94e4de294107f17bf53a74caecca2de691ba9413b6abd64537f620da7bb9a9d1cbc44346fb173e2a262ea76cadba8d521b1de85c8600a100c37869da276605dade223a1e9008c858b383;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bf0536ca47484339d40041444e5475c1e0cd4dd152626395be983a8351267c89d4093c6bb8ec3794fadd4eb424a7564b01782066875f975ea811f98c1df8c29a72f4b601fdb60dd84d20fb5d1eb1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14a7a5ddb1d92ba1d7aa7e7ff96f7a31d5ce80fa553bf482957310a38ca859863448b0cb2687ecd8669cbce516f38bf9c5d55f32d48b612c7a5ab0e949fbc1e3b518ef9c460d1b22afd22b5988f66;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1147075fdcf2a7453e24b377d6455f800cc6742b3b6a2f43e6f48932046bb2b3aa67059ed477d3dd10f3c5b25d94b3e6b3ea19f6cfb36e03d648f7792909bfb7fb590fa489abfc56001aef1d6814c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h972dff6c531d8eff0723320e72bfc3d7acef0e1a54ead139a86bd752f2db9f1772a3b4dcac0687d10802ecc66d57914dbf961b10d1d67ba8be2db11e1b183cdef78b5f6653bda04c99024e782ebb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf0abc8ec405578fcd8c7561167c31736743836996e411975db53fabd4cdd262075b987ce5beef7bfc9fc958d9dd3b02a3862c78745d06b57e0f7ca8733f058dfa22ab8e5eb9fe3615838ca6ef833;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1db893076a141ea71ace7829d3d6edd285119f390c8928802275cd1b2d449510c8923cec089057dacd4c62e7f4a1c6885b96e7af38b3b03ca6e54d21fcde42f56e897ccca7f12f65a8be167efd9ab;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h37343eabd2e60208af476691b6e03323e888d431f7ade538e4c16ca78d47aa3d3697d86d114ca5374152aa9bfaa050597be273fb19fe1f4fd70ba617dc1eb6704ac11400365e27ef8344803978d3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16b0cd3236a3d6ecdfbe23ec667daff994f51fe907a962eb5dd49f0212e14d492d7462121447b245517185fe3a51ae1cf2d229ec1e9df6e455839eea1b202f769315e817650d4936878f138111fda;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcfcc43e9126cffaefcc915787836670ed34391abda436085182d385cf1846585c2b7ae74401dc0f5b42ade1b1abe31e64bb06fabfbe8f63276a44ca4a97d05da85aa2ee3540cb946c2bb82aff799;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14b773b430c70cb3fa6a69cd8a6101084b4cc259147ae387525f79922b1e27d91928b065bf5b5defe6dc4e6f7648e2fd4df214176806f5715b55bc74057d5ae10c9a23e574533f34fd0eb3e3e77c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he93e4da8f6a4f9df7049f0ad271c93b2ab290f54b27bee8e85279b5d834a7f1a0bd6ad31f41e215609bbe1bc4da04bb251054785fab12a491bf8958729243b1be8ace474f0b51b082634221bd8bb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1acf840a39e73e6c15454a461ba255f5937bc8ca61f2975d603d17370ae35662de4777e0d60660e50183968a09dbfb62bd0dc6cc1219676ac2e90eac4384d67f5f171ecc3ca1c6da57e35d9e11b2c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13c3a47ca86144c513ea628e6a11e6e3ef9e13a3330b95be2494f403540f7d8b57adcec5573fcda0e92e291c8d5222018d5b20403fb2865afbaf67ff6e09265b25e7a48afa89d3c1198f38d61d477;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dad4bdf83ff4d90defe69e6cbee731eef648319d99548a289042551da9366a9dcb6b660498e11890ad42a541f3e633a843adb3b46a7b10ac945c844571b3972190943b8a3ebfcd71623f1c554e76;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1be3cc92b34a3b3b44a014219ae288e8ee38710da89982c53ee5f65d09d482680707d1284a5ab4eadbc16d057c2fcb87320ab637781c8d24868bbbd360b3da13d0cd21b0be1a01cc5e464af86b142;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1947d6bcfc4fb414ef71714b6fcdf659f059311e9f9ac52151f7b72f5672da919e86fe6a1de1890dffa61d6f69127eee60515482376e6f0c6c0483066e808964ee6e6c43d87fa0fb7479ed93339b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h66113b9d475ebb08cafd69a2cbfa2226d746da1de8d4c421e85a0a80237bc83cd5c60e1d2d0329fdc91ae68eb130cbaa5a613cb105eb3a54eee6d5f3c66a2ad88208775508758328f4e571990a34;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h173ed3e4c054eea48b61e367cc599d6ef2eb49923337bbee1767e23f595d07c13799df050a54b83fc1e8faa114a15214d21e343d694e640dd1062f26c400e22d54f78802903e44193563f4cab17a8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5074c2fe1ce633d784c1c85f43a0016db3d4f9640a3bb223a958a7b7012f791bb5419c5197342d072ecad92facb3bf5dfbe200b0a2e7a7c5f85c6980be720a5727478c88483e3e5526a0fc62b835;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd1eaf202f8ffe367b1a38d8338266416f824b3a77ed1da202738c31caf8731a4fcd83ad635e668da8ab291ff368d2323fcad5f0476bf11c6febe2702eed1f966259488732beb6c9a97997afdab5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d9dd29148d4ec6c512b1c3685a6d05b9c8c4efb241f944d800827a1835f06735508055b322831b18035fa60c4fad629549e4e956beb40e54982caedc8a196ead186ee4f146fd41c4d35e325efec6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha50abe00bc375d9d626d6288d2697574419e5cb57480df0226860a74b4926dcefbcc5e425a92786c51b0d3283a755668b55ea5b90929d4d830a02f38276e5916abb081edc8b03581d09daa650436;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18eae054ce51275476fdb4663d7ea539aa867522e3bfcddb4e8e73e7fa07735b4cb0d3f03dc390b449d6b2b90826634f358ee381a311fff5ed4b6dce7e51eefdfd2cda304a6fa459a632608ab9f84;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a03dead06483772e7661539d3c39a7ba5834b923a0513c4ba78266949553d9ea7f8d2ac7875727ed3d60878c8392f9b3faf6bb873871647c15afac1e0e8e87f2b58e8029f17d51553ac3f1c6e95e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1825e021f16ccd1daa097d2c604bf8b67e0ff08b79100c07fc281c21384e39d643efd8142e30165aac97441dd2c618b4d40ee72afaf90b11b8f9d8cf8ac45e0bb80bfc91ce8326b3a5c92d1b5647a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h82ca729bb57d61026882897f2f3f0889924bd535c4ab4b8cfcea71af1811e18f5a2f13a6fea960e067b04ef68afc6551082afb751aae1d2f409062f4358b2e3d67b02b73fb792abbcb46538d38e9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1757b3ea4b32610159006d2e07ee66a86c4382b16fea59db9345ef6941dc72734281a070e023bf5940113968c3f2e2b6d2c6c242b6bf60e9624e6a96d399c84440f075d1cc1a4e607024725036a14;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h659296ba8c40e09a3a00bd18f792295162f9ec1e623a4911f226154210293c98f56cd0944a62af48cd3bc958c5557a9bd7000a508567323f9caf1001f1d4dc2a1ebd3f1f5268aa52f0aac03e584e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h870737276cdeff586e7de30ee827ea548ce681e79841674616cf85ab452aff6f7a473ea8dcb4c091272dab3b380238ea9e245f6fea7993bb360422e0f451e3c0d13ec0f1e5f7fd6af0d7cf540420;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd4ed797fed31fe335e98e821e103cfdac04cf877ed285d835778ed209f927e531048ae2bdfb2c65d2aa9edc3222158e19619f1d5d0b7a60a9e1afbda7aeabef623ee905570628a54ccaadceb8002;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d7a0b38212f92e8db2909985bfb86b43c49242fd0231bafbbd15922043a5f71f6cb7b9794b0e7aa1e64f92cf91e853dcc29892378344dbbcf25d99fd90b53da66e549c4835e242d63ed99744114b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4ef560d70725da35d4f656f96025a38924038556e3afd52643643b6d16c15ee417ca67d19d4604f641c748a7d33a3e7013e73dae1319ec627db20d1426093c3f76a64ba38ea5bf545c5aca1b651c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cc1fc8de6d8024d1111aa1e07f7ca86e381175fc716345c8cbb857f362dccd7c33a0291b46795a864a4b0c2c684511df0c16c28f12acf633d972c30438c849aaa2ef55c71210b3b7dc3fef576c60;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hddaaa9822a5bb7cb5537ffaf09953d6f51b5d937cc2c31ab3975d44314bb459c0da5e0f375d6bfc3da2a6cb803532f3ceaf54bc756f75fce6c07b37098aafa8ac1d5cb5b481925921426f7b509c9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1739b021da99da3d1dc8cb9230293b6a8ddd66c680c89a9bdf37f8345c22875460a03d3f22c4dbbebc69f9cf97f9135926b2b8034df502bf1811ebe03f946e28202b5e5a25b47acaa9709f5d8c86d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10425945fa5a135bbeaef103d9800e230510fb97526026b7fb0e4dad6ac78df22f7c7698737ab54e721fe8f76b34ecf240c0918d92b82c1efc315fb3d9d16e589d89c0512d19e4af487ce0d1c3e4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c96362312525bda4de447a0c82b697c8d25b6e6eb77bd3a33d728d42087537b5b32a3794e812a09fd47e521de225c88e8b8daa6797a5daf2a1f01281b39b014d0d065f83c71d9acf5f6f45e3c7d2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc5955d713fa42844c2a57f42bc4a69678ed2acbc1cf7b066073d57756a7e935e96134c1eac3997b4cb7f364299216f900888f23d4a3a0cfc6660dd7d30198e56a34309bb44965a97ccda1b30cb6b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb8dee60e56e6031ef45969818669e9599ae077335e2a27074076dd459892cf645625f6f026637f293bcb345a6855eb7407206c90c509d6e9ba4952825abd446d1febdd1437ddaaf717ac76d11965;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e39c02c00a7b3bdf1d2c36907107cc7dcdff3878e37b2c7cfd2128eb761d6cec1192fcf214a96f8da06fcc62e2462ebdba495fb0676225df36d8e79959186ab32bd23d26308de2f6ea2046a1e482;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he7616dce86094ed6f929c03354f50b71a2abe10d74cd2c9b2b447fd88c8f3dd28a77cfe382462a4f7d2405bcff687bad710b2b0f9e104c54609f3633992a9bbbf43a2f42cd98e798440ff92abdf1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15b3affd595b1d4726c73c91b3292edc415228533ffeffa35cf3397da106972c7d1367a0ca9c53651a5cbf21540b6274aa66a6b4f522d994c6f30691d5150b34c6699a3047fdd94c99734e4719d37;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8ff34dc26a9ba1764bb4009aa338e542a4947cec92f3cbe927f560645f3aa301eab8f6ec1cecaaa8bfc436f91cf6269d6cd073c9a23c58c31905f76b7381b6033017ad7eb7183893365b5393df8f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h52fb2148d2bcf0af690c0af22d6ca34fc7a7ee4904adfa9808a628737ec4d9578da9606733d764319fea1945a83aeb5db60f47a9a0d53dbac29ec0a364f19b034a97bc41de152430a6768724c033;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbf4ac558fa4ff81e251e07aa3b0713c8dc9ae4f43b2018ffe9b8b2ce304a0b15cb76a82ddfe928e05dfee48b128be03ca5d5892dd34a97a52e2b7db17a70515ec414141ff7d8b23d7d3b3c35f1e5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12f65214cc72b5e2118b3c0bd54842583c5f93ad38affb65139ea4f5c0f0c5da188e95f13aed3d8d36e63322c75d8f1248c19da69ffb87255f62e6e0559b7daf60e948f68d989c57ca6edc2c8f2dd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a1eb4eba7efe23aff3626fe9e279d827457765a76f41379951671c180624d5223899dfbc9e5752cc686f4e44a5b007c392eed5034cf087b921e78b30f0d417910a1ec00363ed04768ea580d9781c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12d66fe3d623fee755e6c5d48120ee4fdbca8960f4ba3f131c3251369f84991136b16c2b56fe5b972a3280cce3c30fd33389d47d5e85805af9c5b49058e0cdfd609831feb1aa326b1e4cb5a3755ef;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h31f4d867a80346ef1da73c956eccbb1d16dc22cee36630da95c61ccccdd3a93fda7258449a71377b473b47ba2a3e95d1d7e6074205a6200814e9dd683d39f833f664e28031efd4f52455b7824541;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc5ab320a50c9fabac2215392798ad1441ff37b89acd9efb33063ca74d8f08581cb5ce57e60a61edcd405e4710175d086abcc05d4db237258e914ea79f6dd59711e438ee52ff1300686b54f9f7bf4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h22db293751a29f4a5ed6b5408cba3aec2c1e440e315af201ede622e18474b339a405933d189fdc88c0215c75b1ad5013848d6b1f07228737feb83118c6ac81d484586f76790e87b95c47b728c491;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heac2757d08209bcce01fecd1e45e99752b2db27879b20f6f7905330c11f47263c8ea3bb4b797051e9616327e479dd8adec872cea8b08743b3c10562f590cb47b311dfd27e0e9778bc3d4c5092c29;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c13a2262d4a7a32a54ad91445600497266530b988c576e6dd985d87052ca944e565b771c19f315cd89eae4ab3b2bb7827d7d277893a0300e6bbd3f829f91b57184a363c914ce746c7d1dded45da5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h160cc00e41f234d0ae78d3ca902ddb8f6049f9db9fede85a45611274b36cb6965abbf6362fbda928a089d0e1c89c211ded9aa906f60e20f10931d36f2130a743afb59b51cadcc0f81b5a5d7adb42;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b229dbcd714777ecba8ad72ae034579b27f0d5a11059b2281f3b4ab5faa92ff6a41dff7999b9110da37183e2360ad2e4ce7c508eed0b25dd97352b09c2217e5efec36380fb83e6c80d67432556b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc0de64764011805eb15a96ac08d1a1f6d4043fa6f816ad0c67b42977dbc6af36b0a5c482e6d93c26e178f39e81ec2d1adf2bfc808592667e99db2ff1da85426cd0e277e5aa7625d23faca2cfec8d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h148ba731d29dfd5d87f43b68d05a0305e93b6a58481d885376a6c3e0391afebb69a577365da7b9f921ba7c235315446dced0bfec8798fa8ff3ac001e134b29d3ea5a6b0ea4ad0cc83c63a97b924a6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c49dd82e07d9f16eccb40962f729b60b1ee598b987f417d78e69b4a082d64abef96a8043c74cc3d3e76d508138008b2a58d8ea1f4be3cf824cdbe574ec0e592c205f9945d925b9f130641dd60f0d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h70b50e9d2881e3d74412c86a3e4bc2f4ef5abbbc3cc6754fff0a025422d1640743398a825e3e2dcc94ea365d625f566daf0f9178dc6168acaf8806fa806009b4e863a18821ca4bde64b69c0d7dee;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hffbb4dccdbcb0e5b7e966404415620e827637aa613d93cde6f3256edce5e3388db251ecb4712d58f795fb44e80d9f368ada6469e765dd02305e32fe3853695f3cb56c9e2f53eae762e48cbfd475d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19369e6b4298d40a95f6dacf8c6329f81fc94665e4af3669eae5be670795bedc666aa7b6d9ba6c3b5e4605bfb9c911c969616b9fde22a963a9f93fb70e0216dfaa586c41e8eee54e04d085a8049af;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h739675cbd0fa67cf2493d26b80c9d61ffcbd12b2244b8472baae0152bb14cf1b40209cf59ef86bb309e8af99ac4e349375747ecca440d687222d404feb0a8cb44426e1c7c964780613b1a8a449bc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcb72e515a82d4e25d6bbbfca7b48bb913623cc48859ee6c3a1ae4de28c2c39135fce710a9087be8190c0893f9d2e0de4cf98ec6feed026544ee1161cfb6c4b4098b0716928dea28b43bbd38418cd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ed289b4529515e37bb262f41bfb5060ee7e11fbec7b642af04ba46cf664851cf34373201d391432dc61015dd8f912074b150fae43c7d7246a2b92115de6dd3ae8987c5051da6c651f3def9a8df78;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19af3a9e8aada49aaee1c8486a62271b12d14e77ebe35a8fc1b18f8c0956c7633ad80ce15c95c86a70665e8d8922a44d0c4c9a6d2d7bfa97e8a67a827b2242916371c33c0ce0ef95fdb01a0a09007;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16abb9e8b2ef73c16d8b89e1b58eafaef6d2158d0fd016dc3eef838d7c1d4c6b20a60270c8e65cd31f7a298b1fd56f6357e25b6a68c77e6981c16ad0fd51a90d41ea1cdcf9b7c46ea36f0a7dd1bbf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h277b306e60ce4da08e79113e237522df3daa1735e07c9b308f3d9f215d743bab007ead0025dbbefe2a82a3fd7c08765762051831a5b2fa0a70accc8c06f5a61dfee6bfcee0113c40cb0b14a65dea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10048ee8ab89120a1c2c6892000fed9312cb087c0977ae0a357c0b94f02e6335e388e374fe9e88fd29cb96c7d80e3753423ebe50ea2c0b924f8eeade7142773ae8dd76e8a1610f23804384fb0273b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e8d86168add4a6f1c663aad5d2adaf369fcdb824f40823397f6586c22bebbb0ca21735a3bd8a2dd5040897e005a4f948848403f22770c1f35cfa8bff70d98df3123c8378f119e83bb640a84345f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11eaec1b1986ddcda2cdb8fc47f9d1cedf390aef1efc3ac65e741308654fb28e597e461b8c1d099e5e35ca7c227134da97726263adee58bcbc6fccd3d4d8d3b189cf8f4509101f6875b65677f9b04;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h64686534f41581320bf24da71b67103c57859edb17a6e312be5e9da939261b37557c8e609b1aba03e86b7db74b9622554b39067a829e7b70bc9b7bfd255126c7e9c0d8bb22df0ac89e63cd89edfd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b01c25dc532b8a087aadca549240b434442ff852bead0a7502603023b0e71481a32935d35f71b1929c9c548a30cea55c446d10cf6c2c3d092ced2f8d22670c5d0e4440f7f7f70ced037d28fa7e64;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3bd0c16ac5ceff6c42a0069c317d9a8de3ae120b4db9eefcb2c67005e4026d4742049bb244a90b6f079d35ec91fdaf314244a8c530eb0b7fd1eb73b9607eb51ea8cc45c4aeb529994e4c8d6e54fc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12a7a2e7019a088683aae89f154e0655d0a69fa70a52a0e59ac7792f60b06cee3fe076d70df399d0d29b2e46dc277068d80e5bdafc952cfc68ed78352ae1a54653d3170ca1d93ec6504766bf304c9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c1ae22743efc2ac7e5534eb6d4270b1660bd57e152a3106b7e2477f442311dda3cf21dacf057fc609a753737086719ee8f0170214be83ba10d8ad0124ef851562768a386d84e0b52ee8826d1f6d3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dfb005cae466e52a0e39ebeded5268d2fa7d97c85c7d19b70d3d7cbfc33ff89ff6a5d8c916b4e787b724973179282c3cf63e43a87788f32673a25ed38eba9552ab6913564c9160f68b5e1aced85f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf464d1bf3624d132d5f2be0fd46083469fb74fb83e8491051b5463c27895e8d93bd9f51f17688fd27f1755eae6f17ff0bcfa95ee8a628a2e1d2eac5420b396ac63e2496a028655a4b86c49ad6a71;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h189c1d352d96e8fb4d4deffc08fb3093f1b20e5d8a931b363256a4dbc505631a4feef4afd3266df2fa7ba589cf162c9c2447bc618d3f4c87d59303a05782bf8084788c291297dd19804209105126;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1435e7679d8d5f8cab034b76cb200c4bf427ce8a34910bb290c08f744c386e28d991e20b6d05a6fc6555940c17e8dc603e9d7ad2f613da329c18a375a19ffeb8221fcc7fe22beaac95546f8470014;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h47fc817020ae56a81c5c9064b02c829c647bd367d979e1e7215a1c80b4b84febf94037c8394767d3e8735f82831e6edaceef88faaee80daad57c4a2af024538374a18f95bb7e8da9f9c6832d678e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h157350e929cca79b911b3e57be5a1b5557afde6d20dcc3b21c29f2ff428b2ff4ca5807742a60fdc3d8317bfb1a3ca5cecf868dc2fdf1d73c2c4f451244a30b7c7b28578a001c658aa7c76f6c7b4ce;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1561aaf75a027111c88beee93513de137a6fdd6d592a3e56ab067b064d4d4b5ac322073bf1901df541f3212918a6b85e5143110574a00797f912f010ed2b8d7bd748c0045d2661c041c494521f86c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h192f7e5f27e94c676b9a599e4bd643e836eef35a78996c15b152382c540aa177c3ade8c0c3a843b4f2d851eec4b45f0c4e57b77aacf8475df93102ceeb9b9dddf50c0e78dceb29582dceffb959bce;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h118e43ee54dd0493714928241b1d283626be06f3db841c62fa5df52c6687b8e2ed64c84a44b3ac2aad8d17301f5380c83209ba1e71bca7825ab6bf8181d665fc83175bd75e594cc90e9a19527f4e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ea0fe7c7a6f9bc61ac091baea950a43d59f8c689a503c939ffa47d5c7eef33d03241f01d6609badc23c8f54e5e3f1623cc9f29bbeb386dce94291009e3e76f57092da8129c92958206ac43de6a99;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h80a3fb6c1437a18d97943fb97602cfc6faebab4b6221e7edc405200faccd8c3b845e84ee7fca281d5cac719f56cfd68eb1dbf09b22b848e048b54cdb71127d768ade3f41c06772e60e55affa0eb1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4e1c2dad99d77dc811b11e79da098bc1e326ec7016536af18e9a43230a2ed093428a3bb550efc67b43943aecbde8879d9191dd5dc23aa562429eb783432016c054752eb71d69f8c1f180582917cb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heafc2f396556dd8a2d637598eaa6d4496ef88153cabc62db8acace4169d0fb39c3d86d29a29e036e6362c4a73a729a57bd89d57d2147fbe5b7cf12ec2a3a6ae92468833142ea7ac8e6bc3e522214;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8ab799a747d513d6dcdd90eb98474cb2135d1b1080c673c055afd23499fb9b54b76450c3d5df4f47433db0181b44a373dd5c770d11908286ccf1456d2e6a0c6258827a213eea11e72477e1610b97;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h92074fa43c0a10edab279cf2a5f355d32d05458573691122be6c43f9d1d5c50472124378930512f6b83eca82067ff433e4cce28c285c4d5850ad982bf3bdc2858c1ffe899723719240866bf90d4a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16df6c336e0ee66fa0db49915c87d436c6716bc184e29a86106907c4bc37e994613fb764687b7f8a110ae8b62abed7d8ef76589cc5ecf4528ee0ba2cc843881f1673f80728cdb15aa090d7317714d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h718994ca8d92e3531271eb68f51ca7151c3be45855b6e12d59b460568db4da79f232a458903dd39d1ff87cd459a038abceb8f6f80607a462d15c205ed22c16a4853d3d32f6cc578d78640557d6e4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h104f1b259ec7ad3cfe7a575f65dfa21687ce5c92075f84617d468a6d96249524d27a4c7d7b7fec121af658c2567649891f7059b2a3c042ad2b9adad5f3e901e86b2223f950ed220ce08b4204e32f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h161b9213a30c313316f5582633aa819dc0d4630f9333b7ad4ffe08ffea5ea59a2e03245065f1ef750be21fe756bf5e64f6fc47806930b511a9b6ac7623358602241ba29c5a3b71d5998b30fac9458;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h198dac96efa39b14f1686c5768e9dbbb7175aeea091f2e3c3806b606903f4e27ee5726740af622f33a7be84fa95253038442bb15813f9a775c5eea955831a86d2218d6ea64378c3187aba8d606e31;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h173fab2f8adca6ad6d2f76c4896890741dd8a739fc9b38bd2f0583ef7200c16a872ab1e4ca5c189bc2c4ca1ba1a077db28546e573b1c0f1bc4017930138be90e39fee9f3188b9855a1e91011ca296;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1febf8aea415ac266851b494ed6cf499c4a54d4c57a81eb3f3a6e0bf5ecfe5919c8713e8120c3aa51f57f8679096a45313bc941c57d3d0b8f5b77d6b86fd5a4f1c7c585af86380d415da10109c31d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eba7efc0027a04c1ae73a45d70496dc013fe6b14ad75b804455291c6e9de2602d6c6311a7029c10cdad8fe45cc5f279c9186e7124f7f7cbe3b4bb9272ddb225d20dbca165d6053b353df062a6c71;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16eb6b5a1efaabd153b4815fc220e20dd5019f547246eb09e9947d6909b81e9dfb9c5da260c74e7e94b0c698916846bd30c4908bd38cd4c917ea533a12b1de348a02eb83654127ff0312d820db543;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b39f31157413560c6121a7ed1bfcc478d9d9a2f77282a6926fc5bfd36df109fc16cf7a2c9ff94e8eee598c197a57e575de86ea14770edc7e136a6ea46528cf1f2df53b4fe6c4d75107cabd671e08;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h127d4912bd299db4c3e3701e0f2232c7d476da7da06d46a0e7dd0f022f0cc9583af501e97ea10626a837ef261ebfb912612715df44d24f56940c1a314ec806aded166f68e495910dd2821f3fbb5d9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h98a8cf824243e18ae17c70a7109b6454c4c7ba760fac100e9c68322ff2a14e5125b348d6579200753b3a182b0711610eb60010469542e08f80b6ac4ecaa9b83bab60dd03f282fd416a53554757fd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc388ab485672b90a2c28bcc204a37cfece268363caae6509b4e60203e3a96bd0c6d2c1fd3d1ad90cb8c25a0b3f5012eda41f37716dd7b8f5d116ef8a42d884307eecfd9d01d3149734b1b09efb25;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2eb6266253dd7913a78ef51b5d96f5385900117f4a5346c277ccd72af1756adeda9488a4d37faf84e266becb5254fce3656b47b4999eb63e14c534603c228e55f3b3c5a8f0d00f5daa4e17db8cdb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbd34a1c730604fe3149b52351e90c8dd227062c6670d873bbf31fcf7d071a0877ac1a8c8471166cf833301e966d11af9221a1b85a27af78e855883e20f3c435f0a66f03353d6fa60a41bcc7fe45;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10a7f49e10211f04513c2cdbd22d512add317b7e1d5a7d237e41a7543038a2fd4837fa796ff49913a6f59cfa46cac1016ad6d2683af27d3335b3ebf9a1ce1416c6b7acf4599e4d21546dfe7592fc1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb60a6572b409019d0c66680d3a48858df4d69a4fd2bb3bd8f89f890be6e979333ee315c3d9e19d51b531999dfba9ce3bd84e89d50b945fe807a979ad05e0bd0570fb1367574a4f57552b64cdab3c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19261ce36b93b97264be55e3229414e6174c9582bd7e4a902a9fc09b5730b65fb9fb980d93bb33a7d18118ff8ad22324e6f7f736dc78c8a07e22dac474e6907b7e1bab7f1d335b677beecb162c802;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10f748ff7396eb3b4884c72bed807709ed3bb84c268e225fef9a5ec144c9728ca508f30988666674da06460d3b54e47634f1cf8ed090a6f058961a88be06e6fa9c41f3bd4bba90cd7ea4b0937bee3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b6507375d8acc30d557192a335a2de1b6b5ef64750743e40f03a9ed6010f69e9558d0742dca4b767ba74aa168c8c0c9dfa246217006f6e328a4d7806f11caeef8b954a3bf765b4a9882ed05335a7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7f8a03115e87d4f805aa7b64dc0f8d9cb9dbbb1a7c152222abd8828316f98d828e48b246a3a313b22e4bc152b87182a41508cb97c43b9298fc459d8890ff811a41a2cfcc72ac397afea3917feb97;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18d3721662d24e670485a94abbc54b440ec60a14e83cb01245ade85772ce9f3831dde7525ea8084c75205eb04fdffe632483cb2c9d166888a767a003118db3114c408078e220b508c3b8596e7c09c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf404803fd6f81d07fb84b0241df19b74f032837f6e06bf44a847ce54f17af346c9628433a744db3b96e7724abc4282f64235a5d903d7075b4e725e071f93a9208cea880ff78b0087e3be868c31b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16bb990029634229cb99c7764d42f4ec79fd97aaf7985cd622b8b6848d95a2dfbfac7d412feb6676641cb2ed6818788a075950338ebcd8bfed072929bf7a06774cbefae295c57764ea4df288bf53a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdd1bc2a5fb1bbe55295cafa09849d58166ad39feb4a5def0ef686d2d71ff48dad62225411adc616c9fff119d075993b2f9a484f1836b8a2320d48f628451b037870c74a72f29efaeeae24ee22bd9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc9ad5c83cd005beebe7e9127ef049fe661d8c323c44001be65f94ecbe750c0fa62edccf310080e4aa7e99feda9b85bd65bc5d73a6ac3a8cf11b6caf7c47d9e3009fa3862d1964bb18812efe0192d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4103dbcfbe884cec5f878a46fc660f5e9706d756e92e73582426768b944272be552a48ef73b01d5fee662457576f4083f57c92b16919ddb8553b7a90a523eca12a003c711722c790b6f612905756;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h737e974a70bab23311627d0ed59c1de6a4f6f95adf29e49ffd691a6b772d6625b5c5e238860c6be5581c5ce13b995333c8efb109f96d887a420eb6bc8c75b232fd79a3c595332706853d975189eb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he936976a2d848d9edf144c974f86b7141809fef0b4d7ad57d0558988ac8cd3bdb3be7b094d626391987a7a641f53665aafe2057421f8eb1ec31396f7822211aced43b08ffc7cc711dd8447c43598;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1043fb673b3ebf5f4800a6626d01928d4d57821f19291a6f175ae1befa1be77e9fd0f8216d7c731234a7c7c54799732e28554370464555b14820043a1a3bc20e1db6a9d85bc2591d5fe675088ad48;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4ce78498031665e6f038c75a730e687175b8d1874cc6de18f3544c76ceab1accbb6b180c725b766e2a7a91b5632b2cb37d1fb09d086e27016e83a7e8f0fb0a967dcff4c3f5070769ae015d48c373;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12285e2e2845aeca363cdad8cf5d8d2508732286efa345181d110cbd6f4b8937ab2fe903af6ba2ed73286b95388f7dd3cd443cc10f27694406ac7a7fb564523200cd408fb4689fecb7b4e9bf28043;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf9a1ef0bb8b4be057e24486bdc14f8e5de5cc433e178ec8b2b2aa2ccefd060428ba5611420ab1d00c0079197ce1ba46f6b1e75d2358558adda376c379831f4f62fe74f67e608adbf2fafda709b87;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h648ffbe5907ba52812e8ebd634fd7918b8e713e1f8c51cf0527ad39bc5edb633066b74b787f322af42b17b03a6252338859e34149001cc9761b92b70ef5f170e2ce37ad32c352092bc04d9c7e5de;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fde2587951293c204303abefcb039034405c40cf3b02e3e614322368b47c1debcdcdb242d02fc96c474bd5f1e5ae75f8d57dc1e2943bfef74ebf9af1c3a04fd92c50df9fda11ba4f4665a645b7cf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd66fc0343e86d8f247b309a592a9911f765f10b5d70497231513a626e1394221f8fc17a8bea57af5174b3e04036a7de72094090010415dec36d6d031045a7e023a856a38404524e95500471cfd5d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdd2ba4a8dffaa8b734e3f103ed3d28052ddce3b112073038175bc037800a1a0c4f4d461d1daddbf22829bc91c16f72060dceb6460277397bd21742abba593024e8bed7ab9fd2ebdca51b990838ec;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5fee5ff1682d939c12d610a5c0d8e1c8a04249302c5f549a7ff003216ecc260c5827840aa48f180f1c17e11a4296bc1ac55b675789451ad6bb4c7dc65eb0c656e3b76d8779622d3b68139aaed3f3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f14875982d4d3fb3832683622a7a2464764dcffc8b106ebb00edb2fc5d3b78943020791d3ff7257fd3ddab3c58d36db48d237431e1281b226b1070814023dc0f97c801f33ce316d95bb528d79192;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19a78aa5be35a04e1bd258c28b046aba24e98b7455699dee56b5b010856b87bdcd3054f958616ba7ff0b236c0854d3a2d846a8d79a063da1dfc2d75681d395732a2828db41dc8cf921d781f83e01b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10bed6454b2e91c037330476ed988a10ab308ee2f6c242cf432bf742ac0c0da032e74834e90be35de2f8a92e5a7345391ac506fece1cca3ac97bc8b630138d49a0d4d746af57c82b47f352467af88;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h177cefcd57365aaa6b433cc86414b2cd9daf35fc149afb6d7b731768aa6aa388a63a9199d42db8ea89131b3c43adffd4e031c037134f6dbf1d47f6a5b89a67f653061ad41b53f48fb15e2b2e6101d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c14b3bb7ceeb59550e06fff1e7d2588d2f705b7cc1236bb0f44b71515eed7b755a302affcef45bd8e1fae838294e144758655fba50c92278a625b79e69b8d343a1d459d2a6cd429258636eec8cf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5bd655bfb23db39926dc241ce232289b8fa2b2c90d62fa305dc21508ca9d46c12afd9df997e2e4467fa5c80e7cf1a8446f4844ab5385d386caafd23005b4091e468670db424639f373b1bd334a66;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ecefa039c345625d345889c90b57a06b7a54611a9c675c7794f8cb7e327cd1dbf665247c6f0590814ea120e7b77b3d4265d33f93643b64fad9dd041f70e88bb6df404e54ed8effa8d27f042ba397;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c5cc6d49dc06369d11f0e1f6e80aa899f3862026aff16a7cefb7ec1f7749d7c48e0df57f3d29faccdc6db3b54e8f37f49f937b712cdd354a55f05966fcc9486557ea24da879591563b470359fce2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ff58272b9e46396c421a6992d6b0d6ede93e578f43d1161859595bf96de6e92e0248c91f620249ca83d6758b8317a9281772da6c478632c65f3cf490347f5fb6836b8a5da417a0fd221718c8c19e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hddf8635e8f7b3db83319b38b987f6844983e0c9e3915c8b97dddd23c338bcd82a52afebd53ed0dd6b1382fdbff526d858a7c4729517d1fe7817a94cf33b8e8a64a08164328ec06248183fee3f03f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdcae7d5b36112422bb958ef642829c5494ff0fc09e0ea16bd527bdec7a53ee3749e9639660463135cc1f7350e59e4b86f4ed0a2bc7dc82645b639f608e4af13d1400d073db7af8cd55dc625216e8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h28af2f87188e59e1c6cfe8099b5ffc8e6abc837e67cef1f6e86685ac08c5bae8ff796690635f14a39a631be34f4868266511dc6cb42f3426fdebd9f8484e0ffc20aac3e6f3636630af5fdb6f80f3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16e3439f353a4034315bb1e540bb69a8662e99cc48d27f17e996608dbc5a5c2a5ad41afca34ccf73d9f9939ac7b9c59edd9c2149e33f71037f5bcbb2713e096d65cf4e460b7b53106b74f53833313;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h576f28e4a3053a0b07fcb6703ae8d68d87e60d7f9f5bb402b8855e597e57bcd2e287d88aaf30fada0d8557df333c205841fcaf7ca332d06503a85d56eee6215f9d399169c3cd15fde89877aae715;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15c7f058ec0830a3b3b804e40787fa0287378711baa064bd789352f801a20ac45b6ef1d0d5641d877dbb5c27a301f88da3b5577555323ad09818cefcebeb5b794b72ed5ee5521d6af0bc526774cbb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bc5c355794565d3477404e37d766ca5dc0d92b2f793218179535dee4839e568a74360d9b392ac8ea16ea27d1bd66d35471008b67156f9ce9cc21ab7072f6c6b1afc736b1a0afc3b76f4ba556c4c8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdd8413913fa27c5027cb57ab2b0a384eb2efa33585a3688e76f3b07d86ae2e30d6fb37f6bb6aee44eae43e64034c12be4683d2d1959124d27654af4ec50f475a8fcf3a64c3e0a5a8ac1fb5b786c7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11395ac0c72b0dcf0951d121f9986c36d570dc75b3b0359f951051f2a947387184807673521a4d6d2078b0c534f3c724edac7818f5688c5f43ef5c13b718031cc67d3f6fef8880779e92025a6ead4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f07dd8cf215e7fb53deaa7a8ce4bca9e579d0e4329ef04b7d9c55078fed613d2bd2162b997d544a169888cb89ed01363ae006264dbf6e2bf1dbd40484130d00973ea5e69eaed9d1c50b6909ef46b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10ca3ad406b3bb0865d2c550f8b5566cff0f6c2614f898a6e40947ceb5095adc026f5a7669a04800eac9d0ea052394e451aa15346e10d281c21197f8f8c6329a456866b943f64a9b9f75e7e5e756b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha719c7dd1b146e261f8238d5768a5a58e337da0bc5b1d2fd81d19cf94bc41e7fbf96d1ed58118e29e79cfedb82f6c02ab28d7fc3d535906b7c31ac6125db5bddad54828789348202613e4b3b55e6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fb4f95c3c20430b2a03efd5d7417497faca400f73fc6ecd2c3e06e671a67857a4e062f0750c2b4b000cbcc5d3bb63294a0c68168342507e9a27281a6ef433196402a3e92f1dfb3e6e41b1492fc65;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hec024a5f338e5d10d9566724bf9231e0dc74055ee8c93c246f87a9a24af463531eb535589ee71e181a921fd55f4f813eff79f527e5bc7b828fb898cb16a8689cb7c6246d07b150d886c29735609e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h196ec2cc81e2962184c0668db624b28bb189ee008cb5445cfd120c60797967ca2a43b718d7320fb6276335209bb9cd2b676f73f8e775a1dec546b5ed2d580fd5783649ed62da5512f348816145a8a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b36a8cae778137b869d10dac3c24e292f975d2fc56deb47d4112443290436d0fbcbc834c29fe73f558e2c3d3a6c175abb726b97d392ad9e75cb6ee27f7c23d5c8759846f8ecdca97627c3813d4cc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h548cea857d2d516acea2b16260522f38c9c6ab112c6884379493bdaa663d5151fc854df7db0bf247a0596716ef5b0b9eff6d15dbe4cf3dbdbbf1eff6b5517921293d0a1318ac8b2cf5da400058c4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d341023cce0d6cbd93adc26894ab629f42816bcea1dbba22190373e54a88c680249ae1f3d533a12b294806adfbfbc92721fd82a22b2396944b6da846e140fdde67df7cf1b048620701773de9154c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc8f00df26139d7fdfba53d957563ed20f5384b8bba92c9e9ceb71f1f553dac2bf7dd458bb7846ba80bbb2eedb7623ecc2f40bb19a085570eb1a40272e2542745a5607ec6d9ae91385054f3e0d542;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d8738fef7b5316076d8681f60b246da88a3fb2f9a4de32a3a02fa3d41dda3b14b7e00b263c07fc24f718480b9c9f9e32c678b29e202176cff10b9f3d89f538d923f1f1a0841ec15552203e9b1195;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha09f27290e451f199815c10d33d4424a5ab11fb5f02b12fb632913bbcf008cca3f4a59f622b55f7b443e8342fefaa0828fadb79e91fa084f77cd599ccdb5ac0247c29a3c4d5b4347becb95ff28bd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18704921355c26707c1b109d4f841dace80c67b466e93681348d7c647ae807111d7b11eedb9c5d85aee0181300c4cd4c9300c11e769a5e095ec5bda76f4cd4fb6440494ab8ad17c918dfb359f7f9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10f67ab16c8bdf165dc9f879a1e1515e126143c7c8698dd200ef0d6e2aac9699f1283bf24aba73eed787e83b6ba6b5047972db23aa18dcd46852d452c7ea56253ecc9b139aa93418316512a696197;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18af81555b41f99d6001a54cd7c9815ca528b4acd6731b97ccdd53fba2abb754c034bb8f6d7ad21a3e8aea2d0d5a58b70fe802b3cb373fe3989e68361a9de3f177d95f1ce489b6511c265c733a1bf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a2f4789b05a672c768932830b17f4c218665b98735b12c951587612ad800c47a1d5db1ca2e424b1222d2e2c0436cb53bb0c39a73d1739e57f5fcdc2214f046b339fb2c17af9af5be18206c141cd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17e047b050f57d677f3067c0c42bfc738e2be8c549817ed01d4e2ca69c6c26b4993e0708edf2b54bfddfe65b6ab8b13da0470e9737eba8faaca2cac36dead162ef492e2d090e1ffb5a3af833d7cb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h149f56ae5da5aed5c0ac0ba26c47396f0cc794a7fb8f2d45eb6dbb89c49e022f3c0dd09d5e2c70cacac96c68184ccc9539f4a8de7c9294384f35a08d53a079e8bd1351e6446ecd6fdd51bc638f7fb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h57dc843cce325452d16a1b652762a533ec7ebc5d85261f9624535a27477e8fe3c2b6148fb1fd174b772d31e35bd5b53bd1e25ee401afa3f4d8e60b94773e2e086461ff3a1feb006271c03db33401;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c4784db94f6ecf2dc55a933c6b3ee297997b498f3af7a445a7d7319f79b002969de8986d45d690023d462191bb78821a80d42251690ea49d68716c1e5fdf7287fe29654446d2168b8d0ad7fd21a6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h37a36ca6ae4a31dce47d5ffc9416341f2e155a2bbb22646c1a2d639f379cfae7a7e7a8f73dd9b0ab1fb6b5a94dd60c53c18a73d4a35dfa449c55c90ef8a17dec8752e7108b4c6d6d7c1b4ed329ba;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6ca62e01ccd97073cecd1b5c96343bda440640abf64c7f869b8858ccf80c3dc5cef39f87db5c15c9fc8d8c8116c2164e4f23fc051f2a85213e8d2a83602ed25cefa047d6764d6e88a6d97064c1a2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3f13b02a4a72736c2160779db2385c9dab3efebb7d8620830fc5e57c4cf252b5d911715e730922b8911e3aecae6bec39a884ac3f2ec374c7b530b0c0ba9984bcc303d38f5c02ab79687c4214b041;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1849cd2e0a42c5ec2b6faf1b215960715c110f13f86fe7469592251a12472246b40a0c7b16f9c3416bd6c4e0a653e3da1f0a445a7a2cc61b2523526a0c944359d670678e53b542583b482defa3047;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b26d0ccec8df92545baf79fa2847e5ec081685164d543243ed452e8f2ae8cbeef8c1dc0015a872c40e3b4b11a84880cdaf630e53f762bdb2869ec792cb17604cf4bca9dc081cff01d2303b9ac991;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14d36e689dc495503ccb99b2d1d0fc502dec2bb585dcbcb583c11a2768a4f4379445d0d489a149d6ba497a6a4ab8abe1caf837ec4d0ca8cc253e0b05926081f290c611ab8f467f4bb5e6b5b83181;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h394fdd410c4f0c5257ebee02bc4fbb61db50bb4b64bb6ca5359f96c57f7caa244e411eab7a750c3f04c7e0385e767e9a48285701e3840f412dcee2e298fad2ea8aa6faff6bf7f2040fe19675ad29;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7ce661d2cc79bb4baa05a47c1502b204d2837d5747258ba1355f75ec7043465c692d782f1a50b4968c0ffc0cc6771302888f91b81dbc609564f96a4ecaa58fa668dfb54e6344ff8c10f7c978f458;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11af7adadc024dbbfb2de52e0b5948bd5e6ea9401d1c01fc579d58b357c3ea0712771bc1a3e49146c11a859bf68b9ae29a970aee8c7d08c188817725106e9df0fd3c8b3cc0758c930810137478a07;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd023a46fc424d971d8cc6a82fff5a60b73c924277d5033b76bb257fbb52e0f0964be45aef293963bc606f9672a415bf9b7e86e5fe76ed7f8e19ee875a45f42a4f7f14c1e0a383362eb05ae5b4559;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h147e9b73b1bc748f177314c268be560bb836148919cbd15b7dd32e0b4d43ead2dcd939b0329bb98583a455fd37a152672286b016465f222b3f9b1685904d9c3e97f6b75629c9bb14fdc9e73438828;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18e9f8cb7140ad10b5916ac1a2cefc10974360019fb1d4736222079dc3f574c743a54d6050d6a0d6edcc795ca7235bda8d835262cd7b6415981ec1d5331f599c84b032d6315d878a6570956b5a492;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he3687e2547800c4c5890f8bb16ac64bfabfb030dda3b170d8642d43c1cf6d96dd31e2e5bd6a17db8fc7018b8d8eb0d32f6e8cdd8f28b9e36ef9c552483d1486fec9046ad2be6ccaed2275c3c9818;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12570a9b895e4661f1a195662736e863c26ee91ea1b91f573422320ecabd0b501e19cc812f902cc3726aa050215f6196408a57e6c84b7111050d132c3abec2cf79a6a4a41c01273c78db4eee45b07;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hed5a05a5551a9c22b0e225c1eec227062d2f5d768d809f17df55d7b166a90484ec4f48b62a00dc6aafe09e3eb7c13667f84fc6b2509cd4dae232fdcf27609048472b087b6acaeffe5c6e4ff1b508;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7517eae9500ed6abb07436494fa2d0a9a0e65ddfb9ffbb37c3b39370d14f677aa5441ee0247ebcd6e29c8eada503017ac3d3fd2fa073acb52452ec018b8f38178d7327233417f9740a7b2487fdac;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc91c5e61e3d3b2e941db0dc37fdcb9ccd3fb0f78fc6cee592191ab1d79b5b83a3d536e4e2c36bbb3e46dadc8dd8894c367ea013c11801274200e92bfa866041347063fd0200078e02117a10c6758;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a59f0859d6fe9c2bfe5f2e7ab557ac026e8228f42d1466c7f99840e84cf4e6ec6b8abd09f77861751fc1f09520f6c99a7373e8d2c6dc0b2dac7f810c441a702c0d56b94ec8b8807f13eb7a6699ee;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1de06f45069cdcaf1a34365f8b052f826323a3eec141905940ce46861b524c55b1e618ae2f3a4f8840ba14acd0f2ec14fe77cd33372023a52c867e3cbb2bdd8e6e4e471ea9cfe489f078b133056aa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6e580c1b1b42123038f0dbd5d55affa2332b2c23e3ca00e30779f4fe5f062df8d07aa89bc7f91721fd8e05a17795ed371186c0dcae779e248d1537a3ef7976c7a06ada3317bfa3d90efab2dd80bc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15dba64842e9136a10581ab1308c08ee9af1a0f49ffd577033b415439c85ec512aef9445d2b1ed0f616beed8d1f69bae5bff10c4edfcd50086ec82ef2573daf53f00f4d58ebdb85c0df1bec7db56d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h183f0d62558bde78a2724b5c820830a52b3e875c0aa4ba09dfb8b2e088a9a306429b7c7d4a054bfcd3bc1834c1936c41f2b975132ed08a2d138168fea45dfd6f04bf2ca74111b65cf0465c000b019;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h63fa8acab7ca651cd91b9a88fe9f5563324ce3666798cd3220cbb4c07f46829794ef3548618af006308b91a2a85ab3f546cc3573cb4e5b9e1e00e0e6284d2fc5946dbc0add2d46292c5e575e5c03;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd9be4dd38cfd199cebc97af6b1e7b4e426966a82827f9bbf921364d9945bcd8fe2151707a4eaed7aede43d778c13f46fef25a4e93bb78fcba7f3265912330da91859240fd060ed3af60ed08b5937;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2881c054f8e052b984a90f50be93e4cc99c662378eb53befcc758d1dab5e620453e4941fab5440f71cf45d90b61fa5683bc5459563397111c7e26aeb366bfc797fa1ce37cf832b14cb8042a37828;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17129ce96d2ab97658af0f1bbcf5adc8d4c8256d5a72fcbbc2055035b1c3cf7b95f42454c38175f9afbf9a25bf5ea6f0fa8bd9755c7391f3f6bf2023e6a12a9d405818199d84004940b0a018c02bc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h60e2ea7726569e04d577d4d87b62b0da3c3b39830f140d9f3109abe953b699934e1e0010956bcd357ccbc8e325fc2f7dc2e38fcabee382b858c5ccb7088ac84a34659071ae315c19a5fe38563399;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha3a360da970503be4d94f7c84407b534844446061be7ec7228f57fcb84fbc79b16f5e388312ca0bc3a62cac71d01a10c2887a2d309f38b7b3adab04c21f25fc85cc4a9ca9d812034ec0b7fa96ace;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6b74ef58929bdb627816cf74fb97835aa312da8a05751cdbccbad7ee47a29c6363705dea41f4c4572c92037b1467c96d965021300a88b186f7f46ffa04f10a3463a2f7b31702b78eaa9fd8dbd1b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h932ac85301c81c35b2420ef88fa2c0eaa0f2596343255902d5313bb103ebf4dd4ae43bd4c0f8ab81789d32b47f1f2650b4ee96dfd1ff635ab8b057e26eee118ca067486ccb2a4be872feb4570f94;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h86c3215461a48b921bf64ce4bd50f518598f4dc82a66551b598ff95e93980a762abc3411e62d44eeba3ac5e8084698cf725b2da4c0911777fab508016bf32d6903683866c22e31dcfd5d46eae53c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha141f616398162de5d384b04ed53dc23124db6bedf9002ca0233ef9676108d8740dc45ef14b2294c43bfa4facd4651db702faba39ce0df4cf26129ef1043a32fedbcc689793f444352fad2b3ccb5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d14ab4e253f20aa97c5826e857dceffbad83c6a6684772dc99428a0c275b8f577482cf8f4d58c3b248c5cf18949d58664ac80ec7a0d3eab07536a5cd45d1260392985fa71717f046ae96f3753e23;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13b04e6153c59f58b2d532510bc62b2e46d613f2e3bdd0726b4e276b0e1203395182235aadae24b71ff7163e7fbd1c1cc2f1622bfc2218672829cebb1a8f7ba71206f5ca58ddff836305482d950b8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16f6e467b64707ab515d28ddc0d9a8c1cfb77757702360813deae4defbda005b716a25e52c4ee3653ce57e53fbb115d7d22c1a7d8110e028370030113f2aa83a989e54315aa9fe03a6090d7662c27;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1637f951e79b343ad645d9ec5638b622753e43f29808be303a5d1dac8a6bb4d4aefe40c060c4c23a2f249bd0debd366adf31708e5ba21847d0631205ba6ea201fd2f3bea1ded544e8af22e9a0b96f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h63180d2a46e07c022521bf340157a85c79bfc32f87ce657a6f4984a72a5383742788107c441a904ca5b9bcb60144bd61449e45e171c292859622d4a8fa4bf52ce2e2d1c7607351b015078f152208;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13863ba336ef5e42d0db5c9308ec9146b00b023223b74bb0b62c0333758ff63a727514e2939d6137dbbfc6c8ce37835f382d64327e0330ca97a285ac3c183e35c1cfc25c486aa7d089912d1363199;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8d8ac03779c5a6715133bf69740fd3eb6d2002738bda7c5f76befde228f83deb42bb1612bc257344e614edce6a4ca89c0c3014b32f58499c606330c658809c6bfa9809e723d58dd69696cb8fdad2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3a17d190ec46556401c2b0727d68149815b21d4c7d3ce1f720ab3b75f73d711437ad3f468d0cdbcb29669863916491792d7c987463ec012b5f85e452ba4f47cc5f20aa1058e7df3e53fd56174f47;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haf6e19361149140458201f09a26c4945108b426fc55b52aa0901eb8bbf271c190acd911266a6be7787abf78dfb4057b0a5917c30f5d64b99e9b29e8ab2ba0b77d818400a8935b62494c4d6754487;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ead0a438d2ce9ed2e1db9652d5da68f4bb1527c7df3e521f2592f52ed53f03837d4ecef4bf2b1c23a043df1d3b167b5823bcaf56f1f68c89fa2f7b25aafa5b38375e0f42f764ac65960da8d6196;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7b5e2b409a9170f4c7a3d9be5864454ab81a2dbc455fd5c8853a1b402eae4eacbd67504cbb2388850a91284efa66d9937d9195991e05675b4ce2bba40941557f2f1d7da12d65c94a54039fa9c7ca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c48f2c91faeaaa39ac40b121fee56201cfb198ff06bbaf30e9d1055ef4a755881c7b40445fb20f97d33cb98e40fac1cc039147d4eee879cb63d356144fa3ef9d2b6d51a38a295a7e6b3e4a7b603;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h70c20bd4982aaaf1abc3ae23fc58e145b2f52abc231b986bd393199ab08ec327c81dff989144cb679a6350fb1e08c9647e90d49d438e99ea079df7fc44bafdda5ecf26a941f424cf5af72637bfe9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h175eebaeb2506f67844880b8a6495d647155eae0a32c3cbafdf19dda09d13508c610e0514f3cb9da825f49b45a0488c6c9819e23d4009ad8d92d6302e8121e8772175d6879984f1f4838a5a6c7c84;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12905a57b7a398995bc9c4f1c69631b7d522e3ea0c4092dc5659daa281061704ab8482a2d7aa651a397f68b266a3acbee7a3839634b3eae8eafe9276b911e371b90902947918debbc57a3e77214a9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6ea9424813158e72e762ea740bee7dd47a0bd0e2260164cbcd7bc63fb35d80a07ea1ff09084197f54538296ee697707a5321440b2dc50ed4e78978abd71e04d9d6d0f4ee6abc084b845b325a8cc5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdb8de93fa6857b3fd40ad1973efedc9dd17429de9ee3d2dc12217757adc97746fc7a8130cbeb8573fe67ec497bf583cd67018e2a5a83ff7874742bde27513eddae62b65732a6557136ba6653ae49;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18dce2071a424efca8adbde937802a1a87d1a4bcfc599515fbc7346418fe1562000101db8c56cb03da096e5c1ae7d680494e1aa40a00d3d98ad41636b66dec7eb76eb3e676a03a086b9f52128b82b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16b1cbf85f62e315155743f09791f6735b72e748ab3c8c4bddae5cc97cfd910412c6f6ece1f5c020a98cc78bcd377086d8179d25b3bc24e712529d075caf27e99c1ae0a4831210e57ae31c7e54649;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16b6331ef176cff628a3d76767d2baa884ac500699111d705fcf822a0d5fb92b8c5be54279cb9c19d4a87649a798ed56c63367394d8f03d802fa6a1b51eb5387c925c305af16e9bb0485c263d7ef6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a007da149f5e75ba58000997aa336711f71989911ff40dad0d0b0f511a38513b8a65d42ef63d8fd357dd7114acec724949bae21fc909a0c0ee7f760cb76e29781c79ea5cc7cfcfcc33ab232e165f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3c8f795ae2503ef95674cdfea3c1a795be0879a9f59c13f5417a9073cc3033b6b12c876c4d12aae6a4fd165b3c7216dd9cc1f63dfe879a4192296912759b5396e75aaaaccc286c2a1131dd8b9802;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5e5956a4ea97d6b43691514d5420610c10ec63d5357d941a17a8657d3fd9e53c28f9b34e0831777e701a6df6c645284910d62d5aab5774d7319a74822ee530b7a72f931462d6215a8f1ebc773b07;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h37830ffa795299cb09bfede215bb56a2e300b2fbfc7953911241270b178e7c28c2388d448b677538ffdcb54ab348f72cec95ccd831c2c3063d63edd7a2766c3059c7292bba24c4264215e5f5b79b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcccef658f05afb2bdf8e33d2bc2e329729ffa1f82649d874ec1838fa6c75d8396b9c26d9d612d264d7ac9d29d75fdd7387fa255ce9b9a821243651b0c64ad693ea9d7e49f5919104a587e7cccc3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1286861d3a7d97c88df088da345693c06c47a6e968f9f1d1369d20901653225e29fbdeeeb8f3e6a818356d0501491d1d682229ec22b376c0ae15357ce0675d515dc6eace86fd42ee850b6b4379bd2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h282f3cfeaf4a810778a3911d3b82ea853e0e66f59431d2be728afe4c442f1dfd92ea5191e342063925f908e2ee0fc9c18c9dedc3be1deccd86a24316f7e6ec6618c680a73dfbaefb0ef2c69dccf5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3bdb013ca02fcfed5d14f0d3d236ed93aec6c79f4b46bd635ef14d6903ab1ff0b2ea0b77c68d1dbb5c6fa7f6f63100a3dc15ccb79ca0360482739bb961bfa1e373d5ad040111e4d5a4ddab57c421;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h56d702b7e5192a787d7f04c6e6bc7d75764a25293941e194e7e865fc81e1b03f5fad879590555dcc0f7a761741e6ff48e636a0b2a7f3b4db99f651704a14ace5a5f4ac5c33ccebabeb971595a855;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdfa82025299cee8ca8d81d92b4426aa2ddd58eb93e3aa2e3f40c6270044e5f55df26609968cd3ca92c8ae05831da973191e2e507c42d48152ef98a0fea58abebfdc5e9c32fa48bf1cb97a0af3c14;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e35efa6e9bd09d33747e76d94774e098f31a0e8698f7d7bc3fe6fe7be9fa870bcbf53fdea06a192b4f9c072398f032b89b506cd0e55d8592a1a8cc3c7017fa6b24b584ba9fb51eaef5ade9afadba;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16d012eed3a586d251a461a84e8179b080674ba58648fc84c774495103cda7e79808e585dee12229a47ee583218342e8510fad56b50cf35b1c6a1a284ee390bcb32849e0d67840c05d2018369e749;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1302c6dc4b4af858aec3ca1bbde5575928bdc70ca630fb85c5d41faf0e979287491002c9dd4284c96e4dfbc6be86c11552a2178fdbf735af1c686c4747febf187ed5e19a70dae8863d7dcbc6e380f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1952d9e4ad2ce98ced35fb56b3d5e62b2bdd7dc7ba609a337cbd3cb3c506e90b7d957231fac4afbd6b6274af5be36b9fcdadf62c07a58be53bfff4beeedfa5bc9cf5ced448ecb223bc41b7116cfac;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h121465a2a0659c548783be2927b924ff69f622c1e41075132df8c5148d194e6828a1897e89f96a0ab1e8b760c9e5b31248952114ea306dd71c70d1ab9dd18bb0d89f60176cb2f4d52dccc9a602daa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18019aae3ea06a4412ffb25d2cfc63de2aa6dbbbefd3465e98ac4fda580c9aee4f5cf0880a02e4cff33546c0db48884344f9a0d97765e75e1110989398efa1cd82f210578f4275955f62d80c7f9c9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2012bcf19978cc6446c38c64a8876160ce35873aa1cb5f47a1cbe84f419b8fe107e8cafe0a6e56bd436a489fb5909de1c9d9e36963786ad17720fce512f1d10370a39330b585103a0eed876d92d1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6337ecfb9c17ead39d10dbbdd8d0e41e0724208c93902971fe71c8912fab8a48685e00e78fdb2bca120e5c6f61fc2707935dbeb289b6414e02f17d137b17ca54215a88d3240d777d8dd3f1931bb9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14bda66c0d761347c73e5d6809be92691fd46089d73e045f28ac59e05dda326150f6b3f855455749e528e80cf6b9d147ee0cfea4b0334e93eebf7a9528643c766f4e71f70ca10fcdc9a16f0017f82;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hda2c4dfc5958f70ac6e4a1bcc98bb9264dc28f62fd9188ddd3b39834fa02c4f1605b40c5c505aae425f5cb415d8942ae17808721e69136eeae53f69ed6fafb54db5db94b48fe22b9cdf2152e4971;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hddaa0d41225e087b3009a2bf2844308e72ed64e247ca01c2810194a983590cb0e821880c140dcc5059e2f1e9f0b7f28180f41c0b1d699bc50057ff480c8c9326d4e265d05af27e60adfbe29de991;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d5da7729da6dba41dc0b6d4a7a048f17f994cac69261f9e2371931993c25b29d98b65b74bc2b4f49bbacd9b3b34932055d3ab0fc76e47561daa07f58a830fea836102da01dbe3c5a33d334914a4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b15d6da548d8f148f52daeaca19ca8bbb3f041e0058fc15e6d0f0b59a10f678db9fb334271f48259212cd2d6edd13f8d407d59ec37b8b7e4804abf0b369e06b2449dc8c0b118349d624c083bfa1e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16e2b894a80c3f88b676a91c10b11f377aacaa2e2d555c3ff90bcef01031057c6c3f9af0478d1d2abed3e6ee5ce5c14fd36f583adda0a2c4cddad5b4e2f3d2fa78cb7fb39b68f4d2b2abdb37719d3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15873b24f0b40060a8728fd9fde8b736c7dc6df3acd5db19dc9c1121eaa15d1fd6154b5f6548b2a4d293def99c1c5de98bdd5c8b36026275478090e907f5f7fa3a0fe4f76ec49e8c7a5d77a9146ec;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10262aa324ebd58e20247ab1e04602b436eca2209eef34a8b817092cc1a44e3ac47c84f2e420f5bec5262fa3fc35f75874b50cd6f38c3b75340281f55f8e93ebfb42c45cf9fcdaec2c961c1f38b42;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haaa422962cb6127ad6773a6df1201b5250875b42e712685b8b5fd89fb5d5e65a45510cef52c5d8a8dbf43795b978bb9ab3d63278f85d43d34cd6140e22b8887f83143e418e4a5b1edf88c858def8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h28c2ebc2bb25fbd6bcdd9f982477b7cd7da8f863e47cdaff9ace11ae907a351493fa67299c7813aa88bd3398705b5e8c446b03122a38f0bb6cee06184c7f5f757c081590f295b1a89f5cbf994574;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h118ae23962be5420b4498ad550781d5b2e372dc043a30a3590790f4346dfdb934b3575b8a800598df8046991f7ca93463ee35c0b3c94d32499ae5a0a4da8ee19a51738dbd512a82951a1a90b8bee0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc844756b23793f6edaa12c59bf3c2aa936f541c683faec0c37e16222dc808cfee421bbae379f756778d9c25f5141020edebc17a68d4b650782e9163b8a436dbf7d178661e8fc42ce2e0d6b4be259;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18049cbf3b75a15740726826120eccd3b32cb7f50701016441e19594bbc3c318ba750e5ddf1336dd6fc91fc782b70c053c67d4f1530199b8b76cac67979594c4530dcdafc0294f69915efb265e824;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a95019ba1e0f63edc295efdceebf987facf39d2c5cc81f003f3f305f604c3b3880346ed3a9a7ce72e1f15f05a2a18379e3f13c7fe0c4162d9f60e4c2b7605d6ce05d2d667acaa7cb2d5a151bdb25;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h102ee806e1e86d32397fd690a3b02f2235c07d75df21522e319bcf6e4878df72920bf2768c048a226b06d4aa6656b5f45b730408c5f79ea54bb471dd28aeb62781ef7bcedd59c2bb2f86976f6dfb4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17b99817fcfe550a51bb6eac52f2468e9294094bda794feda679958c21056bf2174942465dcd093b391b88e47b953357967222f0b12c4e39a86a3fa135bc39db32703f3d1195e5da5d978d188d7ad;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h191f2cba9169b979ad15b11816ba5eead0b3fd5ab2d6e4e6ed0962964dc282c92807a49b649660a4558ae484b01d6154886672d24c7dda9b3afcd8f922ecc043c78b12105cc34e4493aece016752e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1be75115acdaf68aec5ef8d3a7a36f4e8665cf875f4e45be984df2cdf4d2d30d474de2b4772ca06b67d3c845da57add3d56a2edc7329de11f5b04a9431fbba96ea39490db966b6dbf9f9fb4434fdc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12d5a715699a071801f6ca41d3142319aa718eb9e1d3dae38d4e5e3db4d3c8cd88284fc8861e38b57c3dd92593952b112b9c2f000c032ff5d57dcdd395eb292da7827a428a5da5941e04c478e902f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he32b6430612bb7269bcd51d2a888c73eafd36d87ad42cfcc426a88ef280e929c1017c4104374599145464832640296a2b88d98b4e0813307f091f11257908682b06ffe1ad6367ad7365a4ae28a84;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h95d855b222f9dad906d7854b8993413af5cb3c9b18050c4d9b5ab47d5ba96512a2a6e7c50cb8d867d2e2d47f2bae5e8ec52786e88c4af213578dbe38e126e40e4e7f2d44bee493c24076d7f3623a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h124c45645e31c1d5f1c3c830012c7f1749d253b5f19fee3ee78d0468a26c107104fc23925eac863c079b47521a868ea14bcd695f7b9a36290cd557a28bbbccea7e71f8166f69af03c5eef47f7ea22;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h99efdcb345dff8a66549c2bd2c430dcc3b4f5784aef65e72e131eaa901672188814f57973d224842a66340bc6e4c528029ec1ea7680c69441e5392dead54a426caf66232be54e2cf49d258c31d6a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha0d9832741b71ec4d901d28129989deb22bd5c1448750e3f51114e50179319b4b86826b8e1980993425159507355f14b539ae7f7effad4fd7f4917a765dffdd04e5cd612adbeae7af6dcc2e1781c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18ad6ade38a1d83e13db4908fa353eef25b0e72e22be21a012c358446703bb75b14a80806862c8723bb35c69f1ee0d73d22ace247114b1bb904b046336d720d8f93d3b7f045866bdbbeb5e386f7e4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18cd26a3d8eb9c6909188c47c6e671364920940530ac980d3d49de4aaaf40a94d415f834a1908b404332c3c4535b561a99d48db8715fc26efa16e10acc3e4870d4a89d55fa0874d688242f09f1974;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13fa3deb397be8be4a276af3a4b4be7ca1035154243e1753a8f22c3dc64839c7c2c4c80fb4b9609db07838c04529c310454330c7ab48ce561668eb209a3a567cf3137d075102486ad49eea4b3d5ee;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11b17c4b2a18162f00d10ac82a45900e9db6e326f0a927973a00df1bf1569fe729b99640c183b82bf7a6aef76d4011c021d45b2b5532d48bb8f430ffbddc144ff6de18fd683a99583e8af607cea39;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1218aaee378adaf44be5757613bfbf669dda94d4a6a9fff3c5b9c033e0f1d77e60d3df2a343bf5940509e296a74e9616e7c0114d408772542d24be9427399a4b294887d0cdca5da526fcddcbcf70a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd089966475f8a627a25ff80bfc646b9792db9c2c9d0ad3620205c3f7cecdf1799a01af9e49dd087b513f7cfd42656de65cd256133630218ad0bad5f6d9b1215f187742dbc70bdca068b98f0ad34a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h133b92b15d8a66d1d317c1896939944dd3070a6a0091f8f50e5ece4ffd619c2a0a76e8c51c816e515abb4a96983869089d69e615a855923e4585199c4c115c021b951759c332b3ffcc442f2cc83e8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11bee56782d4f46f14c0cac5007cc8f5fc491f65740960d805e1667117de698982a19779ea8280e80d828c72e8c4abfad9c7d189053c897b06d42d5274e7f9c5639719d0fd646b480e31778e4230e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h793ed57ba80668bdcce657d47b668286d5e41e92194276c9b0bd114f7e7116b9e0df9e2bd10f2882b0f995f0d6d4cd871c41b1f43c3369695f7221e036735c17c8edf4c136b7873639f68e4e118f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d41e7c8fdb3d9ac49e65cd92369f8752e858ff83a8423e9bd45d3136ddc50fc0c5847dc235579d3adce3acdf623326ee53a11883810504a786dff7eeedb2fb2949e38b08bff87d4b2b2aeff6acf2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15773fa495f87218e185ed0d08bd7985c8209569c532522baff49f6a99988102f073ef384ee938d9d89e5aa18e0bde9899b4e2228dff626e92f42ddfa03ab3baa331b07b583380321c708526e5e1a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbe1fa5fb5d6fcc2060ae5675953c53b7ad4ed4c0cf8fc743cfeb997e8dc065a19fcb154388f9aed6c4fe30790adb44843ff7b49fbca8a88aebb8217c0e4b16cbf8ed91a24425c8484768c121ff3c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7a691d418188cfece0b22d2a3ee41281b493247ed67520e5c5dc5139221f6fd0fb61b1f53fcbaeeb2e2d60810455d76196b282787be420de53b40b063e990186467de90dc441d8731e7fdbe01679;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4e443862e3f72bdee4861c431cbbe1c8bb4247603da5ff8489aaa03805bcf24a569157f4c7ba463cb38fd77e70031833710ea189f67af86d79ac97da31ecd052f9b377af1a440a0d878db1064a80;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3cbb30d3c2545bc3ec4a430bfd7db423e0d54c7679864b5f2def03971d790bbb97b620720dd354dc972b411779c5d12a98cdbc4216b4f38ad382b5a92086efb3ec7c57532e4156f1465f3877ef4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h120611606ab7e5f33c0c54d4438afb2402b159521da26a600f0e839d1b5642ed0dce9ddb67e6eed4ef3f9006ebce15a3be49292b5c85f3cc22d100fd2f8b6b1000fdda35b347d9217f074f673bf4c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h173fb472bada7aa5f9c7bf5b011ef166e1b1267441a3bf87564bc749ce8cf6d638cb54c4b93e729bb7f0bad519659f3227bb83df30faf2794ca57545ad9a5974c199657aa0768a2106f3b407226b2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h595b6507e08a39c51bf64db0db7a4dcc4603fb39e49e295326fff79bda2a09fa6571c27f47d1ec637ad21fb8b3bee326c59a5b97c0e1ff7ae0238a89eb5a37d48136bc24064d5478ec9514917bc8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haecb9883672731729c8221bb1f64c7c7aaafcb9e6a234ae29b817b77068cd4ba3d61f2c71c030857b6a14deacd440baaf853ed14f088e576fa5da6ed91c85102712a8dd2241e01cb0b91dfc96ed9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h394c764975b26618d4f20b2c6590ed575036ba076fc5b7e2b2ff067ab5986a15d13430d494c046abf81817675e2f7615c76c853e2c2de8fbe9a9fe4daedded9a5c0b2600f46a6f2b85bffaf315d5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haab0ddb75f9a86dc323ebfbfa009a505a42b68c0b93a2a4dc32fa0af7ca0da3b929685f82fb77a57cb53dee9dd21528e9a0092d9774ae457b15df2e5004eb651206701320933cf4c5e95c7a544b1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16a223ff83942d6b39d4846e4768004eb9cea6984bf6cf33a1baeea38bf7b24fe023613814bd48127ec5ee030cafd17b5ff555c4d87bef96548d45fad5e7cd05a0d5a7b64aeeb5f4e1ebe3591333d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3bac58c7c0d5e4752f5c37dfdb4dcf9f5848c84d931bae901a6bdb2669acd11d9de0a7dc4644f5f6f6f92ef83f80effc88588b9cb24024dd6882553adc74f8eaa2dc35a2fb0df38433836af15eca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h816db7b51515e90da8c8af507b28b1c54a5f9e82554ae1a97c4c654bd20bc4d4cd8f917133ee8345bb0bd80a55557da20f4fc7298b279e5062b9393f212bcba13215bf945013f6b3ab4398349b5c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3e3b29f92d5ad8f945df2527ea3cbb0b95828f183a715876757ec7400a2330b3428b71736e07893bdcc6b5a1fce15c11ba3054619b4504fd4c982d573fcc47fbcb4950964313d58d9aa38023819;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dba3f397db7d23bbc4c2786c8b18e58364552e6304808e8019aed5cc69b0a7f67b77d850f4a902f372ed663313fdc672bf471069697146ff22d1536578385cddadd836fd1f35136a08cc42f8dee3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18593c7f02bdb1fc52c9829b4ba0ace8de6b7b0576d47565ed95d62eba4674583d1bbac497d3a36f2d2c3ad8d40f5507486e26d000d70c166d30b31fe2242352403f5fb7043135a991c405b985c0c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13441c7befb0b31ea543abbd9375e752434c234ebd78a5930ef96fc799cdfbe483fda7fa7b854948503f20dcb34965ff7176c47723e74a46ac8b96becf95e9eb213e8159d35142c1e35f9c8365d4f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha409ecbf2cdcbc9bfe8cd6a1e0e57969017352e87aea20673064f1f795b221a2fce6cb23006c0795848865168fa0e5207512a4d483af815ef099376e46998d7eb289d1141217c41c66dfe62a8e52;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h474b2ff2f8bf34c7c2a007c301b7e3698bf423c3af818409d3e7eb3d7983863377e161383c75d56b403927fffda57ab62480f322eb4fdd240ce6a999831c0771c60f484c4c67d482e8875b24f675;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15b25dfba98a249bfa7eb6c9c17de1255e4891d542279cd9fd50bdbdfd0cea9a1706fa3100c9fc85d499e39c41cedaae3319e49cdeca1d4b5fa31eece865656edb8137aee0497473fe138909b585a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c462e2973b62725e9ccfe8068fed7715df41b6796ee178e22fdafb4fdbd5819044b1d6e687b9877d04ea6f51851607427a5f9b6f3de342ffa9b2945763664ecccbf1bfdfb0230669fcd820fa2a07;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c7c6d09b1a69214db6bc438401fc7a65c5cdcb24e2c7d77fcdff84ea3d7780d7100fc4fbdc86ccfbde42c1d0608f368f94db3896772d77122c1a99f4a12cbbd2f0af3cdb710e099cd3249e314385;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bbfb383649ac568b2aa19d215679f07eeb514883fb27c693c880ca1f9b9936d89278432895b6c0bcf887adf928cd976ce831cad1bb47ff715e74996e0d28cb9d7292793b92dfb7f17e7fd1b05b31;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3ff427b5f1e00edaaf75058a48c6cb9454eabc51647729caa32f0874cf951a63711e62709ce9d797cd5b0b6ad63d601556f5497bed65af5b584d6838496765463f41c80ecc358def7aa590465eb0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e5151610a01e743c5d217fe710fe6ac39de9d2ff45b70f1f4ef2686f85b68f4115e86337faa3f1a46cef1fe369f78e9f5493c54cc1709c704a84db557b5fce590bb113d5bb953dafe388449e505c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb23f9687472442b775ba509ad03e94a612e7373434290166df771402eaa7c7d44037a3b8fd6e166a5fcb21e9111d0dfdab56760c00321acc21cc26ece12aec86c0399551a82103c87080f7b10c49;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14ffeb2b6402aedae2d1639269b1307d4a13fa5e5ea1d35c1fe95000fb544ae22ece4a3577c0b6a36325bb13186b53662d883f567eb6fc6b33e105935fbcd97957bcc675675dcee7f0369903e331a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16262a9a920e05410180865d66d341397a4c7c6fa2917943e887de375d8b01e32329e90a18663d884727915a373cc5e707333eaae18334fe8b4e93b174006e094496cc4fb85fbdae326f8afd0d062;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6c4598aaa998b048d8eebd3b28525e220dfa2e9dfda5d6a8d9b92fdd64fb1050ed0bdce9b7462ddba6406c4897eeb52fe492708700ca091a648230b2d4e692408ed69812cc914bde3605058665b5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ce575dc5a093b9525ce466d6a9e1ef1369281e63a79ba03aea3afeef791e8c5cea1fda50045f8d01cfdba37a8c0d7970ba76d6ac332f5776eb3ca9ae66d8032379f349fa12a0023cef81a8e8bdef;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hac3bf269595e2a3aad8d82e5f9b901a8b790f16f961c88d25f23867329ebe0fc549fb54d19bfa386ae461c3a19910b222add36e07b6dd9d3fcc9000bfcdfde492560658044a9f175cbeb7623f14c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5af73ac1df1c8badb8d976f3c6c02da923d36ced3631ba31c0d084a44da355326b85e9952f940bf1028339e69d3d99fa49ce29a0fa862386e632a8b98db5698902babf727527f25afb455d4c6ecf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h37996565cc00b67eae1cd399bdb2decb2b4a067d5f46f2cac72bc45c6ad943b64f942621bca2318df42771ab9cd11a4414ba65a10ed724f0e0045dd2158a9a5277da737b783d04251684baa71370;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15fc113a2e3c36d63c159dc48f5f212727139f5f964a65d2c32d9dba7c4d185e2e0b6372797f36b6168710d8d4c52c1d220d3d474a804387b688da4f5a99172dfaed8e6a4e1d09d6ee2bb567e8013;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17ab7d5017496401cc440f41a9663365104f31891716ed59c54f41a0f7819e33266ca3d201886e2248842f5006b4502b78724cdf9ee933719a89d2db1f7c09b2e5ee122a21e56520c0408161098ea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bebf78e20aa61c1c464c1f67875407a62216eb6941b8416b74960b9fae922561491a27461491a8106f17828b9c08ddcfb7840f1eac1328df016b4dcacf014612ce52f46d5527103636aa2678ccbc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h154876ea5cbd53928f582dd3df5cb2fa8b60f9daf4edebe4dd66d380301036dfbc1a1a2ae3f8576ffbb62602e89262a99067dc68cdc8bc1d0d136191c6aff4e28dc8b1f6887de9b25a68a6ccd3d43;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cb1d4f0a009849f76969a4838925a88ce9edba6e5b6fe52a649a73ebcdc0f80cf8e49e664dac31a827766ab6deb90de328fd12e904bca516129a5bb5f9f57e44083fe1b9766c5f5c73eff2ead61a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18f66deb9a9e9e345f2aa02f3b057e9152cd6796bc208a50c0dffe0d38412066e78dd0d5c33e7b6e128fef7cb728061fe30f7bdfaa1cde8f4796984f049d7ce6d042ad54edf9ea6ee3b5809b4a47f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18a107833c612d65265b051928ef0aa956589e4f500f50eca0b1545793c5360a0af68167663a32e9ecac1467e976f86a17d34eeda96b1939edae47c8bbefda710e733892fa01e03165398ce2d0df7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he584e42ea083f2dd23413ce14b54beafaa233167519320f4aaaa931d5043cc4a69446702fa92d06e64f180ca18fda39b31358440996311c54488aee4fd9e08d1f5c4e0c5f131ba4e0336d61d1097;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12079694ab05b667095e69f4d770ddbc2dd497d7e6e74e2add224e88b4bb812d24eedf1cfe37b66b4b20bf2e85904ad28a18da58c689d961897b6b5c01096a31a7be30ec9ddf5c10a0e11f2a4cf7e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc048228b677333a96ec0fcf8212875e552ff61741ac819659ff265c8d15d0464e7dda9c60a585e5b75c61c9e6333a1cb74e66591069549688a54202e7b73ba72e8230bce6bafb5d0b433f4373cf7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbbe95f025535936a965e4286e1b362b643f9d200f4f9f5375182581203c348a346943de0087daf08d8a147e29fcae58856b77ec76e2c81325d11304972cf2a63422f328a6fd9e65ba59bfe5ea5ff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cb100a7a36890a6cecca7429efcb3f4d6ed58e6c0fa31b30463303baf2376ac08657c8a1a864160d36e41f5b46d0040b48620c7f5e6af0d7c4c10f6d6caade5d38984527ae5179b51ba71cb1cfba;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c6a9b0d8f6f46f01c24ddf0b6335cee6f9c0e533cbe68c92406b9a88c7008b605e87cb419f5d44b68bd5ef41f6ecbd8df781063ee29acd2e9f2cf227c031bc07a08e01b5a1e1fe6680e45df7bfc4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19dd3a41269ab52b328bbc7a3eacb6cdc356f306227c4e986faad86ac72b99a5fd2a513e8c3759dac51725dd4670dd32947f659783cd88dd17f379bc98024e382714b205d44d8f04e5dc02a7958a5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ae4e3811d4db289fa26029a15f239ef93ec94adef95cb3a3221ad35ca2ca217051e48be9a0d2dd2ab995175b71b37b209aeea8f36f7bc60a5898ba8b90e8abee88595da5c0274f8c8442c50f5b37;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9d05dc0ac03aac14299ebbc6447ace4e57faa432c2c7fef812414f6eab97f1858329f74d5fe817e9a05570b35ea354c228d7abdc378a9ebf086f16a007a186d4b2e380d56780bb7f42b81054a4ee;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d5123e0d5c03e229bfedcfd740c4e9511a0522d4037e281b4ad1ff4fb49949251ba135e24b856c919253e457e412cb1ea3cdd5da45b4265c9356de3901c4d75bc13fb081adebfd9e450cb7381546;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e9fb9e88e95c56d6deb919e110219a77d9443d16a81bfee78f66ee3aeb25b23080ff4fa156d35321ca2275bff70ceee4ed15182a2386ca0e35bb4d06f48d56e8e06923cbf7d1086ac50b1c4d6743;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a6dcff9d2764ef0ed9f75c1467000492646c41ff1a4293ee0bc699e9c827afd6a3fdb1de6c32059a40f78bb36e4f6fc206287adc23b197a2f32722537a2d3523ec062f95c7bf1b0e0474da9521a4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h52eb7080523c165eb308c2f357ed2288aee56c29aac53be9119875b2f6ffa354b33b2de04393a1c47cb4c3bac04cdf11e50e3ec47b85f808e8bcad17bc695d7bbc3dc7290ccc6f84f4573feee618;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ebbf8bf09b8da3dbc2811d85c7710dd7bf1d88d280653f1d21c1876a087a90c1bf82d7556ed8e01fcd4163953afef18cf21fe99750f1536b520595492056ee414148e1adfa4ce70be0c463a655f2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf2293bb9755524ab340c6b8886ecb0568bfe34cd132c12ea1a64d0776e344bf24f13a65081327d6e180dd1b6f45d7e7b611085276c2dc9e48c9d89093f3714b5065388c69288a97285dbc4feaafa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h549c41672758671e1a7088445b9a018b97665fb3ace2e132a24b767806a486d7a87819042eb9e95cb2cde0f16a1878db22f637c3a34a36c23818f51993aa3be82670a609b51cd64de0acebd5f68d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ab075bbd4de3c32a8ab1dfe20be09fbf2a9601b2bedaa18be0303bab75c955b08a27179a715b0c9cc9fec121c211384a4389b8ce51aef8e8a1a9ae9d9a3ebfbe4b39e4294bb9f4c948bfe8e1eaba;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h345373fb9f1a0427ca875717fea3e55cb09e6a5a45b4b2ae7e8a22483951093acf0ac98fbe31b23cadffec3554d0329792712b3a50ac0da8cf46316aca11aaf3f42409ca1cf43727f70d0438f47;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1712e160e3a6d66f7b8c368152884b8fb68b871ecfc01d5f07f238d119f94980f80b865cd924cc0a7991e62397ec8a5600163c99d2a0aabb2eb5d7d50c4c486bcd84e2876658bca70b91e94e4ea3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b08d729f6268b4b88b5606b55f0dfabdb98732db03f19bd3195e38524f331bb6dd7d2c36414c6c5a2e0401e67606524095890e46bd72b2482e2c28a368e634c82f5a91f9734942f3dd9fc558076d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h49560d19f217c717f2b6e0d114532121539036356af75044d566b96fe670ff16a7f408c411180eeea4dc921b2d21cf61cdc0366c9bca84d4ac3a57d1e3ec5986b12900249c71ebd3aa2d2e85b1a5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d3ad337c7ef6d20fdb4ae34186b10dbcaf37cb531fc010cdc890516abe5707eea67c4d322c382adf618cebc6cfeaa3c8937dac926bd0186bd5c8dc6971f9edcab302d3d18ff8a3ad086e3c633e78;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b5783e8eedb9a6cc43488ef5517a462ea50367d78af6875cef43c7b3e3fc43e3cfc0d63f53ff2a064e268dc2abc726976db223b6b358295da5e9a7f550bfc669c64998da6050199a1ae8a06afe1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h58cc12aa6837860f26c644eedf5e8013c051a0f60ecc21dd8b0db290f91f515220c02b3c177e4f7d316858f7f25463f45d4c5493f8bee33c87be647ca0bfd1fcb34bfa8f8e6adcf6e6f1e2d8ae32;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb987fcd6e789ec27c4efae8f9a9ef5ec260d2c04a9c80a744b309805eebabec2bc0b2041dee688a9949731ce8af848e1c2e87c5cca7b7b0464394c2cabff28949518467e7c8461c71fbf7fb71f82;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h155cee04995e1056ece43f7c41df559d2ae4986b7c0cf1d70da7504499c9ea5c1cf142648c6d181b73dd61a40c1f508b4c740d2c550ebc2d9fa3464fc80f61220b11b361afb2b5cfd5da302f8242a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b7870304db9f34e8cdd69de96aa375d43adf501c00209b8383d80b7ea4f3b110304350fda3c95f7f488bde873240b59c6c997af569e2ec0501c07c5d98b8afdb03176b8c593f383e66c6173ad3db;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h41d4bf819c7a790593004d33027d3336da7f4052999fe59df1917966f61dc47777c6e825e51a53b64c6c37bd34b378b14a7b0983dac17b3cc989076e95f33e91cbec711d77c3b47d97499239b5eb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h76de8a53aa3c4e2a3cf4c016de2f56505694511df1d03039580ca7bb6f87b029de130c34e325a4f346d043d00175f9e16bdaf1de715dde212fe2bcaccefcd5fcddba7000567373ac97f3be6e05c1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19ff622cf82481050695a71c762003c4772d4263afc87116286358e49778e562355d22a632958617db0dbe070d458b9a5bfcdbac2b63a4d9a253e973e86d5070896f1d9063eb9708f9eff140c1136;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2f4bd77460491d8d06da09ce56bf222bf0c1af35ab68bccb8d7e8227178ed6c4ed3078183c53e7bde104c517c8f7e30758524584953d476eacf0c89099ddb8ea659b5d1e40be076ec2639c068465;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3cc72601019db90a4255c5352b4978cb832007faa241c62e760008e0077e34e57372c647cc50af01d87bb5cab73007aba3e6d10368075bc56d443b7dd3f80837fad36203ae4191bf40caa1d61ce1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd286128379387a10927face96b13bca754245179126015daff3ba1f6ac40bf906ab0efed8dff913e67ad15285ba77b4ff40365ce61ffca6969980630a9894eda12d3c0c6394c56c506eae95d419f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc78ce3881f1f1d5dd8b758136d6983feb1dbb9fc2ea9ace86d3fdca25e17b05c581d5ec22b23b56063e71a8a4a96203bdadd82f9fd9f61484f0f38b63ccc5b344f38b346f28b722cec1af7c92dc0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h455b0b16b3ded3736d8d3ed48134868f094a979c03d2b58d7fd12c2ef56d680875f7f65f94087cafac5a2e7f9725a093a9472fec93ce125f55edbeb044b806d9a2e1815c4fe9eed67fe5d16ea7f7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h172aedcde595f6d073cf17f1ca408cbd68eaae7bfa4a90a24c91fcd81010715a6123af6667e96668c3d2f801767584365c5d4ae962ffcfabba31e49770a02f8b300a2b45a336b15741fe113330b5e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2752eaf85816501749486646e83ea39841d502be835e45e0c1c2f8b008b406f9af8c2b805febd8514605d5fff00d097a93839343f2fbb66d05cd840e5a05879fe58593c8c12dfdc979b7c88f42f1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h973f76a2df4bdf57c8e22ca1c44e0d686221abe8308ebca7e74ce0d7fe207a113c04e176ba00c7450e3f936dca15653c302dea19a7afdd61484e9f5d495e08ef6feace2a9ca0df32dac0b0653af7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f05a395c1e8196d819e33472a26e77e0d3ae00aad8928e4315e0e7cf87eb75cad47da486dd2c58fcea974efaab96fdb58cb9ae25fbba87eca542ee4bd50da537ff60e58df12c654909276f8dd90b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha282e3399831ca95211f4c2ab7ec72b79985e7d4bfdb5c1a9de4f21f793d07b48d7981d08e26718258f6b109e6f0fab9be4e1f01ccd8e05b4df6ba826896ce68a8ddffadd51978ec33497628afd7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16c39af64e200edbb98995c6f86b12431500839c05e913ba44e01ab27b4699bcb0f369345f81606dbf18cce2886bb223cbf1fc9ff712dfc439e4eb2d4e84ff2cffcb1b3b6b94904d90c4309f4128d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5e20b5a83588b8fb68e8326422169525a9f4d5ec45e469013af8e8bde257ad0be288f133732519e47960f2d3d65ce4ed37d261b36a442977b3cc10152c334acfab72dee555ff109582aacccacf74;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf37109e3444484e9b4c9f1b382f89da3fb4db218d34ddd5b1a5df8dad9b1ca6b6a0d62084180bd14892ac6ca961cb2b4e9ca421188413a6277f612ddb5c46900837b52ba92918ac440ea3ce7f276;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8cf7d95210f9f4ac06ab0bf486237054de7ac97835279bac173887d68547df48be6fb2638e2e40a161eb44000e594cfec4da74d2623c8d5e818089fabfbf801b198c1018167bbfe153a183e74f0b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e26de7bfd15261a57e16c2236b47a61fd693fb3da5e22348f356ce8ed59eaf086ea763025614e408a8c9cc4ced5fda53e9e4ff9d3a80cf72597c0407eb0516bc629f1557eeb4e5e7a5ed317af3c6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11ab6494673d30db8c0d59a69706437b6b449d54d2fc68f29d2a57de38137130ff920063186452c13e7dc42103d460d7d5ed5d574697b1067e1b0379f3774f6f502aec090547d96314a127e3b3b4e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h120915619efdf6d6ba6723443ba40f19b0ad5fa228157ffa0e269572cdb8bd9c27874a27660464f783219b6d97c53de6128c07abec0ca7114c7571d036bf165ea86f9d34d8275b6e3d8c03b1041ed;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e0b3cc8b2a9b8e51c098d68468345fa76b9aa3522e9d9f5c638b0f89d8e0f18e933270b0ce9230e77dd659ed0619f06ab8eb254f2382924ff1e7ce05008d75cf92b0ef7cee2c28b3ec285e6b3d5a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8ecc9dbf200180eaf766dce22768d6bf295f3043b4a485202d0f12c2a53e9e47f2e7e81de0bcc621da8c587ca995a779e2952a08ecbda7e4c68efefa225714ad21d0f10d74d5b529989b7b175126;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf6d768680fe7930ab2b3b22bd9ad06d33d14738134dadd188fc0361c60f679c815ef26b443c838678b9795bf2c68514af0d00ebd32b4fb33f8a44f8ca61fd7c8236819620c871fe114c88611536b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12c8d58d1783169115ccfd8ccf1396c38ef78b465a5352ad8b05b409d18b90c90d7a6d033ddd6b1bc475dfd13ada0aeaa4ea8cea32788d8a6771582663093300f791f2c3d5789d7dbab8117677d3b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h124da8f93c503bc444e7ed104821994bd5c37132b0043309f7ecadad8ba3575f634581cf8ca5fe0d15e6812b2b52d3baaebc60f115a9d97d956c60f740e1ff0e1e99a8ef24695a563edaaeeaccc3e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h586ce2f3d52a275b00c542a8b1eb9a1a71af002dd8a7cd74547326785852a6ad0adedba474d00765d33afb783614abe8d615b1b3af1eac67344f9bb332edbb3808502437d43150267f46e6d2007e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hec813766e66f3848fe0cf4eb022ecee62da694aaab913d75346ddd2141fb9a1639f3c1879e5b8a0fa610cf2c51871570ed3a268ed8c97c7d5bb3e098688a5c766dc270f465ccf1119efc9e540ef3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ee73e4e8b08bea4eb89a57f0e4f509c4c2e569dd3dd7fb7ff3421d12c4dbeb0249baa0eda529335c1db0843c6ac63c15a9b9992c2bb5ae20e7d2156f6746839ef14d9dc2a13a2f25d5c76c2200b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4f5338fba78274fc1c08c49f3eb8d57098ebd114d5d5d90396d27c76a95a993eef17f5e51cd1dd3f478d671bb41be9838d398651f7ecc96713382a0a0119b24642b57a8d002418cfbcbc5ea12c1e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a86ae67c49266a0d2a7001bb26251bcfeab9228ef6b7352285b45610d027ef3de1e07e6e2acbe4eec7975cdad1266203d40625225bb8d620fb1d69fba5129333d7c0730c26e7b16e8181f9f0a63e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd21aacb74d9e339cc09a9b58ff6d808a7a9a3ace7c0204c3cd603695ab8c83bcd867c793f8db5a71ef644c40862d0e99a5981ba293f3a6cdc211079dae28064d394a372ff9ddf5c012c4632ae680;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13a0492b6385af07179772ab338ce482788262e689dce7509d7bfc35e818b1f066c62bda2e1c6a4136bbe2d5fa0781512be11b69078b8110ab9628866b6dd8ff693de33c7213f1d2318adfc69c82e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f05c4bb79b7b162a01697aa3075d079e4ada833bc34e58495a20ffc310f0e56b657ff68a344f4188d6e0a7dab2dfbd9c210ebe369bfb513e038aeb329f0b1f7d62ff37281ee68e60775011175bb5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h100206a0993e5dd0866a3fe98c1273e8dd6f34851b5e0719ab3d9bc0628da1d43d7e049be3cf98742363e8c03b214cd5aff9a46f7923fea02dec5d3cab5e1ddf54bca41927bbac087b250ea9724a2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7ca03bfc0469c3a65769856fd540bf07727f3973c9e704b3181400ffbc59cca69d6edec9e36fe6570b6ae7ace0e2d384299baa8d0b5297a37cc007994079dd48c12f89de570615374ef96c2a2292;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13d953c4fc04cdc8a20878ff48a08ce7194e15ef274b3fe48f91cbf6024eb597e18ef96cb44c91c69e3c085744d32fa54fb1868177bd691993d033e1a8c6ddf614718dee6e1affa0a5ba896e92396;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9bbf25ff718f3b3d1d4e8d4ec928028b105e525685e7af7ce9cf7130bb107387233e6d0cc79b46421a626c71ebd4c7252348a6b38236bbf647aeb247ad22952652a27ab2c4d21fa8adcf967640c3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb6ef0959bb194327c40b9cfef5caa8fbdfc5b9880e7b1255d49eba56579b5ead03866f70aeeaad22bcbaebf8902ca31543ca41451c66c3e1986455e20da02013a9cc87842749252394452c50c47e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f8dec88a89581f86205278a0c88dfbd3b8fcbc8abb46389f9ae7c4685e258a58a26a0d533c93db1a0c43d1d4a726856563ca3d54aedad0a2043108306280d8b25816e9303ba9b483316d2ae00186;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6560922e0118b544224293a1be4d7af07991d26601edd25a1b43fe79c172b0c26144787e7bd9a4c34af6283cdbfc60f5c17789a80cb446df19e26c7e831dab454515a00a068f63580e0109553a1a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h158b3210b2a5807108df826ecc5211078ead98cab504bacb57cabc29a86fe179f418feee4a28639a07f38218bfed08657afa0bb54a5f9246944c30368d8bcf10b7780ef36f07dee890110e29cbac8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2e60a10da76370f4bf5ea707098ea7f422d14be30c8f72b03596698d77db907aeb743460ce5bf7921beea1494ba2d02be4f7c52af488f0c1a52d65a4ef7fc5cfd8e9c40e3cf5f49f13512585ec0d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d5ad52676610eed94442a7c299703f5fd37edefbf1ba26d6b872683257c9ac91427ad43b45928ea366a5ff66d6a5e78d42523778b40e931fb6cc652227dfa88a7794e3030082b942c75e5bf5c41c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h95b52d07b8e806af62e9349d670ae50be2ae559199260fa69c1956e052babfce4ba3ab9004921207465b26a670ecc3d3dc44508f30b309e99b431541116278daa77431472fc6c812b85858586cfd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9fda7b48e08366c7f43483ac4d62c8cd6e6b84a7ec403bc76f7848878720b0f0d69691db7ee679cf0bb94fd90667619f8620b96a83075c749596f4fc953d3707dae73dfe32f9ec22e98543cf847a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc29985fc07fe4d34f5bbc88df2114287003f290a10560e26cca6490dc73ecff541a376505ffd90ea019232513b471cc7adc56a002192288bda71eaabd75962fa00109b1e8fde5e17b78ebe492f7b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14b7e7b1d7e76a643ce52be3dec7f461286f69e0a5653d461d07f8f3558ff1faf87698f21779a5f84e1803e37398bdc02ac6768c009c286c13b3bdecc774375966fe3cddac2a785fc48b617e575af;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h141fad0686dedf3753ac845ee982f8f5c19c11effeef1c26b2d4dd4bc88ca68f50d8706608fb570338cc31e63f3c5145b9f73685223747a304a411ac0ceebc9e847cc03ce7da8c6fbfc8fda4e1c89;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h50533459c8f135ceb7a8ac7be0a1f98cea584d9c377d1ab4d69cac24162e39f6888c4e883c6f2cf22e33e2b1891c9c50781af7daaf786b2e4c5f8b3c69a55fbc124821a1d728c3183bd00f181ac7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a26bfc96db790b1e41039289148036dc5c1d99e829da2975f8fb3fb3203061aea717264f99296c20beeb7d2dbb59a9a433341048264711639355abe12c67a3690634bf3933f673ae7d783f4d65bb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aa0f3bf2a94c659269099db6124ff1e15d0db619157a44ea004df1c9f3aa3902399ef5201e84b0ec824d024885f72b696f5b8ae6bca0078821c5be5bd2309c18370e91c2f6757329abe947112ed6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h161d43312769f425d30404cae4cb27a84bdd1c8766c20907a2fb5506832a07c645ac8cf59c44f0165dc435dc44c6bc7573f86dba2b7eb6b081dbeeab5622356b359ebc4ae408c6154a6a3f1bc4e6d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13e1e2cc1d6def6bb77ff94fc389d01c1a59bb4a74d347ab20692a010966a69039df26675f395ebf196ce7e16762d8ce5da0c3fffd190b10b334ddd49f99d8945d3c9231527784688459fc2df5dd0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h119603c9dfb98e17724f443d04ad2698ab1a5f1f11fca9c05249a52b1277cad9fc4d53dbb31892b689d8f20cc830b9351d757e779d8229606a497721db417f0266197986875d44cb720ec658a335;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10fbafe662bb162e8b76c39a09c84bc009da8f6895d2d3645e4a83ccd4567740c62fe873c4c9e992edda650c18c2d7bc065e03394a08c13fb1ebfbf34c3cf2edb04a169b71a5ce12e62dac1c30b56;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h24d8b9d32f54cdb1e5d730bdb930ec7ed4f838c079bcd10479e86643754072f510d678daf3247ab39314be8198084003df96573b6cda070dae9f703b064565bfa0961ed1db9c15d88b44bf3de112;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15b053374f3fd1631e45237fd031c1a4d384a5e38f65e2e88fba3887e48ac6053ae2a4bea75059244fee9265998a59093f104a6965e90f88db2f8e1f31184f0df4f6a52ec346833803364bd4eefdd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fc7997167205b0d5bf8762d3ab40fa41fd2bdcacd1c4e3c04e1ed528ef606e24a4d3e7e4a5232a45e5b5a9994f1110fe2dd30101830927f38c9b65c6ca01f47ba3fbb8d703aeb510439dc940ce8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12d5130e3c01e1efd2a06aab19dbcf65df3d5aa2754d72093fd7b9b2d83dc40279d0e3f94f4eb01e8e2440b78f50af385de5c7f880c983bc76a7ae862e88efecb076ced95bdfc6675d634a0f5c2b7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h80b4df2a1c3211e169e4699204c09da3a605d770b574318c4f4da0a4ff5609b58df136c9389b50f495b009259fc4f23a598261f53021605a6ff28733039b8f04212ea584caf04d3979785749007a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hce0776cec3fc9cc241808701d182232827cfb5128f48b0c5cc13149b8012ce19430db6413ece7a6fcdff8e7c770e5b65460aa981b0bfa73d13b997b989da6e0c2f6f1e571b38975a0c524d939314;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h145e679dc6a9ad54705000a43817f58b5e3329933903ce71b59a622c0dd38f7e83dd195dca1bd78004e6861e69feb972994674eff77d2de5f1373fb8cb4b9513bcbdf87f348188ed679f12ef22283;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h76fd1971866ab808f890eecfbb4b0b479d7ee76488511da679fda732671e03f7aacb4b4348563e6c93b08c87ee36ec0ae37f5340026207151ad3c8e6096fce697f57825440d0f81b225084cd408;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c13da8c610769d38c1190e0113a3206abc6c7cefded5c95cfc5b511f6ebf0c3ccda8de30ae57c0788abdf4d945d171ca6016dd7ca15e5d9a11a763fd9d8587cd57f2992519420a99a6d8b5886d97;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2776195ca80fe1713f0fbefec5d40d7bbbb7f8b223cc86bec3a0aa5335df991421481e7f438b15d6f768162a43cf631d306b251f9892ed3f05f865eb5273d986412d05dd2069922d59aa66bf13e8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb758f01a18f441a5092b6fdbc720ee223dc003151690b39b32728760f6a94cb8f1c9b2ce5e7a8d351024aac27cb54b2af3441b60a70b81c7fe2921411afa02c43603fc1c4b39420660ef36307a34;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17084a921e71a6ccd5aa48c1311e962160dbf986a1350287bfdb9bb9f405d5b9012fb470650f131a4ae9add755232c8f78b71f87dff4d8167a62bc24fb0eb26944b73dc01e2477f518c9c28931d78;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h166d27e151786dd6f1aae5030d4c4796ee0855c5045529e4b7292b8ab68705db8b88c60c7634860dfc7485ce1d0275f1d88258bcbea960c96ab0f2b961e8080e54f21295a24c67183135c60ef3aa4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a682a6d21f7d19ae8fd334f8caf01a50fe0b8d59793cf03e7fce83f3e42711d8064532c10ea0df980a606ca6d2d105020055cfa6ae3097706a8c86441c63140465b9193a594cf5dfbc75a146f610;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d0fe3ce47be7839bcd62a70901faec521275a1b2b97f54a0625667aee5c537f5d98fdb61884313fc960ef3b24dab143a28323bc5016bbe7023fc61203172fd67151e033da4b253fcc1381c943478;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he079d0dedb68abed8f2561ea660609826bb830bb4e41b947e547400324d56afd6118452e41594faa92dc988708f10009fa7d3b47299b54f2ca776913aaa59b70f5367256d53209d7204d1f6931ea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h183020cf91f2abda99931dee7fc675e9b621ffdab073a5ad92bf4df69e6b0b74afcade37bfa71dacc46c374e4d22ac0e6e1e87f4774dae6113ff5fb2175243372bdd28e33bcc0a3803389bf79f63;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e7898a9d2afab7a27c7a3c1940fd61b87492a8ca703b686af2f2d3d1e62a0f93990e685a88d535f63b055cdff01bda3f861f794263afd376158e438e5784140dae2a3f950cbf0614dadac922dc76;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha700e039bab2108b70dd9a8d827eae70097310ce772bbfc708a8795147cab0642041052c534039e43a2bbf3c6f9c0fa4b6a62435dd8991816e7a4904e7ff866ff3c0b85ac526a84a00f48ddbbf67;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3eb9951977dec2fb1a5d760289d58fe9ea85d93971f4cf56578b973ea73cfacafb0de13702bf30a1bd8b31de740309bb00d33b131bd634102557abcd20b9964d5b63510399ee40635324b355a1bb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3b9b87706f8de225ebdbee456f9f1da0670cb95c5052721df2e52e118e688b31329d04d10905d015b953a34f62ed2226eb203b993efe5f9ab5ff49ab8baac5dc529f008bda7f75f2e7d29d77fce5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16607e5dcde66900a6b107ab97599152e4f7e02aa6d62074a2587cb793a8d489d35d073a2b66e4f1da94524a6a3edd5c808080ff87ff983569033c05910147f77f0baa20db15379c7a76e0390ba3d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f8018467121159247304bcc13ece741b51a1bfd0994fd63b8d658a8400182eed0d3a9127aedb53e913f5c617ecd48e746b5c8773aac97059fc9c9e131d439fa4109906655aa62b9a731c5e920018;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d2c4c9f25cefe4ebf60f7fde17e107dd67a908ed91fbee95b36b9b84bd5792fadb80129bd6525ff26f6759b5609bfd8c7131a1d16adff478e695976940bd81dd4f3b3b1a427b2e5f2162ef33b763;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he7a5576364a22da4dd26fb83dc8158e37a881386dfa2497a8eca0cf307de072ec96e7fb3fc9ba5964f30490aa99f4c4bb24b393b9c900dae38617da1923d765099e2574da17af7e0db3135540ed8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1593b50aa48c5e52ee743b8492d37543ed843c32d72f8a02a3124f6306361066493c24c666162efed9850f4123a3dcf278d7d468c13ec9be84d3be3876efb5368a578a275d0c0ba467dfa4caa55b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19dfcc3f732952a395a3155c40815d3844be25ad1084577b9f7625efe75acc3c7c89a6f56158b2635da6a6592e0a02b2b90bec221661394ce4e11e086d44c44360445bee07e978acbf92dc6dd69b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h42e9727763158d215c939274284496d19aa627a71e188e292d5aa41f131a637070f7faf870e631cacddb2d7235e2c8fcd92d32c77edd4b6dc6d3b616d41b1f9c6dc3580f75f442d6d595dc38216b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h96dda3e648b81b394fbeb03f20de93060b617d708ec528955365fb59f0361a297df7de4a8a269f80395a1a05ca03b46c73e61a6b436f813058ef96f59024e26eeb4e9304beda7985f44b9dc12079;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h559d9f01fef181864295c9a94182a7b4b4d45ae5cd10a6b4928580c14d1847560cb56e6c17340fce80809b17a8e715babdcda58a06a024f4a16dc4fcfdba2c401ed8945cd95b76648f49d1fbcbe9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19f4d122fc54a9498ce751f67d76bc300a663a8a42d527ce4acdb90b61566d5f1f744052c696a8270330604a7dc420de0a75b5215928fb5cca63b47565ea0e7fc1f7647e3b8f64b251dcc7fa93917;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h170bd8d2cc70768631c20ccb671db1cac8c9315819a8d93abf401f4b176d68a8004fd4abcd045abb0a11566ab39d52ee4613d616d0c8647297e219f2b595eedb24ac3bdd9f2a9403b82b639505b13;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18806c996a089d9d8ad51d366d18cad78d4564c57743e7808ff21439f7f8772c031d6c523668d57dfbe30759ecb053c7cc81c538b15162f8ae7d85945655c2f0596d33f05c016c42824b3614d33e5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dc09eb0179635dec58ce2fa720dab1325e2cb1e7148d3c8a2624f28b22b32ec8f75b700e1b979489cff8a781125c4c19a7ccab4c0b5596a2a9d421005add8cc698e9c7d19a00c19d3d5ecbc14b42;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h44dd63378f6225b2fb889ea4b621c55951bdf02a86ae0196204e8a9a02ba1fb44deab6d541a6ed1310a70a8934519f66cd17734901b66464b217a65e3c2a85e192f9f19a557a55ad9c27a5f93cf3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3619038f0b8814fc8c7ab0cca9895ed12bfd5b0d52a661904d2dbcff51648a99efd291d2f955a0d14c2e2f3d057308bd138b14a275c1e4d788cb760ff96ad3b0aeb8fb80a1e5bccca3f05850147;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1765642f59eb330437e255991f71854f495efb9c77004f4701aef91d43f2c1b266886f48497b6bea648ae52733b70f5058e195e9e7646685bb88824fe1271b663c09e63e99638eda58dd62e2c9807;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18f852e3fde0a46279b4a9d3408d07f66741709d7fdfef2cb749855330934661e503c72558912362adfe155f676569c203a807e3f608dae7beec9fc7d91baccdbdf0fe566c4481f9b58981873384f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h131ccea093ed62f11970ac43ca0302718b11b4f67bdfbba62527d97788f868f35f85f108ea0a5adcd78a85ccea28ffc0aa8544ee10490d7ce09d1f4ceba95cf1425a6b798c1b89ef477306b1f9cc8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10e7b6fa19ddbde3db2cf13c1ffd63eef291ba2d0ca377501dd0f080f6c38baade6de17c68a098d40fd27e2f9e542a9b40a35c0cf887570de0678f70fc688dd2a328dbde918c76af4b58a4b41f8b9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6db0d4f4302bc5f4400fb0a6b9c906088d80a6f57b2806ea45ec1fbd7fc24ec3dbea167012f1084542ab44271009b01e8a60ba67a38d91008d1d7229d73b77286aae3f221bb388acda3bb04e3e7a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1acaacda29a43dafa46887461a9394cb95e2c8a059e7cd2dfe81d86c062b9d8ce9cbf83b35c5b6625fd961568c388b049013dfbc1fd6f6bf6693fa0bee90b8885e30eded23e579947f30bfa0412b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb57b7c04bb43b1a5512a390a747086ff9e3ac51166ecf2cccd088e783c61f98e7f04881506583e87c90c6d81aa35f6fef07553dcb8d7e6cb85fadf0095df26ccc5ea069f71accdb0af8df6a088a6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h48777df2ce47214d9d9ecf36932f76e6151d2421f6b7dfd3bf95a74b892739d4a4bc8a641811c4cfd6fdfa2adfa8c0030b08f1635712a5144237993fc7e9171e2ef3be332ec05b14b887f2776d89;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1132fb08fb0d47a7b7dac28cdf72ebe880208b0efdef890e1e80d084bb01df58113b0881634d4e30e385430df0c2c3aec92e0acc7dbbca075868a774d494ce955cf7932f58bb5802c8980b4a01b17;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1abf1b069a0266c4892babfb134b2dad9181440a064bfde4c7b344a5f4247d51c7efcda904b3461340d5c741700a1877ac5d6bf124ff985447b00cd437a97710e951ec391bd2a8990dddbad83d3e6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h390674b16a3deda770a280114671f3a7d199dcb90bbe2e4f4aaed0fd32018c43906f2c8f02b63a27561813fbd033bd02dd906dc191a7ba6b920f2a6f29d07d126f6882f0544e88aa9772c032d4a9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d67ce7597b7dc0146e0a374da3ee9eeaa830bbf658f6fe1b0d088883d658b714423ec458f77d4bf510871b0f756a9415d717f324d950d03d8346312119f1b9544f6a647477b316712e658721969d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h674ce50f4dabbd3c1d0c4e3265966cae268dfd8611e911eef238b5d46c770c42c95cf3716a31803b15cee6e0a2d5bda75743289be150d13883c42aaadf3631d12a37655aef430a65cc69a82516d9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f59c660b2a2879d6aede898f629acc10498c8277ae6ab8a2a368864b76f224359713b4a2db7e279ea14062f5e94b2eda1b15db2e4879674205934c0e7afa54841aa60607b056df115af5d1b79f07;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7dfb20a371dfd59f546276849ac598b0bfe97700104bb1399b417ad5d7c91aceb69aefac562ed4174693cdf737b36b9a0fa6b818539ec2797b8e7868a9dd21674e7d92069165b3d93a58c31ad23d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h963e41f2f50db97ab809e2bd7877c09a506596d578334b868d4fe443e37c518a1b56bc708a6e9f6a2a90d0250015adff8b8e74bf043631f7b87ad133dbdcca4c2a358850a2e20016670fda5e111e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdcf8de4ef3a136bf7addc5923f101e3e6a6fb968b4e3b7a2ee45fcfcf58114e6bd13397984365893d52b9eda813b1efe9c6effa0fcb971f260bd9e7d2dfa85817830e3ccb2cb3ed213f5fd7b1864;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b554d05edfea5efb2bc2be324e47c14f7d0de1abd0cd85d8669a3517ae35004c228a56491d03373d98fe5c55ff3938e9a88ca6cdc29f37698c5f146c6b3d31d452d015ec7b25062961db3256c4a3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3402ad6deccd007c4eb91eecc55ad8984e4ee552cd63375302c1626623069b7a3e2a63b4e56d8c0f3f41b1526dc3ef8683635c3eeaea7458b38200df5f002229ee5b25ffff76ca211cf00fa4dadc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10e85c7dbcf23ff6146b67642b37fc18704bd7a7351dad7d88e256e572860f51271a845761ea6592e52ad69a9a6f8b11c4500d815a280d03b8c9e202a64b76361000d0ed8ae3b28a8f03d3cebda5d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d9c602027ccbc8f83e18c80343f91a2abc59ed718f93dc8bfe16869fc4b4e9dab7e3f2cbfcb62f7a0fc2b647d6a0768080ee1d2d6049675d1d067c0bbb0baacb7186df5b39f8d78fed77f552db3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18ada2d25abd3002b66c7ad333e5d2e43f2f9f47a1c8f6ee2f5d64af28cff1431b247b542b26bedbdb3e837ccd8cbe3d998804819668e3a776366665ec27d53af9242d3b05662778c65657076747e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5c1d1383f07c59085aac01db8a513eff8f79604aefc4205ef59e2de1ac8cecc517704c684d6bc137fe18ba7e353020553da96f450effdb48a1a96ba3b6371e0f94a0531809749dcfeebfdfa9d00b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15e9421612e03421bb61b595a4f4384370481bcf1aad25d5a8b018baf3cb04ba2c80b808e7abc1831f0fe6abf0902a53fbaafa776dd4762cbabebba2cd49ca2739d749317ff802c541ef62072e9c6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14506f88f64bca4f25d6ebe171b9b14fa293287fff10ae231eef3f88ad1b74c7d3edc45608849953f8fa92465dfa2018e61055cf0b5e696b8cbcc6ff825d4aab90572563455b565b5648097505b26;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf402d7b67a94ebbdf857c37f595c1817e9d0869c7a409819d2af46773555509f90d8f138d445c38dc441726c5fb8487ad4836dc5738169cc5ddecf29c402e632595cc76ff8e127ec55bf6abec613;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1301c847383258095839607ae15add9d172f9991ed34928004a1621ebd36b5a86c391bee53f9d7b553d89e51631ffc4bf8471263949d46ef135ab2246e967b72f0f67b3c08b17425f758604033057;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h136538d868d08681386ebc7a78e7c8839abb3a4a576d28f5ca5baaa1bb54ebddb47ff0cac1a9ff77184af5f2dc6b69571bbd51ff45d0bfbd6bb4468bd29c6fb4085bb1f98de65b89a8f6c47e63709;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1edc9e6dc466f43585e20883fb70f929abfcdbbb27701cd3d10a1220fd042fa00c9cc91faa2e6d574d0bf81c20e9ec32b1b64d659ff10fee354bcab3585bcb40143b236e288508cb1083c4b5cdcd5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2ed5485d23b4f194f2d7d5027dfdaf82e3ecc5d05502a4784243dd49f98ae1709e8cf1b01614d8c0f31c9838d44f31731fdbbfe3b0ab838036feab7d7581ff0030d63eda24ea7efcdfab739a9a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h107722388cf45c97ab27ad35501ce3d953a310cdd8f1169d2804517503e57b813516849617268326ec4073eb8f1e55b544afa36757d7faaac4d3a1d183f6d3ec8604369a12bfa7dc8d9c5020b2469;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h981a529c143fbd7325722f4d0ed89f8cdb6ff16216d532fa97949b865ed346516f6c98cb1def6a0955a9c555af87431cb2586ecb0eebfdc67ac0799901a3e2af6eafb8cf5c5f25d6a64e69086256;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7c9801d0835833fd13bcef0ffcd5c9c2c381119e7af904f4af0c881f30edcff42834f896d74739a150f61d3e8f156fcd7f39014dfcafc42fb5cd4194ddab1e73d192ab46fa79b6e9c99121df6923;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17f96f0e1b153811850fd59defabcafd314e93309381a9904b7faa50a8cfc00b755955ec43c6009e94c907b3acd966f693b8fd8f76a678ea4fc95cf1b4e7eec8bed0888fa9910b1feae3d7aa4a578;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hebeb081ba482017f9fbea7de13d51a4d5427e348bdf2b4d8f1e827eed4f8a54d12997ecc2c1dcf41570d2d200fc443fe6ae82036b70829844053273fd1350c5839a4a6ac4f48703e68c7c92b9ff0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h790cac9170abb01369cae45a37dfd8aecc93eba969a797d953be4a74faad97ffe98b92cfcec197f503447e39a579100063bc32e25261133ce74a4a6a4d82a3195b42ffd77dccbbfff93fff7c7c38;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8660a0277d88f5ed277685385cde96393559e3bfba866bb02049cfd53fbd1f7fd433e6148d4ecca3ae041d5c536faf6f28aa208e01500471c21b0563c111bd13d1f1c15c6310f0b1d7b498ce03d7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dbcc88e41e5ce33cd64dfe0a83a95bb3d8bf9a32b9fdfad6d30d9fab757915fc77b417c1e576db9494b1a91fe02f0a0a56aac9467e755d2af63fbc0670ede0cb5494a4072c42cb81ccaac4aa8576;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc23cdcfe8bb6a2202b1c8f35e48fa63910dcb1d14b30e76d02449dd02b756ee45261434a59d91318d522d06fd983bb3e0892f8ce460be0d9ed554b55cef90baecf67461ba993d3d753c7fd6f2e9f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h221cd1ab40370412938b4f19b6297ff77d672fc67d3ad5da697f5c2843da7200bc644fd3b7b717403469c9192c6d95a7bb7baf4c1f5103c9117b80cdd7f0fe23d72ed93e90861969be169d1fdb45;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8cfde3a3b5127a99f7eac0eac4d8d892be11d6dd27325f3eab12cb14c72de421ebad513e87dc617c39db0af0de1532e138fe08ab6a971967758052f1e5b107242ff2aa7ff2f8b9e7432ec41d573a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9ab4ea83439446298929ee8fe24ccb26a65f681b31d184e244684de7efd5b2404c55fb9f6f0e8099ba62d228c9cb967833a4e6da6f13769f2922e2867a000fd89d5e5d4b3e0c8d287e28914b4c8a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bdf3fc0c9d52ce2b031c70b9c11d80e3d8e1801c130350c494996da925d021bc4fe4efad79edb746f1e356e1cc1e917c9aab972aaa671eb09ff7b3c45f029b3a81630a9e0b7b2ab46b4de1a28f2e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11c0a3466aea5ab6bc742dfb61805338eb5db56853b9f4a5f250684d9f9951c820788f6bc8800e50022b08c2d4093b8d627e78f99ef112f8090cfc878864af6ae3e748e2e82959600a946becefec;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1377a09cf6d3d59d67da54e8096082dd3485e87aa8c073977538e31e689f78bf39adaec55012d136422e1610bd786ddc9ffa51cdd46fe2acd9f3a700ea4451fd04a038f732e0226e4b3cce5d17ac5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5a5106326f8b4fee336e17e8f0b125cb43572995eba7f0d96812b877639eb6fdbe246bf25de1e72e7819912674f0ca6112f0a92a3c1e7b504e618b10c97b2304e12b8a6028f19e5b7b4e5f59d784;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc18e23b5f70f4ee44b0e15cded3abb4a89a50b226810419ef9e2ec94fc87f81235a6c87f684fd0d560c0759afa6a56284cfc51b5773f11122ceba20c62f3108237111bcf932bab5ff7627d306fbc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h40e2b59801118ae600b1362fe2d8155fec27d7c2f8d74e325d80db0b6a88c64add54f16aecd24635afd2e446c423d22fd64928b562d869d72afda60c8cc6d9eaea7c88dc5b2d15a11fed8137b673;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5aad5f36739543ac5ef60551fd5ec6276e5e003da43290d24c077716b1d8140c76749523aaac044aaf6d9f1255712e5407727f8345d51cd3de5e50d7dd6bafbf2998f05642b61dcb4599241753a7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ad66c446f0c10c9db343bab9927aa505d3fee0c87280ff2ce580d77e8b8b6f9d3950d92ec2b9351f2463cf5aff77d8ec9af540b24ae00902608df3ba53995cca5e5630a20f0af737d1ca7aeac904;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e0b43b38a4dbc0fc893179d06a6e83056e6229c37651cd5d3cf4828fec5c5a1661d8dafe724bee7135bd50c0a81f6389cc7ed8f73aba56683c89689f2a1c3f39edbef0b48cdb0996c4ac9ee4e42d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h25a73853e88f5c2cabe5ae40b00bf12f4948c8529f769212acc1f9f50f125d50970525f30e8fec6fc9e37aee3f380681eac91991d15bb53e6b246226298c5341467097cf790c6aa17170d7c7101f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c3b23c6e39cef01467251d0b7756ff0420c4e774c6fb49f274e0f3a37af6036f639e6439a7351d83f5c3da23c5af7e7b4d304f13b13b0c806630481cb569c5cda5d82d865d5a6163efb0f02e095f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcc45ced03d139d5a36ed1554a7caa0d2a4788e8eed0631a65fecc13819e8042ffc6b4ef275d3fff3733fa701144e32621d59ed5aa691de68b8eab5feb983089b8c8ecc061c6748f3e5cb22f66e97;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h86ef33197ce9a82ed8337768136301144223e10f209d4f5fde49ce85e4ffd6c6ce6177e7c002e97c36e81f7ea88754fcbdfdf93bd2e3652fcba7d4cc78702a8a47b160fed6ef5bbbd1cb658a58a2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h49eba76259acfed185151f22e47d054389a0dbf3f0eca6f7a352dc91d7a94c78fc88498e41247d74ca5b4608660244f9ea4b65958b8ba505e82b083ea4497c25e8ca59e19fa66aee209a63f328fd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15d65b8f7890f89de137deab2bde621bfaa78b68ec967ef6c85622819479287c89befb02cc12a7af4ba83cdc48f98b7c560de0114eb95135188d620c337bf3d4a556943890566d1341fab16e8484e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d33ecdbf5b1288fc7d4e8615bb29944cb74df027b4653d1678f92c632feac28251bfe57fdccc524693b1a9873954c7cea46d4c311f1287c0fa0bc81116b3efe045c1fee848ee534e4742afc6e1a9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ba615f7d20fd4902a64eb43887ff53782d5f332229f127ca9b400992c95e14211225727a1a251573dc839e7237302248987c43bf5996efcb7a3a7d52dc14438e0a3dd30699d117a78dda42512456;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d0226e9b0e36ba29d4c06e088cc989082f5f5bc771ffde707a1cbdfd65c593012edf04ec2a6f6954d06bcf2e4bfe42ef2ed0a3ce7d4dec1a43f98e9e631d3866bca137b254254f74df55660bca0c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h346d956a471cd944692df105ad91f149f991311a6fb7fdefae31c77e876692419b068dcefaba6e91f16d62494a8348cdc5017fc6c27fa9cbd3560b7340f7e4253dea61f693c9f4682819cb156b3e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbf0b2720c8250eb151878dbf16a26d9db2ffcb0aa4e6cf34180b28c5a928cd42a790d4f1668d42677c6e8613d37b1274d8edc2742a6ed832b66323ff40f4f3411f3e1886a5d4a51fdddb90fc9e13;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hce0539a84d25ab7b37bc031f197c00e8530ee18a50b945adecd7b992219c7065f6c007d7aa4d7b152603288f3e040ce1ff80674bc64446b65939d7e784e10d52504e3c681c50586ff91aa37c6c75;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc49e227a2de3b4582c55566c1235fb1235bf0333af9512c4effdc657f6dc4faa674ae12f9540dbfcef6ce9e742c4219f6ac6f3c1e458a9f99b5888bd1fd07fbaa4dd4f4d35fa53eb96615f2d4b42;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h124f5b503b7001053014d886595355f510fef646652b0ac02653e6550e8abbd44036a7197aa284f048413b5581873c10f23c377feeaa59402798199590bdf26b898bae4e0dbafa2c869906aa95564;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8c473958800399e636c71c5604c15f8702984b0e9abbcf98309374f3f67c80879c28a0c37ab83c04e234a4b56ec553a204e69bbbe860d6dcff198007218f7825b240c50c9990a8bd5d3678804e58;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a62edee3fbd0194bf87cbf10ba9768a9318ad9ff9945cfc6929a7f35d696742ca66b3c1c5a02645f76cb10f838335bada8e963c97d6a4862457412ad89d6ec084fdffdb7beaa21b236e3a9d94f98;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19fb9302de21377050d6980ab83cc721cc08eb1656b8eb0ae29a2068ffbd5a973c0c9fb1f072ef41e1971c9e263e4d2f0ef0470d5d2e58099822a0bc300888add6742ee494dbe5b8ddec140e13c0f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1caf4b46f7e6967a2293b308513b0ae3ab37db25af38d9bcdf454dec33d98ba785d39c47c852c04bd253216ab8a77b3ef2b049242546075386f1c9dc7b4b6c4adef913b24d95cdba1d0861229324b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1581a569aea081381a0b2af71e3a27e5f662353ee155931dc9b99e59b4ac23df653ff65c44afd485b234dd29e43cd895afc56e05b7fbf6459ec0cf28f71777d84b8eab835c0c52fe916ab776fc97e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17f76580e578b86ebf070eb78597b30fa9ab82f5c44dd0d7d49c8dfe39d2439da2c078285e0e2dcf8d450b8ae1f2c925d54edee7ecf5bbe1a57661a5cc48688bde49b15a5c04d64f56bd332569a90;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16a7a041d2381b6835cbc272560a62e026ac977c71809d8a00fc1621b67e335a31957dc092bf8c92379aa2f1ed792630b5e1162d3d7fffd616bbf6de5481fcd3a4478aba7412657c334aa9ccf5eff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ab46ef75b68b32176d4a54d24a51be0bcb7b6c48c3edc5e63a1ffe5789ac4c0fff201e9ecf1647609ab4d8d9cef81e4bba10dbdd028048bdc452491177e1688535161624a67f02f7e5d7cd761f7a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1837c53af5498a42436d23f3b7c3b0fbce7ab1b690350fa5272c1f6b827c0432fd62d16da949ba21e9b2f9c31dffa7248496863575e655db56173e11023bf35f92605532fcd6ac70267a5cd22675e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a1b8bd4451a08c1748d38bc9a445b606e0d207c34615ae30059c887ce3d0d0d4d772d6c882f14ff40e256cb8b9245ed06558a83eab146b2022a71ca44ba28c214197edf0855a08f778812cc24823;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha18a45cbf404cd191f5eaefa128a378ff717bf1767338f3e623d46ba472012ea4c4b747c49c41bd11b39e14185fff54ad0905111fe281ab7e1245100488334915ee09f7a9a3fd614c27a7f943327;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h298a6ae2926d536781e39ff60c5a1b54542411edfe4a018ce32c47724c6c14b4e6e9946f1d1c006582708abc05ae84bceaca62119f546b53cddc06ef818d3004ce89cc9c194f8534d15f9f1d6c90;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h713e83af0c4b444b7012d8cabb346545131e37c1d1ed263c70ad3240c0be7d64be56db9447b2bc1cf7d473b2564d3f086e5907004e7035bb925ae8a882131ae63f816c85bd1f8ec7cd0b10ad1313;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1500b3cc93b24376dd0ec2631248e7dbc0d17d067182dc7cd7ce42c06eb2dfd410ce1e2c6f26f54a87d4c0f185fbf7608d96944ff0365ac11361487dc9aa8918f0a31f06bd6a71ef0e6fed40ff412;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7d30309f065f00c93f5d293abdb0bdcc25aa02538b19aafa40377a012728df8bea68acaffb5892f65afcf8fa64aff2c1b015ebf6734d9d15e57543b9bcf7d344a9361069092b322e4139ed21905f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14493e0f351109d9e4dd0912dff608c7b64658c6619be93f8345e0899af27f2bb3b715a7266f4a23313ef536fd247b7a3a1b51af77be379319dcda4c481769b2251b3fe6709b09df5d8dee4ed750f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h845539d574a1dfbe96073163f6a1b11e2fe28f6cd5e1550b17ba1059f02296563dfe8638c6df04b94641ff35f90b69d80ba66707d7e89c081f803cc261cdcb1745b10452a098985426ce9b5ae59b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c8a099ac8dd13336643f6551574353f77043e7d526782af6cc6113e993c4bf50ebef094d0e9f1d1d77b83759d0a254d21161591b9f9c53715068c6baa0ee75c5f2221f76dfbfddbf1067ab4a1b41;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8bb02f7ccbae40d9a544b3230712117f86fecb4d0772e5d837e2097ece8d44029f8b9e1cec88c78add4d418679ed55706a05643ae9aec197d6d272fd6778d2f7060f0acd73d31257252daa132f87;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16b00bfc04ac3e9ae85f3d0e9f9070c36e56751e6611efed08e86fcc7a0f87bb7d673cea577abebdb2e09e86f2122c91fa1ae7b5380c129f0138a27c25704fe73df4c42303933eee966a84f82d570;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcb902dd944cd3d5051620b94d91be4fc745b707b422e1ac0b7237c99b91379d52b1e69e389ded4f63a4bc047ee93849a7c9db377554207b7987b80c5e096920bba6092f9ee84c2f8164a28ad9b7d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h92cfcd2017b7dec898e11c34ea044e59d423a2daec77bc4a167b816fdd6865ede6a5936316967308be84a607ea92cf10699624e635a6c2e321f99c6476469bdd44d900514bdaa8f064c26789aadc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcf04c45e0635aac9883d661f4396adeb7298c08e2f40c0346a913fe8fe871c43df7a949064760f69d7ba3d3f854985ef3380decda55c5ab7fd69d63e7b2e4a7ba9c369c752f03eb5f3c0050174cb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h110451ac8bcee8d0627cedf48a8e3d1fd8fcefe604114a88d616876b8fd32dea6126443caea937ee6bfd0c5ea5fa05b55b18db8daeb8530ef3997b406175a7b4c1f1af795ac4f4b54964074a89bed;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ce0e1f73028294f58505e04f979a2647877b6c4e3150c7fe0debafd4041939357c7877662612b2e93e06305d7420dbdaa8e7bf5d35e2776256627d0cafcfb038ce588e6514543cd3ed41fdc1bb5c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11790e14ce3048390c2fdccce607621d021aaba7fadf50439c5c05a2493a9867df9968a63d7722e426651041424c6221c624306d5e76f7f1883c7f0bafcca961e0220fe107c188778a1486b14d6a9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h192b8e2cc4bb62a0ef238e9f028ab894c628c84be3f5767bc80ca8f6d06f38c14387a3f956de62d88b7c8e07a5594e8776557a053591651949e4200c829d7eeced5bfc50a33ddf9aef370a3327878;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hed5bc56c758ce3b7dd0fe5f293cf5aa42b6e15b89ca07703627d2e47651e47c6f1c3c86a51aa47cdf0e71b7c6ccd5f09e90492d6d7c8e71cb3490685635225540bf0d0888d3309cce2a4dcb669c6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bba085e493fb279e79c1a2b4fd9706d99187913894264a7a60273a0b56ca0872300689ec8913f2551e01eeea455112f269a0c6c31ed4729f829553579c52464861bcdf3ff0bd9e729483130a2649;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a2ead5cd6a93f5153b400b1a790eee9e8b7685f06ffd4084c7046934434e79e0dd0f6a755f2046bcef9f88864057033dc1f5467a460f10e22a43b8d1b4bcfa4ff64ac5d333f12f34a38eee90723e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbefb1159d693e5fd44a9cd35f973254af9ff4023fdfca97b29d857216235c67bb8e9e7afd8ac48e6f6e145f589ce0bb3bafa9aeccb003584b0e4eba23d57f7a1386bdb6e38c3264b484992baed51;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6c07bcb0fc8caad700d659011576b438b7a767c1dc0f691fdc6e2f34b217f5b4750f1e8bef8cd68c440556b5fc5b5731a6a1cd946ca92232ee513c75b308a6086f640861788c241f8b0000c3781b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2c9ed361ee6edbf4124d3ef332beeb0f01ae72474fe90f37e3b932567fbae24344b1b5570cb4d7fba020b1c7cb1bcbf52b88b2205940605c792affe621b10f840534b020b8d46b7ff692f25c5a25;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc42afdabb7c687af8a8d954ec4f79ca0ca3b8a3b64b409ff067b5529929b4907d51101c63ca46460e1e0ce0a4e0ddcd823f706881f64264ca99110846da418ed4fe3b3a6960718c8a99091240789;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h96bb2e1c1321d3866f21cb250b57a0aced7f6bfa36f1da9254e52ede31db79a1d27d428cde8c2a11b8e56bba35e50f0a8d46b73f9879dee06c80b97307c436acb9471a95d1f00af3d35ca5695560;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfe061e11e1ede5f6e0be365d14b41f3ad170238bcd98ffa06e52b2f9265ffd04b3f1ff3b2267c5465d9bae1ffc8ecc8f6bf3e97dd915912d094e4bbd162946618fd73e16f21b1bd3b4fae2bb4342;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h58f54e9a97041f63e4a5039e1df37c4a8533a648fdfcad237b305de66e2b8f2f282d575d2c90e27e244de9ae2bcf1618cc2feec31be5245394e013b7f11f595d5bf218ca9e3d3ac3a09eb763fbac;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dc3b83ff364165e397ce8d6d949eb5677a63f8d0c56a2113c6de423f31713a487a10b3b90a829cc6752a1d32c2d0e2829c97264d6ac59b40f250842234c22d6ade1040ae04e8fa26239b0f4cf1b1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6932ec5bd7a234b79f945176f4f7b3799f13643ae9ae961c5b56f1d90d2e78935f5581239f7c25d9b3412af8577fdece92ca4985a906c962f65d57bdb0538190c950200b1509df2e133979f4b9a0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18b69ed9be46ea91dace27090da0f720883cdc8e43b2d104225867bc1e9d670c36a38d8eeffff5b71a72a3cdef8d2a3604883a42dabf46fe417721f601098ec59dda91fe121a7214e5f61722effcb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1062cff91aae4da6a091ff39b7fef0d155ff591636b8fb05f06d313990f742cf180750fc06e234931bc720be9b6a5fc3773b0aa87a21c64c5b47e56fc20224760fa55314f7db6e06fcd2a0deee44b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h110d548471fc7925c6d3b6411fe3438094a1260e668ddb1be0877caa92584043a31594449aff3e6275bea142eb68beb7b4d672c0f80c1b69f41becb45c23024d65ee64d447beefd86e76aeac9cb6b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8966c58c5b061494d9f5c87a1d77033df7ae35f837c9812836bc2ecbc66e5596fe76ceecbc9711f994baebc392e3e8daa65ab8a19502d2475d3f21431446e3da42a28294425aa232b89a4494d344;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a92ca856fd600baad392ef4c93f05ad61a4a85ab2be6197911802da6bd030e2e5ccecec671844e0e232eca503ff4432a96e3c439d2435f68f551890db6380464fe1f14e18ab5c4f52da40f98b4f4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11a047c1b774469e7af594f51be8b6c8223fbee219c070fad181558e2e1b9ff6864ed013cb43a149b92fea1002d1c896c1e58e5e43f48579cbc60972f9732df009180486948ee398c17df099793c7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b55605ad54d8c6f1b77ec7422b1b9cd0bc821d6b1b74beef21d91aaa9676faddd06c319e490f562b5c8f83f8fecf3face46d749aeb7ccfc2cbb18f9064234a7e2f330ddbca440a61f08153101d1e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17b8c9f5a08c0ce56d5bc3f7d41a2c74463309a620617d42ee99c5632feaf3240f99431c9eb3d076f4a237a3921744ddaba592d62bff951aac86e7953b9952d85213c586e725152d55557128fa29f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19488a2c3aed94c026f825f4fdedc48faf5a29559ec287d8ce7f73e0b16aa0916851f4f5d85ad93d8087c8d10b59529170ebb89ac41caa68a790d757fe7838b91bb963b0d503cbf494d6e4a512672;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcda37c96ae72c73c2c0dd37e58ec3ff9f1b331c892353d0a6b8c2b40467ce193ff7c823e17767e2ef75bf7c50d58eac9e177868dfea4098c0e85558d37481f7a22a3e5b7024243d221c7cc059b64;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a9e30d7b71edbe23035eea37fbe406d4df497ef0552f09b7608b3c895a779e9c818feaf0dc7633a16292add60e433bdcfcd5bab69c6e3a1ecec59c17e9faee380b3e9d74bf6cf137d2633c0e614d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17a02bf1862ca1c0feaab23ef6e1d1cc89dfa58152784407df878c1c947cc3864302c58b726428ed692dbf624a4d8117613846aa940cb696169f18da7830d0ae23a96ef6da5727d4aea960631b6cd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h103c9203481d908d72d897cd660261e41913e293c7ed51c15c963c3392b20c20c6b48f1ee3c5d4b40dcbb0ea541a450fa5648ad8ecee511eb10c78cf95c8ad8dec32e220021c85e2a9831ce06029;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6df9f6e427289c43dc046d3e2d91a9486d24338df96b972e3e48afe115e18907399b8ea00f68954df7f0a0306fd47c4afd6c455d26860ed770b80170b8b29caf4e8291de0a4aeb54b8890ccc452d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a01754b25e990f8e3f55d89e929c92261a0523804dec9d009e341cb41d8539d72ae5933dd08e7f620c3e7f3fff5b13bbcacd0f4cce7f40eb8752835906c812459a3c7c71be346ae2d925f7aca25;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5d8ec6374cb6ef5c3aa740a9b19ecdfebbfb6f5dfaadc68024f25550d8fc57c6ab60a2abab5a6a7951d1315e95a707f758c49b18198eca3aeebf79b8204193c093dff6a2e06997c8f92855e1345b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ddf105f071dde8796f15859dbb6adeaefe02923df1dbcba2024a0c1096a8ba1c1ef1b61207865586c5244ed3c21c0d3bff875e5a10bd65199fc0e11ea91ed03be9a7b98a98297ff2f3b040064d75;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcc00d302f38ad8e46fa540de6ffab70febe84d05824d6786fb9baa8537b1e5a8dd497bce18ed625d93d50bfda6676b863ed219e845118bc781b81af310a4838f95e232b2a394bfadaadce8632f24;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a6109d57dc8e196b87d2f6687037dbec29818861f87222bb065d5afb168e2ba676e93f71cc606a7bfcb5b77aa3a0d7c7dc091c9a3ecb0f1dd1213d92202d575144eb0f84260be3a55383e6aeccbe;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7ccc49ab8be839eed090714ebfdb5c82b1b1a89fa8f475cb488adcbf4bf4d3f163fd9994319baf8d198912d2f4c63308c01b1bac3ca3478249868d16e3664419b8268a2930b01a7b831a504e96e7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h282ba797bca7a25db8ab87454498b5d746afdc79d39694d4e4d6015f16a5c7bbd34132868c09a4e67b12a2d3ff8f019b4eece76cab109312142356aba8b55d15a4fdf917a6d6a6d6593d7b870ef;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h101c64d27fe35fec2f78f1f597cf414073a41a98c285e55106403db78c97e2693484ae9abbeebe11ee3a47e001da12d8bbffaf4f27bf4307c181b41049a019a7c54ed7cf5a6f42027b4bbf94d6778;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19d43e62cd419784ba6172f272bf3a6ad16cae95f538ce1668d41aa57c6b6de93f153f6480bb31a649f8ad4e8193c5f1d8f8f8a096b1c5fe0c6b79f1688fe6a6ac23549600aab7e726d42a1267df9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h112d31f1f5e6d6105825e30d4fee69cae2799e964bb29c755386a268adcc7c0188ff4301d02eeb7a546371ab6ed49832237d64b40a1410d3f3149234f81551131e92b33b976b8c57595e13c6e7860;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdec078069713e7077deaa9ce53e99b250090bfff25aa7ccd5c6a978b32c687df98af66c45ccd623d52c83d71fd1f49179573831bb7f3361162d750f090ec93202b68fa443ead07a837437fd93c96;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5b3ac5838d84f7f3e8c92e8713c9e9351ee39e76b8584f23e810b038ec8cafeec30227302c41b67f1986bed97129001f58210f026c2423c5f6857d6f5dee901f247c9be5df03defde767d84038bc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hda725659017bdc94ed9cedcb1925b5b4bfe28cd99421c19e2be661474769c5926e250da5d76bb084ed069f88d0ada539f6d07325155f841d0ac3f534213212adcf2e224d9da3ceef33e2b79180f0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f1fc047e159fbf446eb57247ef07efc7be103e57e1e6592283b9ae5e2d4922ec0398967e710e08a4629e2897765f0212c7413a2ac4dd8bc32075a9531336d783e61c7f599650107e0b83215c0af2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h196c8e78e8afef616fb0ac1fb01014317b136af8dd5320344499ccf0f2bf5f70cdbc65a820cf5370358a22256645eff0b627a010b25626e255d8b0b0ea683cd5b0e44c7179c9816388df6a4c39805;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'had1acc5d9fffd1f7c33ea8b05db2fc2de71c049d1b2b816cbe0162cf084cb9700827429cd5d227216f4acbecd2782b3fa33c7df38873eda107150762f9a8a42ab4de9153758bcbec72062c2e5c19;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12a78d8485a56842818af7ff073ee29dc94bdc54e3f58a0b72622e3f187978b3ea33eeccd1ef01c46634f4f17dc268068dbc6d7694243ead91847091ae32a6eb9a53bc9c960b6fae6c41dc7a80eb0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfec82dd07d4856a8d498dd528429578c387f290f91bc17b1564b1df16f4ae89918ddcc1a729402e19067c168d73a8ee08c6f0270c5ded8083cfb7eb96063aa301bb9ca8b9ee95e55f221d6ffae36;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd4ae1291560e17cc6a8af8e9bd1e354d95b4fcec5c5541169bc2018b6f5f9e0a87857a519dc729c0005367a725fc7369eb67612805ff43165b31dac90e121d4e529a97fd53234b7170a48476d99e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h274f4a7050da23182b27a5bd5ac42becc9694db77c4c583a6a1a868259a4d29f1cf143497566b6593c60db6e64bf9f134923854c388f5d34a0c4b233da234304757534be86cf3aaa2afda4423d2c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18ab36f7e519641aa9b98f29d4f60c2aa08f4f3b60841c496ee51f3cb36761002696dd70c4ecdca580f73e96dce5a3b05d51634544dada826b761a703694c36def170530846b036a7598a52e5573c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hab3a5849de0471c117f0701e39284bf4ce5e07512610a063e00e5957b4ff1c0b1558da907e045161babcf552146043fe76e83a7167b49d7c8c8ea083cae55ba6fe3d6bd32f671ca88318e654be93;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he1a4162159a31ffd86c70fe5b5b2bfa92c7449ea1e7ff60254e11e4584a118518e863c8e7bba491a43ad10fbeb580ea09c9515ab8861aaeee4ad5e0f0d8470cab1e12baccca37deaf4887153958f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4ca89800b3520a5e0cafbb6f017fa13fc9f34ddc935ae85afcfafc4dc44981dbb706ed4dfa35499f8aacbfe17787226d634f0c4633c6b11b0b0be368863ad104505e7be12b53ab5068e61a07e4c5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h445bf778faee769af959915ded4db761149d25083d65698b74f12acd620dbeeb7cb92eb4ac3868f288979d466a7b3fae28cc9a6700e79dc2936fe9ab36a770091b595fb69c9e284f977c22a943a0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16439741053753d7b70c6ec658d9373f7bf2249cc872edf17dd7a5e89e8a0f4ffff263f1641320078e5ade6406b76d0c60145cfa20643343f9364c891d65172b67a82c5f5e47d8cb6d4cf533e8085;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11cd1828aa1de342e0cf79fe401fd6752e5a8db247df638e3232b84aaaa23109d3894fd7c0d847de87b52779c7b47bf84482a6fe840f89279426457ba3ed0448f2b81081e3193acaa7faea12e7f8c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3304ad124b3be36f155807037ac89816cda377b7f3561b91c53bb62112babc5304309ec0417ff07c7a1f74ee5a600030f1628a397cc063d2817ed1f27aeca2c898d105df6c539977b20e156d37c4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1606e15affc85c8f5edf94a8803851b2acb3d260c0a6be2ff5bee74b0842d6a7b0ef17d470b945bcb6dab3885ae29cd92a87340254ea716020c9fae8f76f7df697a8e69432c7168abc6da3dcc16c3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hde49425afadf8d0f830e9d1fdb17eafca79d33e548425ef01b25c13a2b855683b9542a1988c64161df098115e278fa7324de3f55506dec043937d5e9d1d7b646992a6b0a2cc0115f1cba9c298d50;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h186e371386e120b145b7a12aed052c2f2577209d69d1cce91fc9609c74b660f0822e1bdd269057a6d47c726da81afd62fd731c318f9fad3e5a0c1e334be66d4fd3c7fda5f29952d98c91138ce8c2c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4ee09e272204a1f6e943a07648231f8fa7382a13d2a03b43b967564d1fa3d60736d9a1fe2e678cb85ade93395760fefc0cf1964ff23d832eda5c414a3cf613c02f8b48656e2094abb00ae0ad1328;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb5b092c36c12b7499600c3eaf8f0bab72e72653d4fd58433758c5bcc2bcc0b5cdb2f0a7415829294cc8213e45503bfb8d85ce5432d1462d950af2233cd7822c01cb12de44b6a145202286443b848;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1107a0950bc97f6addbe28e4bfe0cc798e3d2f381bb4f6bbc5329646be2e3dd49007e97cdb50083543c31257c8dde4cf82338ca6d05f5b8eaa09b1362e4d30a7c38c7c133d6591de7321fb9a5451c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d586abba0e84e583a0c17770aac3449f7175853097145c9101c2e4bc586cbb8d4d3326107b3e895191f1fd02e6b368066a898a50a8e54b90243e948c50db82659b4b053ce6daa4584bf95dd17213;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h87ed608782db81e85d018bdfa79306a5cdd7565374b4ad4988772096dab6b043b3aa918705a04c5446fe2e4a49e3e268f9536a0cbd84c4e876df7f1811e1f47adc2c45063526da284c096b359c4f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15309f9f1cae25c0c8e6db01a52b8be3c59dbbef9c716d74c66e9fac921390747d7bbca404d3102b9d4f5b76bcaadfac438ce58fd7596bebfa703699dd27c7e767b0541c9a537fe7c23456c6599e7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10f1f063133d2ec07cf128033150cd3a01f970f15050b86bcc80d085388b6accca9a4f6af340e244ad36e812bd7e14b71951c9061b3848c7f34d8f4fba00baa7b8d887f5e80d8915acd19ee1e7103;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3c41d1a614cb8f3c3826807ecddde26da6641594372bc4db81409c4c9eb233a12ccfb26e89b8ed4b031706a5c86ed00c13c0dbe8ebe174201fd9ca950b4b7ccc9f2f4268ba05714942a37806f063;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hee03f0f7970ebe06aa59506a50714990045426898967b18c59efe4e8190bde86dce40af37f30f1e4a3388f2a32dc8345d2d31bb2c8541e70455ae11859219a53c3edcdc52553e696f6619e1d2df2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cdfa79ce3c8cf43b6d043f79b8742d7c9351c664696de65471266412db82b0d3f2e972d474632a35f279b73e8e52f64eb268e06492a0ffe89a1bec69eed92cbb0b6993285e71287fd80ab22887ce;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a1652257f9ead8c6dc4637c019ef633f27c3e7a0672f253a3c1c2a6ce9a0e40f95cf8c1cca59366fc817c40e7f3f3290dc217d135bdbb27dc2abdb12783ce6907d0acec0a83e2fd8a01086a49ff8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1586d4062e13819289bffa6a701327515ce59cb3e8c8a39e86394bd673d36e409e24adbbf6f696f12e033c6beab294f55d7344f3c78fc26e73647aaa988aa0a62d4ca4c4c656865773873c88ee11e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8738af74e588e7c7306fbdb8d2c35bc7f3f6bee8bb8ed07da76f81d43e01deffde553bf2a6ab2311248cd89f0999eb41fa51856433266e089a8cd1dc121c0474818c51ef8a5234e69056fdaa2240;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1076584cda6114cc583e1bd7bdd9971d44c16d9a60e5cbc5de30265dddae222d5387b773e217f781ea7eaf28c76fde56590d616463010938dad037e259746af2cab12819b4a4a7888a91b203df3d2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h918d992db30b9e22820dcbaaa63adcab208f993271c80963fbd6b711ebbcf284bbab8a056f01bde064051d9d729176721f3bd90f41b6139eb1a0d2ab4f5979d6a1e1fc23eb7ef6544c5f18813ab;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f4c0cc7fe0f7c0335195954a0751071e8f3182763c20fc918e74048095582d58eceb043303498fbed295d1a72edea33557b72c660f55a91c69a34690606871c310b9dcabe27669ed6ea17e36e368;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c19d2b8c3e9c0ff5ba961ce840e6a363f5f311a492505ca9b0412bd84e5db7af3303ce673dc4b4c52021a56e6f1174aeef42caa4eeb165a9b2c1fabea32dee38b46d636db19ed8b5c8d206d8ddab;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10a85180463400d275f75e4dab5b52fe82703f89f5474a19538808449400386d230234cc2e37f432137ff0770fb228f56aa59e2c71bae6bf045588a0f9b8ff40161cfdb56a593d12f3409322a691e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7c5bfb022125a59240b9e6e1811d3b9e1d790ed212f9f5d8840045956e6372cbbbacbbc265cc71aae84650a898c69f0f1ee56f78d32077fcab95f43355eb69c4fb2f79c4f3aec210c4f2a510ddd4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h189085a5e4a77bd31f2eb5c23be87a0506580acb89a346c45521b8df51eabb93273ebe69dee098cbc4d769221311e00a5e8e94eff225900ba889d13922b2cca7e7930347141c7b48c50e0b779b866;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2a85ad0ea6b3f17b1e1e78a467025e34898f047bc640fd512cdb5d067474fef58e9f40de5c6c380f87542919d839b9fb639123698103b9b416deb2edd5c00a796512db86100061132ba17cd00086;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha80c1fe9e512e2daf4410d85d1acfb2cc41f31102c99f51c8b907ad95b71e7534f1863ef45d5dbe7e49c6d5d60eeadb30128469f6d6ba3250b170c317d3e71d7709dc252e0577d02c4d5439c95ba;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbd6d679235c7a55f12f9fecdf4580230f2bbbd111344feb41b9aa9bcbc471457fce6d7ef2ad1e84d800884a36199945ab7f2c0f2c4140798428c9fb918deaaa75ba45e1953a2bc4d28233149c6f9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ac31a2b6ecc2304b4bedf6aadc7c12b750c5d78fc593ae474c86e006ed3889e5da2f6256951b81096aa8e6a49562c12c2f7fbb32db7b3b55303374d97b2bfee8f42f76afde75caa71acd21bb5fde;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h177443bb0e9be8073e324067f88390e10d93fa4d1df28e72584649a8d7d07403a9776aee212c53c845e6ac06187a914a0a1f82a6e3d70403ceb24449b0062ede0e68d71161971301945f027536ec1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hac327f44d0b0dea61b3b9ebecfd22dc4bf05f2b394481a13d6a1296ecc0fdb7eed2d20645aa754e9562bd751cec8d045b612d5ee3716e8cfa47cd9f6ba6f51769c9c0f4d9f60a27ccf1274044526;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1065f014b8f4a6a16c58c40a36e83f20d3d85adb3af36ae3820399d1bd7de86046e2351101cca817cb380d4b85dc5a748591d4bca780c96716af64408cbe7328f0efe537f77a20c879ec324a0bbde;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f3ed5c39a1344d938e1db6772a450179ee79621b518be22cbbddc1ebe26017bdb19f7a3c55cb56d1780932422f96468292283d21f2e56fbe98b0f466c6533c6741f508434c8e1fa85be9aa5800ad;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h180fecdcf222a4cb0df3fd3bf5715ed834edaefa0f9fc7d94ac6daee64d60b87a855cfd58e66d4691a54dae06f93132468e698aac25e56a5ee42495fd606677486da0b16236613e69a4d4e259c8bc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd2a333e7f23d460a53a00436e7ed100e05cbed54a1d1b90e2a4fc30b6e6e8a38a3d3fb777859b7a432bd2702330b41d3dca992a96b9a18ed28301037e1b5ea45af79754e8a3ebe99f402bc86570e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdb3b9b24917474c131d8c125f7b766ddbe7217d3d0fc6699816d630d44ae4e4a4cd0390d9cab32be05be411eb482efaf4da65baa5f019123b25f86380ddf5c6b7cf5364c6fcb7a8b124f106df64;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dcb34d59ac216a2bc5f41bb4194b1413a65ad3d940cb5193cab9b263a1e0f960dca6ed08cac7ca4fe702a7f8f38839c0f914b10b5c21ab88e45449f831bccb56aaeae57cc484d09bb8370316599b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h31710df0f811a11e3e41f34b78aad844287e98614433d286a304b09c81663e8f5e079a202a1427d5f8e6e0476028659c5938d406f180584a5c12d80c6672f07fcb76728e58bf337c3d9315ba7835;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb00272a0a66556ccf9b1a4045812a22da37b0c306278239653c8328af8a7f7985cb6a26cb065611ff8fb87014d72082fe801a098cdc1a489243df73d3016ba7f69eed0211d13dff695371391d3b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15d0cc20eec6260de82ea2ef9d8908e5d5946436a39293f53d1887d6c035cd5b81dd42da03c7c8b90756658e28add9c1ebe04d4a501eefe96c2d9c3b9fe427c36642c43f6acfa52864d9db60a3f2e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1902de15ce6d4fa9707632d1ab7340132673a0e26114d910f5897d52dea9e799203039467630d6fd4f1b854d8f544b6a0e4b1ce058953e782dfa745f92ce2493d1103c50c7a588ab121d5c0bb0f9f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c17b9b68a2012ec4a0a272c0fbadda3af9d4e97655c615fed961f2b5c4771e7735c138305d0a8ec74dadd09c7eb110038642dda7e48e18c6f286b3bd79d37be34a2eaafeb807e970951933b4b5b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f104b12499f8fca0dca92a299d129f1ab5a176d2ecddb901f45ab7b771e73e673f84afdb99b14412a980675f6b83dcdda9b9dd69513af95b48a21ca98c877a55bb6f3aa8fa1bd848e9301e44f4e1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7367a71feee0e710295574ad083d7855780e2261fa9dff9eac788b126ba89ffe4d8cf0270f00f20899ed1a70aa00a8c1308fa3e8a126cd173e9f6e807fb6251cb03daa912daf2964fd9fdb7a5ce4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h197b8708fb5b11f0232728a6c5341e09cf6febd5a0e5c8e6dc498f295b6d068c0959ba97dbd3bea6f032d2a2d09002ecf0740fbd29f9a2878d2333e505874d5f5537d712fd53d173954e13d2e10b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he1f1025fb2e57cf74b4facc661fdb57b3828e493e57f439be3858e6e6f8cb0cfe3299830a21aba44023aaea5b745f08d7bbbf8ddf5d7d9493ece514c0e213dc9fa738f6f6bc5a157a9411c6c5c7d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h67f8460b448f1fc244ca4617b5636d52dd4cd6a076d798217bcd43d826c30a61ce98a4f07b1be7e8fd8713c136afa36271b9c29d79dd076070d1815f47491d9d36ee1759c3be2b7b19d52ff981cb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hef33022a8682dab030deecc67e2e9031142c4cbe7af55791f85e9177b7c38af8bc0a5b406bab02b7d67a953175640b7b7397289e0554cb045e15f5ce82f95ef00661da408b0ff2847489a694fd7a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hafb4ca1bd1fcf2928732c9742fb1dc71006ac2cfe6289fc78df13018ca93538793f7b9c527e0a11203229add5edc275a5ded76fc4a57979bdcd24759ddb52a389721ea1977e7f98a6c1d79df29e7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdced6cca84954ca3425ee8d45e80a689e225ec848f77a13d3574c1af8ee991feb42dadc2fc328a05e883dd2c4a2cbfd58367bdbd149718fa9be5386523f3ff33886efa05cdacb383aae1e0dd4380;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h164b8c1b19b1ce912dfe028ec320621e6ade08da176861b13aadfdd73f3e0fe31a266dd5e72c3a304f27c48061af288fae97fa35d119a63f78ffb6f6925c83b5e6bcf51b6035b2cc075abb9d80442;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eb2cbd2baa1f22bff08f9216bae97f6631da206d836df9fc606ee07ff4e516f8df934fbfe0decbaefc3a3a3d35c130d94080d2690195a5d2bd9177f003ac9b410afd99598ab2526265113d3f9314;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ff864787d5611bbe473fe237000db73b89e6be7fae3f01476a5a4a16e1870a3b9db6958724ed077b2b1f84e2410a81ad5628395994e2eb51b7cb0b6e2b415d4334d93032ec8de9672fb94688b17c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7c1109cc65657c3252d63e3d493c8b6d88124fd482ee66ff5d26f64a5fd6f4b4b75733fd5f394340383ae699ec08baabf192dc25d8e99c13b3c2271c8d42d50d62cf5142a6d50ad3bd2769170549;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13ae58c069eedca7db9bd97eae556dc201dc6ff9bba7fbbca53103fdf5f8e1737a160a1f5770aa1fb0d58bdfeafb943d732d662fe7519863c9571e6f7bb1deb466a19046a3241b27e7e11ccf47490;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11b4d6f56e086cfb13926ccdda62b2f59b1a2927ff38b9ab3efa65b44642ef1c9f337eda6a906d986eec9eeec229c5bf429b35713247a873fe3b4562f3c1385498206f94ba6a2a9b7466304d3bccb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4d6f2562b13c68726921756ae45ee1ca73cc41f3b02d946cff7b05bc81fbe4f38b9136d7d3dc232bd214e5f2f212999b99ad5607b0137b7a45382052363dc4c27d36c9f189e6f0c059d9347b1aa6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4fa62f293f089f0d2a6ef0121c979874d464f850cd88dd8050a7bec026bece9b5a86d1ab7d33688d86b69aa3aec4580ff2611685a4af037864931a0cc743270c99aa5024e894373e55c46518ae81;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h362de6b48dbb6d8a0578418655dac42b65a7e1c303b5a5586f1a698c1fa9e17f9fff7237306c2e054e8ccfddd5d48f639104d3b9cff89271cea1fbc1f3e1cf800d0cd49e285d98abd0bd60fbec0b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h907ed8eabc631253dadb49c302c684f176f638bd2bc9a3cd72c0787a3c888373511229e3406cb8fe09fdcb216712b72d01764b24dbdf8d372983c20f826dac185fdf55be3ab9988211af1a0f4790;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hab54cb5f1d172934597ff1212866940f8b61790d7c351b3101cfe189d1e62db1f68a44a77d2b4579dda2a6db105f2dd74da6ab0aaabebc9396284e4b02aea18b056ace2181ee976a1bc4d442b7e3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h76cf6ff25721692ffef4661cab041c13253b70b6c3d2bd249a820ce9e233b7d7b8d8bec4dc5559ecb29d51c16b7324be307b0eaf48d0731b13a31a01317532759951b588aca7e84abd9170b76934;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b9129541d3ffd003cbaaa06d3cf6f47f9e113da62ca9e7c981feca7fcf3ce0385a1b6c12f97b8467e8059dcf7e3c753643c5a07d000b31f6de10d41928ce13ffdc2702b04d6d31ad5c9f0b914998;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14558fa7786d380949d1070a41734c3901e3a37afdbdc9632502344050d86b659a3ad6189164311e17c07c540f840fdb2be5bc5e21bf806fb0fed040fb2b875722b6839c7301eb645f16877d51e1f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13c57cb076eceeaea573633da85111ff6fcc0e12bede14bb93047fbb6e70b4dca74e77e7e30622525d6fbb82488509dcd83ec05aef6934bd91c148152b2ebc2f69e8ca1fce5216ee3220118dfa7d7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2e7f96744ecfbf0cbc778537e9e067cc471d219e4f085cf0f1b951306e94904d12a541f99292ead78e91253a254251f8b200a19f76f3a302312bf1e31f869107a9766ca2adda3afe12ab6bc0a7fd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he5a546da60d1253ed1f4d72629d5c1de0f327f10c7479eb9cf32fc2b741de0aa745ec19eee6247ee0fce3d403b77dfc077344473148b63f48ad0b2b009a5314f411846842631de5c539b2fa8b4f0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10bc04416cbd75a2a7bf4e747001482822337f3537f3f1475a13386a2db401cc3f1ad11e73061e9552231ba0049d1b53ac663f8974fba93aa3f386ef3274ec9271682488fb389e609e9a6cabeb23b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfa670270ec3e3f5e25ebdd29c3e27fc10afd0ed4f31e21726247e315a40e81d9ea58be0efc1c4b8e910203b66affb91e364edbd6b062cdfad9ac8a18c7178b60239805bdfa0d0914e7d0c9cb1182;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h84a1e44cb4706bf7cec15f1e707e3d21408c2d5c4663303e8b1a13f065a42c5a2e7ebae65c4c0d4b75d302be79307ad292a01d1ce9a7f61110308f95917b082b7ae1fe72e04f39425e36c21457a1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h494732354b1a010554da36c4ee76fe0d1eac0e2401452d42671e58aa175bf3b0a7ac9d6b822f4062f6e1d3dce0a3f63a9154c3df4d4a32828013678c1b5d51a416298b9831d5b029634acdecad10;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8ee89a85a6882147374dc263dcf22287318b45c344b31f4a20ca03369663a78220e3c1919e9269090f6b9590f3bbe4960d5ce69ea767f4b5b013531948d8f0b52059fc6b65af74ca4077a3ef94c2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h455bb141d1c678727d7b918c95e3fd1ed75a2d24f4a834db288b46331b8dd40fb55868c93508f4a3e0dc30ce3ad3d0feb5991a67282385174b30c83954b9d679c582efd8cd83452f4064e28c7321;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16ce0e1168deab2ba8c78ca8f3702758bdb26fae78affc36dcf246d8dd8e576aec4f1cfd9b85723ac178f980f11d3dda037630526f96221f4cdb274c6329a7d64cb3a666625727b962dc59ff60f5a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19fe95c71ee1409e5c1d7795bc12de43a955843fe1089d3925b0584d486ab0a72017de63770a625c29196a2af232d9c1e980655e7fd403a588d68532a6246845ea383b2a3bd35931165f72d1396f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd7b3d14aca5f2d56479a62743a8c767e50cbc88277530a7a4c7489966cb039feb7c532053a3d17002e512222ec098b5d704dafa1c35c9850a8dd88f652061b75e375a81adf522e441316f7562896;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h124667629b045aec0dea9822498897af006e2f6237ca2b265b8c5ebec42f9c01d6189793bba31c16119e4b9e2011ac61391d44d7ca49b2787749d966b0392d7bfe4abb7758ba004bead025bc254fa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18d600b839f209b5fd2a524f75eea728835a040999eb68c3c48994dd961b832feaf4b2484a131ef65906763b59f4856c5093e3dd063457a4cc7a8e852e16e9c1da0dce5876ed72badc839c947674a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h35916c0d74081167492282425fd483745578e47b1bdac23e994a646324e578d9660cd98653709a466579e50e10d591706402685bf40fbec1bd78bb8d1959dcc4499c916123a4982394b55d7a6f8a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17195b2c22c806c295ca84a709e9ccc4cc1a9c5fd0351c2842b4bcb361f9384c4d2386fd44e124a6b5a24e72bf06f922512351bfab96bcd82d904e9085ffd976977850e3693ea670a21a985394c53;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc254fc7a3b2075f93a2e216eb7812afb8d02849315d8e53f24ff78f9a31819cee6a9273dfeebe5bc4bd4665a1fd20c61277b3de439e19b88765ecaada0dc7670fdc84ebfed1e78fade22bf568d0a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bdf3159a2391ba650e1dd401d5c80789f4c324cd6a7305e3defe12cc4edab0c3dcfd29a4393054e9d650d18b51a1a0257f03bd5527a0a40d243db6bbe64ca7ffe3e3369a856d651835ec737a4d01;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc38a33f24d18953975ff2a497a399cd3d12c32fb6aa314ce256008c3c3d1a736bbc0b46896c6ab61988a88908a90648fef9b04bfa2b6e56adc9c8a9edde33738f1b7580fe5468c77fc0402ab6fe0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4b49fa0776b305290c86cb855ddbb7eaa1b39652d58cc40a713c220bc8094dc02cca4100bbdf3136c83926015ff2e05f5b84aff14c5b6e9053c3c418f6308de2853ed7b90dc6eeed08764fbef72c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd6285c8e0d8371a961a3bd9cd87508085511287cf731f750e3c503a0f2a043dd75fc164ce5ac11378151e691d6d5e1e653651b284b3ecd6c95b235b81de6beec02fed2570f92a07c2d174814618d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d80060823b5368f0772433edc090e090f66a49fb0cf90115a636a331ee631f6b4b22f82e550151a3fa7b36bb9c56d05a268ff85f519893f080d81888abd913b09c23f327f37b7af4cc4a25c9ba4f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1784b374a9a93f5fa8e8ba4670f9a3a69e349d6ed12a23bbb19f153969bc0c6a3d598b245cba8b253f38049cb7ad4aa2899a4e0cfb21cdc91fcef4892f15db778c94a84d570107c1a75aa871734bb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb2312d6aeac2aa61958d1a40ab5239b61e2a87541c909224c7e737c73cd1fb8ba188e49bd9d14079cefeae40f182268ff6d44ce04a107b6cf4ba416a316b8ad2417b669e69dffab14ba623d99807;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h43bc76b7017020197e3255f339e20fb807f5663624ddc289a16b8e62dd6d1fa6096b070364106d3eca99f561ffcd432417617e6c66e42457373f5ce3633d232d1def833c581bff649bb2f7740959;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6a44eb278aaf0c352121e6317332c21b12d2f1d02f30ba76f5f91ce2fa6343875fcc4d35c169525486a4aa497e5c6ed983dabb35e9936ec7a8ec0e4d6ef0881d81c4128efc9490d6d644c3334444;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf64b8b62bf418783d3afbf21717866964bbfe2512b231f62d8a1a8ac0ddf59b81d1121ee68cb65421ee0e7b8a834271de4163a216a09a57d927c3dcdeba38e97f713daecb23146b364c822b0d576;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h145d5f99f07d6d41f75926d7a15553ade171b16bd4a45e538e3e74ce7a0ac0f1a53bcb7a8aec3a48a5f5f2ac986dcf8fc8cdaeb7d07b866cf876273f16dd4bc0de34dbf235c85c6f7bf96dd0dd7a4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1029ce553f487650cb07b11b737aa01f4d356e0a0d21eca54a39bb58648d531f065d89125e8c7bdd351e48289b0d0ecda2359c72e59d83b7db77d7aa1846236119d3a9217551de17f5507a622eaa5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha49db32b821ae2531c69ac78b788f7c9c025cc7366dd8dc227095585a39d994e5539bf2a089e634d4c1beb59268d1716297178d801876573f58f1cb20ca5859d03a2db4cb7fc5bc1d8ac231c3590;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cb304158a4404d4c77e7a815939a8ad6f9e31737c558bd42c52a7c0b0de609c0ab5185fd71c52cd42a5ba700d96b782af247d8611279d6aac4b6e6f3921f3681e3ee5d8f86f00c425c58f2f82109;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a9d70217b5f9383fc6ab1ef2a0e4adcf9af449bf2ac88808b5f7d9d5cd1c9ea32344934cec5d857e56388064a33c081b3b15be2fff1bba39cf84d009a2505a878b45b08fd55707e5f3a254f44bf4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13478516f85245aab410da553b0e57550e5aa28b335b83b6237860b4b3e7f3bab61c291f380443c57d0655a9afdbfd3c31427a7d489fa5069e9440af8984ff920ab8a688c6d22c0569219c63cd29c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2cd7f92b383b158956e14cabe646bebed12abefae8feb0609e66b5ac5dbf2d8a539bad9c37bdaab004952ca64b203b715f402eca9cf06f45d27d72f4acd437cb0689b279cf275aa4204e7d13fbd0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16e35a75ce39d343b4f03c6b2758c14407ff5835e778dba7ce6c04842787ba6f7d2c2230f403815c382ef8c31c00fe2bf24f66c2183fbc0bcb4c080c988d3a99631745f2641584176dd947ba5218e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b2b00ecc51aac89239471304a92aedc73cb27b761782d2ee47ad8aaef97578eae5fa4c81e433842400f1881d75a3fc33f40360636144ad15ea7fbe7564caf8eba32bdd170fca8aaa70ac5432f68e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2b15251bdd8fefca28a07f564dd56cf5b25bd41db6051d02f443cc7d8bd848657e594d3788c5aacea67300d879ecdc3da0e47dfa423a444c819b290ae7b1ea9ebf36cdaeeb3c7ebf71bbe962b901;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h41d96d091087f33c85f9a024c01a730b8a509316c8a74e61b22a4674085af1f26dbd426fe51971780854d357d3501cd86afdea962cb814406a1290f51c96c53e7ae625434d85157a123e17c284b2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13cc0373ee5899c6a553ffa1561d5589890da21a37307cabf0f84bb90cdd7465fee4c3d2f10d4b2edb15b40ee7a59cadd10a6b5a234ce577b844555101812049b886fd1fc9135c06570a32b892bb5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7934215467f4f2f5df81c0e635b11fa3a0ac76687940b14029527b97729ca2d5471b146b837befc48ffa1a36a6047151cea0b152b951b35b5242e5fa4e9f8d2aa3671daffc34e68615ca9a90ded2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7cebefdc36bd935ad702b99399bb9cfe6923ebdde3df564f230a572a4a6416c473c3bd5cda8fab0c98cf83a0a0b7fc160d513e0cc8798faf563948d9d6c11210846e5027cf773b3e670292199cd6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h136218359707fafe85a719f14f8e574ec31f9cfd1147697979073e8baae6e23001ba7bb75e7f9e3a4c05d9a1256982699b924bda202d2fe9230bf784b2764f820f026e4132883d67435b956e37d81;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h171ddc76ea2fc91727abe53320e5f96131ededc784228a85c589192e37d5bea143f39b181fff684b33639c0a088fa3c2b2d41d62375f76569cda1a860b9aa66c2f457b018fd00ad16fbee1fa5d2b5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hea7e0e853b4041144897a31620440b31d7726022d5fc387d9be6415712744b370d103873485a6a7ca760f1f7bcf44de0947a84d49fac769fa70e3c82bb9471a25e6c974fd4de45a24e70c6fd1127;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2b595de1b4211795141ff4461e62b3ac00a86ed432821391ba7af082823ddd895685a7ed4e4f0a0aea80f646be2441414278a03d1714faa5e17bf743ab444302661e0107e9ee17db8c7fd28e1d8f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1958002144fc11f1bc72c7cfc3282f1871fc0948c338ff1d9d94d2e244925d81fe4e645730d6ea886bd513d8c94f145f615f7340b9378fed1d86f5c98705764cddf6ecd7651e5b3936fadb66f984d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cf2b4c1cd96ef46f8d568365ebe018506f7d71f1b6d46220494d0f8fdc3aa07132708de613d8ccf67e7b7180049cab30fa7172ea9164a7b8c5f93f7b66477ea84bd65207dc986fd891c6f73a1fe7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19b91d8feb6e50d73946c418d305240fd2884757c9d5aff911e79ea97f8b7366bc6cfa73a621762034e2ef7b623eca1a9fb8f8c0ba34ec8982c4467ea8fd59b222976def8e222ac210594b26ee315;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc42e49debe7b90836837bdc10d6f3aa70cfb5fd9c532e60dc7effdae837c9238b6f4373b2366c79c2a365fece299064e7782cc7553f24469e2f91c4c024fa9b77c3cf1a9e2492a33de1b0b25df15;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10546dd2ab521e7dd467c3d4f2d2376017635e2627c35d32dfedc3592ccb6943e56408511353079ca87662f0ddc05119585d136898b732a30275cd180a0d590a3c75b25a4889e4972bcd54f05600d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13a741ca7c20a97c3722eaefbf6da3db9626f42541ec30e7ad1b7f98e00dec9e0e6350f20d4292665ee58814851124c4106f847021efe9135112e826b2e107acf6ca0245016ae1da85439b0a8abd7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c566ff4ece3eaf49394b6bb514b1c3406d6a450b9be8640464a043a247fdc01bf4b7760e2a8a8fbc89daf5e7dcf3b5d7e8404f73c33b2108ad80d3df3d6c96ab6fe0af9bcc8ed8c5bacc40fbaff9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13a6daf3cbbbd9e8488a6c378d64b40d34db5ed8c1c3198c9e60c572b1e296a54c7f023e732c342246e4d7b55103cc12a80ad299e02693051eb09a366e7bd4df22c6d5cb537cb4cf2280178fdbdff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcf17651d10f3d7381082a5eb44b6a32aa59b1cc8e66b2d18a347547c51ad00548e91a31f677596cc12f87a7573e735dae8b3f770afa3070f2ee53ebfec4b2e90b219e067b9e9608c982e445a65a8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2e2a1633c59250ce794dcd6c53d94d35e04afecdd3c3984108212e98eb43506aca52d40bd064dffce5a07e795baae197f9edfc9238f888e327896e2048867ffa7536157ac3f4961db41461f290cb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b88c0aa93a2df1bfc31cc0b13f271d20f954bad6f03a763c75182f6efed728a92778ad1ba7242d447183e9f3c89a71a5ff5caabaa2cf0955db2bf7ebb10e39c895ec8f4f51c27deeda528244f489;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h134a1fae97a62eb9228c35d0d102569937a68491936971c52ca43baf1be824199ee7c5b774cd2f788fb22864149665ffe44b3d710a1ec85eb10db0f835861e72fdb8a9882952c8415d0a37d0a8417;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f567f7575a7b098d5ffad3925a723f6ba14e1ee56d9f4506f8cd1b5332135993cd7a35c9f90fad745527e5324878e4b590a551ccb6b2b19f83d8b00da9d04b03b1d90dac726ed2a84e8cf24715c9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha95ef408b3bd5ae1312663ce2704af36dd6eae16446d60190dd42fbf2f105c963a89d183cdedb8b0b1ba53b8e801d9368a514617f86f9b1823f23727f1812abcdb2ad84bb2cc155225c4f161ad5b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e229903fd6bdfb2681f4476083b8ba6b7bc5fa0e1d89c92f28ecdfc5d7bc3f7f2f6d8b18d6595dfb2ead05590133a64cb226b418124195770933fe1eae162a3a67cb9621967e85c98282657129d9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9242279dd4678ba382aeb016a84ebd3bb3591c8c42050b3b8938d0b9a93b8ed3aad7cc4dfe707457794edf2f3a37c237c07f9c54b029b58763fe7cf74ea613becf644f226b5b46613002a34a6e9e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1736ac0013081350c7f7e50bdae36a7691a1cb5e45362a23f37d4021fd073b3b3ef323e88ecafcc0f963a1fc0a031b889bd20c94a4bd5611b3dc3469f9746748a86f64bd2a123b6b63ba7d7d1757c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h30435bcd0fd434dd6e968c76eba6a1fae02b68deefaafa648de93595bc14cae87a0bbd59f46d9f4a12641077587184f569c322681ee0e313c5a97dbff179bec17e489a3cdf70a284471c4e64fc36;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1146ba92f98dc57f8b976a7160a10f8be71d69ce7f80941dc86e9cce45db31aeb9cefe779b553f74471fded861efe34f3aa1937181c95e4c1e696f7e34ccdd5baf74906fae75abfe4cce164564bf5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18c3de67f25a4accebc9fe71e6451dab91b6e90ff0a370e5fdcf62ed38018ec27ee2e233b46bae2ff16aa943d652a44737a7c3d5c7d5ab58eafe4392d165f0287f51257edc83fcb10cc35a977b6f8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h183f2175145c260137c787b2cf0487bb8c4d212d06f26a7f460268c8a6d4e39d29e626f0724d5272c8171c169acac173d8d586e39c76450bf930dbfcdf5aac599afefb2bab6b3cf3d1314222b8e8b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1931db149523a1e7c261693c5be1fda3350119765a59b2b231a747799ac2baf8d1329b1834407f9b8c7f5fcc80ee372b7617afddba197c5b745d40c78df5388567c122a71b3259e836529b1f3a81;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9565ae24272c8df3cefaca02dc8b40b1140da184b9ca442fe1a68fa47e1c0ac268f8fcc37fd0a2595a4eef5da9f9fd8a773cf88cce085e8574eeece40cb71a0160025a44997ed40ddc74867d1d6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h189a19af98ed83ae62746a558fad5c8b4e50acb640aba842c0a3fb7642124c343252e2720def0c781d47de65a063f2f8982442fb20fac7c4f718b30146f766418795d6f790e38e760be0af4ad8d77;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a6aad1f56ced5d2778ca36ce07f747da3d517aa87c82a7fb89aa6003dfe4ea9ce6a67a7d7ff35ef682dfe222e67d8070d1179bc00a7dc66a94457c35c8a333b6d389392f73dc38e4d01c3a11f79a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1582b138b11b23354a4d127f88a4043811c751ed6a7a101e5c191404657b1d990da70c9980a44f90c133ccd847b2895a85b9bd6da3ee1b25ad5d4ebba1a6fd2285ec47cdaa3af12de54fd84fdf283;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd129333f79ef75bdc04a75c007e1a255598db816dc9e418de52d92b1ac7b1009304265c605f93b10b65d8e496032f49f0e87360713bee27dd49af953568e829eb86bef72c361010ade7e5fb9a6b6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha0285ca6b97b9acd4586c3917725094eba2ad11625c57c5cccc4f86ea9617a38af5e0d66b6647eefef1c80a605adaa006afb977ea65f5303b78384359f3e0151fbafcd317f6f7859519ca0727016;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h149f0fe4a65467fc960e16b8e7235bd22e90e951807ee4d9405d7ee277202895ef0493dc56af263dd6aa69507fc90fad5a2d3889a29969a9afe7088a2ccb364acd144023f97dcffd62b3bbe83b1d2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h193ae0aef1a8b55b1a3dc89a9f8aa73b01ec793e2cc0aaab5d36bbc740a65b11213a1236963ee6b63d0748463dbe70afbcf033dd3f4499d0026c1bb46ea871612df48f9772ea7089baf5520418163;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aadc892cfce7e0b898f4671e4f6e20abfc01078d8607e9cd60010ceef9297ba595f17622ab9eb7971d75d087bb1c56c46a6698f5a5873902420cdd037d82fd9a016cc68941a8225665b4b66ffe2c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d42e34d7a2a58adc0c2f6e11a5c6a310798e55889bbf670d5d81ef6db44f2d256e1968154b2639e6ff9bd36da5644cafd158522f6e837f09404bfefb2209af9850249578730c8e26c1bdd94322a1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd7ba43e1343b46369633b1b8e984261894511a4bd7c4b52002eb7e848c25c8af9696166d02e519519c0b063ffd91632a46f31bb71529a74c132384be0d326b9a18c81cde0268766c4fb531b792e1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hea7232c2c7a76eaa0ac21693fab0ca8ea16723cb2e4971a11fddbc84ca4f45a2491693c8f003a7dc0fddcc5fe29205b106384e3e381b1ef5653a615be968d7f80acec6aaba289bbccf1b8cd0a588;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14828e75263cf7671c3b2c4a579f58bcdacbd28042342a3ade0536fec3e55941560c8d911dc0f0fa19c1c5ffa2fb2d4625456190e23de820fde917190b5d56c03e02c1d593c8ee7846fc06f15dc54;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h57da1827282a227ba92176f1dc6bc048dea5d6b66d0e73eb6001469a99106a30644d014f0be4077a9ed706a1e7d9e9b8f9d3975d0a6eb7236c61c3e18c69a4f2a467b810a9610c86ef9c7631468d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbe6556dfae71530c95301fea1da7430a9b8cbcb1ca89b98e814afa50484e3eee7cdb77988b9c4b90c0ea0db929eb3cfea18eb238cc836c94b587392bde8eb7ef7b3af13bf741e11cf3b360a137f1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f64c9f5e6067e6d06539be82e507e7fd20d5e3bd6e04de92ad20e5a14b26e1067e3cd0e2df2ad247105dcf595dbeac893bc2836194c4be6b82246187d88f76ab3d32dd59809932c8d45a3374d9c2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2614d5668d45039577e29cb3c86cbf7825d63dba0438f6245617599ef062d564e1b2b91ccfbd4f4dbe853ef957c3b242d778ea1cadb3ded8a368afe96be58c9d64feabc8077accc5877a3cc494b5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h71b0b6c61f0eea0c3ab9888d0732ffc6fe9d9f0e5d1d413846586172f8c21373b731d786edbb841d03b1bb0ce5d9453aaa155d9376457bc00a287f4a39b5ec047da1776198efc67219f7af0a4bf1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbfa7465f30e354b2092e6ae1d5bdde4085c6d5fa6b24bfa1aa7985586ff71c5f9977b16387e7da577dc5a17a952341f01a24df9c042159b5f35616dd9d5eba2157d8b0b953c34ca50774989b91b9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1893ab071b2b413bf287412adeebfe5aff1e66de1e8ffc6b8a1bb6fbe9e49601df2cc580619c382e65f0f1be93891e55d1bec3c31fa9192d8cbe8294483e7dca146deb16a44488387fb60aee4d900;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfb6a3609855ea787abff888b30d4a6a548ab40d16ab904e0d93d78a11e8721cb0d9a8e2b7044c374549b52a468baab9d592b9a4fde388772b371a41b54ea22d82504c88b0071bcb30ad4cf36b36e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h198eed54a91287cef78f9591e499adb2c077076a24466969ce236e041213ce4acbe7bd170cfce2a6ad3b5380283f1b7789a378c2943be81eafd2a7b9f88318a822e596dfb3687d621abe7ac40be3d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h91158f007a2e30aede2deb880e4dab460b028ded7ddb60d990d5d66f5f5de59e5efa1dfb3fa31892a6ed8ea7292793b0a6edf46693075e20820cb5ca3f9ac002461b835ee2dce0ae103d451af750;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h576f1b0be36cbdd7776cfaef84f9e887baeb88523f0ccc8a93db641166a3048233239971968d1b4c26c6baad2ae1c07f402c8c5ddb76a185ca71f8b5a4c66ac8712c77895f28129ceb687845197e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h80b178d22e12035e9818a5d6fbd9442346a64e831fdbbe0ffd4abe87da1dd4cfc086faf333160ec912a61ec7d20dd8d84572c521a139aa01b5bb6e2d8af92336ce3aeda412a0f13a07dc45728bec;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h127189d5be586fd3ad3ce44f7360a0a8cf84ef494c7204f53406c9539270ee682cb9b49f9fec994dbefbd536f642f0aaf132b73c1b0b7a90bd43739576a7046e0f926e1684c1bdfc101aa2930b36c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd5df25dcf0032c83c55ef465d43c4605f667fc20df3fa0ec280adad7bd07b0f5b16e1132826042526750821345fc63ff3abee7cce4bf423e3ada34048be38564a67d372a163673fc225b2c859534;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h101b15dc6434296db0e8f5f1388af9c9f20ce49a89efbffd7fe6550738542749870342edd931536ff6b86d57dbe8611752076f64a7505881d125ea6b1202b9cf64499b0b862aa5528efdf0abbf8ba;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1afe8e2b1aad48d7f4ff4ef3d9bb6bb506cf73058a8cbf647e7e3adabf73d2ef88d6317e8a77992a4fb1c14541b33ac7486c2f95aaaff2818e31ab4dda1ff30ead8379f33d52d9bee290c6e257f24;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h172690b4e1d6bd5a78ad3344c1f7ba39955eb323668244fb3a8eaf71ba83342a6521787265f624d44b917458703ba5b8833ef909de3d4af3d6555e641224881843ccd62422bb019678ee09775ca10;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9515aa6e06fec432bcf976dbce391cee7f242963c4ac6be076509aa83ba2ed2b6ddcea75567ee1c9af603413fabfd06b512b3f646b72d7bad5428b4026e0dfbb0c8c2c0ebdff078739c0921e4a61;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ac4a125ef8f6c036e8be4429bb474869ebdb7eadb08683b1d3fbcfc5fc471ec2b39d8fdb4b343f7460bc3b93151af78d09c25f0f38694b0e463b0386c553eebd6f5fa851595cfbca062444764feb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5fc90e4220828aa34b63dc11ee4cc1409ebbbeebaf58b9c37be416ce2872915bb8029649570b5d866926905c3145ba2b79eb5caf1a3893b8d30168bb865744b70a45c7d31784f4a12e83ecb43a8a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h76dc24bbfa874705301f27b524183db00460fba55ebac226dee32b30fb2d4ad7d2c611274f9cc47f83b2975be414eaa24e99b0022694fe13c925cb95b58a5cfb05e3014caf5fc773e1230144340f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c9f8b42c840c51733f4bce2d39f074f43e4303e4efe571cd65ede187ab5ec50797f22a150c1896b2616fda55a2168a2ed421ed01878a90a6823355725a1f09b2e4064665dc848d0bba5f32261081;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a35ea74eaa0a9a6d017a86d1ae4e5da58e44e4013323790753dcfbd954c15d39dfb1a3d62c450b10f6bf3fd77fed7c9cfe45aa1ea25a9c8fd09d62c1d96c1df5619db8423b26f1a3ff215e8cf935;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h809ed09499d2382580981502077f674a924a0ae4a5b1e8e4aaf395d2abf64a73a232d3bf27328ea45c9ad9060a014e50387182dcb03004e04e23b509808ed0f5e4e43b29702bb8b6bf1057083f27;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2483869eb21304278052e1d2800f1fcf83101d7482cb4927346de54af563b4b419f9370d40fd8cf9adcb70120200f9de8f56bcf8e21f1ee653c90ffda295cc8bb3831cf42c1b04ef08f5bd07b8ed;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2caa09d735a6405e4493ab9cb2959d1ee26e14548531e55b0cb24d67f567c3d2db707ac54cd2a3b1b77eea955d33e37b15a27270b08dc64b2c6aa77cd0a38d571dce8c9ca87b265904dadcfb7eae;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1646daf75da732792a25dcf44cf65add65a431dbc00c6f4941a23d391be950d2c6e88f96b712d178964e911f633b645fd0dd5c6becb6ed89e705a4e6d77792ee72bc25c7aa421780b6bd8eeb4a080;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10fa447d8a2e48f402270e15acb242c109d9a17ed0b03c297ebfcc9d4f2bdfcae58f3bb60566544d4710e1e10b5d6f0aa12a7036b1c38d966ec5133547829ac181a15f24f10add84732da80114e8b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15aa47c94743f9cf2a3a086c3da4b724568b777dd9152ed779a42d51be501f6b101cc421f7a8b95f37a16443bf916cfac0944fcc5f7b0bfaa19daf06066889fc62014d90ac1306126b73690480c5e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9d06abac923f114a0bb3c49c46d079a067aa67b85e4ecadd42c799f0f5c3473c25f9642a7586650daa9e30c43a459350ee98fdaaafba35da89920b0fe217a678bf1fe882ce9e0ad23405f056baac;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11c8a128e05d74cbce87148161fe88fa9a33e156166bb4c8a55decdd9ae3fc98837da3c576791e68e34d14c39a89a0754a6c93c0f5879793b40028c33887b46af76031313437aa2895e62dffe000;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he54dc2199590a8d272b6ace57855a892b32af0e3d90e3fe241773c030b9124954c7daa8eabda7dd006e32399f0142da4a10dd9c81517fadfaaacab5b04f834dda1bbded2380efaf0a16a789ab9e4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dc570f3f0625bfe53a354907f2c61f4ef825de74d01b1a4b12e52b3afe41fec25ef7360427a05defc1ab0dd61227b8e3d246d4d4bdcc3c63ab5efd972d24fcbba3b2b6cc4eec25cacfb1d82787af;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdec49224ff491a5fa5d892d5c7fd9180954686b517c49e6597527885b764c8279108b940323f10658adeb67284d45f324e0777879da4de68269f330049e2b3558ddb97ec7bb818fbfb2419b0d972;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16459513c5c912008904724429522a56704684c9d808140ba1df7ea87f81cfc55d6cbb469bbd28b818651f081154845605dc15a47e1cf18db82586f10c24e889a219a9a749ddf0394a36101a1c309;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19cee93628a121c0048daa12e832cc6babad16e9c2b0bee37325dff073f9ee59d3a383d6917df737ade729de98033f7022540f2bfd8a855118140e7d0ca6f000413404a7346f103c4f0bd844bbf3c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7cd2a02db2ce89123f66e9c4c0147740cef44f59783929eab8ee9a5119c6cfe31ed477e77acb464bb9298bf49a9e0e1b85fad917c9d9772ed4e4ddc2e27ac13130e40f55ca3a23d0bb52872ea1e1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2d5e113fdd6ccff27b651d0557168c95b9aac864eaba6f99e587ed1e37d7c36f004fd2c523ca4383d60c671b759fbc6f46c51771b3cd80a182937776c1dfcda88da713394ac7c0b290d97192733e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heedc0f8600b247b64616076edd1f168455910141eaf35a6299ef947b3117e38ce3adec46e9834eb6f58710ae32066fe64e1670b25a6a18f737885a93184c5f66d38891ad3d6b7394bbeeea22c6eb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9c35d71d7779481ae454e3087c07d000922e38104a4b6053f22ebb29ac4988734514775671df725978c2d3a5d6c48c7340a1d325c20404f0aab62de7b0dbef2fa4bc8f3fd1eaa94e8d6d0fb57ff3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf6f689a36c05cfbd59e37da220b0488b5362c180a1d9ed52549f6dd9bf3791d632b54c159b03bb76f5943bf9313a3e78196d210d9bde39c18c8fda771252ef133a8bba263c743c1b967567dfca36;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ec3752a664881b02c8529375984ba3ffe1c93fe3673974caea7f14894b75cc71ab8ba0180caec67db03834310ea6dcd8f00dd20418e34b770042b09cffebb84f0054c997fc204387e41e8b842feb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a046d0500c7cb3b83cc80c253d11053fbf170fcc14cf8c95e765b6d70e059cc49727fae5a2b10c47cf3f18ea949c33028572213ce4d910477f52a9fae3da95fdd2a241c32933f71e0a25c95e58c0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf7c6a4fb75a9acc49a0947f0dec99dbaf6e1625122473401bfd6b22bde3be8d3543082deea335cd69a07f907ba65b4f178d2b697328de13e201cb848f1612ff46bcd397ffc9a3d17ee0b81094e64;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17f54c40df5797d8b5c7278aad3009251ba93230c62575d32b2ee82669176b16cca0fe5a3fbdc78ba70e46177bdae13165b17c22a63202a5f22fc17a444be678278a7369d15a6db0caa2001422642;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcded9f64418afc396074b0b34c40fd47309c24d558ea289c056f9adbe95bbed7e5687186ce5e19157f14d755c78d754b7d1a89de4b7b3a83cf9b9305072377a31141bd697cfedeff05a1359184eb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he811a7110d4564abb11afb0647049860148c7e7ef65390d421ff2cee45b7dbc4f8579cf45849390d64ae229a84c765e71e4d131952df7897cde020a2b19432ed30ec56cfc36916d3e1a3c3886568;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1727d7e038de5cb15dfc3de91a9ff7e847a6d8274cf22f76bf5fd409dde2053021bdfe1492eb44ac797dd4b0637d6714cfd9e8dbb4f8bddf3c668f0a65d9eba8faa7a10bdcc3510afbbc0af94cd4a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ad1b48c96df3c2f1e699087e5ec4ff9643bf18651ee73c523b21cea9032226c0a9be06ab4148a47f50e41807c78d8ba465e031a7b8551b8db9ba317a85e957782ba7b0b98c0a261700eec8521751;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9ae33eca34cfcf23a08b636d0e7c1efc40f73895d6873ba172a1157c0e074fb51be97a45fcf8d7c379e4d8a7df69700eb6c51db3cbe44f9448646c69579aaffed3e5a1646f0eaab374ec7b6540ca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b7163c9419f49129563d6a2158942d3f0c10db466a569a8dbd3b0d24fd6217ade6306fc88b0d0339379c49bb701816dd8d997b6d9b133832389a271ea90ec15a5173784cd9ed9813adc8d0e58274;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he9faf8bec1cbe157124cf092d62235c3261cda90d146f2b96c994fc80a9f59efbfd67a184c7fb6c71d8e251e1217cde7c4f931ec7306dc5f5e97bf251ad3ee0c2b8a134656ad3c0964ec8224c8a2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13569691af63320584c2a05b5f6f81f3d3daa8f7b1c59fa84b1ace545a0f76d877aba77a00efdcf94396256337717ae3dd4dbc979c3d62187f8c9af5aa704ca676e2e2db6925f733895ad4b720357;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18eff3e09cded9c439002fa6d2828823fac6e87f2dc1b8c87eeac21421d6177096b3b8ff99f7eca06d95a255917770ab5c04e32ecde6d82bb34d5f5430320bc60a2ccbcbb53bd6d6d3b5ab2f36f38;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14f7e3bbcd3e0780517b787d5faebe46626c99916c05d58e6686583406ca9be9ccd2c066cc64cb75531b691658048688dc9b5ad32b24f616d5eb2f4195d1b742e715ba0bdd0fc5a815d95d0f65865;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h411518682ad039b5a683ac04c33a3cdf3cfd0770ed32a1fac286de93794e6227af0c3de0ed8685ba483794ac75876fb1995c9d5bac68a003dc4b78192a542175ca050de7c2455e134d43448774d9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h147542d635adab7b49450933c563ab852492873c04610801cc5306e5fd68f8fc7eaf89f8f2bbe8603ec70b2b5f4e340dd409502c936548973244ae5590b32c42d4c764ca97319c6f65ecbd0470b7b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7cab6083bcd1a30a8960498709762cec8fc78d25094337ef077796400ebc2605faf2cb5c59d391d5297bd42aa3b89325dd58888bc814bf348f66c5909be1dd2f74b5d0a65b4ffef54c48c669be71;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h47d7d0ea815b95164ea7f27109b85816fc758a063a40dae3a15238e374cf112e29c34041cd47246a9f09920bf715743bceb0ba592dcde65123ebfe4c5cfee2733ff8800d403e5c3906795a11045d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1396f70c7770b9d2425b2a1c93395a12dbaa0b8b5b9b1e81b7cce199556229bc4a6fc581a7671cac21bd3ab7960e9c3d5555fa5cf260081e74300fa647c8495d9d2940e55b98db198a6374cc9ec0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h197c4a0bc5637919d76759544659d1ef750aebc6170738526c2e14c63097bf9f41ecb911af9fc2a6669f6e25eae8b29fbc80ad41d5d9bfae74de6d57455b9e6cb5d2b596097330a57cb40c694b917;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd1a0a97220e4b2f87f9f7f3b84ef92e899ae2902c2168140ada0f7556c6754d02cd54b7e2da963c6e86a1cad8c0249679fde2365048a5b66187f3b05644b12431efd9d39582217aa9b58d886fbfc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6dabb04f80fe5ec5fca252a4b011deeea58c4965f6fbddd6c1819ab0bfd476bcc4545f7f3bea8900ced612e72fd0f1604e49f245708137b0b96b4372f6d3cf276d684cff0736fc428e3e698e09f5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcc278db320444702fe00e41f6c8d4c6a8f5a124f06ca9d1694e630607b2ab96b925e76ebb2172bf68ccac993e47b7338faf45570f958b902757b511c7e159f0df2d7bdee54dd0a79486032e0da40;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7cb833c2c7ce3ed2245a691433216304dc9a9c4d17c6199c4c7677e115be4d2aed892e581e28574db6bd3d5a8b487f69779b94c8168800976c56adc7bce626c15f763a78cf0b5ea9ef78e89e6dba;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e2d55a4a50f6bdd417e7b872e1302c9c80478487180161b082e2ce4ad395c1ff25af8e67ccb4fc81e987e565efce72b442ac9e2a69c63d680bcb89931609b4a931c9bb393ff7a059f7c8835c0b91;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18d4c880d97756a0d03b78a4e301879307b9dfeab82645622d4baffd318168b0fd5b204436d0ea4aad7c4bf78db6483d234b5992128037326eff6fe5f1fed4bc550795ce21df14d3636468e2742a8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h180d991d15f44f94ad9a9f3d8c15e28d3436c901130e1b0fda9bb5ddb9f4027645b7ceede27ecb04c0dd05ee5c2ff8c01a5e0aba87c547fcd82f470a0a4c5909c7809d61c60ff8608ef1a3930973c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e17a0e6e2ee2ecd19a46f4241be9fcd7a1b6d23e008a055ca85aa67be032f44b34dd74d7f42f3d89265c0b89a4655ad3f4eb0cf00fbc927c7085ea56575d54dd3cd498f2520620dfc1ebad91ce0b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ac129747f97c48e5631a72520d4405d59aec21df420f5185a69c867f781c3ad061ea4ba06525ebe9cff3b4d83c4e7f4ffdefd8a4621ec69b0f15a7b97896000ad49bebe3026c283a3c69edcd48a6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12640a48cfe6e8f13ebf7fa30a394d3c670b9d0e7d3de029d01944635fc8ed409956bb3b91bbcf5911205b2013d5ff1d6e0ec9a8aa095d71d63ead3ca00adb9f84fc2064b564e458b6b24b149e88d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18d98a24609bccaaa38b5648a9f90ea110cf587aef141c86b29b50dcaf5ade8c6bd5041f3855beae7b515b67b00608b7861cc9a3d9bc414cf7648dd11febf718799e17f4e7ad7ac57242e8d545b5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h85f5fbcda1470b609bf8af2b9c88631219a44f25514ac7d5730d364f2f4fb4db1c3bea187c0978747d583dc0c240a24e8019daca719a16d5a031bca3cb104af5b957ea7e01c87c5867d585c558;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8c7dcbf5b54448e896838cef11be666bfa5da24bdc44df7e39acfe2429fd21fb73174f2d7b29b2891a8cfb079bf50653113a551f19a310834871ef3f99073af8b95b08683068e43edc84e3d9ac1c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9eabd527bb899290bd4063ea5dfa592326d4b8d186396ea9ebf1b3cd662291b41dabb9058ca296e73b55be7ea9fa0b938afb15dce99ca3e6622062ad902d30352c9c3b95d9abab6be880b8f65c05;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19ecafbc9d98f5f593af4f6c0f3842d521934eda97f3e62a376d0a28985b9ca5bb5a5ecff3796b77e5c3785c4ff8cfe4cc8df33c4d6c9b0ae1a9e45192b29630789bf83d4f0217cd05f33389c11b2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7869225ab37546508224e2b8f87e7ac7cb37fe94a78c8bfae6f200b5ffc4b8aeb7a07d88f9ddb3381cb2d454b4c961a949709e8e0400a28b4e76b97ab6707a810bf86cef226a2accd06aee057ae0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he2e8db81d3a5cb38cb70e26dc3a2198d2c9ffd614179bc1055b455a80bf24330c62c56ef67938758b9c8ca5f827a6ea39df3e7524cded75e365f09a1dcf0eee22cc334d41f3785d61749271df87d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c6bf56523867731b86b2e4481a05bb5e2524d3b700f18b10f62b43030bfee8804e069ce0471e32fa3442f683867ee81ddb63de9874b96a23d538c86cc39c571d1da7732bdad9674866a238a48b5f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1702e4ea05c62bca1225855f508522c00843ef10f35e7a1c3b9d78eb7f78b986927b74c578d2b2ccd38885cd784730353697e58038731d7308a99066cd759140704227b225f9841cf90612da4420c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3e5f436bcfeb6768ce261656d1aad06c448403ffa1dea6df6aa3d9693c48f0e8516cd07b0e73c67fc753470db63386eb508a8ef3b019515cdd68a5353605a06f806c80549cdc3682a68f8aa0a150;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ebd1e10faa345cc2d7301d807da8a2849fdb347df32389f5c3d3d2a090b0ef2ef8a6be9cfda0b74ba33a9e6f84e904397b506871aa0265d0d3d335a7e04caa2689e3f1f7f876b3d3e72eaa2ddaf8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9cefcee3c923a2ed12bd0eb6938be167d4a33610f185dd11090e05340f076230c0a50277550638204fc366d75187ccd128a03cd984acae1449b13804abfde4aa3b322803c75e5488e33afbe5bf93;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbd1db8e97aebfdcfab68fa2058beb03b291bc8667f2430d26670174e5c4a376f929e105523dc9a40617cecd943c826086c6774b5f90a670c41cfb243b086b95870d27754d7f5e8242da44926dd3c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11a7710e0d1cef7ef6917717ffed65193893184e8ea13aebc367daaa1ce05dc5b6593d85c5ae5c5e6617c4c2925e2327df84c9d38c8b2c893a1dd8c3299fe2b4c341b5893ea65a10cb85272804a2f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h42fbd0218faf46f99f9375f8c50defaad8abb8db1a754b05e1d36037dbeb17e126fcb999e2e94efe26a596bda11b06ba1775e7ddbb31704c4e0504cbf9c444f76ea142fd3bd12a517c9dc3163c32;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c8ced08e1e1c44c0f1cc520c68b8f6057f984f51b00d513a3ae9c85c36424d5041f18d0b92d2def932d93f797cb48055452f0887ab70e05565d444fc5ce938eb89aba7597519981adc93783807f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fc7c8dae93de063de97318452abdbac3b36be5eb4dcbdbad5d6a0697fc4c2f97187fe277a917fa17d8a0fe2c717667dfec0806a106267643170bbd1833b3795c359b04381a03308cfdc0188e40d8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12b0eeb3abd6830625953ecc712a56a51566c745620be6cba6014c4be68a51306be7bb862dead51f208e195e2e925ec656e658b262ab3112b2eb681d72f2ea6bf8e509a04f06a1fd1722f9a445570;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h77e534054dd84b35e04cf4bdc35b9415a9cd44735f889a086dad4584d79c825ced5bb1fe9c5bf3a1e408ad2a590a793b5b6a5e60e641063ee95d7db271f5cd9c51bb5a93bb68208ac9f7c93e0ee9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14c490f39f2b71d9cbb699e4757f49f7220b40cd44f2531b9c705399a4870f454b51e7fc6c6beddca070fc39765f7f9ce987bf942c12761bd97f57532a1c6fbc424c125eee83fa5d4f353069633fb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc00416c3f62077af11ab61f7d8fe484fc1e992df537eacb477abc51e78e0557c995ba56e9d7855c8aa1e2410b30781402452e247a37379185a56be43eebcfe9f72825bef64baacccc6890495e86c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1517c75ef47d168d004ded2a2659e9d7be454e7fa2bd668f45fcc7b51b54b3fc00dbe1a747b5185ab15b5bbc016d395d839daa9136d46a3a7f4eaaa1c24569eba328dc5cb0ae12f95287d827541f6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19c8a76c62e11a93d5d72ec418945ec6098185ba285b984083f1753f0bb2c4661506d0883a66692b496fde6c7f081ceccc7e544f2eb5280f1d7794fcf3c6a8701bb528f0f239d102d9a342062d7a3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8d902da3338bdb25b83ce4fe0311fdf3dc5243babe829cd0636f29ded6b0b1b8dfaf2b9c55757de5b8d5396ad80d318057b6d1e8c8846b7cf923b8e703ac563d6c1eab6cb8e67ed307bb7851335d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h125bbf17af6afe2f77a874d1a52f1cf5617994c9a9bbdeed857e52b96c80abff61914e74026ea0d59a65c81398d08694eb927966623845dba4d17455dcc315710c1c3ef0f6f64dbc443c17bb8d2df;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13e214c8c6f0ea96e665082fe5dbc33eeaab8a1a00d430daf6a7db625be40b19f2a0e9c99aec2d7d0646b6734b8777d3568fa5df3957060f8174a8a70454abff5a0d0f8a6432db818fb93ca2ccda;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1816d176bbb5d9a4d0c27483289425809c48d18db699fb0daa1398b193c20e2d7ad2f4daa35fdc04b4cc970ce09c64c5331d6a00a8fe9f6a9a1c319a7f8f106736b03f461c9073b03b60dcd5db4d7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13d02871fdbd8944a59c9ff9cf7de7c8e2d050ec78aac042d24d5a183d667047c58bb37fcac8da79c23478fe82879b5ad9329657cec3a765e1db939abaca2a9d249012a372a94738785062d41bb3f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd453537496b5f08b2b25068fb48a24086c5c59395d8bc7fcf7c68cd06205e3ba8aa4ca3554a837c189e2a713f448a384159f466eb6208fac77cee43b97caa2452d022e28cbb6ccfb2d8a193aa99b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1adbd7d462fbf5a62cc549a13c6de5af80528800645f1b9fd66e8fb44412cc2f58939dbc72ac0accb7e8445daeb7cfde5a4f6c6976776267c851cef71d8feee4a186534dbc66e2f11ea01682e40f2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he1b840165b422ecd6df1895f00b7b77fad1e583312eb8650fab2964cdc030367695e835945dc8309a22c107c1c7cbaa2a1f29dcec97da26c2c148bfedc55c9241674ad82fc0b7393e4e787f044e6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfa02c4996dfa665c9917d6478265a8d02981a017ea28aedf9bbed77431605085facba8839ace6c72599d6f32bb68c480e2049d75a706f67e07f090de55b46f24577d9ff1cd55687d9f64d1a2964a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h58824311495591724d1bb908c4dde0152db96faed2d2175775ed836fbf87cde0534d6c43b74c0e5c5b67cda8af896bd621368bbb9f24018df5022da56343c2b4e36ef6ada16fbc1c6e5bb25bbb5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h126156a7ce88fedad4d63aa4d07623a3858e76bd62a39a9edd1979408a9d887083b55ece08c111ecd26cd8905e4111f0afa71251ac6e37fe96a2e6ea6ba8fd06b7d7a2914f2a0a904c1161d9fe271;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fc648c9cc963ed1f6fa4f970169a64c75b51cb6c19902e3525e274cb3c2f53320bda633df31cf9c48d0f22ce8bfea0b2f6a2a296fd46488c6ee674090c18676a310e3ca92b46004d597a1b68f2d1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h709930a248068134116b4e86dbe48dcc80c1e73ec61efba71d097f769f8862369f696a49f4930a9b3b7f8f2a7d97d7c27c60b1620a99e3da7e8174b612020e4fb55095c1ffd1746369858d3dad15;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h140315e17038a3aead2a8ae8aadec944c7d3fee55b7d94f5b5a8605ae77a4ebc149f3e18dc85b4653d02e7c8ad8db07a1bf8bda59aec600b68c96eec74ac7cbdee5ab87eebb35490fedaa2d763464;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h176602638ac2a1988216bae5439d61ab9b84ed01728098d910fb9fa7f27a46de93eeac0240100b33b8e1531296bc367acc0ff808b5a00b697e9a088f39c631d9deb92daa4de32430c0e5e880ebb33;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h23c147578b73726978291babef9a7cdd2f9c7cb609e79df33d88234ebd13aafbbaa5dd6c89f0ffa03640ab4c6169221d6cc42b7ca76dc91da00939a448ae6e2df11e4ac3d80a6bde83d8c992aa2b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15afb7155a66b77d34d7e5cd8e44705195c8c1203e1b605cf6f7e121cc1e35323dca323f7db8b2bfec32c98c6da072bc3640ae246656e6873ad64a72689f1f67192a11793275ff79daf56a85278a1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha6414154d840afbe8f7acc56649540535263a49f95bbc1610af8da47b68b4993ab2c103b915bcf343f7dd3f8a37713eb5acd97bcec8fab73a2ea107ed454d97fb7eb2430bbf373c8f78f0c07f4ef;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha5a73bda5a8de95f53bc831d0dcc516978ae53f809f543ac3e349768258743f6bb8b6b993866510022b71a943ba8d00403e7124032457875d93a01104e1e3230bf1068beb3969c9f07e17bf7df6f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h165fcfca54d61fcd44f993ce8aaa9eef2c7529c7ed031953ebbe51867c00aa651666596cd550cbe859d7b07f6546aa9bc0dee723a770b2ff79db3be8021269ce03964851d14a6205292685283d836;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1190a245d9072cfee7748f5178e81034a97f6f9e4ebcea29faaadac5cceb9be49359ef0ef2aded5f75b77d4aefcfa6ad6eea72506ee392504b12bc0c29e8996bbf8b6ac87dba6a7641612e63595b8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ec1bef8b6a6962556350c626dff0143023e6f60ea26eb08c49ffe0893919e9d66730f3d253c4c86fcef48638446fc5e808139d2ef9c4718d54f62b9e1edeb1abfbeb2fe6ba3750ca83b61b350680;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h85cd6c529fffc1ed04db30c8d7e1740f0114305134b37d3290a1afa8d86a58063f93b425cdc8a5549497dfcef4d55dca243c5417f2d147e99754f31c4839a68067de207b961d2f3827d2678ba558;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13b3b3bd16518978429805ee552e441fc78875440a298015dcbe64468245f88307bbcdd82cc96875150a3334036d9a90a4f63c056a71c516d6e30281535636beaab79123f6b2de43b346376506f29;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1115f019447bb8a9a276ba2fad726935d30e0cb273efae26f23117c7f3f4ce70c8ee5774577e15ce92c62ef60ab230e4e1728e2f4d34468ae334e83275d7aab089b438fb8a000804136cb2907fb8d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c7aab9607d06bf09474c2fcaddb9e5ee2f62826e4ba23d58aa69b0df8db0fbb300565d4a27db417502a7e6f101b7c33dbc7f462c47951dfad3ab9b4376346660f596c37ceab7d01e73e2221ebbbe;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hda9f381da7dc1e70e64e43c82e645cda5e7c1961c8f485b9317e6c8fbe45b0e0b972fd54a40931a7bd6422b13f0f79d5ddb662d2948bd045ef2a084c12e3df012546930935168279ccf7d172e0d9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19b6bc1b6866cf729a1a82df02c8afd92bdbc7279dd4cd49283080406b1422be20ad4c61d93f16d83481798808a88c0b1f75291a602a3bc843077e5813edf3b657ca9e123139c6b62d97ef9a6bcc1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1477488cc18a6a8c8fbe6b52a967d63a3c63a523d4c0a02c0bcff631b5a4888b0c2e086ca15bad9bde918b6da1550b6580c57a58676ac200b269a452453d1e9ffdb5a1f2b61f383bed4afabba21cb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bf6df384c5d2d52f1e3ba1e637836541db3dcb146e44498dea3ce0553258a79209f24d9b4f276b9a390318931026c8322a84397f48a0a635f1e56eba729d2f1e8749dc359336c6f3f2c4d3962ade;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6bd48ba33d43ffad6fc57f8f546671c863853a0f5a9836daf5205c0e92b4040f84b16d1fcde542c74339ad222ce8fe0f04bce491733667a86e9fa53d685e23369bcf753bd88f778b6225b8ce8c92;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h150c4a7bbd15354aa80341c60cf9d1e35dde5c177c30caf2efc17c104e8894af72a2d614bf9801141cf70cf07c4ba9ec46b4c69b84bb7beee221f5dc94f0dfd32423b2e5d2561ac8d471293aa66bb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h49d9db906d0ef4b4515c89b8889183ec58b47368c813d1de9ad124695d6d9769010308c0cfab7909521e88b743fb0a23f8df8d82e2ebebb634c666755f55df6b1b9be99d9fbf1ee54a8f0b1e0b29;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1da06c76cde909073379c42ee1a1ee560d57495ebe58120f91e9cd9c78c506597a4fbff32e97b4862135205f2fcb1ff45269c19816aff9231c2a48f753cd684a291f753bfd24c74eaacd0a8f6ee82;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h670336ce5c6723e010b73e9bc9ce7d58bb9c789167eeb3feb2af1b11b1aab49174643d245fb5a6ca13e1ae2393c06d26f901d5056fd226d82d15138983414f3c49d28a6909362699c966122eccea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12da34e580941c3cab88704a6cc3772803262535e501d5bedc9aba3b400461360ab91a6f3ae8203ba75bdaac82272b91b0610aea8e9ca58b8da8cc407717fa310659f5c5f9a6d2ee2da3e9dc2c143;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6d0ba94a4e2628c1947c13f3984a6809af74751c1d2b8714d6656a3f82aef16f6d11610046cd85944fc8c1d25736a3c7013964486183c496d9282f73f12e4848fd5a1889504dba3a5097a44febc6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc19617de550be8ececbf79d1de201b19ec2353ac21d00a0fdba6674b7b764f4d860a604e503a769c06e9ab3e33ed46042c1778ff72689c69d5ddf67b33ac9a2cc5cacc808ef33041d1b6598d44d2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16d53550a77f3d890db40e93a4de55b7e3dcddb1acfd574e64c36b9276dc330f7cd2b389bd8d0e07d5c1ca624d1ef4c80eabb1c0ccaabb660ccf0b9b7b0a3b306677ef8b7def584a28171de24755;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1274ce2f9893e88723f60edf2936b04e394d4c4243ad34c0659bc4228532bbe5f60f1a4e7107a5285f9fcdb4616777f9be3ef2bdf3646adea8e24401469a5f6a85bddc0f7e9198f02e9d80bbd87e7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7bd2317d91090e8a988085769fcb3abc4afcd6bc4e4ce147a74249ab159c802226782628d7430ee98ab3aec66d6a51271be3da4cb482cdedb1f4cf9d90b46e0e7442c9dcc052ce904dfae0b8022f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha20cd4063ff96544ecf2c9467637aa5157ae7e5217b97e6c86c4e58d793677ff0e99f13e5024383d5986fb881c4473d487963c1bd646ef6f4aca3548107b01e6fbc78fa0cbaf145c6fc16b2d113f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h113e9943491576cbecf6316fe2abffc397afe3206723084f012588c3300ea3bcc9eccacc7ef651a27183429687169fdfa3eb6fdcfa75069e65d455c5b9ec795a003a9d9d76e8aad0007ea5ba6c2d6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h177981a9dcb2b6f11162d1888472cd9b12820d69cbb17faf423f04c06695a11b9506f8cb3858321522431ddf92560f5af8625421ea27307d3e3a80c45eeff12a148a555552456900801603c89caf6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10dfec1eedd63250a0ab10ec68df783c89c210b2e7041db2be4debd293d25967d997baa138508987cf79d39cc6d1587433fcfe07022baf33d04d40ccaac191fe3cac1e764e235530373d8a9e5f12;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb44028a6e7279cd85802810716f823270f6c034e2dea92883c8a5ac3f4ec6344e50d8caa74d3c0d823d48e3e710fd24a574dd560304cd3f888e1635d7415c2e9939d2d015163cb9e742c6c16ff2d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18cbf1f0e79321ab5d5ebe4e6bcf1d88fce6df0cb8ace6fe56ec9c4752c550e8488f7bf63d3b89ffd6d2d9e010f911ed75e9c024a34c2aa79ed61c3930fb3aa8a78d5fedca7e93412878753dc4cd4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5b7cc36e091e2398cf737db8db453dbf2ba2de93ee5b373aab8b0e8787bf73191b7c95fa381b77ac8a30634fc1f75f615c05ec0394bf4917af79b3216af1d6b829ccf5348a1e3c971338db8e2db7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf587f797553ae4a5cbb4c7bc5c9e97be4d1be43473545b11b1c58e1ac7d7e87c5a24e402261796f1145d14dc9d4a3486df1e77a8b4ee8b4280133431c5bf37826d5e139929c657073fd0a1681904;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h57024873db011abcfff04dbb6a243a6b141d4e859fa7c6c725d4a4fc05ae1f33f988d0a9d9294767e3757cb3569bb2aca902a710956ef152b0a66bc44f4a25e71a5514ddadb500500c144e350cbc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c48218e852f4c6db4bc7226791e9d7df91708ac29d6445c0b7eb0920baa80a632984f3ab925636ac1971109261dfc485bea64a7257cab29a0abbb2bc013362b9e3762d950f6cdba25deca3e2536e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a4bda493840fe08be2bf0adeb4873b7d7edec7b93de6d42fc896111f0366abe0896733dd75008a1517fbf0abd183b71adb62d75ba7afc27661de91e485708d703309d51262743c8c2f225c1f1244;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18da3162b9a2e3ddae165b5c28c44a58f56ef7f10e5a8834bff0d7781ed18d5a1497856d7205005b5a5031b888675862252bb2ff9baa6bdd7639997e0808456e9268730445e6bb07092deac8e7aac;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1babe02e16e9aa9a2848cbd1c34d6540ef5206501f6070887d4d77c074a63b562b57a6ace32d0551f6346e06b7d610386482763138b473ea99e877250ca60a8595f2ac64565e363bde1c3db255138;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19b153ba60cbdfc416967e1c31df2b47d9f56c48d872d9d5792d960e729f80a1d069547983d9178407603d4dda0829b9ef0cf940550298f5d8fb68fedbc2d9b0facf214b0d18049bc4b564bebfc09;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1797da02454f1f28857f0880cfbc689cc653d2b6b0220b283f03dd420daaabcd91a1065c0f25ad1e19f7e1a36d33d583ff78b4b644bff7d0e6171a675c495eeb039c66b261582781aa620a923dd6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a2dd8d3bb46d454b5284685d8237071476ed8c12b83abb82e3da53f94d1dd47c76a6d85dde6c5c3d7ec22be6e12a0606f5297da6dd8a1db569a728b126b270c0d14dfcaa269a4d0ae622bfdfab0a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h199b1169ebe666b38d013423b7be107db9e84fa2d41004ef08832bb88f2b9336698f86e201a64df04f903805e7ec5d700ec6326a6518f5c20e6542d7bc56a01911b9047a4b3fe1f4dbdfa7235626f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18792516d74640466c89674d7564b941ce39cfb8fd77f72ca24a689a702a7e6ec7a56d211cb842d08393a22a43d66643a6c6dcc134675bdaec0b69e3eedd1da00264af19f107ba6b7eb9a7da14933;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8990aed7a5b845f2dc86fb6b76924ad4d201fc8b496b06a4be0441f9b71648ca5ad42de6d87c296c31c8a843481afaa7dcbbec8cac27b620c540845d2e2805774f97426c6da9a168bf794e173e40;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5329563addf5c288b9a3362a7cc1a436061dbb12de7c77defe627dee63c639084cbfc69bd33f72480b3344fff2b7f17619babd945c2346f34c701f867eb5069e24d9596d36b0974e6aa2038815fc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11d968e1290cd346c15691fdd4899fe556886790916a82d7a419fdd284a904938b184d2bf590ca735a34f0a3b1a10fe15c6f9205c823122fda2b276d01f41b4a62c5f0338d0d6e921912db8e64643;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h895d3789fddf3b046b2bd5e0ad67566e492db7c0b8e12d26b84cce7512451d410446bf48629a6cb7d2ea1d4a95b7856c44171164be34e9767031ac3a3e4ba48fa480366d7b9045ff6ca4fb7b876a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd923067d2b574d3af079ce9de4f3bf58370f481ad20b40beef07c82ec9d1a9ff34678c5c3daef1dc45c78d057cae4d30ec257ec4d3ffa55d66969e2126c35cae15fbcbc9f6ba3cfb0c77f81d0833;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h87cae141b58301754cc1073947d93613f26619fb2295b68edb35c575ccbe11ce9addbdf05bffe186be530d1ae16286ca2b9bfddf95575fbee4aca3b99012927e7339a799439abedf85bf4cb904de;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17f582af088c8294076c05cb5fde3b8087d6fc0950c90c365d061fc34a6b4787dcd292730f660e44ed6e2e87403b8d3444abc78e10ec816a7e047ef51c1fe586c2771f3e963494df1b7308e26e471;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb337f57efc84f992b88bd1f394f64159345145110eb7f66dec6647615339c892eee21711d014693c75f2a2fd2119f583726b031195dff876a54d255fa793b6605cb7bc8c89ed4248836dbda7f4b7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a5043eef50610c02e8e28ee5accc03bf6a1f4d7df569bcef7035546d3cd5c525e959f9ae92eb3f5b8960d27131b6d428ede0aa34a4123531ac6df31cef6417aab2f62dc4e911f75cd8d40b12036f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14bf67c7b9bb15b742598c8c584206f427244e1b75c58bb993428e1adfd608bf45ff3cf0a51b4ed54a1007f78503e13674dfd4b48176dc7bc989bffa9fbcbf619beff35f3250787c679f5dc8be878;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h84995e7c6d2a6e8b8df5a61dddd7f435c01f5603d3a2fcd654be8dd25835d6d59055b48868484831e48b84f287f256a582565ff55c0ba5f4f5a51515eec705b1a6bf64a569ff09dbc90b53a6a8a5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h44d9608ccd75d8ee738dbef8c0398059ebaabba2c397edae811bbbd1ddb980b0394c5e5079a4de124e37b5be17908c2855dac2151d137e9dbea4ada78f367a06b47cee7704348fe1542caffcb618;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb8f5c20571dea8a81ba76f36fe2bfd1713b662c6597b42f0ef22092d60dec560b5cd61fcc817c781ae6e8b321149819fb0dcd841d76180213bac6cab75ef1399eb5a1984bb8a02afb03c897d27e6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcb3aafbf9d25bb0a455a47fba16171b2037af29d4dc313fac3f6aadcc5c00987e0d30633f78b1006bad7df577adeb309dc27cb588195064d88584dcbded8e2a72f8da611ec2897630b8a3168e78c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19d0af142a91a68f4e8903b9d4b8efd3a64991339149e9f66a1840be9fad2d0728373350d4fd67aa3f64a684ebb7480fc1e821175d4c24c8d8943a1561629812833d04f5bdb0b01e828d3168dc2a8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc4f9c73e8fc4b9c4cb7a71f5232af180b78604ad5eca30ddbb2963196bf11caa6aa73bff350807574569caf81360207199ebdd88d7f2363999fe3b6440b3938e635c40cf7542f13ae9775c47872b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e027cecad6e32eb9e4abd610bb687670c3dde2c8b2ce8c7d4c43544f5fa58fba1eb009bb36a556296846b18e0e53f6c3f710c5a715aea03a4fa052a1bf32e2fd23870784161c0c1117588e542f92;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11c60d1928623ebf4e47e6453b661f382396dbe3c9287747233fb407c5caa684377fe44b3e6a2f5b65985371c74cc5159027ff8bbaa020f62593a26b7d94b1e231e87c3dd45e8782e3d45b34392cd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19ea9153a0402976bdfe57b6885b472672f0bcf59ce0a411d3ecdc0c214a23cc98813acbc86265c6e5f15677d99abb72b95012c5aaa188e3f7e578f6e4468d71e578d5ea11a04ae7dedaa79abeadd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14632907162ea2c059d54d69a61c193862fe52ca8cfa78ffb4521bb7159a1aefb861b73fa59002f9127b72ef6900dcc527938c7e2bdda0ee1598e0af071fb129ac50e1da473b30c80e2097d5de1c5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16058acbd2849c50c5f5163d298935751fc452527af20398d3f11c8173923117aeb8b7689ff8f79b347859873ecf8ac672a395d0498accf9693ed1091c574623178306bb1880099573d5852e99682;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14a4cb4191dbee383a0b7874dd9047f1244351791a56578f3af29cf39a0cc227f06ffeacb34a199f0f181eed391ab459f031e9c1335f75d0a729242cb30f35961cab2493655dcde345c952b7d3f34;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cbc811a233a7f5bd7fc91a19d879c8bb84f858ebf596b87276b6f1b443a1cf09ee167668272195c246827dc55ec9b18c35ad7bbc0b419796a70f72292846998843b09721a61d29991b7f95cb717b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1542ab3faa6993b8f38901b2551cffa3cd589a0252fb0cdbd0b650cbe6562b4492b0645442d66c99027c94a280e6eb56713be3f6f27d20e0cc58dccf5ddd45d721cacce2a05bb3c04de7f3341ab8a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18f09c1d690f52d71d5c38cb7d7d233e13230cc6e560c96fec5ce519612b145695d2bfe35e99f171a8d8963ffe81640c5291c3e9f1f6cb4035ca9b916a23b6213b17f8924260fe72b44722983e808;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h250e3cde67ff5e1e92501363d071b71087adef9c140c287b86b884a41ee0231592812a25104e3c8b65d17c87008a8237f2eb67cc9a5197adf10d443b29c8f275a9f2b05d6a75cd38342e72555427;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d52723e363ae2548a16c7c0cfa0de452a4fc42c66e96e85499439f9c2accec9870cf8d11ae6a53ef1c412231cf72878abcc3f4ef0d94f70618038a6b1a1ddb6e8c95b79f1cdf7b62e97cd27358ff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h114f8e1c0c4b0110733ad5e7e0e639378b183ac85befd2a67cef36e4c221af15f9effe40ff6ca8038123b1f1185cc74f7d896ac8aa6cbe51d628311d127d1f73d27c7532563cc604ca0a4672e405b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bc5a2ac35947c3f53591911667c9d01216fdd652a614ba2d0760e762f958b764d86e67c61f3ad243804ab495233541c4173ca3750fd92bd653fcdd1fcb1656201f802e54d9c26e40bec99f936320;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h87e9edde4aba6e9e73b9d16858bc307e37b49377cda68123144a33e6141145861409358032ca7d58e839c08a28f6651e57ca8cedcd589e94c592fa0d07df9a7436665560230f01fd07e024c868be;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11cc466e8ca89f0620bb803c07e722a612543775d2c6addf0283d28d7117789e8bd08798656a85cf03a1b4f4ffa4ec53388389158171b8c2f1598b90aa5f1027391f6a2a6e98a2c23aee5ec128695;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d4fa5af9113d00a27ecdb71e705570708f2f8066578b17a7ec8313c57e686937d1f7adf6c486ebcebd1f619604f478d84a2d959953b7ea69d0bf5700a879d26de71b78c85690f9bf866ef75b62eb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9ed8a3c08abca82f3d3bce13fe2959dba5bc9382d5d13b5cbf805fe18b507ae35af1afba3b9459e50383e33f699343f65e0b2571bdb2c4bd75592639d55f581e8a100fbd6233a445ba35a8b61271;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1db1801694bce661315504fa817dbae2b0c569a149f4c34939b538105ba71bd7a04543ec68f100db54d7556e7230a833fef11c871e94f4a516932969c6fabcc7d44eb70a394abf346fef7c7e81d87;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18c87fd72bc7f3a04184d33ec5cb7919d33c5eac6eac6900cf4db6c7f502cfa7390bec2c16dfd9d541d46db11c037b99716def80a059cfe6aecd7f35b012c85b4301b4d01e71e8322574860830701;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6e2cb42b77867460515be8f02ecc79bd1e8a813089324a3b07074472ee40b3bab87335c12eb862f5db4cb1897546e8cc925249eb2a090aae8ca7d84e97c9ec0faccac93e2623ebb2bfbf59fa367;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h149dda47c362a70ee5455bf55aa42f3142de1efbe1f7eee78ca36fe7cabd54f6a72d99371d469a2655f9bd712fd31466a754e92596ea81e82dbaf7712b06b577f9dceed62bdf22c9522273f135853;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1804c820fe0b0b712e4de48a75dcd5c52a9097bcbe91b7f53a83659841a68b958f383e00cdf9374c47f1bdc10a01762438b1d80b51c3ed19d968e0499f84e7648ef85bd64dde674b92f9ecf661c7f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h61fd4c7d8080862950d19f77d9e4522c4db38d70e1f593978c97dbae747fb6db43248efbbf59fd29af16e5e06fda6125d1ef899e58b808b25a1bb928f0428cd1ce31cb3b383d1bc8df7433671a23;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f486e0bac5acdbffc8e4d9c97e4cf9135a76eb3481eff1726658b0034f877cf154ab98c78852695b4936b342b7412cc5bf257d33230642f94fd43ad2f74af16ac0f85b18aebb2393b76b0af1bb97;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8d31f871947c7854f821da543dca350f2f67cc0bbf08113194dc0f893b8c29ef8398488549f058c00286ab01232a7e0897c0efe62766b4bc23bac49bd5d7a8b4f2f3fb955d28fe88e993ffa265ab;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5bc4d689f19f8f6fa79bad5e6df284f71e428fbaf803d578c733f7868df188b2c66d46223c473a25ee9e40b332c3c679027de66a4d22969bc87df098715a243f04d3ee4e201cf27ddc116b089421;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1027fca2d11b85108568dc2c2ed7918a2102effc27f435f8e50ab937200d036b4ca93c62708e0cb0cbafde13bb72e974396ebc5eedfe8929d2ada16a56648547688df08a3853f82d33c35d814f99c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfece858d8cdc67ef85cbd6540f604b499951dcbfedb08670ba2ee30ecaee231867403378b528728e7eb64633578366b3d306575c78bf9253c5ddc489936ab2d79b4d123a121170621bd448121d81;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1222f018f4d478bd0ceaa14f6c841d5c624837680bc27f87b5e1b10151fa33f9abf34a3bcea81f9afc613cf766ce8c99d93e5c9bc242f651da38025c8ba9d351fda7f975d517c398894202a4c6978;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cb3b696115769e3038ae8a432375993b2b5f7d6cf43ede62165a5971c7e59035433da2ed5b6b40e22c9e28e35be1bdd1f3a3f9b501bfa8dbe8f774bb2ab522de005dc247d5e10e9fcf1061c19717;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h516ddf7bca8d3b00018e303d11aaedbcf357ae9d80c52110a496a6e09bec3aa641cce6d9d3f153b4b98ef9e745819fe1c91ff57a5f00da6784ff607b76de84c9f41130dacda0551ba7b4f535012a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h31f866394010c9fede72ce1bd8b66c55410ac068252122a86f6d7e381247af5d6e268f65d1f514c06be0e6f626972fde33460c46bd2674492fd69458172714f72f53e5bc092d1b00d5bd8eaa602b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2c69fd10a6618a4e1f2ede562aa8c999dd4dbbddd2bd84993c1ce287b351ea63c9ded69716c15c7ed1ad1bbf9f6f5f66477c9ee49c1b50a8d9ff86b8cfbd56a6351593881d4654f6e6f3ffd44b68;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f196f1d479e956fd2f7d1f1977705a65731d36d3247b9c519ee0abf9690a36cff470c9dc3384d93a9782713c5f60c2ee16335e09b01bdd8a67af9eabc77da2187ad70c918c7e4a0af9ba5dea230f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9d85117d910e3dcdee33cc739e955db96f177ac8780c8b6fd0b5b8b2693a73e38687a97e5354e7991a09b9f9dd2bd69aad788de67734e3f3a41954195567041c10f02e752c99dcc4c4069a865803;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h25a1ac598113856598a736f7da8a380dba629edec42e953c2151249dbe6d90059644f4bcd676cbdef4b004f6fac9044c473e6b60967ff1efac558a6bec90a87212cc5d1740bbd23c915e21122d7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h23e9d94320e3e9e13667c98359cba9dca5f5f58229175c1d622fb3bc5975acc8119d733b839fcf40bf44097f31946ba843ab34a382ea1fca91df78d051c6ad393a39f09c9b51379290f81e7041d8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h780777d9df229ef249616ae9eed51ffc813aa40ed9d1b9d11bfbd0600050350e67e3a7dd6fd25fa35528e9f2667acfa38da4ba2c29e7bd6935882e3daaf2c99d01b8a5cf52a0d5ee390a4f67457a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a5b1544aae3498cd3114477f9bfc102779e5aa2f0e3e4cee9f48fb958e0906ff625e09ecccd9bdcb65222c47f17b7dbfe5234adab2249101aa0ad7e119e070e963e48716bc86e2ff849c1b23a8a5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf95f44f8e46563348379a31c4043314ed79d109af5b5f0b680be50de29cd6a38abe9cf9d81a01082ec321de1121b40aee82f350c10efcd5074300d0aa13caf323b366a929e7a0e7dbe9f122f637d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b6d000de813850f44f5d384fc81133432fb79ebce13f10d5419da9c72319c03e50978c1a9a8befe6072f81acca9e796a1fd0c1a38d8fffb17138b1fd65cb8662d07c76572cc4612961cb6d41153;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16a1b6780ec16927a34c53da3caa84153264ea1e8783a3e9a2bbd29e45771bbdf219bd1a1984fd621172c27128b7ee4049554a2be7a1949aac66f18d24fd6814795938ce39d8464e3ff091a957150;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h685a05192ef13bf94037b935e6d1abdf0c38f2eab592c2aac63de4e0e048c06161c9b3fbbae6b94756a2b4ed6dc603f0be931272a9befc878e4903dca5e40f480f163cae5edfd736a6a14036951d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2e1370170ed86e6c3e5c4ba5ac53bd8b4f9bb0964fefee71ae87e703192c112aae13bd432b90ad5f146df728fc2be612206efce1304b171abff9be244681e91ad1eb6ed744b238e45064e3b48c77;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h118fb08fb7fc07d339826a9af8829039814be7659b8bad320192787200ee8ae0c661370d05f1b77c043592852c9560fc9a3ce01234e67d81294450aff28d0dfe35a9b6e96ba14b0785598a5687e41;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he2c0d5f9aaf1e9a9ebaf0dd32e9a47bb60ac319bbf8ff90620c0d822c8c409aeb1e5e72f2acde12edcccb80701fba0e42187ea67ba0f0728673f0e78125b3088c6c9f74cfabd4dbb17a9545cc8f5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1767a5072960f08795121eee737f9db3caac8684d085de76f1d89591c538031943468a08f17a36aa6dcd1f042965a8fbe43542f192c2f7539aedc335ef059c7cbd348f1f7e6267a536b0656126201;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h109c5d490adff680ea6f280a0f9086421f558ddedf237a9969a64f4b9ad213adb62e884d567a1348861342bb7e918e8990d0ffe177ea68097a4b5164cdbd904da60a865d4519405c76830391e5dc6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h165fbaaaecabf6c645b77f0df1fd114cf41215c44aa8729719bf847d8dcbc67cb7578a49d3ac40e0caa323c0cccf5605fe728369ce68218c7821296da519215d28c5b97783d82fa4dceb0215ac1c3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1102e70f224ade11be6872dcff5b76feb7136d98b0a5e7925a3d7ed826e8b9f56ce957fbf15798fdfcf316f2be3c22c36250fe2dac36b32bdcd21ac9666f7bf0d0c5435f08b02fa1ba9ec7603b7b9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2cec871c0bf8ca87f4526b19b9019e45e8cf9b43148ea3ed392b885e1e42cdea70705c5c7152962aacaa88ecc9bf051b34f90c24e012cfc057b984f1b84ef0c22a56f5bd80cf30ea7b01e224e3ba;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdbe562505a77e5dff4b273ad69f10591ce626bac2ce5923d3bb145e55b7888e24b2320e53c16acb3d45b62c7a18e8d321c1362d369268dc5571fe9e6e0276e291a18bb82b39ef50419a04942be5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10eae4a4bf7b45ad22847faf1e1ba10017f612ddef7ffb171cb3847440b57a9f776ce372d28ce0d0fdb0264b90bc4e4e0e517a3585c739ffd8432a021d293d959ecfcd3c9d28d9ba206bff526a25d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hea38f4dcaeceadf5bfa4280a9297b3ae80c9234de52cb424d93a730c635bcae5fde50a14af651ad95bc91f40b8a452a17a6aedeead2134db2928debbf376ad30c6e3814330ec73c2b92ea9faa282;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1953f38eef75594e5ed1dea40793d732300f7988d577aa6a7ed823bd135eeebfed4c02d7a6207e6a7e0480b279f0b37241bf96e0dfa8d42d33ac2cfcf672fc1d3f2737f8a71f79df9850437ba54f6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he5aed36b9f728a67fb17f696fe03f8fbe9f464c112e0d43ceeb417e4304185951a9ad5296dbb4c6d2f337fba744308e0c3b5062d03cced0a05fac6b59d7c6a67ef401135013ee0e635151a2782b8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h161d7fc309aa802042f6b940603708f0a5700cdad386eeebced2071e73d9a647a9f4bd3a9158ebacd51390c635cc0643a9c24b083b2b540932a59131226b510cdc62181b3cb44cc2be255d2a166fa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3364eefbfc53b84bc93316602501a999ffe67abc6b5bd1763e1a511f81493e5d36b0932b6d3db246f6b32fc319ba8f4504425157cc6b85624e2be1c6a100a42832605e259078995c95ac6efcaac1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3bb0446303fb1d8e651510a419afa67a5bb6fdd47c3e0ea6340e25cf186c467e666fb15f62bd908313d26a8ff306483c6df52c4894eff1653171f45a24bdc16e75263af62ada7dec0864b41836c4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7f641c449beca6e87559304c263d8b8a4075e48edda62efac11229fe6ca9e851f72486b89d52d3f0f6415dbff8172876fd89912d2f6902590a22d413e4d5d6a69ca0ebe31a1e10d6a849f59b05e5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc557edc5bd152a23c10d0620f54fa47baa51dab7293ab2103d9a94f538c17dd3e120dcc453d441bca15bedabb992bd60a951430dcbef6471c000a059e0227862b8ab7f35ba098a37558414edbf56;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h645787fea08efcd2065ade071bd2656679bf87795f62110bb77340d1f60f9b0d0ae45c98690e70938dbfa4c7d8ee6b21ef1de944cbf68f1102d3f9e94a09ab544e1aefbde5b4a3cca96f344c8343;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h85a3d5f0bbb9b46669af1f433ea3035dccd4c5ba59ea25cd6d205897763b861032926b711d259f0da12baa23d378ed73e42d5ebc371d000beaa290b5a63df9abfe9b1b9750031a4b87de8f832d13;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19acfca7e0037a90a4b3b4a8ad1d9b157f992ac3c94f7d47aedc74271dcc097d937d1017d82583b578d75016482146fc704043182644a17bfde5826f6ec12533dc03aa7021428dfa7bbae96c502f4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8f890ef7d9943cecb5acd91ea82051174754e4d1c1dcd2a1baa5b3bf5e68e3af6514ad98ad3e26203561b9381a7efd36e25b95c76ae016f362fa247d37e2c988256fb4b6d0b242371b75fc1c7fe6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f5fe8cd94edf5989e73ed421438417bbf4155ec4dca0a020360195e175f134aba5f111962117b0145805cf473445f52c619f284db3e6d5b212d843892aff6f541bfceae4e5860fa3234c81346108;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haf1e2d077006cceee668920d4e133b8db246bf71458f1e5313406b4d293c5fa57d1e0744181e18f8d8d5ab89337698a7a62a97de3a7a32d1c405eb81f04879fdd67b2e98ef1e4bc1d81c04b87422;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haf3242506fb2e42d6984c6706ef95be0311c5ba266eeff56b9743225875627935ac12718abfebb9bdcce1feb39642bb66f460297db7241b1ee40af98362e8190138c1c3cf6d36954394c53f2bab4;
        #1
        $finish();
    end
endmodule
