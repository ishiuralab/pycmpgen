module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [27:0] src27;
    reg [28:0] src28;
    reg [29:0] src29;
    reg [30:0] src30;
    reg [31:0] src31;
    reg [30:0] src32;
    reg [29:0] src33;
    reg [28:0] src34;
    reg [27:0] src35;
    reg [26:0] src36;
    reg [25:0] src37;
    reg [24:0] src38;
    reg [23:0] src39;
    reg [22:0] src40;
    reg [21:0] src41;
    reg [20:0] src42;
    reg [19:0] src43;
    reg [18:0] src44;
    reg [17:0] src45;
    reg [16:0] src46;
    reg [15:0] src47;
    reg [14:0] src48;
    reg [13:0] src49;
    reg [12:0] src50;
    reg [11:0] src51;
    reg [10:0] src52;
    reg [9:0] src53;
    reg [8:0] src54;
    reg [7:0] src55;
    reg [6:0] src56;
    reg [5:0] src57;
    reg [4:0] src58;
    reg [3:0] src59;
    reg [2:0] src60;
    reg [1:0] src61;
    reg [0:0] src62;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [0:0] dst63;
    wire [63:0] srcsum;
    wire [63:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62),
        .dst63(dst63));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28] + src32[29] + src32[30])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27] + src33[28] + src33[29])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26] + src34[27] + src34[28])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25] + src35[26] + src35[27])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24] + src36[25] + src36[26])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23] + src37[24] + src37[25])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22] + src38[23] + src38[24])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21] + src39[22] + src39[23])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20] + src40[21] + src40[22])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19] + src41[20] + src41[21])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18] + src42[19] + src42[20])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17] + src43[18] + src43[19])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16] + src44[17] + src44[18])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15] + src45[16] + src45[17])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14] + src46[15] + src46[16])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13] + src47[14] + src47[15])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12] + src48[13] + src48[14])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11] + src49[12] + src49[13])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10] + src50[11] + src50[12])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9] + src51[10] + src51[11])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8] + src52[9] + src52[10])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7] + src53[8] + src53[9])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6] + src54[7] + src54[8])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5] + src55[6] + src55[7])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4] + src56[5] + src56[6])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3] + src57[4] + src57[5])<<57) + ((src58[0] + src58[1] + src58[2] + src58[3] + src58[4])<<58) + ((src59[0] + src59[1] + src59[2] + src59[3])<<59) + ((src60[0] + src60[1] + src60[2])<<60) + ((src61[0] + src61[1])<<61) + ((src62[0])<<62);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62) + ((dst63[0])<<63);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61dd41f50ffdace5112ce0e18b0c966ef311ea3f32472d043933cb4a583d8e337ba18dee1d76ff636ae76ab0aed057b189dc791a836306c84762ec1a34d4772d334d4ad0553c5b0ffab30b45ee7febde591fac015d600f19acb3de6ba3b98cc810e28cdf74c77093f8db0aa07f36a1f7e6e0487cbc2a2a745f391362893003ee;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he1ffdcc08ca59b487014a52d487306daed31d8c5a96dca3c332f26e584d3198b8304ddd5102bf15a0f8f64c70629e8b9ad6735bdf3fe7e002d5d1115e8303c972a6a7306a6e61b0c270f42d299ff7a534af8a76b9c9d1d75811a12c64cfc79fda46bfcc7301063b3c3957816db4148d79bea632021819ae6099f21366cc52a3c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8fa3dfb593cd736cc7a7a7376af7704e749e150082353bc52cb75d0b21d4d18b2ea16148b8cf4a2d6e65a8fef4a3a1afee628a7ba936daf67a65c33e31980c5c312a436f34af26eacb5c11ea15a3c08c7b692e2de248120c63f26ea6ff9726d022c53ae7119a60ed168d7c1164539b083018530bb7619d67ded169c1b1696aba;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce8cc84c2a0efdf29a2495a15440fb27c4a45e928adcd555ea2742835f2eb46bc30d6c450108ca982d29e1f165d81592b5461a6291613cb6d776ab7d0295008dd000e8c8520bdd580bd439d2d458a612377de1f1d294b557604a7cc4a1756778b953dea06064a3e2779b8c171fa65485dbb6cd3a16bb97e1b7555cb3d12e14be;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h823b1dd5f9f391437f3476f8247358cf2a306709be0b4b0f2b04fce3c597ba20d92b7ee7fe0adff9145cc703a7af9b8b590b089cb05edae2a68b2755b737575d9f6e37bd668843e8a03c2c33dd357bd26a9bfcbd3fe01db204a757a4525f152bada78f313c9d2977aec739173e467e5f58edac2e89e9b7b6890a16225626d35f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce09bee533d2ef2056e53bbe6102e6a2ce4505b0a8ef969796d75bc8b6c84b526804dfbef6549dcbda9d89e4683c5e9e52025f14b11958dee38e72a44bdfa5f20a2ecbc524e716b181790e2c7ab803fb542c62049eaad4f14d97e7ed814cadd50a4ca0487cb8dd9e462254eb7dc38ecc53e62b4e00326eee7088658123529555;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he15549c2534a220a85ad6bcd25d49ba4327bf207e4aa96d2f0227b69354bdad89a858c90cb2018d1117427796bf08cc9e6b528c9416d3c0b0b71585aaeac22fdf1246d3c70eb7ae7e5beabdbeae20a8032d67e40c9f6cb2b54012e0b494644f693c6a57bb0ec4b204ce0e3277763562af9bad72043fcef35508b8109430b8e5c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb3ea7f21da75505fad7408994764c3e2c7826a056c421c3c02764b344b05e3b108f80f827f8f3936b0353dd9d41cd312a87ceec14916f2d179d73c88b5327917cb3c44aa2540f9f441b273bf472c2e60a4682abcd44ac1a5e67291ea471f0a0032a2aed225b6905309532b64d27a20f3ea7ec31d70435fae7e5a3fe0cf1103aa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h964cb5ff8a15531d7c45129c28565923ddf3adc4e568241d66707fae0592ea3e6855f1cc54e4a0096d8c02141d1b80a8cc512479fd51c977ee14f8b80b8f53a695d2f21e0a9cdcbbc83fcb47475bee91f7541b024daddb8aa6dff6fe4fc1c7ebdf263301224014bfa0abfd1b1f1c49481d71ef9c4ef8aa9621fc73e0fafa6fd2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d0e79dbbc3500fe4ad7348ce3f7a257d9b0123952db05c3849c6fbfa329f6a679cad1a7635758355e03a670b11d367b920795393599b5890da1524e4f1e5851c4115097147a35189b1f5d34bc0bcee129b50e7b5bc784bdf2ec9d90babbfd5deb9eae04a5363bb25b7c0fd76a6b6bcdfef096fd99178b75eb804a7502ee04e1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3dea11f63be1481f0da7ddb683c6462e55c0bfdb1e0d86796c77cf80ffac6bc35f87f9d000c063505fb32f98b2125f95cede77825f5ff3c111a49a7dbc22922d9ae53c2e5f32cf63edb54b06957d1ad219dbfe4962191adb0ebcb81cb9fd95ddf9dafe1bb69d26cd75dd7ecc3b0f62016339b91484cc118ebd9f95f77ea71f62;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha05b992951718502f5f5ae3d4c85d12580d574a1cf8253de5a9f62531d1e7562811844abfdb85bbc4f3e52c2759a413e4212663b0fa80024ece8334cc47c6bbfbde90d90a5f279f626ff8919ff00e708a31791996392549380118cfd757e88800f13f354f83fa1d0e2a85351c491ed76ebc32724b9f0abdd3453d668ca8789d8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc161ca3aae078f2181b863eb23273aa0185d809df6dd7d5612af77c69c57d2c20854bd38f5802c4d6cd155d30bfbd2ee36a0199607b9c9c7b4e74f0f8f527c8814777bb225f86d38723f634d591814f93cdab1f1e156be2b2f0c428c78513db2fa5799e79d1f78fc053addcae6c1163693aef89cb5c5247667c941820ca86b2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha511b9fef0447c258a9ddf3b8d9416b26a5f07d72874bebd1ce41186426e9783af77013483b300f83222f3f6d2beda0a992c95f58d8c87461a43a8aad5d6dc282358bf41bb266eaed7d59f2aca27d3ec21e75ac0e60252d4a9e8801168c30263cc9464f088fb3cfa2d65712f458107571e0ad314a84be0ecc8954f113d540837;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ea63bc2a367d57aba33b537dc03cd7e09b35622fe5df414e568debe093723048630b45dc70ce945aa5f2dd1aba7651a3ae82fac5df6f935645d5275496f903ef298ee252c045a184745dd56e8627603951cc8537633ecd9bc16953e37674b2c1053dae1ed58f5fad046793374301e57fca9c12e2adeb71a085776ed32173658;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he2b1e3da247186abfa833382e51907c05ad956f70f4d403c54cf97e7955d68c1f16ec69bb9ac4d248ac13f88f58ea3df60fdf311b1721963ed6b5683b4d29b57676d183d35fc6e0ff95e84384336c2791be37a76a039e8e9a1d909cadb9a33e535d24bbf0d13a60364d1b226bd50a110053734a7af43b532a1e9d73933dba012;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hda56bae4af0f3680e1d6ffb4723b65164d8971d065ac29f51b77536086dba084ae231fe56982130da0b501289ac839febd7bb5b80afd656004ac47e0f30f6a5e35a904aff40733f65fc26261ccfbbe389eb4387fdc2212cfc5e7ebc622a80bd0b20216eecd974125d54475694ed2cdf552aefc03c80e4a48805ad485fb0a992a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h92270e70ae6145acc76eeb0340ede051e9266d899e391205885192b63e63e989d48b60a0b05d6ef3f405ecbe572b3d34d46a1b8820c7dedaaec294034db04407510794210d582966beb8e6bd20f4f01027a34121f07275b299853c1b1bd4f036a475b8e9a89f724bfecd076dc965687ef51396275894e83602a4eb5fee3a0e42;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc4fd56befd7d3cbb454dc141247076c3c2f0f2327da27a7c8ccec782ffec78240e6697223efb65fe2d134e7723c60bb2c9bb3e373eedce0c2da5a40a491185b79b24ecc80b89415ed5d30887e0218ff1465c78c36cf6dd401ece1f127e181e84bacb93a021c4572d390025713bfe922940887dbf07097d545af4a30792df8083;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h33ddb0369aad6a59f56c09ca2f8a51f6d70e0476fa824ee47e997a228a53e2627974bbbe4fc9d3834f31a0220b5bc7b815f16254da5eec031707a5cf343570a41d62485f52d7d2a0584b48b2cad8259619737235a533cfb6695ee7349a297696303cc34db9a76aa81883240f2e55486f4e7ad0dbe4e175eb22717cc65e9d80eb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h96f402782c5c95dbff65e4dea6de403e95bc6580eac819c47998aebd486321f208a99549b76ac28aeaf37fe7d6eb82be8bada69fbeb91c7176e7e06bbc9e6a4e69b84078eeb8774a0a4891b482e1d9087f3f469e6c577fb01eb7fc963d6b5539c1233e9f57552c50f4095fe356ed529310c711574f7084c495f1de767d0b818d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b73d1822b2ba8de263db973da64cde7dac97fcf77c4e712242c69ceadeb44984c0e991133f6d9b83c2c607dd0c7c16a0268bbd12c0c86b19f4893564ce9f8248e5fc4fdf11781f50d735e63493b9795a47e0f99ce4e6c03afb292cf46b0d1089555b7ffd0108a5db8aba29426b032c3e7820498659fc6b9527a58a0c586d2bf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf15064a582543428883c072ed284f441fe45ee174ce715ec2f2549acb273135f9d3b9f2eb53d7a4236eb3ecb9a9f558ad2f36cc604c74cc2ad87d0b01941a70d5af49bf29c8faef40a7a7614847696974e1cf0f6a32abb4a8cd41a377b1239dc75a21ef6deb531cb4fddf11ea84c28d94333e0dc886bb8b552473359e98be513;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h12ea61f05619cfa69e1568ca9eda074de26a80c8be724951126c80a2b9b939faaf7ef59c61f774d769bbe941ce1a3ef76685dc5b38a42d51c6b51d93e0a91f06a27bed0e0a2d90779cde30192b1b9b05da545e081433e63d8d62362a0921501186a2f0bf3f2410955e46282cccb89268d1ca2358dfb721664b4312826d8fae29;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h566a09d06ba6bdd65288db5090fbc0d9bb4cf912c4c621242d9f285adf798c5494c4fead9780b9b83f16b38d501afda5709c556a4d6ef2ac770fe259305508ba91498caac76b263d6c4a318c80d40d75cff8893c8cf11913829718c19b82d8d74d543851d51b4fbfb07a921b422e40b2fbca8a76dda818e303cfd669dd192065;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6060587276cd877eb15af8c9f98c9c8a38366a7f8a7fce37a2e16698cf74762dba913cef2b97b3bea3940cbd2297b1c316143b10730ccbf6ae14ea80d799e3140460134292054d9b81f142ba8531bd80c536d69a76b43ccea5b55e79c19f81ef5e8e832a9728a6f92bc970dbfc4c9f93a021c7ecfd2ae7814f1debc0df1dfb4a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2377251bb9c3f9b286ab7c68bbf291e43ca121574fd8e5b6d9dd274568e8158a32a0bee16920741c9096b6962a1ddf2b1ea28ce0d967d6a757b426fb215aaaa95cf011dbe0a7e74ee72949f9c8a976a4f2117dfea02831081c2b2337b8e682200d7519a4c4a16d539376610cdb8fabc2bce1b88b100e34ca796564b296bebadc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6481799a377912ba1955a70ee7d34a33d621927b3d4658c4dc3a8ceb0ee542fd1002abe00c953f085995e8d309147bb1c8a2e038c9d767e906e8d6cb65c039935250f97650aff82294c8a5e2cdcb35eb007720cf38f8805111df979dc071da036f2c62cae7cde4215f49e453658265322cb9de1af0636c0be50d482d63807a1b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h973d72d6ce7fa9506a9d830a99ed7484b276093db400fae5dff8748ba537c6272b7aa5a95c7e392fdeac64faaa28b4e5657bf460ce981cd80de384cfc854ae0afbe1a30f2d08133ffb6736cb37c7170ea730e081957b7d287d4d17836bddc93ca9acd23b85020c9a0eed9359c1fbd7f5e99d9e941b71e71500f9a7ec3f47e2dd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h43f3dbed144e35a84003445305fbf83234b3dafa35d02249ef1c4cfb11c5ae42f4fad264cd5193ae8730f4759a935c6335c02838dd1340f5e83e81a7c587326d29339368b189344212629d3f7c95e550f3e957d0f333f1f296f93230a48eb79b726a0d4670dadac8973d35552372aae6620fb980efcf69c65bcdb7ece1b7451c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd8676b923ffd5fdc771c87f324adb36512c2be55b81268ed5b7a35b5f1232783fbb135f5d222e8708d92cf01fba18f7a43f5d3262c438d4d89627725a517e7504cc1314db8a4d2c4d55f666b15439bff1a0a539165cb244b2ffe830e2b44ef48227ee7f9b3e6c9b71282f2fa0915bc03566ba7ce9675f0576b94ca1af0cdabf8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h376057c97205182b42165e8dd2f06fa8eab05b3561bcf7c0e28bb7cef4711b77145569f44dd438c591c0ff8fe26694168b2df0b4d4eaa0c8931243ecb0dc214e1eddba2d2e3e7ca85ef0cf726eee71c7b5d6b76f04719f7eecd13487f5d2e6dd55566051314c3aa8b8e5eb17763a84e94ab4cd7a200ba0871e6c9d6da67e7125;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h65a41f39de8d3c84a9f0db02d9e99efa882cdb30326fa741aebca19de4a4dbe96ab46784a89bbb72082164643c101ba6d00567765449428b1cb7970d970b099aa8accf8ee56d8315eea1dc0b2c7091e6b3b57a333d39811d432dc8fce13f94b473bd8bf87cf24b4aadee56e219dc3fca3ffe8f1fc8c46632dfad8490ac0f2fe9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha3a0fe3bedf0890d482208b5b3768f0f59cb107618ffd9b382a3370568bd71a50e2cac8fbdab7da8e5338b3dc29966c26b487ed5757bcfd616681ade1ea6f8c9b30f2a148c5d9799a81bb1e052969cfb23d1e2c81cf18ef4757e4be0a7647c85f8360a02f28a3c222388e7914597b78c471f347301a173bbf1db771e37d557fd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd174073ed6959eddf056f9a1830151cbe8b07218c14c61c7131b03349e076b8cf95728482f3643ccebb4249ca3d6faa529b67444dc733805367be871877490637e29f23e4316b4a6d38ce66dcd007cd035899501870a2caa3c5f875ed7becd9aae12999e72b24f5ecf4777b65a7e7160b5c909d47dd68c27404622034a5aa2db;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h68b829f393511e01961537b8587d26d88547a606353a2f1653bfacbfb394407b6bb93b19729bc654888118b71c73eeda25c1b6e5e84e4bb66d7b8e3edad1d1f6d0fa92f314103dc9105e611d99b79c5f92d26336a51ef936123da771cb6f6253f634521948a287e35e83c74ecdf104127158a2134c362f80c3a3898634208fb3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6a8843a1af4b1a1a0079ba68dce117648edc3b9c329df1ccf050916340a67c4f02f33511ff81bd6c1f058b16da7d9b9e94416c2c3be58d2458bde3b500a7b7355d5762053b840522ace188a1dae51e9f8bd89a7cdfed4ac0ea3b98ba3de823da5a7375f3eefb9a33ec6e6bde55f517b7b0aaeacf6748995b7445a12fa4f15c09;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd867353d31938d8ae0e37be8fa1f62d541a8835ce3859f56c9c0bd52580c87860381924a274e8582e01d7c914f255a91c4482584b93d4262f4846b572ceaf066d93169adabd82ca2a420dfe5971156010f4737eac8d518bd20adec1bfe55ba1d5724be3dbca4697632b6cc5bc21dda181e10f0f83749cb463400231faa7fa09b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h799b49adda8add1249c3de5ceedea18886fd9826da5b70c57bdd9770d1634a193c6793af1431547390b9f1f470aaa75c98ae39e80fce99338d5815f59a0dfe0884f9d271cbb357d3dd46e78d2213539c87400c7c02e9c027aa26fe10bc7fea3832e95b7a5c8f358399b2c7ae1271288204f0bb7ac9b9672746fc07eba1cce29a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf2bb129a6e323450d6c0b6eecb1bdebc41f4947cf1c5b47e7b616541c532020548ea4e03432ee378e21ca10132d4d5e0fd90fcfe072752f51b12267c31653b40f270219ff5736492734c8144d1912bd20ee98bfe89589d53d0fc37a3247eda5c7e269b66b7bbbd4c1d07bef2db290a5bb9c8e0140adec5c39383e244446ecae4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4b8e0746897da30ab4ab660dd655ed03b45b51d7d84ac2ebd03b491363a5f97b15d75a48072a28ccc6517953b52986fe131512348e6f324cdcffe33311f242b6d15587519946ba67609a134c5f4e273d7cb5e1251d541f9f0ec84424876df24c3d920b3438a05ad7392ac3598b448d670f458fc57cfbd746aebc6baf8d464b9a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h20e8d4657382cec304144ea4cd4fe063b18972b5bb2af1731f89dbc98f447b3a7cf09f7e4eb57dc8c06bb0987e0a14ff39b9cd28fe56d26a87b57ad4500343c6bb9a7ccc5787ef0ef4cd6fa9878615ef4aca92b6a3c59fd1763fe4000291e35a9ca131579fdb97cc91c65091c668a03083b382663b9900b3344e41d9c2dca1e1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h49a77faaa9327fec46f20ef2f10f79ff14dac104c20f37cc026b7f8f90d518124a474d80d55fbe0d044d6ff7d05e7b7af3fa7acb51bdde102e1dfe4c40b4327514b377cd00064251dda17fd6a3fdfb309a732c0e6b47f0470ecbe8fb6887b95c7bab37eda9a765cb3ce9b1cc7bf3af53f3b7a48f881167fa7f42289843998bb3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdfd1f54ddf8907d67926193e922f2a05d292c691fbdf6eb7dcc646228374a42d9f90d76952d777e498101662685282a890f2d635b76d72f910a3ad914a2c9c595efcd59301866524e90b616e288a928e28d778326332c618f8e02b0165712ed485e4e0b0120a6c3607fac97bee0dcd54058b2b4691ee662d9d9be08b4fc71a13;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h98d2ddd7737f141d441978211218f917d0aa26c03718e0ac9ba7215cd18ed7aaa5988122ca1995b1667f382d1c4ebdc90ce0a3f0da4694cffaf8c11dcca942e34e0d92a1866dd6357c630b679ec7ce26b81d3100f63468f67d5d6e10628764c5b746228f65d014a4d35cbeff9e99cfe864c6a6132f93cb4b9a4c17a27352311;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc22ae0395e07f3567fec5374b50c487507f52f349183ce901c7ddf36cc774527638870b3b60aaa814dcd227aaefef9e0ccbbcf6476ddc4ada404e7c0fa32e04ca99e780aba0fcbfa8806a33dafecc75b3e2009cde863f015a9a2b6d7e6947d89bd4d67fdda1f5b1233f2e3443bd1dc11e01a96434e88bcf9afef14be26ad928c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hea7bd97c0a7b1b38138f121d9c67f49a2703529f1708599fe875fdeea83fac3d36e90b2c0aeff1a66a3baeced22bc497e32c60cb6bb23d103460be578c7b73403dd62957385725eff447e95bf10448c305f834449e9ecfd6400d66290ddffa7a356d3310e95c0acbb2f062dfe2850e3f4c108e507436358815380bb1886dcbbe;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13308c9a76f6cdd84608d32b9ae82fb4573c28df75f580afd01223221f9b41916cca7a52db3d0c822064b973cad5a0346aea2a0f6899910bdb4af1cfc8f3071d8fb4f40afad9f21f17d8e8ecf900120df061e9dace10139fe3fb4f7c498305b787199fc24a09845ad3ba174dbe8114c92cc02578a147f56ba7ca421ad1680d99;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9fab13e127db1c73fd9601b4b0bc23b71aa85346a283286168954193a78d8185bfa17165b81e8e4b621254df953ae7f1d144e48094f003c05a5153f6823798b0388dc325b66d3bae2b15bffab0c7313d156e87e03aed86eaead796968221c4f2396887afb042d35916aacda65a562452eccaaff867e8081d4a20701653f2ddf9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b471f295cf5df887a753080a3ff33f7208366e1fedf537396db2a36068fc17ada72e5248fd0930bea109d2bb9223e09d9c3e3692bc7e5d26edfdf2d490a794efee6560e7b542de80ca64919567ee6090e3256f4446eaab6e16c75ace0509771034399025d1d96c147315ddb00975f47cc2938cf23a3412685041de20811e68a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h42ccc9bbdb73469cf3f8b017321486363b30ff49f0991c0cbb26e890d5fa482314d49066f9c084451cbda114336528ed3cb235e886c669939a660153015a1d3723ccb30cdd846453fabedf1e2a507303aacb1e27bfc2e3903d3cbf839fbd9191f29ab0c65a06cf5d061dd29f6a7dbfd6393977815a93264d066f082cdf408e46;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h64da2bbc97d37cc166d774e3eb3e21d239330791c241eec765f14331f14846bf240ea619e9bd90f348a677ba2dcf1f76d11af0b9b227a6b17604c36a2f1e9fd67d8a8a1a636779e4794a3ae7aeee629f251a5aa582831d5ede8e26536a51a5a5ab05b58e05accc044990e969a5e4d9564cb3402eb4c208b60a8ed81661a04811;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f13b24b1d50833e5e82d93b9bad459cfe626f0a4f0de1ed151b1c10d56745da1878d4d62fccc24adb167c6e75f5d7cf5f6b493ffb7468993cecbba44ca88d7a1974ed6048e09cc97adef9bc74acfa768c542b2ce35175540fbbbb4f45ac877e38f06bacb4e0b46696561f60277ac6b20c3ad2654f6dca51494214c9e5382ef2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbe778d22a862bd1ef02111db8dadf0a6b70d8ccad5a87643e7448779128a837e7006f2a16119c5ad01cd11a0a418fc4ea8b5793a675df7c37dc501367c803463b2298d4630c0f3a2b356d8a400e3d2761657b79ce966373b6f636ad31b4c0e4bf06a7e93c4ccde92e3f32906ae9220d924a304ee4f6c146bec436e731a123399;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haae67d20cc10ce77a6d045df969f8f67777da50fc23cc965750fb796c0e5ed011f5b8ed476ad0472fd3374a67311f143b7f7d7f4f13018987a39f31014bfa2d57719ae9ba9d1b1d93a91320a2e5b08c30187eba8e8d2cf33159b9b07ec0265f3b8a8e94eaa711f3c87f738f4af6abf4ba553ebfb1e23d55776426a4b08a5a75e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h98a46ced5cdda409e45a38cd428d1d722e668a5f693d37e4bbd9a16344b5b688a19454d4cb7b8d57b35050207a6ffe1b717978c6826abded515907b1069f21fe2ffdc305a54b9c41e762d92f7939e6e2123cd60abca75cbbec338438dbaf8d55bb85e43a7e9d9cdee916fc02dfa75c0d4cc137677ed9ec8439370516413cd30b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha35a1d9ae5a674f0b478ec7e76ca51c19019f2c3a16402b9d35dd618c321e0212f127fb633795816a3bfed99c4ce3b53870ed660925a29e44d7ea849e4a68c1b52bdf4d2ec2c7359f15c2d1b7f03b4dd258b87c218f788f9cb84905b29b3c229defe30a9ac87d7a2d8ef2a7a7ded57f6a8dc9e4f68c69f251b3764f4ddb18a48;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb65eff408c3cb5b4edcc08e0b5e5b46e734920b112d4a5dd46df8ec89228296a3f0d7cfd26085f3b99c14df5b5946bba52aa349f193bd747031648c07060a67170aa6979d3203f82a8290ec43c0e4650d6e4e2eb1b3fa8010d837490d6233f465845cab8822493202d4d6b80afbad8b4c51a78e5888efd9c7a80fb0f04124f2e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7c3bee29f519cdca9a72ad676f2052212ab271b15da69773d7260796e14c0e4340fc916db7384cb10caf2bdbb6006e1fac459c7a2be5b633878e409d0939a59abe1df9ecb0892467d3faba05911f200403b0b38eb44fd3a76c5a1b2006047bdfe4d098be7c89941521832a2e23b990a2f2d070a92ef527f332c5b834a86c1c6e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9a5ed0c02470de764cf26f2d57479f1a00ad4e98219a4ebc0731437136ea223d768d42981b1818d5beec045b8eab87da499d68be796a093f38695b5c4ac2a9a561d61cd9b2d9753c5451b7206e7178463bd78c60ecdc7bbc72032b2a250f626b90a4c02dc9803ea10ee5f60c244607bcdbb98c3fef679a592b6932b6e1518572;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7214f3f8b0e5d29cb6da2bc830e0cdd12c80f07e8f04090147ae5bd7628273a54c3034d40811d40bae9c405aea1f706eb7933e31e9ebd3f58f2e57c82cc175ad200b8d7b4d6fda9e49c5347d5f371f8a0af6b030a61031f25ef0776c87747d44fd1d97998ca355bcf70895361d71df4a0b53baeda844e7c2f9fbaa4ea800ef66;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb984b776da46398a9f1c186047dc9f5816b9f33068d9de5fa77450d04708c9362dd84f73e4a23246dbd3cff1aa8d74577d7369be4ce1f9e7e6e6cf1b583295adca1a61d92f9fddaed014c5b24eaf8f39a0e80c53f6220151be8fd14985942a2078f193bcc943f37875c240ae988009185896cb5dfa1e354716cc01fb63006beb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h89b943bcfe2bb1607867730a370e3d049e67bfddaa1fd0f4a87b867396db55345ef330c9972adf302276005464213afd68b51b5597a4093c63373e60bdda2b5fdd5888420ad2179365275de47eab5ae96c5af36a56d418d92a3961d355586db57b21855ed9659050f9e865323216a6a45d06516efc41f4bec20e4674e3b126d5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h66f994c529eb4811d821c3c217b22b828a44248707ee401849cf8df9af6a13d3a8c554786b76d313b00f4d26775389c3d12f946758db9097c5d1373bfc4810f6ee448e39089d99aa3759572a0a30c2a67b2ff418315d761ef7c7812072e0ac6560ffd08980f8eca6e6d339f1ffba3a25778bce62dd5258eb3152708942d0e813;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9ed646b4c155536f221237d5ab4bc69fe1eb878a31ad6f80d3ffee7522772f2af6fb97b392b56ed13f455c88a30828e051a46aed8f7fe9feb2504853af4edbe4d15f0ae8e9557ecb18bd8ab316b7e095d3b4830236098d39ad4be6cdcb2d7af32f8ff932aa1a9332e123794492aadd3b3ded3005ea07d757c4ba9944e25472f3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h85c38cf34abe77f237a7f82d2610dcabbde35396f52fbb5f0d7d96beaf50875d5f34af8a22252b9ab841885482439928b442d4638bf33543d6bfcca8947a7f6d7141ff9e789e2aecb94a558d665ca25c641e02bcd3b41d8544223214a8165e5e50b0820ddfafe49e3eafd3e532766ae06d211c5b982cb0ccf88fe4a2a928f607;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hedb8062b9816d3f2ba55bb04fbe97dcab665d686987999ed978ca2f9931fe2cf9262eea5fc6f1e87fb45f6673bd9ff61685bda9f852668c2da848b6f8ca0b981120b811b2fb60450b7745ca491852bd916248d4425367ec154368bf3a9a8f77b02f9da31eb302aba7dd93875577cf919d51eb97de74627f0a0fd0761d40921e6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h851038296d8e25815ed54b57c8de99051b7be4dc7e98dc2bfe0e4e1e3f3f3067c1fe26c35c9e197297fbbcb09232d72f02910f6290df476be7c57c311a0e397df98d5b1c79191f65c3b1163108de2745f281b26c15287d834ef3116722b48fc365d9488334d4739276dffe8390b9f91bc28e6c61636a827b314bfa1d190c5506;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd318579eb3603783f6087ab32ab2d217885054a5b1b4a7c8f8b8882438c4d0c46cb8bbbf2a7f425093b6dac594d6ef187186c9048fdd70744cd8502fde8528db9ee3e1ad839a57e6bb3d4050d47ca2e0ad3bfd67cf8fae39551c8bbd19e59043fe57129c322892ad26274a7f7059acc694250bbf6eafa1f0c73277aa1026153f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb618100cd2872cda5a0d2927ed8a9a8cfaf84f2da4ccf0b0614f37cb69104c696ff16bd7f543f80dafb63c9360123f6d9ac7b34456413d8c12dcc30e61dfba2e5323314bda850a9b46502371c7318486e5b90acada6f0fdd79475aad5ac5e1b691536014b7ca4a1c9bd53ad30cb86e303fc3d66c3c661bbc0eb173f567962a10;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5e1d06e7907bf0d4e803c037cf1c25466ed49e483f0e03990ee83058494350917a62ff24d9ae3ac7cc1179e45412d89e6868d4ee3f9f58d3c7f90cf7df84f23b08d90145d4653cf6ada53b4c0f97d7a21ff9036c7b025c11fadf2ba7aeac2ad59da6bc64d21d209ada582250f60eb3f9b0e064ba2b5717d28eebbee72da6e3a9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8ec564963fd291df7ae6ae12c68d9f5cfda64706c51c38a8bbdb10caabf543867c485239d2e2662fcabe2a90ba96b418ffef61e5244310d9628047d13cb39699ffe545c12fb1510293f61e53847dc6c4bdf5cde2a88128dcf2b1c448882c23f9278bb118fa1aeed709538e2333ea37c74b23fdb77a1a026342f8cec0131d36f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h742034c7e45535cd98ce1123cd181a11cbf4b0c4b9a9df9c418af4ce0a5889ce7cc366096faccec1b0428d1f7a6d2bbb8e52206338924e4f749129578a51cd8d2d668b47bc24e91d03ba462a77703b08836e53bcef262c7643cdda2024be30c613dd1dbdeb8634a9bf86baa583a0e2ab1f6c3b7f6179cc048f908168a128e7a1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he0b40bdfd15e2868bf1c930aca82dedc7bb02f27881f6f4c4ac54bf58ddcd0041fa4a3d1cf401e0cfd2b75abcb6989e4d48ca511da535fb55a6317a34135bbe9c2dfee054baa3f231764f8db08f83c61a2ccdf06a9aba3be8ad45019151f009a388d4dc9bbb4d4fc6d946c3219843311d655448cbe739c513fb3c7d11dbb5fbb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h812b0f641825880543dfc304b835aa3a8c36001bd99ad56b1bf5fe7e8365a8ca1c14eda55a22d07108dd1dfcf58b7a9425364e163c1006bd670fd54d149b12130f41e64d768cbb8249d2058556355fa24f2e0246166e47979b90cea4f362c58af08b4de0169400315cec0bd814c7b3305bdf04272086ad4d134f7d3a5b621940;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd473cf881a3367491ac476843650c6f383ee55027fb107a23bdab67d555e7750412ef254bae89d9c9476416b2fa6264100d02756bb1d652024792dd22704fd73d2e8ce6c40444b9b86137c6960afcc0c324fdfb3123426b3e4f2981febedf9e20fdcccf1fae96076c6fcd6283545a5d0a2534197960d7625e2c44d591a0501e9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h31d9f3b9550554e153dd4409bb54c96fc65752a7633f2ca44b83c5c5231bf695904c6369b4b18952c86773d14b95eac404fd8408219248cf0e8594ac1aa5b506b675a3ed63d169cc2da5fcb8db7fc8a0279f45ca2d65a15f4a2d0cc7ff1fbf047b57eb5725eb4c332ca6da8a1d007fc828dea4f55326df02289c9cf6c5d8e9c7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he03a2eb87b88a1ed551d9f84302fd84c12ee65976f88a75d25f8b8b10ab6ff6b1afa50267d60beb9799e28abc9dc2a0f0175e5d1fa34e279d34de6f41ca779680cf3656869aeb80598e6fe493efd3a05378d9931ed5a46b25a87a0dc2c2f9f036171f0f58aec11799e1d02124f2d78a77bbb7bb4e207ab198737c3f4bf4a960a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd1edc796e625969f9cdd9fbae8a02773b327d0570cf86617a071b96df624b78694400c8ffd1b93d4cc8388830b408766e85a27de0619ad81fbd069a37c0f79d749c87e7fc29ffa07b9bc2085b5d566965a7926d8e2ce5db043591c84a7b6b05c1b57b9c2489031e58fa6046ecab9ee514bd704eb0e86198fca2b42f2b782ed35;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d21a983d00061b49ba71b7c51b220641b0b7cb3a9cf70b47d9e4dabfa010695dbfaefe9ea864b6d73554f7699905d4fc97ae2126605d9c01ee14c0aac50259171c61c35a7c8d4bd20da9ce2da6eb68fe21cf23a79635e1dc7e7c52f0eaf46fd7f6648b3c138c24263f3459cce2e9bb7b027754d17d423243427e19d70508804;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd8f3d34584217478a5b377d37d4a4741b1d7030a44f88a7b78339e29cdfadfc4a7a7802c4fe1e077ee878df5219d925d10f05e9849dd995fe14de4eb4752ebb895512f500bc8a4c3affc977fe1b448e688455118a28884ad00f183f679c2eea52c1fe1e35a5089ba7e591a1b8204fd7d1637dcc9346f3255cdf3d93c1776f3a1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7573da648f6734ae86595ed584fc2b053713634ba4fad3cd6c14b324ed6cb1ab06256f647a1aa8d4d5f816a14e74963cc88d36dede2667451252e1438af882bb92cc1331312c8db419450e50089b60bd30788ec8d536fab2e8fc1dfafccf0ee17c35bc844e84e33827bdb38bfb31251bbeb7cbeb8d05c738af15b41c18c85978;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd9333c6e65ceeeb5d307dd2c58e8b6a8a65b58d93001aaed483f4224a7e0c329eccf5a62f6420f69cdb8cf49eeafc7bf1fd156337489880f70bd91a242941fa39c0b5fdb27c04b5e19a3ecad64eded327379c587fcbaa8d7ce1e8a497250ef3c06b5fcb5186e032d8026e408a8cdfb3a6325d940ee6caa5fdb759209181538;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h11fb7f40ff591a1c8fa5db9a558cb1cca1094bc1a5a6e15a15a137242f7377ec06e1907a4efe26a4b3aa33844f26886afe301386bcbda1a8ad5ba1b2b3e1ae97f909aaf83b076f7ab9530ab3ad9e0b36f309c009cbb09e46085fcbd64c507e9dbc075f34a3b80bf2fae9c341f8dc367bebfb59cc0a46e33dffcc03d6a9967232;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1f24a43aac92d512f6812436b56317ff849027dfd7e796dbabb58d17dedbbdc9d5bb073ad20ab82076e7b2d799831b0c9804a10ad18ef3083ee53463804bcb26a658bd43de39fe564604b66e72d1aee37af8086a8a284c28051aab9376d26206f0f015525421e4a7daacd22bfc85add9b5df762104ccaa77dae3f0fa61e8f6fe;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3ce65e551bcb37bcb55c209fccb031aa0147b9b3c06a3fabe6885a2c8cfed6beabc7d9f07d26a94c005f8842230448807e390b008e77ce2d49cbc205b96f257191c912f9f2a38ba89df6084da07c7defc9a298db5e383d9567c501fa06d473360c63b924a0484a182d2850254083c05d8cd18300645f56e3410dc3503c5417d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha0143365d656929b8f74775017013f9cdc22cd9f643131e1ea93529bfe2cad05e0d8715487f1112475a5dcc77300a8b561b8c50227f9656fc9512fc2c85e9403771a6806e05e516645c80a8d1184da82364ac22008351d6383a6d5e1d8d9f49d62a207d056ebf44a0bc4ad71cdb6d085521579450b94b89364dbd852e751fc2f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97e30555c00f8e2e74aa4563cc972e6aea2c04a692e6927fcefcc878e64d99dac2598dc467b48a89d93bbfcd21dcd41c74d48b3640ff89fece82e9624a2ed533f7d73ddb64f11d2a0d1d9186d78387163f1337c717046aa828f533df9e72ff71bd5407779062233fffef53c54ff7b43a80a7e2b96111fb80a86e1ccc8b82cd0d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba1a65ae51a18d0256129b182c094bd0c44a2eb6822cfde122860e28e9804308697448c518e1174d842fa639536602297960754ba51f1f0fc032fc6f82e7f05d4455bb147d9d657c3ef3745cdcd180f61913b00c27d96af5d30aa1f13774e7d9490b812700412a57f020e93f31a23a195840cdde723297401bc0d1c3d10dcde5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd4db329d5b0ec48c4618d31abcc1c147a8fa9e8b091dbfa117c38b7741e3d5d8573ee9465bdf4c3239933a226f7934cae7134e9ed6fb9e29157495d4f4c3d61f05182d2a0a5d27ff4fdad7a02f1b5a945e3b54cc6dcafd4edf81fa8b95fe82ffe46609471dec68897129694ed692676ed0db757b0c3472a0c69bbc6e70d2756;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7089a70a8dd93d8950af3e58e0251c7ad915e425f058b5136e43489e9cb8be78bc34caab4aab145dd6005070d9a28510f25de464eda6f29cc2b0f2c0ddeac86fbe22a084e0c045078354e0e26ec33fb88fc7def1dff8638f4924fba06ce04ab49238a34c2c4d56fd2307c0e873df0c3788617e43ff8b477bf87a65f4e22afe75;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd34805777cfafaa3dd1943eaf21fde6b403614634c1560f8f83f6f3cc3cb8b6ef6df43a1f692606a74df7c9d65ebef072cea8c131fafe8978c2f7f59b00b9b0f91cb1dab408432a8c50e6e3806d8a63a0ca909097a2e5acd9677afb6e91c15d3a1a00719f9c6e3358746fc9dd2d81f0c1f03a353ebc9491c4dbd5c5ed7686d02;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc2a0ddc4ca6413284bbe2f24d28e327891f112bd013a789ff847bfecdda90ae3dc5c9702ba1ece735fecf52829258830a7f71b97f8aac0597dcb3f3cc882951603b8cc0684baf30b817beca65abd0a5b56e3514280c727b15bbe7421bae2d228d599689c63787ac671e7fbaa804ab958bb47515ebfbb585c49281cfd62ab88c2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8233c4f8a4ea15e3582c79d6db07b2b0e7defe0e091b4e05288724b3d8009574b9c534f83ebc49ea01c71acc14f85abf5528993e584e7f9a0dbc1299b86268893ea98903f4266a3cb03b990a8473089e1229420d522720a7b1690a24c221c3c5a193248958698f0e79c9704520ef2118946bda7779dcc8647077e297406a0c42;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h854263c1ad990df7cfeba33a8ebe91bbeaaa2eaffb590aa2be659127a42acaf2f05cc95d07a8f9007936922941958ed6c5dbb548d6fb503a864cc6a355fa1a9c0a0ed5c1bad854005787d02940953d5f5b466f1e592126d61c743fc0cafeece0f70ead2396cf9d02e6d29c94749ef64c048dadac652c595d2c7f6cd348baba60;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h51e6b2f6570ac7edf8f1a5ed9dc77a0b102332d6715cc177d7c49655a72a71e8a517ddf0da31566a205024aae4c313cdda7705e262257c3d4a9daa78848f2adfa439be52a479e8e9efe5ba067ec42e1584f99131975829d25f48db377038315fdf6bcdf5259fc88e3e787756af968f407da6d70aa47d6603820251803a39017d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb25aa256a7b90f0ac9534f7f7c9aa85544f6f3f87a7589cea6a0262cbdd21fcfab3db1c85c302348b05c8eb34e10bfd6b46d387abd9f844398d78bf5b199afce2ef1f6c5892b14e8c082b1c0bc6825baf8b6c8650edb7b1d7bde35feffbfe74ba7b9a34c1f405bce5085e7b08bba4687d663c69351bb2943320c39447c569c0c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c419afe65b17d65fdc732af6fe4f10cf442d6404e1077c31d6e2988c4d3ead14a6380311df1a14cc163e58664a04a44e7772e041bf9bd8e95f2f2d4138dc3fb9c08a24f43ed1a130891219c34c6240de65d03c366cae20f3fb3654bc3467db98d0cf2c865315a59150a9664fe95a60faa709bf488521202a7409ba039bfd393;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4495ac09e5e84152b37887113e7a67dc6ea43dceb96375247dbb4239dcee705c2a186f9d5f24f4aed7c1aeb42f17d6029217ed7d0cdd2dba53b4c5ea0c329593a4f8ad891f5449124078d451d751baaeca6698f5d18398bdb2228cebc183a140ff1ca49fc08c0c6821af3bd1fad621d177923299e20eeb83dfead939de97c993;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he68717d89701b2c891bdc1c2e3b212af0e82c0fec2b7cdb7b52ee79e6a44c6c7c8634039a4d5cdb1894e95023add06315a5ceeb43c4dc1cd54154309f9e30084f29e7ed07d3eb7e8c2a58c8c14dff26021a86c8688a54752b9ca4ba27eb2fb37cda5f200c85f3dc2923fd61e7c9d3d887b4b4aa66a4851abdc20db9193dc8fd6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha304e4e14cb81ace6768c580ae1f69734a47f40a9ab064b80afea50c1dd1792c1455c021f05259237efbc26ee38f5bf51509ee622f7071bce6dd5579f46d87e46e766cf2caa84799de560546dc098560aca7e91486e16a3039f7cda1b1b99dd2cf64fd60f845b21aa2ed04f475bb3a8ff363eab6c046d1e16063a9c4eea22c44;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha7e4fac3faa8d984ca8cbb57ad82718f139a509bc2cde68cc9ce6c45548a75ab63d6841cb9efe20e97b3d955471125d26f91c24e07edaa697a04a5ce17e57893e6dd0b65b7339ebdf9e6653d66d6748dab15ec16f39937a627c57173452da421f87dc2048958f8450d5f0fb5573be71f448e000a3a78223f7ba0e0d1cb0d913c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8adfd2d67390654c76ba0d77083272e0e97d326f5b12ae1656d71aa7a114376a311699f8783f15131d5fab8b35b31818f14398712c07818670ba30d2c2ad2bed018396611ca301f259a228fd2a1728b46475a459b73c705cb6334fa3eb09b85db6428a10bfe8f30687af3d2d7f2ddd77c98e4cdc563320e24c23c3a635d57a84;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h27ee40d2154c3618a921515db6f189fd378074ffec2b1792a77e3ea7d354368fd398724cde46d732117fd2cd17d531f757bcda1e11590e0a5e68fae3af774f12f2fa44a705d3f8dca7c1f2da3776925d04d801b7c178dda4712edaa44310c6aadc491b5541455f90a68e37d5f2e5b1832df3078e8e704012a562c1a67542b11e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbde7485b32dc6ed85c7a928dc55880c9cb73e65ae58027b9bf175104561928683ac59386bf032fbb5f1795e74625c6123b7809b5c4c84d858d7b24efdcec1788a3f8842111fe8958c7ae330935472db6fb4822d1975518696209ab92e5b67d40d73dcfdee976bce6e86b8a6440d27bae0f0710d58e68cc0a27878910c45a0f9c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc1fa5316a6c6dd04f5b684be915b7e5abce29a5f0ed25a42ec8933e1b115d443c688b81a5d9b475cb157aca630a88ad9c8aa03a61feee6cefe0526e8566f6f73cb93a3ad226eda13fadd7d9c147a45c06df9244cf04bae25dc08b45eabdf1e904b08471fcf8399bbdd79d62c26adf0441a6bab77fb3ed8e8577e2d81f42c21e2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1228743a9205fd6012a4e6aac7ff129ff2400090ea73d79e3932305fb3225d16247eb797dd8277bec773dc23d8af5a183c161ee8872f2a9590f7589af8576583f0bd6bf69478fa087b3005b1e3ffb7d4ac89d2e4c43211ee4d5ad390338240d020706c4cd643ad4792a307dcad8bc3a7cc888546564b460b806363680109db8b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc261b4f8be0e92a48c50977c339e3a87943d0b713b7a238f857dca8d7c4638d54f3178576bf17a7e78d16496984e9e34e8ea2130ba0bef1b3bf14eb211bb47a8852099a13f144b392f6d522d68fa992cfcbd5451325951346e982e6652df7199fdddeb15ddffd8fc399893bda12820287880c3bbb12d9b1d70ff298faa7e881;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd32dc1edc0e71896db42a71f74818230a4a2e6b95d7b43dad4a77e6c26b8de476f32164d0fb5a1c87cdba912d7526c633c58e48ef7119863c6732ae8a8b535ea734d5f62055a6bf0edf71b01d23ecb350dd197e2062e3234bb0475276c3b8039700bdafe19ea2c718aba1805aeea3c4b69541ce2cfeed3fb60cb1fc7e12c933d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdd1e1dc6aceb7d586f33936a5ca1888b634a801d3ada7b21b4d051cbb4736cba982f290d3ae08ef82e6dcc88c84d3f8f62fb3febd4d0f2f45e5185c48ca6a9ae51c79ac06bae99a8a975282255ef81fd3a6f6ec783bb07313eeaab74618801205e11f78b6f357f6d93f92f2cb1de797ae21d955c9c24a53f69540bdc54430b14;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd45370d9f6bf65adf2b0643853e77b0a5c87e099854b683ca64e5571000f6367d69b61a15d0485405df719fd7578139f3259616a2acf776330b61950bcdff5bf57f078382def93559eff481197029eaceb671bcfc8b29238fbd4dd500ab562a28855d6e6b03823d2bd0d7efb0e137c129aa5c22c8af07c323fd1e693edaeeb7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ab5e12082ab4a1f4ad86321c735ca300b84289df65b266cc9602bf025ef573287e46c07bc7850a42bc070e0a182abf9059b955ea399d7dfec12650ec949956f59cb647a815926d2b0f6657b04b570f347dc2e9c3960aed481a79edaade25f1a90fa7d3ecf5a3fbea13d415219888305bc7b1b24e2e2eefddd00af44ab238bb3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7697ae818acb7c1839d336ecfa53c328f5019e5fd486820331076daaa504b314382be22908f280e3e87b12f31d3afa1e81735836e6536cc7dde15773e5963eecc3afe982dd0aae6ba92540e39a6a5a19dba05f11b47eee4002a629d6fee3623833aaf34a5ee096ef249f0e953a738059a971b8060a10dbf0fb2bf5b994675a2f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb2df0aeab851c5a2c45f3a577881060071d105a3b14c51662f8ddf9926a87a377f1818faaeadf0200abea6bbc083438bfa6f0942cd099cc122ac37fd9646462098aa930bc2255fd0d051e203b6748bd36e4c43e1cf81763d4d751be7915202e632e7007a9d55cc0390f782ee50204ec39c6c5fb83397194c6a2962af35eb612d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e608deb62e2786e1cbc44382dca184cdfd9dd0779091cf44bc2867ae78e727f05fa11a942850ddf6975a5abc5a216993229041299efb3fc1fcaf6c63c11d52204e2dc3d6c87cd2bf0b385023b248d24a9299af2c494d0c2a694e499f7e7c16e7a7ef16100cc98ac44adf87b4549cc9fada8f8a55251f603ccd5870472d250ae;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h66470955d34770ed7b6b552d598596006174198bc50db2dd9ead959bc08f4527fc49ec5096f899d7eaa2338ad528b506d2d35cef395fb48c602d502997a41cbecc6d5b715585c565a09e465139ff0e8c597af6fb7346f28909a2a64ceb82ac8a463cd00e789d788d419c65d51e52d32640d66f711d153a971b5b0e6885a9a856;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h79e4f7a7fabd93a873fe1df977327e1f632eb164ca6c2a709492ff4ad82ff536b777c9b579ea9cf9e596815ad26cfa38bfe206ea68a3e54c310348bc0987165ebc9bdc4e47e60b963aaeb83cc77344419ac18e3eb20461c7312331bda9067d581c5116c1c8278c4d33728c26c923f62058a711c3443b500ced34d3eab45be4e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had0feeb0b69758949c8f04ea13d41dbe54c377df0720fd4cb53b528cb630a975cf0e64530e4fef32dd30d71c0a9e8c42dd4abf5b3d55e6126cb18165623c8665b1ff522913a5630b4b1e1537e4e209510a1b068f3f1200d0670ae315fa5722a636894c79ca8c236bfd4b4c884a5fbb05bf32ec35a82a558c6ec0214cc6aba6a8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hea97fe2df7d5d086e1261ded4682b4470903d147aabd4550e16d39837a7aafdf741ea7ec3ed92fbbe6e595ceb8b1e3a607b0157156485bcf0c986bdcdfcdeacfdbca7d29a37e20121443025a5e156f3df0a8915d797e50927ec32b8acb33a7bc2df53197db5eb5aadb7af3d02ff75ec715bdd4f047dae68a6b0c67ba5bfc84da;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2659b0eb74e74b06ada36f609c600cbe252628ba6d6b5342100e2fc61e110cdbd9741c86bf4bc79f2879b82d89914024f7545cf670e6969068d7a4e4d8356b06c5afa57dfac7fe841ed4277eb1b8a52a8f7af9829b411475a1f3c27918930d772acdefa7530d2d94976d0abd033414f3bbadaec0d3c8cfcffd6e83f296a9e68f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha112c4ed2d539ce476994efcfa97513e8d236af769379e69dfe14f0f61c4cdc74ed253ffa4838fa27528f15bb2b4f7c8aff1579909e05ef6e247041e3c31e5aaf338d743c6572be3942f9fab59b68220992a68b82bbe066992ddd7c0bdd981ecfc3db9532f07975483cd63a4cb26db87cc45b978590e0f2a6c8509408ddb354;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee290e57c67cddd1aceb225d72cfa79a97118229ece4dcb43503e23dbb599d3f7a3885dfbbdb498f0fbdb2e6ebd4e4aed98b567cf60e7306bd25b520033ac13014870e637fd68d4f64d52fe3604638b7f27d600fd0f2773c918040245a2e8ad8d75bc38ad26ad4e65fd20677cd0f8a3d90ca35d32e9ff9a0a7d9d958c6d5de27;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcbae6447d87a0413603ccdc06d422c56ed7e11aedf5fb97ec3c5c9a5afe765f65feb8388bfecb676675e0d13ad8a20151ac3be1653f9133a183eb46902a641c3b52c0e9d3fccffc895eb283c17478751d2652c823268eba79ab1a3ecaedb7b5d78d6a3fc034d07bd1cab506cb9aff34599629c207f3cd74efcd7609a5c8ed5b1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h158ec81a41c449f3c12912eaa9f090e95b0a33c028ad8007e985332cf2082d41a5990893ea440e0777e283442587ae407f0c5216a021bd383f0a83de42de7e847c55bd5d9b64a3905cd92add4e5f148df384d362bfa2afe5edb567f9b28637ab196bb84e7372f4fe4b97c2975455f4aaff484e7e178724ed0c6166321a976bfd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c6f71da0e22a86f880976f46a85133074a0eb252a5add64731065d818c082dc0e4bbad2f39ba80e458e75b1c6c62f8f03550ad676ecc06c08c6865ab0530df15e78ee5a5f26c2c2a9a88fd9ec2dc340858dfc855dbb4fd4e8ccb8c5be73a701e9039b803456317e23b0b1989531e02d2d8f3031c2e9a89ecb6d3922e482d7f3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h386e91ce690096518f6019babda1a2705c5e8b6c6e05af56a9450363d17f19301f127813bfbb3c62f13941207e30bb6156c0545145cc80c2920f0c053e7346214b44b9679727963aa7ebcbd4aba545c3007418705324bacf361dcdd4d8030fc7c873334ecad89ce61221b80cebcc80d2ce512b1b5e00605faba51d22ad0b7493;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4624c00a6829756291f2552f2af71a3a374a9d21cc8d3dc9ff8e7b72878ece366bdd6b92ba001580a689d54cf40812650e59a11321f5f0055ffef5161c70edd1887fa4d494c054d25646833dc987633e311b0055ec48588d59e64b62127261ac3198df844022470393e8622f5eb7fad47df303341111dc20817d2907ffd42461;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3f30b8abc5f32446249ba520b71f25d9014376bbbf505287102cff6fdc9ce2411c2042b3acb7f5e14863b36a632dc233883f8b410741479c9355f49959d4bbbfb349e410a3e3686efccb37f1e321bf9aeb6e91ba77d918d64129ec12755e83bdbd74436536a7393dc061501a92bd964f27153cee4b2d2a0c6aa3aef5ddf721b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9857906f9382ca18cfaa357e90c1fcf80f2619d7d61726511817f343cc2330561816f9b97e19427db473b69a66a4f750cb907a0bf91072f7acc34c551909956883e95a70e4dc370181cbc9cc877d0e9a03f7af4e1d8dd6b589d1d0df36b2e06cd4e00339564f442848be7b621eece2895c1e805945f1e87a8788b16f617d3ff;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1eee8aa7d00f140f6f5c7d7c215987b1e3a43d353c2be80507f0e607e92c93d4932254c49271794d49fb2cbfdf6ec37e3801654301e4bb3363005757174809231905ba7aa6131bd55e05d526352341f50e1d022942150b10f54715efc4abfca980c27b42821c19298b85c16c95db8978be7c458c8b8ac77443572a3656179bb5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he1292ca4319704504e2b501157170c29555eb65245a9338ae78ebe685882fd6bf9360b5db1dc444f219ad5a82e74a1b039b11c01971d266e4f759be2dbbe6907686a52996b609deea5249fdd0f0116225bf3ef7c9eec4a9379929de27a28338d6dd0d527de95a655fea08741b5710e07daec0e23993739290117efaeac889385;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd6095feeb52178b25e00945a1fc9bcc61548bc63f27f1737efd66d06706603abdd573164e337080f31d085cfb68dcb5f77574bd1164b6afca31aa0f54e4edde5961ac0c63dc561e6b6e6bdfae0c99ae0c96e70af8a81b5a28bf2c3d50261dfcb01c85a59add711964f4ec0da7c69cf0d9674f4dd2165f718920aa9f90fe7834a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5fd21c704fa26edf87c558661660d075a8f50e52f609a92133bcade93bad7abd16b219ad3d53de3d547db22ba0c3bd30d429d27d4f4935b4959fd7effcb6e6e69762aa19e495b96db25d7fcea4046f33ab2ef1859d8e1fc59852b7ada2568ad3e3e8c1a80a6b33d26610a71616bf5a4d322b01e4feb547364bdb276b48a3edb8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4364c31d95563a79e4027ab1695e66ef690d8f226906c2ea9e9d003f6afe16eb140f1153359cb5271bcc58cb37c5a6904e1ca143848643d56cbaf2e0795dfc3969dab2224181c149fc4c3a31575b56364db21885858b0bb80952edfa9776eda8bc3ea43642ac4bd0d9e20d689e50f1a379e054a1c4898e4400b6fa01b69f28ca;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h70c80a866869e4a2cf0fe2b2b28ff7a015111941bb6ca25ba8f6eb552232a679caa604975b962a3454deef03771f7903abd8a067fbfd2900ec6c6100c621d5eb18382082d76a619fbd81dda68a51f01972b221475e21a6131c7e894587b54fdae1e3edff20ba1ff134c990e0dfdf29aa7f4e305158b9df71c3263733724e833d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc312aec6f24fd1ffce88cdf595f7d8e1a9623b76b814317a553f69695401972861b39bb7544e4e1b1b507fcb1c56497dc65392f72da8e78ca025bd430cdadd00fbe67477b234db3a026b47d15738259b20086ad19cc2224192c65a367413716a8890195582e09bd4a0a7b8304723abe4c78ac9d03e297deaf0137dd403f4ff06;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hccd9a629b4d5271218cdc0b42afc1bb03bf9cee3316bdd931d99833fb0269c062063f050c0d17d5e0ffe46a830cba8ba5d4d64db75de4deed392133365dfc3ec320e48909b774983675bf622145825bf1d910c2aa6375e1aae83ba59c87853adebc007256b14b79e494f70b5a760f02df05de1fc128229c651ca40b477bbf5c2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha9870741a8b2b7d00516f32d04c3b1d6f4c721d91c6cb99e1b506e2d17f2318b2b28f85aa69d2047f334a3355aa703584533a4fd3ef139be84d8b5c88ce79c0fcc2ac47dd90e7058f1461e1f1fc11e73e85955bcca6552881ee5a37e79b5665bee175a7d9ff8c34b9e2537ab0e4df433429edb23226d54cdbb03873e973f6880;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h578d05b6647046bd8f7ffc4b74c1f3170d71da44fca85f00eb0ebc2cdc7b6b012ae397a54bf0f2e7416f3e0f91acbec3e803c3d2e2fe45edece54fe9e0b718f350a4b5515b6f8c824cb861984fdfeee3a06dcab0e2ecc17ea34f03b3182eda13bd0975869ab534873459199901abedfd1dac4f3fd776ee0ff1307b3daffea314;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2a6a0c6558f885bd6b9f4e78a5ec46ff8991920c8098800cde51da9304f56281e6f31ec9bad85d14bac0167045ddce2574446b2192deca9725d30c68a7096a9ae8e5ac6b1a102f36a51c747c09eb01114669f151caf1daf6f68377d68b0b38c4052e060b03048284e31c442bb0a2d4f196481d66f2836005ef0c5d4c489a8350;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hae147112ae5970622a9ad27878b02debd24ba0b75b18ea3dc4b16dd79e75203c4667d8d6c828c361179577f9b8d0e7a9dcf7ab3e34a058b872429f9669f7311acff28bc3486cf4b4f42669008526c5044b7dd5bf2e5fdab795c6f1d110bdbdaf0de215beac26e005772013e4a537ea91c4dab18fd59def2a5f76656a9d69bbbe;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7ad999aa0b46033fd6556025c636266fc91a6c339fc1cd4d99543070c3b11e5a3be8daa35e3816d752f81031cb0ea4f380cbedfd45faa4445d4b9d957fbed30ce5f210d54137a9822437c91c4745a7f62ac879c6000f3062741f26d45e2ac9b968b8c1ca0ed7a72e17941de8d699056f45da266819df906a1fb38240bc9e2c2c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9c2c61bbad29d66527fddea13c80c0f04212e1edc409f301830fd7adb5af2c456ffa65ef3f66c4041238a0e1fe43d3615479ba66316bb784162a8ee675d12f95dfa60d2faeb27a30050a4240957db1ee0e880e6122356abe876741aa5833eb71f6aa5af6150de7728a2704e594ce606c8f19dd1cbea35ecf18b20a1d1d23381;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h41885055eb7a538ac090849f6fd4073cd3a23f492cf5509007cd48e0035d65b2f8a70ba94f336d49ba396acb1157c5998047c7d31a59c9a946c10a5a5349d852b7f937d2eb6605c51491fa86ca689560586a65745dcb03c13ac0a50818b737bce6e7aac857f8217bec0aaadb9acc8ec091c84e4f878be9429805e5b137d64558;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc5d0247d284cd08285cc439e20b05bb0ff05ca19d8ff1451cb3addda1d9f5de7ce9262cf40a2813eb9d651ab7600b6af94ec0050421a1fd83da72a1eaf2510108e71665b2664a54c6d6ede76ccc6f1dbbdae44d462001c004a9b191c7cb5363d1769c3d414b92a05bd036f5cb46a3dcad92d6b27fad2d7d5466e97448d98d100;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h69376467e6a779c9863f6fe4668045db24696e4dec401ede0430adda9fcfe3b83cdb974bfbb1f729237811a090f9ea068b223a9f3d67bbe675c374bb5152860325ad39d4895c675d97b77b5340762a380bd78820b161064c5be8e16032e1e975907de493bb9bd9e33681566fecd3ba075944064b4dc4f0f3239353a4a2100ab4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ca30855a8412966a9a549980af0b2112aa0e4ee1230301be71938489e0e82b1ff2ab2c6a442d2ec4d05bccea358b0e860a93721bbadb9f62f57592637643d32930b7ce418610ccac2e0552dfc74f799d1f34a80a80e2ab0a18fdc9969312fb788edcb0e56d9fded1dfad8304476fb5c9c32a9efda957560791a5b5f9457bb2b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc901d9e7fcc4eadae2a4eb346d5f8e2db1f7b4febad8ecc1138ad93e348ee5cdb147dd7fe0cfc52b71d608aafa2c23f9692a364ea89511915ddf049bb4ba831c9582dfc52661fe779db03f10ce4ff283f82d97a6202a1737f42c86e473a60dddc3912b63048b37da7fc697a58abe61f68e288edd55a5d47cf807d7d90419ba2f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd271255bf736c37b5366a9e753cf89599416cb652c4302bdc1c3f075f473d5a9ba0f7d6f24e42bd639ba92bfdb7fe6df794d96c89029d26d9cc2decb62acb558f1a79b6bb36a91245f024a93840916de31c4fcec8ef4705234da1d74cb21403362869a45398f376db574631e344a2e9f41dab37d07b794cdee0c920669b7d4db;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcecc4a12466c9d8973269736e78b7aac56ef05feb55ffdc0564c4f333c78596d40703ff9f5c58bad57e6395c06a4b316dfc6d84b37b122dacb14f145e8494a8e790911119eb0175fe0a1e4e8b318c95695c8c8f45b749c2c1e43600191d2fa729bf7bafd29e4ce687e4a61e2fe6b51623ef570f6045b5ac4f90e6093a93018ec;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73d336f7eca0d6c774ef9bd7911968a522f1eefc404ee088bff0541f5160763d8107045aa744a9db1b0314c4e97fd254a8ddb33d704383ebe0bcaeff15aa3396ce6da78fc12cfb88267298723cddb852a40eab94f1859ba19dfb24b984185afd015f17e7b71c6b8ebb5aceb83e28a12a61f46ef592f67ad6f8b95a2c4f7e937f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h807d64c32e331c4e0c29b1eed11203166e18db72850fa923a4344655dc532bc6ae56edf664e50104d7164c2ed88bcd0d4484f9dcaef005468a8bacb631afa89c5d4295ec37f38f380934278c70243f2bf6db3f1ca279123626c82359752ce035588753913b316e863f5fbebffa41a2036710ad44b2ad390a929b7356525865b5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h39f7876688d7b20bd08d3f27e839ca16c141ceef3cdd09f2362f379584c1d9be113c095bc17db33cb1a84a104883a9cb8b6deff94da13da81ed21435492fabfbe6bf2d2cbb46224d180081b98fdb2a27d49ac996de9992aa14e4bfa1d4d16b9f63e208fd620e6de9feec89111d7d8e6404edd2edcbe62b6d5af612acc2ff9b59;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hde09821e3bd92eb9ab38ac62d9488df7657071b0c7d873da9019a959538d3815b57b8ca6692a1359a1b4984c8649a18d40a91a6e3f850061fc7a9541c2b4fe71306a4f2c74b2ed879c38d917621d03b45cd6040be15f621922a283e5d0e1b9d7819bd8fdddf9a16cabbc746e6f4a49c0a5d71bf4fa98b390cb969950238acb2b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d59d27f2301272a31ad073854bdd878bc120562e936cf286b2057efc7f7d48bafe529c6e2a810230bff7a0d80dfcc9f52a86523c952252d0764fbb2a687dc06257051c1923fc8edaa7a3dbde1dbe312e1526b9333776440df89fa234dc304335a264afc2674f6552c3d70fe2b21971700a888d81ad4c16076934e92040fe7df;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hef16eb9f7fef34c77aa1961ce31cf571c3e46bd72bc966cae3050741e50dc93315f39caebf54caa4b88919fadb4da23247b3cf41843e7f927553026e96f460d50776321a8b3454cb606dcfc6561e4a56699df3f28d8b82f0999b0b1e032776d4af79b787d91e4dcdf083a74d56a22437ba22c0ad8365f19d548c350383dc5635;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he7187a058fc3083026be04ae123738f4c1b5001648a56a7a1cc8f1c177eeb4a54109384fd7f6dd90a4a25f4d06836ed77acd52283880a47f899fb490c28a29ecb64de63608e623d49e0eba91d95f43b49b43f36fe7c881a009f127c36ce8d322145d7a14ccdf4b86319243d3f0f79fedd8ab5ba2a0c3f8e506f6809003a00d4e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc71e1021e31a8b635a18a2dbad506a429b304dc8c2a2d6b4d99f908081eeb7542824e992fd12502a0f59bf7221ad25c5aa29b98c95701984f9a8651216a63c4673dc866f1a3fbda3067f5a0e9b177c2da11b9871a7992b490ab9cb4a2d447937f57a575d0bfcf66e557a55b0aab475c487d6d545c3dabc2e2d63824732305995;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfbf20a8fa757c544d717eb6ebd3ec1ea2befd82d8ce2e70c3a7f37b6faa272b64e214a2eba6d1a3bdc8d001ac075a0982961aafd9070a2d9295e58ebd8347e8a88c26a95252b90985e8ccec2a47771d120703c4a7d0940d28d0c50999aa2b85a9d01bdeeefe7d131b2246d0ed19cc1fe4b60ee058aa578e22b309ba1f501e3e5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hceb521e81d8884fec0cc6dc4aa981b44689e0a1e49ec07341595794a0b0624930e7afb3020a5030b10f141de0b366d241f22d777dbe2889756bc6c3cebf618ad7d5420195b37967f2467f8a5e8378fc66fce0196917dd057c1f9d7cbc06e3858e294c6e31390296a86d9cbc1ccaca9e2381efecf394b2f0e8bc863c6ed70bf9f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf758ef7ba862a91a7197c4e9f7b13f6a30ec2accc1a89423eb87a4b74dc8ef9b9e03f54d77596410f68c9aef3d80838483f3a17d35a0027d2b3985bb5541ce1644917759f14d61b2fcc11af7656c7613b17cbce7812282a381abb821836ba0479a344584d441b0720e5536242cb481aaf7151a1c3668ff2ab80a468f86d02a7e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haa11ae9d0ce35f86cb5cddd6af4383e77077a67cd48ddb8dee60f00aae3005bb5c76e544500bdc1810124be3befa0c73abf378df0dd0e9203196fc3923a4bd780d7191786a46df64a9b117c5d41ee5269a50dd2e858c9cb3f3397727e94842b36784caeb13aa4a3f76358e0005212de56b6f5ef1d1ccb341ae7a391cd9d9ca4f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd06b24823a420d8e363b7eb79a409f6a917c7aabedea760ca90d4bf73e91f59371eb169310803d4b1a048cc70113e7a1b300d99a2f2e5f227bf08cdcd22441c37ca1fee6fb885fe7bd03c85a3269167308b5f3da96a2ccefcabeb0823527b4dcc2419590407df32874ee5a07d89937e3a9859d0ba9e0da70195fbd995a7a1bc7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h40497d8885a8ee8fef6ef52fa80f674721d3e143e5d605821425990ec53196ed8bbef0f1db237a8deca083cd35e0f3039b8d69312421cbea4e34150945cf2bd8f584fd7b7bff4aacb03b67c28a50f40aae349b3042878d755ccb8d381a5f463c4ad1a875026b2ebe66738a2544816467814d754e39f67c27f94db83d84a86d5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2dc0ac913de022b3f20edfdeb8d3f241adbb65dc976238e14f820ecfb6640a4a67db70d9987018a5e5afa338e03b7f0a864812ba6f472a06908848453b73008affb08bf36502b34bfcc75d09d9feffeb0a60286efdcd69a06d67dd3fad352e2f5a519ece9d4690ba63dda9c7b6a7c8f6f0dcde769ae1acb6f05e06f9baaa47c1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6623d8d993cdffa99c9ad24333153804d4136eb1a5959a2052f7eda9d27628f39f392b0fe9a9391dba81c39291603e486aae6829f8df96cf03c5db56dd737ca3fa280ae1cf2157aea0151c2c32016f2336dcec8418cf6a650ece998ac58544d3ff1ee02d29c0f5f8155cb215cd200b38dd13d2c62f70f35054a249fb21621320;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h55fc6239ca5edf272ae1d52cf8c4fdf0a3c20c70ba43e31ff83aba5b4d0eb1a5556a68447bd7bb70684f2a4740a61d1359e229cca3a219db79caa8bcb8a3786aee10e73a703cd5a89f0d0824ade9404e805a1d02829353911250ed26c36026607b95a334dc18cf5bd0af7181312c2fc06dc371f8c3f4dc3202a5c9f091f41cb1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he973ab64a238a863f2882a7ef5f4f3d16d371435354e49e1dfc5c698b3019f980e7ad8d8cbc54608f8f21ee1741f99f0ae9e0b367369d637f04fcae7a60624d438a24ec7f15eea66e7b6dc952325fe715bffbaa872c9fccbf908f523388e62fd2607758013d9ca4d39501b081ba06d91bb5c4f771cd154b7b15842770bde605b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he71df8093afb1ef1c0eecb533a38a5c5ba1a04f0143838b2cc4f5ac336b9df4caca099a8c6051c3d2a50b096b8518561807135a25acdd50ea846157976e24f2381a78042883172c5fc83449f6950dc4102cc859ef0d2ffcc7ad3d43a1ac5ae9f680bd812c778df492d80715c3a56097dfcd14b6a021173c9cf244bf45aacd07b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6e42b32840ec5e2adaa0185f312c193ec26cb9b9c3f32283a6f9d682b5929d4ee9ce4f5d2c304a6de264293df72e9341a2e90f4812d138af5ef661bd47a3c9746743ddbd1ecc71e91b43c4a31e1828053e20c5c096fb88217aba528ab110f4a0a520b0cd8093945036b7a5cf452cf5b78dde30b4416acc782c0c65a1dc12bdef;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1443f938dbcb477895939a406363f310e8e95325b155ce9bc5604960169c0dae3d9795343ee4a74a9fc273cac8b31e8119e6b8299196b3634492c3b374bbb1ecba1d5707088f248eb1fc2891368881e0b28ec9c33c0563356880007822d4f74aa230bb5cf2fcf7565da25df1f2014d212ab090933adf06b2c01c7ace99acbc42;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h62d4320c469667209fe541a9be21511d83283aa78f103ff372f8b011e5674fa0e986eff4e2ec8e53efbb286ccf49969d320bf102b758900bde57ddb05c10a0c391a67e4260379a80067d1a11244b8f31a3b1baf4b6e4dd8eb3b396d5ef32dadd93b1f8c3fc826358b62eafeac31ac7d6223b0eb56dab94706a3b4296b4e786df;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5766390cc4429dfd60b8845122a4ad13951b7ecd9d6dedca96f663887030a1211d66d46e5333b1290b0ad5bfbf990e9a2aa0f8b6dafca0f72ce21ae70be09d78a923870731b2d41d8b1a43ae4933dd8db239b71523cc5cc1beaf4e97187bbfbf4bb89af9a748c7f09f0dea035d0aeb773fc7a873d6daca192bd83981c1ac0425;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he43d4860ffef2877f72e10857e67c9cb0bbef02454fa53e771fd259e4ef19465ac04314e7335ffa6f2a68179a8f6c2040237ff618469396277350cb5be1a111c9148b03d9f1a8451e0306a4a5a345a9eada99e1a3a18b4bceeee43d92a6859964f3d52f6400af91251eaf609395b8248e9b9d17b7d851695249bfb9cd87a7ba9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d93d1b324af38514fdf15346eb30b5bc5c33584509fcb7002a62ecb60cdf872286244095ad17ff0e7cdce5cf1bd5c9e1d99ef7c002a251e5d9a8728153601758a152b5a8bf62cd24db1f13558e1a48102c590f2a796db347a366bf3c90e88f4992f49382849a2ee25c3f84b2d9b9f4146b7cfe10fc02bdf14c216859749108c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8bc919daea9bf86fe83342375fc922ed7afc685379c6ca7614fe8f5894f71e0dde3e72d79b94a83d516346980b8a814f7b72bba6e7c4fda86fe1a237b8643aade351c02aeeb8e7f423b17fce5bd01f14889ba22e0409279a841b4d7d6b2d61e907a8edafacface7e3b53097dd2cbf10fde2500f2902d1131dc3c3e49c9eac428;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcaa9b351b9ab33307245009a2028cfddf3e216c87c6b031dd5686a6f1037b322a5094cd5f2cc98c5b7dd3c0ba2b43325dba54246f46590affc57f0c216fa7ae872b7a200db338d3f728dd2cd513f0366a2f731c2beb7c7da713798432d1871b5ccf8182417e0760d2eaef3d646eb96932deae51abaa505d91d07ae1b146cf261;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hff617050aeb6a8f4a21fe5f64dd5b2ca531f24095977b8fcb555d6a070cd4041f897f93d1b9e3d95f039bc653a099eec462d48ad532bde932807d881b548cc63841712618507040c0284b5caa85cecb2519b77b56ed31390c2b505f6ad4c9e515da3be41f2a8253b46a0dddf1d59574adf7061901077278014bb3935e65260fb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hac23e9a4e5872d98196edd0e1442454d8cab52970591ff8f51374d0dd15ec04958922090796566094c919f65e90c67b8ac001e1eb42c02843ef0a0700eb7fc082448469bc5b8b56ae0a6c28053b7ab747f5255d4a92cdc3e08cbfb11e10a7261f967f590a2cddbf174cfa55deb82a70b2a7c3a0dd062d58a93ebcadd0f65c6fb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h661d355681e3f322cb17932ffe0353debb609b10139d3235f0b2ce01a032d41653bdb817031ab4115e592bd264003ef6d0535d980cc66882f8347604e8568e022d3d1a3d7ee783dcc309e3a5cc164655b6e3c3ee5a70282d09cfb779fbcb9ace93d1afbd2beeffe972f527f30df71dca0ab99e2c326999f3125ddb2d0af3190c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h56aa1cd8b305ef9e14a4eb2d2ec8538cd213cd3169ce941bb7d7efcd308d7bbdacc6d3154aff9dbadb4d2450356fee2612621ed0e4a8cad3143e1570a32eaf90aa3084dfcee1056fa568da5c8bf40dd9e25cf49f907f0f109ae3d6ee70e27e40d5bd454f21df7fd574b392660c721285dd36119c3b66ea2c71d1c17d2dccec1f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf220a39d5c5a83e50e6380b274af60bb643476da28eb35cb0ddbf2b8ca78d29df764fc4308dd6fddb3c3c5c2853bc8830f0754756dde81ad020b6afea4866847591ac16c66b09f5c24b4f2785f84620f0f1fd7597bbbeece4d660abfed134414f04a56bba41c47481b551e6f685456c8a29508ff748330fe069b5546b159684;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9ea7b9bc76b87515e38680844b33d91c629355af5418a978f7bf564e578e0007d4c308d08f39b2a3b93569d607ebf2e32f770e600e086e21ba67a0ae5716ba21b9a3a9070c9d31c968a4c82ad0f107958a74d76f905084f9bcc1d897b1355a55446390e0e24b3c1944f3da0bddde9a2ac58a837822a6cd38b3a895f56320de8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h78c6a9e74eff80ddcd5a8f4e9388dd78b9fa97e2fabb65b2bbeaa050b671dc8e31b338a4959c4b2199fbed97f89146122eea35cac4aa42e18293531b7a64c4a81a701492b801ee5a0e93bdafdccf30e37133f3e819e1b92312038a1c46ed54f6fd64763a965143e3046cf8250b7995e30a38430632cc289610583c24c8619294;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ad8c8541060bd6a095bee9d458858bd8231df293a76360e21b0ac39e6da8171a1743928ff800449fe794db3549a90378d3cb440dffd225d4fc49fc1c6a21a73f90eb72375c4c4d2607cb026ac3dd3a950a11556aa7dc0bd34ea55a1471edd757db877dfb8183dc4762ad40dba7ce3dcdc0a3db195a3eb64a030b650a9e3c0bb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2be31ab9dd039f6bac69b5947375d4ba3fb605b557af99822c8796dab9599d7cc2f3f145376e62bbfd21f32a20a648618590dd1b15ef01cc1dfad64a4dae3da81e4f61542f61764cd53dad563f5372065a521fa00d9665ca9175bfef7c6052d5b791bda87e52c74b7b2913029355d23db51e3cac7f0117f351370de7bb506c17;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdfb594ea2c918ec9f0410391bee372c197245a209c4096561c5d5ed4ef7c490334776a8a4b9f53625af15a45035f7368a9292c0cd65ae682e95a4ec5df0b9c3705c7e818f2c4c48a20ae3385e627e484ded441fdae9366aca38c8282eb5606241d89bab2ec0fec10fdca2a1c1f58235cc8316daa292ebca7038ee759a471e9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h722040d95bd366a29a9921de89953596e7226017982d7a46fcfbd2d60ce30565c7265cbc381f5ba5d1af2661139b9f5da01d3b3e3d9eca4db25e5e06073c2beb5667ef345ed201528a308ad3208261134c4f5c928789fac738cb5fb1d65b0c65ea5fe77092f89664aa613553b1a1dac63f433a5a29085fcb3e5e5add359f083d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h85839ee49c67fd4990ca6c1fbcc19c412a957ed1738304abbf2e5518219c2b44a5ddbae375e44c490de31a79d87293188b9ed2c78a3c6fd51d0b8db7f8f475bf6985fc6cc8d34c7180fa09b70ce661682c5794a5f373057029483be92c4fbd5e94a5b8133ec1238f380e7aab5d1107f7a11b5a2db5a16a271a63ec90d6382c95;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h87a63a4272426c02949b319a32a46895d67b7f80fb822164f91c2319887d8bd5d6eeb0c404cb4d82047ffd6c4b1b5ef9e3dc88c20307c7e297f65dabb48b69378f42f4d599c2e89fc4dfe367ce3818fe2760e4021ac5070ddd93eecd6e2a06396b442440074c668ac1a26a6c3152cfe0d7d2c274951888a22168c52f315288c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h71f9046fdafa288835755d7e878ee8928105956abd2054cde22fb46e0ed19bd0bf0b1638d9b8fbe5a07df2000a1bab50d970b5d97c451ee12ac7a4838ebaf27042874eb3d9b78e6c320065670bb52b52d4d2c9c52521b18edda5a3c002a6355655048076cd7f4fc965574e1311472a24f724b40e58fba1f68f46294379779985;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hede223bff4f9cf7d497987aa503defd8a63aa43071f73b46f2cb9a3bc798ab5c880fd84d02521cd0086b4d0dca3cc56898979b75d413a5e63e085e98735e6f3084c68dd3cb75f1565dd0740a25fa6e8b2abac7c8ab8e4dabbacc30bc1c4e1494b3faf66e19fe0e439cc40014d5c4259d5ee91ca23bd3a88b26e8c7d8173ef3a6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb509790c3ad5e13250ea915e2e343e61dacf1f2d26a0adc9591f1eb4a9ffdb49a1e0255f35e53f42a738f684ce9a1dca79cd9edfdad7118615811952e76b1a2dcd0ab3d3e42c0eca0615c95ae9756a9de94af324fc32a984948a8267357e3d5f94e5f479361a687054d9711b6f8e99af7e27ce3975be8fcbd60dbae88adad646;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h275c5ad1a0eac9a80c65655a3997fcf2872d6f17d8aba6d9353090ccb9ad71cee0c31d41be14acd8504e5941fcdb8bd2cdd1f98deb81fb325a54292341fe5a730bcf219008a5166f9f42494877bc2b1371e52666465731dc15955a06db22e0a0c0769ab5636b4eed875a4b71c30ac6796a347bbea61d069c545651258687af48;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b5d22fde4e1ebfb6b453a09bb1b27272e8ca938f000706c484d979dbd658946057580b70b86285697b876d4395187b1edb64bea4d40ea48e691d6c5bf152db5f0db931951deda635cff6e6529ab22338993a3eda82e174cc7acb83f662c351f1664bf290c5fa9883c507fb7cd0088dc11842cff70484c451582b47f2e8dd86c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h85c1d7753ceb4f4767a3581c00e712e2cbfda79e43824ff09d83d40890b5ccc3fd0ceebbd46511a803e7b449c26da3f9a1db649e70e3a238f624bb5e720939aacac3ac116b0d3e8fd29a7a22c94e01a954e128c3c03dd3ec765a993bf44c4a3ea6ceb346ac5ab2deeebe97e405d4ccff24ca2c15e670965b897b37744c45a4a1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha2409c83e46c33b80b3b34dcd024211116369fe0c334f4482102a3d3f0a99cae5aa0b9e078a29308b7500805615fac8ef5cc0da55675be228ac4fb9ecf9ba4f7b256de787d29e019b6318e5252adb2a7a75ae194ed42082046e5e2340093bfc33126017b32d122bbb4efea15c23fb92a560972643b6e9fc70a8b28c1f4aba9af;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf75dade7ed8a15f756e22a402b9ad8cbca5495ee41bc5898b06e9765454a0956785f77e97895db360b279781f53a4412941473837cc98bc4f2ccca0c5bff950fabddc5b5b3ff1c00dbea18dde83d0b832537684936a4946d190fec3242c6aaa3b261bc09d45da9e066c5ea95e45d9e6fc910332d8cc762b1205a33d68a029a7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h266a1dd3053c55e66fa664469225b4acb871e3509bb96f9b6de3acc109a79d806b749cb466ff79fa87e641ff0d7499d9a7b8cad08bc72dff8064940fdb46d2a9300dbd0bac15c9117420e5e4fa8f4f7b010b38b8b229a39b5466fdc05d8718ad2ce9246163231e4231983261e7293b3a84a6e860d51964459f7a9cd090f2a4b9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd5c817b784242ffd4ebffcd81108bb2afae243d546e2b452346e31549a1dcc5d0bd0a0afedfe964b528033bcf0760af8513d4e131c1e77b0e021c8eee553e9620b22cb09282ca2fcf4e0f6910075de00eb21c4650bd9e21d56f984e37467dc0de6f79d7040464e7c4e03aead1255011b2e112814e806e2cd2c1b50be33835c85;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hec37258a896467208fc631fd70a1e7eacea87dcfdc908b8c8b5b58acc9a9280b61374949a1ef891f0a91b6b849eebec91f76bfd02b4841d35c92886c0aaea1edb174234a076ee50962fb6ebabcabd8ea2c82e26b3b05240efb329804dd961bbfcc4f4772480fcb77a229d837f6473d1af6277e5a0ba4e28ea91870e91c7e09e1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d7821c21b6d0e0b1ea3e20a93c0d70d7778ee95ff4901b3cc86414cd6c9f32d0ab7ea562bdb332239a5409f740845bfb643f0cb98052581ca61c7e652102b8469d1f2a1ece0e8ae6400951c6a9e08037afe2106a8dc881819f03a766c6c6e50fa5704a5582e523d95f3b8ed58433fa9b125ec655afa5cda0629d1a7c4348b73;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6d9ca699383e87be6efd2c9824834f37f1605f233839427599d8dda674acbcb54c7ff94fa2f58b5d573b5102a6b1c6d561dd0e0027c13d6d6638cd55ef056eba7cb9392a5e81e37756508b9cd0490e247311539cf13c28cc63c372c6854f2072b2b041d405dd4d998b808a4c68af6e0eaa40e925cca4626df5b9668abf3d9305;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3b00e74f71e18d97bd68636825fdf3388b2da18a65a5235b135e71042ea3d09a4382b7f61d72db1924e54d315bbaac2c3304fe59852c1114a526ebe7a1d8aeebd38e2147c71f1bbbe4b3aa14e3db655f7781b4f19e50a66114ad3e4971cdd1b5ae1deef2768aa43d014974567b666fb9d7af65c170e5a1d5bd94ad71ec6a6cb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd2bcc3544557e4d55d5e973d538a930952d266fb370a044876f842d047787bdef6a5ee098b765d8c3294cfd3e337430ce545b7fbb45909755fcb6618ba9ac6bcd04d4ad270e677af0c2cf757a6f08a74b5aa679681b8a9813d1cb86e67c75acfabb3d9fd8527f7fc9906f2208cfb3a37cabf74a1377d4b7d352bebb549c24da;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h693d7920ec1e4041971de653a4651b782aa59b92fa54804630e82763ca7c77dd4d77c41050be957780781f83115ca29a938376012f7587d4e8d49eafed51b8964abc26a248b2eef5f9709cf23dd72907dbd89a2b6fde83c196c28d4a010c8a8725a40feb7fca03d04f9bd84711ccbc7165824eb99b59f8d2f2963a62e52540d6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h88a98cae9c7855e0021f4084d81ba7ff7682745ff0621ce34d188862359abe6d5432ea0a5f355033dfa8331dbeb6ecbf52c4c6b2cf110b8670953261790db000a3a53bc98b10cbdc8c78f561b1f5ed0ac3c6c8c1a140e230a25079dcf98aea7e5738234d45a4c7358536bccfd05173eeb092c65e965c5a966bf696a80586dc05;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5adf41d0785352ac320b07903b0d7d610daa2512fbc09b2a637dac2d1abfd16038042a7da6e5df3637429139cacd0f289481743f58de268d2b2891cafaa127d9108bce47d228f6ab31ee713f31ed2b87125edf4cda5a9eeddcacd4efc0468f02d767ba449a5b33bc3b167e38e410784d6bbe9dd75e5ebaf073312e7e9c4c83a5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha97518aeeb673079bd61bf6689020bfca39871ed6cb8427c37aa6d2056d113ce5aa63034888f450a97024c4c4dba14d122f5a484a440292ab0cdf7646f6a041cbf2241365b555cdb4b143c9dfad906013e9aa32fc18d38b0076be602dcab08fd4fa31fc857fc2e016f6fd30dd27448bf3d193fe0253463e35a04e3e302fbd08d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha9d9138f534d2b445acf5e2cfdf67992d24525f9ff28a3441616733b26ff592a42c7086caa24bb09a914243ff760e181e52b22ffb368d9ee5a3bf104b6692e4bccea503a44b50d15aec077fe22edd4e67d5c1da9da7b9c67b111553e97d39282e11118ac698daf6cec558ebbb4bf3f508b2af9a5632daf4389962051d75d987d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfc2ac32f3aa7c6a81357b6ee778b465718ecdae8f3f093d09bef91cc8998d0659f025e0e9f94457e4e6d8db23945b5d2ecac032289388c0feec4bedb2f03c839cef5b057b74555e9672061b120cea3114377fa95966188ec011ced7c7b43cf967af1fbcd1f7821c16a2034ef692f67eddea038bd5655ccd4fbf93f8914340336;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8750cf4b23934a83725268e8ece7334171391d708eabf7f1d98aed61af1a22eea3d058d2c62e0b12e652008e6d4775ed4b2f9bb6f06d4232f64ceb1c07b21400f8a3fa5f394e5d53d3a23b2c4ec75ad9433d0ec02c90ebe1bd4e18b0dc29d9c4c298b6da2aa43aadb1bf9fd972eab9b568fe7855db0711b62c14c2f84bda140;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab28678838a72555cca8391da5e7111ec2e3db1c897e430a69f837c0df9dd4ac39e0b3743f19e4b83edeb237f39d65a86bfb824dff4fc2408e10a0decdf5395f4f45ea0988f866717402c66a67d014f182f1902ab3b62d5b94642fae27e64d7e00425a9bb51cf86a63ed62501acb621a9142aba959cc1f1edb311c19ef43c15;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc8fda6c281144c640ad41cd1576529ed9baac840f54e0ae4233e5bda5e1147bfec378e319ea9e8da525686d227847c45182ae5d897986bfc56c19d4bfadf2b36b1712cdab2033b8f0a6ee1b004644d97495563e29d4642a0de6ede9b942241f870bfece9bb1a1c0ceb5cbd1083074f5023f9d5cfd5b32ee406eb03f32bb06bd4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9c2b140278847d80cc0d2f564aae0ab346eb180f5b5e8c5958300804ce60c01ed50f67d261b7c6b82e401941dc988a2da554055a667e7e9edf2a2253adb41f44f4a5571debca8ea91d0ed8462d45ca559a4650be2681b977b77c50055e0e9cdfa572033f006e978307e2f7f3d4a5c572db6a2f1119be4e360a99566689b4f0c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h34d71399f0c8760fdb8752922908e935f59dd849d27da774c281383a3aa2a747e90c43ba338aa836c60fea8be2e39cf1c1a002e5d19d25cac56cf1f25afc2f2bc3f3a2527698e8e6efdcd0fc81bd8589591d33361ab43bd141f925987910d65722e64301bab6806f93ebd7f47bc63a39e62b7441a136baa6cff334514c7fe5ed;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h43f5d6cd81a317076964bbce26d9274f481c44a0519a19c49a9ea64496276617e97f33d9d62bc5f2d27d78bd2c7f6f0cdf990308744dbc6a14ce98df75390ed7c32db1467b6fe1df42c0c04c3e9997fca11297ab9f241b94ab246cddd8b6f0032ad62c912a77ff328a8e9ba3003cb247ec38a428ff2bc9c47d08c5d6b4331eeb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc0a100292291826c755f62ccc711a9b65b2389aa21c455b44245983a43b8ac7ab480e6b3deacbd21e294c6917e91428e818dad6b83f982500921a2515eda6d0e1ca401a37b85976ea9f074ef024520432e69128e060d0b1c552ba3c6287faa061b040e243423108ee0f8e3536ca9d2d674bebe9d5666f5b1efb0ef5a4fe6b51e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4c4a144d1e9127dc2a21af693d4f7f09de324a7d4a26d8f2df41be0f129da826b4133da57d126c967fb2a1083a5e71c7674e8459af38f54c51fc09615eb3c8cf7465d3fd2f57357a156bc12658605dbade7a5dcd7c285538fdafccfb0753264b64522fee5c73586acbfa38db42ad014f3a1dad0222e6674e3ec8cae40a768b13;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha54b1b44328838bb85622f6b23fa6ad821b4cc60088a161a3d9601d76f5b5e3c3a24ac6606d39b63c594b7dc92a23e67dfc194c218f1c7d1f17cfbdef2b40716eaf9f6796a638d565a57d34c5e06a92aae0721f8defa8436967510d33467d00c7205ee7b1f7927cf685f74fbf70f46512e7ba0014f04943dbeb3acc9e6676099;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8329a8f3c46d99f4c504bef9fa77c3607d008c138cf10ddfcfde95a57c1c2ab159c8871b57329f07e3c9c7d0b8a44a139e8334213f3e0927810caf74f5e0ec4f62ccd87d54113b257fcf43761b0b45805c1a7ccb795572fc693952d937302bb736878f043ea671afc5bfcd5f1f8728f9db64a54e76f19ae48290fa3aa64bbd0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc84ebd61c1c37f5cf89a09707bac5ee365177e166f605550660093c6e3fc955ecd03d68ba6176ad676472361a583197c5de2918c5f12a8c3280fc62a4879d235fec18efc445fd4d9fabc51ca60c7df35958e9a9cef39025d08665cf6aec816710a60fea8b812af21eec3976145b0dd1f02508689a6ca02fb52b3e132f2dd2218;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h47f9157382302415c58cd143e0e389bad9c701c174340a55f117eb51854044f9cad9152c2ac6af6d94e359eb8e7adce10af369251bdfc5225629fb00bb9df68b0574c03097be7c8a46009516825c6969c6bdc49f32e8dcbda37fde60efce1bb4542a9b6cf2dfa3abbe597756e25784b717bcaaacaced13471abbbe8c64091179;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37f198dd51b93edebaa4b9287656aab5168599ed824e0f88b14e4f1447fd2a68af919a8485f79e78a985ea10e4f00f450201b6679677a3ec371975574c7e9700f9ef3db1285b20a30a87f60158e8fec561ea45750c459900b6e8acf942fc1cae27432fdd33c0b111e5e512379098374fbf068cbacfa691dc5ed4035c7b75d46a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4b195b782a9341336ee7b145b51ab95ad3265d4d4b6ae327c0d52b18f69289d6e7234c001aed6e41137f1f5e3f8311030d58d08cd2caf4ab8501fac07bf7d2de57802db453722fdee712f64b32c110c925c13e9165a81041838e8ffc440afc15e686051bde1eb246aaecf30b234ddcd8fd1479585b3d6690da99afd93a042b5d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haa426c98eb79eebafe9f4f47a9037427b82e2be971f9407a79cf8e1d9cb238f06db07094abd86cc78898f6e1c68c7bacf8c0f2de166bdaed1e9074057fcb92d342c8b415b32c5144c7a80c7a98f77939c9fef27d534e8f5ab635b1aa71d151e01b9a0bd90292b14bad9af2ddc331f0562dbbdd4fd99707bbd98878520af90ff5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h28995a97f03fb2b07b8f2dae2d3f1d893c80585f5cb63fbfd16ebf5b73460429ca6c12a6bb03891ca99ab2bd9643c07560505eb990fd030a6117fcee3f1ed265abdccf8e29a3af36493a692401ccce4acfb0a661d36d50f5a5ab0153d9f613369ddee90999555f91721ff918ae0937a1857a8fc654acfaf4c1855d3f1db267f6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc455f1e76092cb5dc4099249a57f07f92c0b0aa32b0d309c5df512052f1de4b6a534c20ea6c42918332fbec99aba1c7a411d5c0a9bd81181d2ff2834b66a534d0fd3800eb51124c488ccfb00123eb88b3e77a4c0241aeae616cbe4e2ac3b964d52575f717a25e4f08160f73f776ae7b5e1104e88e2b0d2f4a3dc37407123908f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd056e1b7187858633963257388f8bd7b55d047f3ece19e39b46fc9cc1ed4b3ad6cf66099926f076b04219bcfeb66903ba07afff3c8bd5af5507579ad60c79bdcaf3c866fd6b8cbf480ac35ff5aab125ca55e4deccb9c9a826a4f9bee598c7dd1245ee98017cd01985a4e8f3b760cbeb5a88064825a316fd61e031c1898fba8cc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hda9fabd2609346ea7445c96a9964991fe95ae6c0ae16884bac89276a21dffc5ded6d0f8e1b8dadb01d815b26c993155bf03f957fd03997a314c7f7bae579d3e9725748d4810bcc80cad1130852eb95c51986ab806523754dbd16ce91dab65fa053322b0a5aa3398b8a81c23c1064766db9c4d81e9ef85350ed78a1e4fce6ec8c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6b6699514072bcc0874433e0d41f5b3e08bc33f5933bde24aa439ae634701a437ae7c9ec887d377cfbf17c8f11360bb35ccc420c0fac575486616418d5a57095ef8e844f33b86b0e6b4b7ae55e9c609198bccd44796401230feeaa0c3fb1eeb0a3b1ec11c14655c939bcb340596fdaa1786c38f02eefbcff8d9b861b50bf7af7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6d08b21d24c843ab3f4fd4a61bb67c96cae70bd431dc4d6f178cec37ac95fbc972c043101ebb94a9369c046fe95d2b48d6463c1acf0eeb376915cbe74abc4b6b29b15c43e35265a36e9c13b95c34fbeb41954ad8323f6762a209b9426fb40487895784327e5b1d4d255550dd86952acdd62270f11ebd3027df5b60454032c4a9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd7b7cf1e35045b3dd72f23c1fdc7e301a87ea2e0973f0f8f5754ca98f8801725a9944d89219895830efe45405da6807c694cfbd3a2d6b19ab82fcade61bde3c313ff2b955724a4f9087fdad34d3d604d7d00157f5461096f0cfb48191d92fae88434b10cc82114e1a2a58fa8a6dd4a153711275d796c388658be4772bfb829d2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h22025ab7a816ad5c653b88976bcd5c8c1d975d97c4beadc533e222f7e992893eab26aae82a4471a164057d17f63266cbc3a1fe0c36906566d8c96c38c5f372264bf0b8f2f25a194dd29b8eb6f34aef0a4bb3f2e748a8b5f0fc533ea419ca1c0265393c7d357c009734a481c8c70b6113cd181c05f6869d514436d84d3da48a4d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb95a70e4609e275e517b2573ce46eac5dbdd4919b340bd0d86d2836d4f1d970a30be44a5c5d95155a37b9f5282196744392e59dca5a9a1037e171bc0cdc9a01ad945650051b32ea67737670530b649a0324a7a60ff59404b0fd5263837c01c0183c8760e5cde17430a961bd02e0d9886aa469ef3d424b61f3bbba5c0ccc8f020;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h648ccd07f3c1c27ed97be94a0cc75d87459b3a3c759edc9536132b01b6138479cc73807ced18d08bcba18ff08ccb6a5bad0932f9da12450abe44859a64295001739221ec19fe0317216f43cfd9e404e9c6118d6dfb3d844dee999b7b6a9d840846ee91b1a3dea1482a77c4958b696d54dd2e31a0070a635c21dda3f901126809;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f4d71238659fd56d2a52329b0efdba83732fb8b874100bb69254ce6542a5f26234981e16c97b36364278bd1d274f77c60e457a2d6d21771ddc48fea4308d019f462b01f2139e6e692c13e3eef18613c18d59a630e792ac1ed998bd998a2cc44e8220eca4a1b9d0e5f0e78235910376c5498c3dd354f45c1f281da5ff0930c59;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdd30b076590af7a563ee4dbe4090d969310b593e76ac5aaabab59715180fe8eea43e97da9158b80bd652058c3d97605b9a19215125b9c69512d153bf666e9f8217f3f1cfd3746ae29c7ae721b5477271b73c6ef00130ff0cd570e76990c8b6526c2ab7d82700a3794077b5bf5dc0baa8ef14738f6dad0476672daf4229b78e84;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7a0ec297a7b09f4a5633d73c40ec98733bb08c2f947aeeed1e63563778ef6dc071c24bdea754cd2b37a49f9d125df3bffcddfb664402aa54ae4b6912e64e36e7bfb704f55fca6d9e18fc13146251a4159d33ea2015875579a4f7be11eb2640d9981c36cfe1e8618f84060449ef3647b82a638139f889661081a8d0d279116ce4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcffc5082844270c76b54562c386029c0c313c33a109a8e89040d2e3100e917ab34616e9536142a538dd3f5941236cc6de4f128418dab44b437b68ffa0a068ac007d33b2b26872cacf80692ee2559a4a708bf47cc1aae9fafae4336c7d95a52800e88dac4d88f7d679a86ae33dfb29d6e071a7f5bcb91cbf02168169fd4638fff;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hefd33d4b4de2b24302a017b7eadaa9cd3edf6c8df61c168cd2b3f6f45bf0c4142b33e116563af1e5a60e09a033f0e8bd5d1c66cc5074eca09b1425ed1c55e27312c21d7e701ef6d8a17836ee97efc72cf266c5316c3cca5026631b1ca48c417498b15e15e672e5243b8329b99ac3fae4e3b89bbf2bfd9f5b1cc70183c89a7b3b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1e3497ec1bf38bda27b7ee97186ee402f568d0f3cee5cb046180e58448cd8c2e0c61bf1cad4476f3397bee85eff950d8d2ddd59f46ce6e01fa9eb1a3fae6d023fbc6c063a84a3e7aa5b09192042c987c0479ad272be50c02aacc3cbec6f5ee169dceb2fbb75ef516e2ce6eb4ef281437ae3676fef4413fa8be444a5eca95439b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2fd5caa7b32503984e2969d717a21a7263c39d553c4a9b83cffed41c5a2b69324710fa0217759cac9abfd24a4b0e1d2b409d1e0830aa3d1799ae50663851a3578bf6f29f2786e1d5253e21b5b9411855159f9c9919cdbd25122a7763a9c2b9462a7dec5cc170d318598a8ab5fb0a610af4602a327d929db35d455cd3173eade0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e6fda62ac15d2b68ec509c8532e9350499ff786d94b7aa584d19ccd71aa2ae72603514f1b7fe897b05b57896ffe82384f03730776f47f0e6b9db7077b234a11a6df947d6a6525b42b5a2f10465ab788c2264fb359d6dc67ad7dbc0282ccf81869be95855cdd7c5dfd36931d21d6332264cb81a5c3b888db4e28e11bed8e19d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he34fc8ed54092f7a5b016a90b3d732423820bbe59193164f7878a331f7f4238fa701c9009ea865e2ba7f91c8bd66ebeeefdc5cbf5cb8a829b1ff405983c5ee391f9b7890934dbf79bbb3cad0ad55e7e94275f7aadca4bfc1803701869db3e91bc17e72459f3d4445f717367d9601c0a79249eb8a17f286cb7552e43c531ac3cf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd764e5951da3384dba84cae7a4ecc3eb5c8ea5284eefe3003e0b98989d3bc126a2f2a308ab621982af8265a27b19ca8146cb98e7832294db5c33e9c4777f985cb1e10714cf1c468f30940639ba51c0a5ee998a02367bcb1093ad86e959c6d08c72b865a1625f7939880dc76ff3c28053552bd7468e9db37426c3c6efc728041e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8810a0f815a9c4e0544586394165c411c1fed6083b3689a4d044c88c21476d08c99b2b20b2c8b550f6b4ff9243cf6a899e7730e86e8556a8d8abed89a33afd62c1a179a87081efb7412d253150a9a391d523b259e8b1c36e29a338759dbd66f1b582d5a76f17a023bd4a6b3849eff343c499909e45a420adb9c7743f4a4e7735;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h81fefc8272438b882f6c23b65a46358e399991a4acb9e4765045235382184c936a97f5650f1097f7aa7d7b796c501fa589f74c99b0d552de9508b8fbb0aa292b589c01ecbeb9989a843363848aee51e7ac5fdfdb2234e5a4909b0ebe7d4df1aaa1139f17049d82472b8e789806d5362143cd1ebacabd0c5f138ed807440d0fb4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h45542fc2da53cc0e90a76309ad6e7a5add6670b4a928ac5b2f19216674f6f306d661b17e92761c38bb5d76065065d969479283e981be804606c8fe0592d67359b6dff63947b6568f12a0897aa6194ebd772c39d84291bc746b5cbc80ae64846df58b03b96b133d83793378b877c19b57882137cbbc08b4f36dad6762779a452a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf85fc72f32478548d5e38a86344484ed05147407b448caf9c6b03078e4f0e987a39fff908c01450e719acef89f4c7df6aa67e9a7273032d23e7ceff4992f4126dbf831588189bd139dc718f73329995147b008a1ddea53efb4c27c4240f3885a60a0701af1cbb86823eb095b55653f9ec36fdea6cab9d7ba2c605c6c31b6bd49;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1fbbd8bb8ee70e9faf2e2524a4f8add21fa3ed0238d9b8b4137dcb726d3f89e7b0942c795a6625ec81f3117396de37d009c2690511c42c69103f65494b62c93199eb71fe243824f0d720352aa253d76be5055783097a206483c2e0ccc23bfb929d58a9aff018f735c23fe3d237e111841ec1750f805089ddfed57951c68d032;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7c546095c33a71d7834e27b7a784568b3a52ef6b69919496f6f817f176ca050d4007954ab73aaca6ebd75ccbc6733855432837808fefab110e5a826b8edea6aad129661de7b356037f95becb8619967286e0ff13ea757b04cb16b145d592999a48326f51b21c9c41766880870dd08b27bf3385b0f29b2b9bda4d5a622961bbce;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h88666a9582ff96a0f4c7082c797f5c9762790c5c2fed00255a679eaa1a52b1b7c6e849ef6a39675b3402baf414fc32f98890764b9d07814e1dbf9de9195c4acc3032dc4113549490a4138b481835d92c106c618336560b41c9a8f4593b358e2f0cea0b57cd2ae401efef6effdc0fabb48a501a917c510bd4f1c13ab913aa74f8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hedd26b983283b1ac57269a24529877fb91cff542a6637a473dfec2682bafc3669b2f19f29916d9039e612539aabcff9905831b5a5b719d4a42fc7bf247cb8f6062804206bb6fdb12d81c7fd800e8a36dc83fcc33a239f411037ad833a8a380ca4eaf975fc171739c317e734c61568ba5f99539a58e33bb9a386ac55dedd4a162;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd841d64b38a4b7251b219e9fd7b1a44b6461ac39ff88a8840e1ddb8181c3e4b883b908c5cc19244809f3da580f7da2b7d9dc0386eae82098c73e1aade4955e7152596af8d40a681b7e4a7a1179beec6ac48226a2c3fd02a3cabe35570118b1f51c92f0666bd1b2758705f154e8daddfa80e77476a1bd4265fbc137a8d7b2ee2e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5f320b0a3c67633853b7753c5edfab51abd059932b589432098310f33a548cefd2362254ae83407d5afc810952686b3d01ec15a9c8bcf0518ac17982feffea3ee1c92ea7d205a8b087ae80a1d4b9c92584e944790c655b7f759e6dacfd9559d52ca3cae5f46c6ab8cfcedd5607152e17dd0e53f8cd6280cb7c0265149a90f8a2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5721d12b75197a5df94f67ee6ec821d0b1a0e57d26f4c7386ebf9df265bceafd19a65ae6c1e71faf83fc7d453183e267e462ed0f5ff5369c2b10c1412839ebdbf2f3c3ac8add965ad71fe9c9ecff5fc5a8534d70386449e2fda271f9084381b58fea6fd7a823bd92b6f721ae8c273dba64c913dcdbe39fa642bacb8074fe7466;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9225196c09242eac2c5e450fe0bb5aaff2632b870c118f6f698841572dc3bf81bc589fe1daf8e0791dd237026ce510613774f5c00145224a823174f3853c04c07ef451c55810a693f9033feebe37f8fd0a8ce2019c1aa3b7fd198ad07b8e38dfde3a40e2f4e48dc4a32fda4d1749feb5171c4bd611c3e5f2c775fd839920352;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h832a6b8f823b78c8e64d84d50f8f8cc68a3090d8d29f0eb35ce9f7cb4d6d1cc5e2348fdc36eccdbc7c1282950d0dd59be252d92cddbae7e64b32466d714498215d931416c79f9f822b747807f80cdc1d44b1f051ee845f50866b36bf57e77b3e422cec5a8496a69f2afce53082766a8cc349b737bc23054ebdd0773fbe73b53c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3f4a2701ff506e402e0832429c5a4ef187380b62e39ecf13a1aca624a51fabcc15f6a29649abf81ddd77f9735c4a5acfc55404c942b2d5bcdf207b583c34b741e11104f98f0f553cb9668fe21a1ce337144fea52cc2046edfe34ffbac2629638ae53711dc1c9fceeafa480c65da895a67b66e5fcd37c18d51c2b156229f67eb6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc75b24591367fa24c17780200a16e0ca90eb9ec1f1459d05408d317ba87047142635fd3eb68792204cd7391fd058393f38cd5d58c9ace0c863c45e5b5b6d60bee0af885f56b30037f89a9b431508e0282b5a467412969cd58a10db281b333b244fe4a48b62e82b7d1bb04e6a30602b46617637ca8830bcfbe93a5b9d23d2a50f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h329046e932eb4e3462af1fdde6161a8144f7d443db4efe749ad78f3bbdfab27654b89a829bc9d017b5cc4c35fe764c6a126ec6fc96b002699ec98c3b6af5b3a69ddbb5543ecf4dcfa92a6e5318a55ddd8a1178ad2010f2af945b658f046ec8a2cc7053e01562441384425ff04de04235be04dbc78245b7278e790ce6898ceee2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h98be965276c54df5663c5003696ff300991e33066624b63925a54a547a57854a304d101175bc0bcafc2c8ed6c1834e6f590bdba1ae4b099b39ffb8a9250a0ff1b4195b21c25ade44ee98307ffb59ef436a06ece0e494dfa0f1534ebf5a6e222e85186d87af02ee7c44e39419ad19597da37fce8fd28235815c0bc62054484420;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7dd6bd472f9a75507b6b2ba4b4bed1c21e696cfcca6beafec70fb0aca6fb5224d4fc5c233088bb1e51d0dca004b1a36f1b201689572c482221e4c3166bad06f51dad1bfd4414b62f62883bf7ecada37e63ba55f693100866b16cf9bf938fc5fd5616be419af9e127a10a24dd108da198c803b75b49be177bc00c276275159b25;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha27c389d2c6e7f676b7df7a36c7554a9ec1fea651a893090819869f01187673d5aeb1e9160e0ab5fe96723cbb519922aefbb7388f9ca5bd40d9dcc5fdd5967824f98d37c6b9acdd49a06f8535e3287430bd014370a385dd987d823db8ae14ad9857cd3f5dff2f6ebaf6c78c223fb210f735580869e0ac0455927b3c5b7840859;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hae19e8daeb0b5b8f61ee5634d8d443c2efab4b18d8c4b9534ad3da8cd6d67f2e8ce9ec08b564e4d7089a3a73914517085dd870a693c0f08d5f82f0f63e1e683c7f6e588437272d8dcd80afdffc7c6fc9f735e62943e66daab6e640d7bfe40e3003abb29193cfd762332b9928f32a8938a0c7f6dd784d38b3f98b862ace815a08;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1bd67633635cb6818220cea2b798a42f5c1e4f8452cd6801727bc87e5490ec78b19646c94902ac264672b3d405f6b2e7a143bb820c13831adfd76835859b55e6adfc74f5cbc687e8efe0015c9fac9e5f8962854639e4bf2ca6633003cc3e25a72f9d7904c9c9b4a4729c3f020fb8bf2babf75b2645a3acf592385f91fae7cdd2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3b4fb8feb31a40e657b0004d37a6ebb8aac85daff7e35129a12cbfa8aaf7b1bcf58bcaa59d41a43a56af66d376a6df9c1d47cdb11835a268f5c6a5a5ab59b72de47a8f7e2ad04f65dc73b9c523d75aec9179b11f4ceabfc275697d77cc052c7ea7cf4748f0bdf323d9347a63c3eb7d1556ebe15b374cd59faa3d7cec9fc04f55;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h34e4f409f0be271d1ba60292b760b008b5fa14a2ba055c3ceb2667219268af30c1f1576c686a17c4c1f30e9cec233f1f7a1cd7526328f5b7356254e82b68f07c9086e9e520f4a2982a1a3c4dc2fd2d48338e9040d6729290f53a350b4468f96e6c5b266a77e3321341108fba0ff79ed6dc21bd3794c5a17b645f56aecbf880af;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b833177e00f2f7716bdef813c29fdba9c055846a35f01f0ea30b391c54c202ea6df30ec4d6902db85b59ba0735c8222fcbfb14d34391f395d6a840bc1092cdde69781f36a470c8db80fe10eee4bb2d0ae7b37332b89aab7edcd6131efd60bda27feb786f35f5b62179db02195f65bf93776b978e7c71feca7230a66c0f5b31c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hecfd6330977f2c7b089fa3aaacd492fc0ffa27bdf682941b2c8f435c7b637c992873248af74b4cd7b61f2fd66556f6b7f36d8f4522b444a7404fd49e9a88c38a3484a758c38680e7fd116c93f397eca885846103c765a005533a2ae3203503521c9f9fd0ae2bb2163ed6adcf4fe8df26d52f76419f3f06c55f68251c78108920;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1597c6a551d6fd753a5a67f7bf0668639b7a6ce77ca735cf59a291fba91ecbcf6fd277a8eb8a2dbd9b981dde77ee9d103c60cd3d1fee593899659528e89b2fffa5855357cae382897ef0279543b65f83e99565e14e5977c346c1700be89ebd30f56aaa6b4b06e63890ae053cbaec77af120e6ea78d5ce72172c7439de51a234b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h511e572860457cb44e009cf044fe2eb90e76d5a86f7b1d9daf38e6e4b6ae8e9d4514e78071c1d7bc6054c4e34b49c199726207a4adf5eec77d59ca2914a10d347857a432e944f2f4393b65725edc6d9955dcf6badc9e3d87ad03f8e29e51fea3caef0e963063b94b2ed2379f305350aeaecfc653a13b99f64ace6ddfb9a697b4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcb43bc82a24eb03827c1b9054b5588de5162f207c83ad70d843c609fc0a3dd0b51f2db0aa65f97290b9bcab0bb1adb1521ef68bcc96003aaeb6fbd16b16ce151ec2edd93f03d756b560df80771889d97fe881670ab7e1bda39c29a945a93c6415f64c59c95d2df4afb304cd897334cda3f00e06c3a4b6c6ce22fc081e7ad8fd7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf390386011e6ca0c2a9759c8d8aeb35ace78a228f06413cdb97013e4fa2d5c054a14a3d861ae2539284e984df0a3904b20162421622eeefbf2a2e9f25178fe7da4b97575708fac125c6bbc9e7c999e67ea8ffec2b7541588759c7ea269b8b4079475d72ef2c1d3a89c37805196e23076c3c71b80920bcb3c399043456fb5c93c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h91d5379c4cb6025ae066ba5a5406c6618524591dc3bed279e2595c1c765b3a3a10d4b90ab4d62a74962c3d8a6c26cf312a5580d0077dc54cc25341f64d6e27acd1c76b0a2f5f417cae20e7f3b676394abf0639fb4d2b74e970fa0b798bd90da5413d80698187b7b89ca1be6d94af71943cf7820c85bee4c4fe4f2223fbc4f1b7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha3731f0560e43001c0256442fc534af78bf9315566c5299176d19c354faafac5999070eba38003db55da8a654d202d4f0112563c210e87392715b61876fdddf52774ceb048b7f858840cf75926d548318e5fe5f2dc5309d48e68069a0a9ca44d3afb87c32616160edbe4b153f211358b8d726c123aa5cec84090d3308d9a1376;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb6ffe749514dce1f2554e8d81c8e1df2c905c429b73e83b746647bbd578b84361e45e907a251d06055a20bdb831f6c5972b0463b35ca5bfffbe8581a8fc4e7716b91bc32fa9bb11ccb23a18ae0712f93260aacf03d40b7e2e484d229d3c728233a35ed9c9c9cb7448945309999a69fd661106afa2b447ff8b83f708f81651966;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfc55439cea5597dc645a975c5f4903227e95f5ec23550c89d3e65e2ea356ee3601f3fc53fdd271bc9dfeb749d15a7046d352304f5ba13ce72342b47cdcb9a91986061883cc9ad2868abc728b284938b5c7d604f956f4fd0561fe1e2605bba409b2b716275d836ac535439deb9f14c04989711f6a8d3898070ac4c8538a16493b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfa96d6f73c09a9bfdc7d88a6dfba1c9f8e09d66616226900f9657bb1aa844acc259bc9635cdb6ff151235481cbb9874f970e22d494a169f61216f3bc65ad3d5ee78f70e205ca147bcdbbbf0b3b52cca8ece499dae15c4f6f2cef6829e999aacc9833f39f7e10d9928085ab776399c6ddb1ad164df644dd97a35bd81e3705f272;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h51c53e2e683efb1fa3ac01c740d03e6483d414e977e047dd5507ad98149f6ff708ad2f3ae753a21e2549621ea9dcb0e57e678c0547f38a88b792cd83bef8f15fcf90fb23e595c4ebe52a7981e51052fd00714ba5eefed79c9c868700b5887f189b1d717e5b53e946009a56818cb3e47f52df253a6bd23ad9c2e8a5999e74414f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7520b7a8b87a32d8aacf071ad80004582531616fc4c39144efebac3a99c7268ca60ccef89c2a73de27f2322ca7bfb7dc98bfb947816646ba872c6c1b25097194c116d9d6b087abaea922cd50b1fff9e8121d9e9dfc3a20fd0de1dac82c977cfecd6ad2471e167976d6d27b09c2a95af7a57f3661a87203afa39988e4c6cc71ec;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h53db62d91667eb93ded8ae7645a9f54f198388a18ff2c6c4a2aa3929c8e4686d67cc59d862a24fc6e25c469256ec3eea2ea578a9d7cd14812378a29fd2ad690f3ba72aede32bb0a46cc9ea11f2e994321a412011a83f2524734933647908d15c1cb70631595963c18e4d71bdf267691bc3d80897f4113ec34698b0e5c192d40c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hac6740552101ea41923f4da3c4c7238cfb88bbf1ba3dde5b683405d53cb051ac7be1cc63ba47bf2ee4cf4c1b75334c2e9f8023cd2c406793cf5ebeda36606f7e452689d5783437be8ca971510fa895cdc1f531f3dedbbba5944a0367c79b9adda055193749f98e0ee06fa5b75682e9120d1cd9c7b05787d3a71c10de528b479a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9c94b5565c006abfcb584d562f708d76e74a9529f850ac291e452191994e933a7ba537183a82cedba7706b3daa148f6550edf710fc5cecf60a7ec683021938db4b175d8007ac72942d9059a56a44e008958509b27a0fffd2904e496b9fc54ef3be0543a04275e0cf086c485d82b443059632d7c79907866b5b903db018f0b18d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he8d08e7736a7b5b413625db68872bcfd0bfaab367dcfe14c84c8962e48831cff5a966ad1590c2fc9f132d0580b6fe97872befb5cd5410afc435394792a40b868b62f22ca5d4745da9b3de75c034d4aeb493cccca7f42c9c37611087338408d26a07593fb7fa0d718fbd81d18cfc21767ff5a26c7732b62b6915180ffab7799a2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hff08b5fd7a9e02628d61a2cab19f73dc5666a966c160a9355246c2db54b158b3f29e3dfb5b5c34a6168dbdfaa3c1752a1418350936c35bd82e3b7140a5cc800104bd50d98e5dd3a5f55ff36db0ed3a8b4cab3113ea5ac2449052cf7c462ed081cb026d87969a61a281beecc2c55260a8df12efa00e0de559ae469d30de7619f2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha857363268d011131a766172c48b905406c9973cef11e649669317c5fccb8828cb50624caadd39087401a9c58bd26d4bf227f36e5979a5c56c7475bccab3f150e76bfbda1429e52bf118cd221fd4ed5af6ad74da01f9de9466e61185820510fa0cc2287e746a075a14ea122151e84b5819faabcc7a327172e907cde54c16d732;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heccef3ca65b2d6e426074e5873f143619b9b077bafd005ebd6390beff2a2d51cc7fa027c3d0338847b81a871732598cc6a161e7bd4305fc4951eb7db04be230adc8a8d4723a8d3e5ef12d94164e23b82ee9afea6532c340f489fb725358ae03155df070c853ab1fab21461837a43412c2d2808081cb1afc30a95a458a71cef49;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h63ce816120fb1326e312d6b914a2a8d7c4167c8c6af1a0e18cb89bc9c4c74145299032743136a8daf0562cb76fa0b425f62410ef3acdeca33983d9161e388ceab8a88a88d19e2c1f427ddc3d62f9a1c57b30aae969dd53450d3e58d989b5ee914c627a1f710f289ea0f9553b601ed6c6f67ff39d5c55cd59cc783a0814baa905;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h39b2e3fb1e475505dc0d7947bad4a6662225bfb742d938ac0980c19fa50d4047cc537501488f266abe2da4b222feae49939a06a6fc7880aec7608a8d4aac67ef52092ff236b4d2492c528dc010a86a89b5bc79dbb6794c9e33bbad81ca03d34bf8eb8421064d24bc58d8b995d6deb510b474ae742c030daf451c326da17e45a8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ba3215f49a580edd89cbc08880cb0ad5fdc68cb03a2324e6031bb03eca48f2bff8a8e8b8585ddbe4b335b9afaf503d32a9f4c34696c6ec041827d6450b0c04a7acc7f851ada163784ef9fcb74ed79ad192404501013cb7d4af87221fa846dec83046cbbb5c9522de456fe5d97f03be2ec5138df1e92e96a48e08eb749c36076;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfad23963ae6d8251be51711e3f5f4d3fc4825663318e5b93e283c0ebf475b276fd8b9a48cb0cc7df1bd80ab026b7e76419665ab30920cf7ba6ae93a2ec89602c03b5040187891e5242ebf27d8f61e45da861aed0abc9dba00894e989b3440b07829df27726a7f08cc99183fd19b112a6ee8fbc4e477200e4b61038ef9cbd036;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h394e13af1c3463780a0f7a787026c19c1108178b3363a75663831746c2fa24c72b5c9def915c2c9d73af5575ccf7d2071e56a6b604308878ae188d49c444acc6bed817f61d05a8a07ea0c4b4cf149cc1a98e35024191d191fce9e7e41b92defba6b81fe3e4b0fe4d77a6faef32af798faa5b959908811e62fe8eccda35aec6d0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8fc88ec9f1073a8bf7fc35abee1e822ed39ec7b7798c08312587f4294f370009ff11e068f165be7e238ae10e96e49c90c1c14245ee1a867cc2b855a90908872e7d27d8a770441fa54eceb92668784258b773e55b5281b044184e4ba701f2a1de3512ecf8fa9294e7a833a6db6c71c6a2ff3dc41f3a8b3f04af7efdaf428f8192;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h869f2afd1fb65de7cb910e0c8f64b92085ded204b217ced306709ad61911fc8b59eeaa5f276eb4104f6e60fbc4f606afa8dbe45520c2d0e2ade79d9816cd176f2caf097486c9e03de534f064880ccc1b492d410997524160eeb75306e4492975e12a3724d290325fc853beb9df672277029c189ac7d15d51b86c3b69f78d31e0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd29f5767246f941ee1f081035e87039a71c05bfd8ef6d7a64207c50d28d821548eb8c63cd15644734aaee9996ffdf10bc6ee4cd3d883fa445c82469090e22033964d3d2655eea41b920d4f8af191a8c04ece13eeddacc61260e4c3678ac260ee7f9e3322eb2de8bfc6db98a63efa6a3610274c4256a7eeda6507c7db91907dd7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h36ca46a6f7dc0cb04bae9ba10b3658c8597700ff17c1e55e59f5d9849c4228a503b816af3be3bc8ffe819d10dd264931924ea63c0a1e88927a891abbc7344c22f8ac7948e815d01372af2477abf80f987f68efaec193f3d59f6dced88e80fdda27d9dd70868fdb93216da3237317232c0c808aeaae7e2781e6d7fcbbf774a85;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h24aa1e76d3bf21676fffe445b0de347955cc5c5e7001379e19c1332188ac3dbe99e1b3836ca6534098e23a4757baeba84b06afe40a19ef0f67329bb88beb758bc3c81d1b900b18dda982787426fb946fb55e7828f27121044a5a8dd460540014987cfcfe3432c0c9ec0c528287450328b1a62434167e67e0ddf79f7818567f1a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb106487859b1168368cdf6f58b6461961db5b2d32f39ea8413146448997562541915cadf97d4685b1c1a17640caa29b56ef26852c8ae3e7fe11cbfef8da325bb3b0be78028d16f75e690d24e5b7fe1d20a01a713db24821cc184bed95477077a6758a9ffaa53dbae8fe9afab57e9816c9879fdb338b49eacdf9d5eaa12c60f18;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f2380820cb397eb3fd614fd3459c351fc9fbd5c8737ad68a647a63c5c4804f4a2ca0b13961b5441be897310cb77561ff9b174bc499420e6a43a90b01e0043e465b76ba3a51bc383490c68481de46a080996ffd6db8045533a2c930b60c605e4ef654c59d497a439873fd34914a6b76b7f44837c11240e244ecf80f303d808ba;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfbe4dd34361ee34f350babc4dc1ccd53c009227b6ff8021cdbe64f2b2d49d6c1301942a8fe6cf64f6b5e85ab8815ca933685f7f36d905e46e0baf0de821bc4b849949d6b12e41f79a1fb3c705845ffee523db28acfec4046a50634cc4d45fde306feafd51510e87fea935115a2e4354da415b7bc5df55de174a04544d6b06b69;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h387970d1a7fc3d1b2569e71ddadfc664b7f4e46cf6d4d7383ec77ad0f9cf079eadc461a015e10b9ffa6197aac7c845631dc2e8e30f29507e56c2861158f1446d18af31013bd8570ac48f006d543a992f8a5e6615e04b1a4adaea5aa089137e31ac16b508d001807b837f1f46c40b0d690de0059c678a880b191345445fa5dabe;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf1c9d0dea87995dc258ce1e5ceda9781b900eec4a78097a5b9a57ef847ef9b9a32878cc7e2f9fa72895e9a5affc7dea10f7e554c87975a51d4566176310e6d6644680c5f116a9fbfb14bbd434e75f0063821535b8c6348ef35a9efeb05475a58fb55e6c1bece70a75d4db2cc2da10af4d2505d64a2164337b7f98e82b634c261;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haa78b78895cc467886d264ede10778480fc16b6c63975ea73ed9f87ac47ac6d37a1afccaf399e1c86fd4cd98b1502033b6a5f0b55cf561f34dfab7d7829a774a5ff24672b24d58e83a5cba07505ae50eff311e30a20151196c62e4d99562c34593a261e7842b2923e1e4b1f56c5aba97dd77c6daee7ee1b5f045313b5f13c84f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h29dfd8a4f16c8e6cd16d96f64532384629c8c485d8f26caf559dd913a6b331b2e4233f5ec91be088a353149e8e849e483c79322f193fd405b25326169dae0f4f5ce1ad4fc480a6c7f4cc6324596f5ac52dbbcd5c5d593e1eea7c0624bc844e3225bab668aba227dbdcb2b5fb4b0ae62776543405b69577e8b78376ef75b2c02f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2678a3e4a9043c618505202861ff8cf51febf5dfaae0fc7c361d1f96b2e5a96fbb08921589809b1cf2f645597044ca734bbacb085f28bc309ec16c70123797f95b679aff5862a49826562b1190b94b6f68565ae00b8372e326d34bcb8759f60ff8d950515794ae9290a51a6170c2039b1151c0fbdd7bc11bb904ddbc8838a40e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6f0d2fd7fbf05883907c620c64359fe484ca5cbe21b1840de0e01958785a3c9d9ba092181a5d3b5229219415ea9c7aa39d07865324d39be5963f8a67945978c838f7d190d41063608b3f41f5ccd02abf68930bdabae32f64464d1798e9eafff6db5651661d076098b7d48266c18bb4e92b4dc6d8219778c1c2e45e1eb1daf699;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haf8f133e330ae9bd0005550b2981db9327b4ec348879bdd2e7bca29972550b438ff69ffd5d41c81106b74218c85dfdf5c8c165d49ae37576ea3277da9938b8184237cea2a61b805753898a740e7b9cbd04150d3d5944aa66b2913d1c3e7da39e2afe5dd373fa167a83865030484894723ab443ffd0de9baf433dd68b81069682;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35a389229edb87ac7083a181cb3d3df631724534ff805cd96f478b5e1eaa993984eefcafd75f72a8ad5c89e49587aa3864f7075d054b53194c425757e282e4476b9c8eff9668a51afa49719ebcd7cdc8745b4fecce0ac07509d84660bd661a97ddf0e3eb86b8070a68e84a49454dca129d4613d58b262f6d861b1a6fd6f96be2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9a3985cca1d03bf696c448da17fc6ab9ec33a9b36df472e9bd04c068eee2111863ecfeb8337d4c1725354baf62ee70d62371825322ef3356f97180cf7ad721bd4b87beb86295d36edc910cf94cbf0039d64cd24a6b01bc4c8d086090090cd16cbd310e2edaed6aeac77823a5244033a969207e8ee14cb8eee873b541c2b18de8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4273055913aebd7104aa9ef6a67f10dd5046ad475894c26fbce18106359313fcc6ca10b8cf954c2d19fbb56131f2b18e36f0adb702661d6bef644e7ba09292b3a19eb80dbb8f705211a1bfe08cf6ed8e059677e45b50b441df57b370dccc50d70ee7bc5eedfea633d6cd7eb872af8832a442b43e57a987436c51f287518a45e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4dc3c1bd5544953b1ab1af7e0ee793c5a9c9aed8fa3a2f1513d375a766e40912e2005015d8eb6d725f760c1f24016d79c34233fc1720a880a27361ec62e15d22bfaaf88985d6d5ee45ed9fa1b384292442986383094cc6e57286b0af46719d74d5f38cf82f65d88cd3eb2b8dcfecce7f1604fa5ea113a786811d1b22d407617c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had3bdd8f917bbbed391fb672bfc130cacefcb8db54e03b3b52f1cec17f69883d630641451ae05314a0be280ced8f1c285990fa65322e66fff2550815740220b9719edb124792b53ef9c4472dce022ef11703cb022b83fe3a671a4c87a76b14f7d3c2a92488907f2c27d291effdab476c1cf3f6378d582a634f6b29fcd185d227;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6cc7258aed9f55b9e5091d83ece878f971ff2ebd3cf3906bdc8037e95011ba2c41aa61b85c8ae68cbe5218eab78f120c5d5c72e4373c02e8e534d2f72e9db5a4a61584a177879ef589d17dd302a11265a38f5c67812d9d28b9981c386982e507a143fe016a8a4eaee655d92d21cbbcfe5763abbe0a02628e7bfa2c69133ab229;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha7da38cc9fbcf76ac143b21e85342f8f5673eba79554f8949fd740bb9c08e50ed4f7de75c1102781a238efa7be8d32ef3a3f51e57b473dcdd4cdb659ac8c2a0ba4fdca5fdd89aceba3789c5c5f571e20de46f9edaaf237e8050b27297b1e01d97a64ec6dcf0f9031c0bd403c7bd8d9fa512c487778da14174ad075506e6facd7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he00fc3ad92434e0382454c16cc2e1ce008ec31c3b33ac3679b06752a6e53f78a5f0bda5c40c7815e87f978b17a0803a1ddb4ad40d54808813e7b7383c9d70ad3888d4f4e5222f90727522d023206b649efe8c0238acc68ab56217b12ac6a96a522174c39467aa27de051b1d65a3ac758c605d89ee709bb028e870cbae3acd62f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2035c35394589119fc7d024f162370d2629f28e38cb47e976522a04e7bbfad2499940aba463fb72ccd23ba92406aca8e7e7b16fb103ef17a30d3ad4fc05bba0d4df779b005897b03323aa630b8729d477cda4cf6ae78fa0bfad3818e054224a65881d858da26b949015ff5cdff5ec468dea83e3d4bfad07afc9624690e12f4c3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h38939863a3d283576f54b2f8071b17c08f190a62d7389554cc297bd5d27ec642486dc95cb0b4dbbd273b9a8d940d6b6707b172e8f1c276ddd7a4da23e0a8211a3179d4a694b7286e1c2dec8bc10a660caf92de5ac45bef20ce9a195597c40c4bce8427af52aa53d241a55d44e920a2bcf4723ecc2322d3bbb5fa0fe5a9eaa1ed;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h91d4ae5341806a36590b4a0b8f786e796761c477e7fbbc1df63b8c9b5f8a2f01dc083f068dbee7e11b14d51f509a388282b77e952cb0ed9255340d83252c2252382701baf28f1737281ef42144fcc60e365ee0b8388a95861c673715c9048579e6f067eb25cf5677d5b2ba0a48fb73d7bcd274d7b00d76bb02908b25cccb30d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc76400b633a636c92e54593e9067286d255dbb4443c179735040552afc01fa2e89b0c1c63843bbdbf983158adc746c686f5748a95cbf52b7b4bee4db71cda7a853a29bb6088a168c32a6701d2f69a7c6f3dd9e09b083b8effdc02be4cd584e7e7ce90c902f5a0c46888dd0462a45ddcbe1af276d0bcf916bd196e7ca02b1966f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8fa51a72ed132de8a72e41fc65ed8600ccebc3c3f264bc68fb2950a29266d390134601ca8c3ccac161eeab9953de9a8dc4122c88b5bd32a986b5b12625863f0c990fdd6f55c6c3405d7c2d24ef5d2c07e4f742f3b732ece67ee7ca4627195e63648f96aac056c63ad6b059db055676e56fd329027bf429544bc6ea79abf000eb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h78dab36077a61658ab7167b54e8aa2f57790fe18e7de93d4016c4dd58e40fc8a74e5cebca182731749d2679630888176cacf9520a6371f4bf7bf95864c15e22c0fdfd097a9d014ba242bec67a8901b28ad622331e548cc721870362cddf04eca9f7126c3394fad6f3423914aa3db04aecba1ea344007e2b1af1b74422b355611;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb95bf171a343729dc57682d131a453f83304153a3846bbda47216f4154ab8bac90bc68dff4e7e8166ed7be7d5db33a67d3fbc6a2475d690b6a561b9f611f713f148a9b77db5b5a46da3b8416425e38763a1d2a4688a53808a90566794c1399289f1be1fb2da0fec600fd4dc7fd0071d1d8bb4294bfdc4f2c7d67fe3a4f45a0c7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e054145b04fa7f9e88c61252fce89cfa669e01946807344f72f0b335152daadf3a2c1ad483532d03ecb9f7777ac7a7c2f5eccb6ef4d5fffb6d42830bf62692d79d0a710a417f7d894adb72eb4b33c19c1f7aaea89a798bc5271fa9951d5110d06c82585d58e9bd6f1b1d74c50e09e55e2b7d1796fb38d3d83b321e7bc89a020;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h52af9463a95b362ce5e9515aee3eea7aa1f2d4bde53af5ab80fe792aa14c61a49577288d851cb16616d89a74298703fb42356b660f1a70f3f7fabdcc1a834ab3fdf720487fcce40dc81b9adf1de17737b4d71168cc0e1f986d00d7613afc0c166de34e32d343054b7468a72b7b5cc809f67b604ba7b8b3943caa685e157acee0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he8b4a2efee269018b244c06860ffc101055f3f9cc48eb87d4fd5dcbcbc193a398e9769b8bacfebb23204512b96f5f0fa084b48b75e9988cf9fa1c17ce63ba7a4e58a35a159fa4eebec638a2c57291b224c698aa131b6b62915b00612b2e185924b9b548407ac52ba87f11d6318d279f1c37ceea81d9b8f5cdb0576df3eafd8b5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6eb7657123d9410203e3ac673a1f9f6328f0cf97d6e7c72ffd79760833472c9a0288398d8b5691d88fb5f3ce75b78a91769124d5cb5db88c7b2ee7ad7ba334b06617892f13ddbfa8422cc63e3b9c30bbf21c39ad5218878a9615293f4b86c5f9c50bf0310c75b1121635853f1de0c9bebf429f274f53543981778d3d31f21f8c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd42924f9bb787075d2ccd14d91079de29407945acf9e774b1e44bd7419a40e0762cefcbe1b32f1782e89f283f3294f7087f9bffc6f709ff5d230835255aa22f9f96635b461ef4ce07275ae45bf4ba48d602f87042482a065b94789e559a21e61c80d54a8194f033094a3524c7c9fcfdc161d7744e8b0ff59d98cb81d7e7d0dd2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc88955136dce2747194f4ef503f10be58746db3879b0837009a8a7331c8892e678081f61e4e38fb3200bc8dfb3bfbe14b2bc9d7fa940d24393ba4c6ef4d88b66c5bfeb569786bc85b22c6693611bcfa7d2dd496887ee6d999a6f08c864aef9a6e6e9e387572d8a1231be8ab68fe27f0f48bc7403bae3a89ca2abc3ee918b63ed;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8baf6b9c1481ff7ea45b181e6f8fcb814c76e4c348868e524135b35e23993a6fe9e06911d7f8578b664ead8578025553c6d1c6d822cbc3b99c4beee32ab9c4fa13465489e2fc828895c47efcbb77482c26abc326e5ad6029f5b9a4e01a359afa1d0e05f2070a42295b64092d6013fad7d79849abdec92117ff4b383583ea3c70;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37e494baf28bbc780f95d4f0fc6a7a8bcd2d951af5c9d0f3bc59fbd113d050327d8e131f82c20cb56381986bc88e5fc8f4ce3dae66024e2bb9aeff0acdb50b424d34c6ecd102c58986c516bcd9654ea455ad4fae54464055bcdcbbc33bc0534c3887fa4d089f44838ea3aba80a64d459d6df26728537c8035ba61e177bb9c07d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he6294d48bcc7405c17de367f13fae2c4c09b874ed0058281004a047427bb5a537fe8dce3ccd11bee5b29bd65bd248311b85d2d20f50e32c3b7fe1c7d3e77b1a13582bf4730cbbf4dd539d4bf09f609861baf0f1d3f7ba12acc7717e9ea750ed2cef26811966c7d44df8ce86deaea3e84ee987643d56519b49020d741f355326a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb03a34a486f5a132dbe1a129f413c7b842255ad5a5634fd7257e33ea50a83c6aa82c0462990412aa8c77120040c709b59e140927fcf60d333247faf6b3fea14fb0e5991598b6928ca6260c0c8a04a948858e15c24ef0522588e7270b403e2f78541736b487a69f725d124f9b713d042a25ebee849f9f2ddbf400291ca17048a3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbfdedc618cb18b519efc92c1bf8f7b138aa5442c1511908ab1a367b7c88b49a63e377e068d8600b7e649fd52007a73fbfbb0212fb15c9fd9d63b2fa4d90b5d53e970ff134fbf7e1dd2089004959ab5e027c326e58b076e2945e2e481edb211feaed5025efb88b4e7f07ab7a193ce15fc2e19cd3f2f424a3f35558ab460d3e757;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had2b3ca28bd79366ccd2fdc480f2e6a1c253aa7b37429e56c7a7d5b30e4c7fddc3263f21aac3b348002b6481db14ec5b540198798bf1bbed731dd6c57c7620ad78fa493c46a273485f8dcdf20dfa8393384251a9e12d42213382fc0931c5ac8bcf1740e5d6c5494ebf2a6dcc5d6b908e95f73e5b651431f50ab3f622741b6904;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hda0568352d24fd438be73f9d5b129dd78c31a60698cbfa94c3e746320a3ff9548d612e3f1bf63da91f4932fbb44c955fde979de4222582506ba8fa723ae0dd91ad531860aa76e44e6f902c4aebee88874ba32881da00971d93a9df74cf1ebcf78e225251719ff9d3a827c202f3ce64d8ea436c5a884d084f4114e8b295e5b6ed;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h845f2c2433c1819024fb0265a68a258adb01cfc722d1b3d37c27f2edb6fe4dca9c9c2496b37167d5aadc92cd0441943fd0f4e88e4ea03eb2ffd90e180561a700ab6dccb9160d3b8dd0443a7bcbd4c3851a0102931648a89ba49f79e48f8f00d5bdd2eb4e002a7253669c9afed57c6ecb6319243a158fc183f429e1998bc82046;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9a41781c0528309fa89590a5e0f2c0cc1a002f94cb3865b1565c45fd24b02b9fdddfd0883c7a6559b1a61f7e57f3aac1dbb8f6db8ad5f5f87a692fdcf64db0a0d79b779a2ff6da16c2103f8de44069e9272d2ee1d0101581018559bd518bd233907daba00149a2caf3abf6c65ec988e8503ec425fe5edecae1ff6f357f0b6676;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h49392b8107aa17dbcfce5e7fc4567d368577b1690f88266d7247d08498591b9e9989b00b2942fe4faca5bca3f170299a5d7ecd8e5b7f67bd361408c451c367930ba7b96f797f53c804ed4ee54e52c0c93c5fd1aa5b35774ab61f0bb8ffa0ed6b0a8efcd96e37bab09d0d7e7c732d9413552b9cbc45aa6e27f1382e3bc52ce4c4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hda0e62983fd77a8b965172c5b689d4de618eb30a4bcbc70960cda99a14e593c8e4ed12329a17f588f3ce71823fded0d32452c6e7cf20b00760764641360f033fcbe8b6a3fe199032ad5962652f7da48f9d709d3a80e54d8f8418f572e04eaec34ad717b1146b315c5e78e239f769cae5010f584f142f79a110a8e1dc0dca8220;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4b31b5c396a86c6b044b5ec8752ab716204648a4333c9734b6d12f86f3f30f6e9ce95100712e2f78e6ae65f28b5b0bb1a5e2e68b1982caeca59114680c0b8ed301e49ef5e0ee62bbf773f2f7cc3b590225b3d8e4cb907912ef98415db9f93a08aa2aa78a61c88ff5c35c5ee0c3ba8649283ed1a1f6694ea538f32c067f2efc9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h536dc7e8ba05720d6a309d3b21f1bc40cfc133f83a4b291da3d4dbfe43f48684d797ccb777dfd6ba978b1421c3d1a85486601028be5a56641630a4d8db15e26b424e3e42e2ccc77fd677724343a38d0c63096921647cc121c073a8000b3c6ef3b26e756cbba6694e8ce537f9135a3c4afa2a56ac949b80963aef05a182b91438;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7a9b5a54a4a7c2516f1f2014c6c482b194517b7d66d25446fe7a090fab82d8d96fd406b122d81ce9dd020b8cececc6481e33c5bb2c77336f31841159bb91e91881906a889a2bade155b00748326d64a6edf365c66480184eb9015c63422da298a82c34a65e433e202657a617afd3f0c9cfa81e22adf902f7100ffb8a7020d56d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5bbd5c81f4f0f60ea6e4816aea0190c336e781979d74ece8d63a5124a7b6debb2242a3376d8aa433f3909b71269312c5caf97628b7a752a74273b81c3ec9ad8fe5c2ba155f85e4fcc4c6f945e7742cfafddcc28e650503ddc8c4817113b86db1e2d887cc78010caa77b6756d1eebb5e36545e6df9dd556f455985f0af8c19c6b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h41b235f226a5b6416d5683098e9ea7480e67fda6288ff590fd9fdbe542042348da5434ae8f6c189749d780f2618e5e0e1dfb518d8526ddda3245ccae9a13184c670ae41fd40072a4cb133a56ee7dadf02513850da64f458c3bfb0e4cb8a8b06bb10011f26bb1695defc18374a217bb46d79ec7ce067585db0fb01a1e0810e7da;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed18f10084224fe8c1c2edb575cb0c0fb8487f7b72e73bb0534044d52b869f9428b988235b7223c9ee48b675dfaaddf750e3c750caabb14de737fada48dcc7b1e991eeb4ced14e23147f254e674dcca990f50b3f2d21872de251d85418660a8a0242d4073679c02ea7e029ab7482afcd94c3106bd67b38aa011cc042d7e0dcf8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2720b50c09e3db9981ced8ea510e47227a290feb00418688ecbc6ebcf76902a8ea773270fb3a764dc9dbb320ad8ac1ad40efc0eaceeb5d417c091195cd424fa60b9fde6258ecf393f199888c8d0efe6e119a3b3d8a3934ef81d48fc574f7e96f860a076eb12c6755252963e49d4e4c2dc9a9070f35b1ea8a644748ce0fe12a8c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97917a3685f79445d1f9697ab74f7ae426ce2e187655f15200d95de189d947722081deec7a5d5cb403ba251a3a36370648038a4a5a7cc5657f2ca072490436bb1b8152779d326c478352b334ae56c3d62e86713891715cff5269ad1731f83d8e94d10fc655d8198f0c053e1387320d7e09c8cfd853ac2e62b96299f790020193;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'habd2950551cd89f17ee600ee7c84f24a16381673aeba7eda28a782aab4c5faa7d65fe3394b46126d8db05c05c0f5fe65929167b4bdeb2cb4ad76d10d980f1f41831d57f0abb8cf8411db727d266f0488244d17c2a348f7be2abefce0d3f991b7b4f6154c2b1fa2232f2a3575b1b6099b758e18e9863df11d7256cf655e0da712;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h23d69abc4883c5daa2cef3457e8c0ad9b551c07e8f150764759bd76dfe27f6db07ea10fd87accf482891bb630b7f8fb1ce374f33e20218c63079caae427fb7183c981d358ab389f104c00d48c9f3cb0508bb425904138ff482d9f3306426896c38dc12cd787351c6980943e4775456acc102f53063e823c3882ba61e3f3a3ad6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd784cd9d47cd85ce8a0827f2bed7fedfb4d9d785f1fcafd78be181319c8c6b30c4667ca07dd886144991fba5b68c8e44b9c16829322837a2b642cbf6c046bc79d250f2e7f1f109c358ba58901f3cf520cebd382db80cf288d9b0749bc55b2fa676398f73b7c4fc0dc8372c78907ac7588a26e37658880ea4dca41b40ad030751;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he4b24960c54026ed0e15598675183d9e7931a5e4fed6d6c14fcddfd8a9c2f21f31eaee4b9b25599128ec36153a7db70fa94f63b9ef8eeb1c734186efaa8ecf4a33cb76cfdf57137380ba1d6d9d49909de4f236ecdbfd9353b5ff2cd50f6316cd1d6691c167e04c94efdeabce4cf98fd00e736c5a8e52a4016892385f8bd2cf59;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h32c3d187085e84ce2e0df86d19aa879914950fed8f444603df370088de948b853fb059fe52eb6b66812c86a05e0a916b561a68c61d03d557a572557c624cf0b95ed6deeace96cc9673b7262bae9ebbc31c5af8add0862c0d4276ce98e3e1693de727fccc871970c94323d68831bf5426294e32bd9645b1a1c6c5a1e3b53bae5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbdb8407c327a2d1ea5ff2bdf5a702efc426d20d46ac36abecdc2b1a8610a568f4712fb780d1341b5ba03e30369059ab7be94137ff5199f43b52481c459ae543a26a117e612d08b326d3e1020d9c43e929315c8317c0d2bc572bfb01e64b412a35688a3b1e464f16fddd84829f140d355db2a5869a79f93a51a654b741d9fd53f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdd2cefc759aea461d78d803e920642398558d2eda0c40d8cdd4f4199deae23f9f6250d182d64205a0d5a78a0db3992644ac59fe3fd4975b8e57a5911fdea1ecd522f33900b0d5ce8a9b5a5d1ed7d40fb8d0392a964c58cf307af9651ce9c15c1017c80871ed068da4e7380b2d16d24450df1b3c814d3b5e237beb1da004fb41a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h89aa47c5f090779ab25148568af2d740906b8428613c3bcd166cc4b9fc14e04bc0a9ca6b094217c442488fe310f17bc77242200280bac03852a5dd2f9fc4721f5d4434b2b863ab9b5b21d163f178d1b3d49848f5c8359c22f309106b1f3b9e8bdd81e648ce74d12f9d29834a3ada37f39076700158cda42e6884efd7d513e060;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3ef2d3d8c8b4fb9e50f382797f9618030587616e42265518c7605f8d3a6afd0e5ba480d18b74ab4f9359e15d5a899bcbd734afb45e0900622229e58aa86ff489614556f0f06183904dc6bdf84aee9543acbfd59e475b4f5795d86c681ede251ab424cd6498475233fde4deced62a227897c71b3536dd2c026408563f9176b54e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcbea3e8cc948531b886101431a478d2ebd75c7696e494141c9c160b7a21487480595de7dccd3b2c082813223c7fee4dff2d49f7fdd08f612f1de1dfcfba22b05a31748f4d6cc70c354a92f787538b1a34699e2aeffbf5acc22a1bbf2e0c8840552709271f2cab414b9eabcff3ae6bab92e4a9837c934f3392412070402cc07a1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd43ab434198ed49b8b275cc72b2a6db1bc9847357f6731343bf3c601b29a4e3c02b5913b58c0727599071cf9a062d9450829feae8ef2be1f6c14af67708e997944d81c23138893dfc16662a397eea55d4409005a1d6bba84a77c8d890329e785399315942090ed69717d69facf527748923d10dcfda05eb4136057154671f304;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he9a32b5c2b3cc4bc01c95c068d7a3d52ad54b1abd245cf0cc53b19114d374797d539908134dbf9c8f0b16ed5158c0bd1acdcf4e12aa9cd7218fa0eaa188207c311bcc53f4b65e10cc84221856b843773bd03016009ede8e5194e6ced7215984e04bc620be0908f16bf4e3700a4719d38611f69fb3fe23fed46ae45f9c55f49b9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5aecef4469785e67a04bf773644ba584d7bf277630b021b856f5beaabb53c4cef79688c945ad742f4c13c798995966f88bbf6496b3a32842f80f49ac502686957db9a681b273b6dbf7e05cec636938377d32fbef63d60a4a87d15b5d4d2d1d5e324e1c8aca65695edc01e5c64e91cfbbeb30a52d2de72795701027c83112f2b1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd07b17527ff0a553fd64134fd02e9b89d0671f67246d6a2a5f72ddfc14b36ebb678666027b27cad719cd3e2c509c630bf7da9accc6d124994390bb11916bf5441997bac3e79ac80deffa3769eddc29f6ca10360107ef6f9bf3bb79faca763cee1bdd3dfa7679abedb8c51e3ef33854ea822da6585c9c2aa338d79a7f5a79ef7e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfacd371761f22645e627ddbee0b456a50b428cfb2b9e43cf5c0418704382aab7629894b62ab12fc2cbe9a407f878ce1f7447a7ef9f02fe3158cb64a2973a59a6516482762b1047de860ecbf18e36c8659f7dc480208d5a46fea7bdfd9009ed42b391b6849b7e42f55da72ec5fb6dd7fcb43a2f652a1911eeaafafa2a548881ca;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h89b9ee35eb36bcad1f6fdca7abcc624e5893faf44df7fef3b475dd6c345f0e71d94105802257ee31df52e388e6e6e6a49087f3979265920eb4a865712369897227d357641376c13cc92692a3002470413d4b9a93b1da446cad2b0e5db093bc3beb4ea044e07f1534ac83d02a1f47acf2112500e6711ea95106cc52d7ab42b05b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb4ed642d5059c43cc5bb0345f2ea752e04876b02b31baaea0c81ddb5ff8e26118112b36a27345658d1e2e17ff6d98202e44751bed0cfaf07163cb1c7af82c66fa29418f33601bfd315e388afaf097956a2e97592890386ddc282882027230becceaea2eb26841de8867f007cd0330d255b44d5611eeeed507ffad52db2182009;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6f02303495c301b7290805610b9659056110e0ff568c282ba8dfc60c5d48f86b4c52627dff7afc9fced6ddc296714c8954c20b4b6b30ff095dbff86d98df64e35e4216e0e7bf76dd30cf9e8462d58986346e0f1ec9bf51d4af3b4afc324faa065e2f3aec4d00d9f31530732d2f56cd5ba356a3f70aa447a06cf40cbb3fdc168d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1775e6f1757cb811c7e9c249c14cef540fac8af094759ac0b7cef98ead04536fa3bbea0d57bcac7a5ba85eff3a7606859006fa1be08ce1f77e5f2017f1429088804204acca1a37704d706b3b5e546407c3f57fb71a5a7593647d950f066d3a5d5daba5b8caff605018ce4e418fb531e51a06c128a73aab05d324fdfa4c2c5c9a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9ca429c2a5250398f7d597fd81251496443c16353743f3197124cbc8b928984b6f9def616524fb20d9aec4064dedde60d01501f8812147947eb184512c89e00118e9e7949ccc32a113a7b5cce342c170ee702d2ce8be60afbd4fc12275713ad34c790e0efe4ba5b014fe16b4dd42a8114deab583ad0fb5282fa295b72064a746;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a9db1d67a3005f6c299ed7718072e09a6478bef5b435ec1269d77825c72184f5d2333e420685e96cb0f821af433058899ea6a05a439500cd354abb6f78ee8c5bad3b7ea91a2c2bdb58fb3e30ef60033ce5812e3e36be6f97c425a71dd54a4b75965f52d8d9187a75a4a9506dd1548b68792790a780e1c4215f69b719ca67811;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e280ecf17723b76216aaae3e75dbba72d47f3c636d8e81cb48d3bfd29a85d72dd29474b3c2f097ff7c88465b3928725aad896905948123dc888f3b644a6eee80934fd32b234c1f116c7bf7df132c32276da701b34f7a33adafd12388e54ca781981f0ae26da75ab9441242dd5e1a82c410d2deec8ded842ba2dfbb2b7f9b0bf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h788ac2a950f6e6832ae3db57937e9f93a01ac9cd66c0d218befc5a189c1ba18592d85cc647dfc7af48de16e67d417fe1246ba686454b7285c4da1bfd8873777bb90d1f73c5838630a9dcdef3477dd77396cd08a4bf29abfd9f4ee5307d56aecaa3fcf97f98101fe4caa7dc3ed0b235edf096f1cbf1f7c1b7e928689a74959b41;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h681e65308b54fa58683b564b1e57f8adc48d1ef71295202832cde402c6482bcf7d4795675424980a9eb6952eea777d113cf7e82d74eb1cf1c4bdd945d02870c6f1d143bcf59f2527ec4f52f9aa9878826ee9aa6ae091041cbcdd3ed16d40be8fde315bada127a31f629d43c257f8903b43c221aca10a4e430e281dab6e654f17;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdaa3a31f4639cb5bd358f82e683ff8b1595c4a520fd15d1593241a4b5966e7aff6847ba2f81e083fa2bfe203a909fcf19845fa4bcdfc06cfee9bafddece521a9fd84120fbe7218a4c01ef9591a21701b26028aa4bf0262078a4861142e23288908bdb524483b3ac30ffed8713f95586a9c519cc5e87aeb40b9b020faa91c6e16;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he5ab47e4a2071753ee725479a31d2151cb0b226864c1730d4597a057b590985574b32d840fea3b88988e5dedf2914efeb08fee5a1541ecabd2eef18aa5c5f02694465363cf31d47562d804d1d579b2d99d2c2fe7a229e5c364d5a0723c632c3fc3f35e53b7922cd3d3b5f7e0cd26341493e3fbb90d929880127abc644ff166f3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e3e07c6cef31239e7c97d6135051706ffd62aeb869685d8c9e7b959b1a0a9a3301d323e0e137f4972b831b47b06027c33ce4a205b823e87ecb64d32f2b521bc0fae58384354c59cad79b0fa0053b10cefc5ca057bc5a4dc1496047f267f9b8926007aa0d43e60fca0049f656d4e7b028af67c1e1334d80c4f9c9bdb039f6ab0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haf52bbabcb0b11bb456545f30eace5b32606a7541a37f1d4cb521dcffb283d120bc162f9121d24cf0a2e97c62091b10e77408e67b01650d3c045a0c0f5c009ee8b35a0024482d4c767d62bf65d93ecb17e68c4d4fbae5677c3ea7b12d46c49da840e804e609e4a986392ee58be83ab2b3e443cf7c103e39edf93dc4fe07434b3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f1b527724d8ad2300bde935178c678db104cb3e046be700d1dd987bd82dce64fb708a9c3acecff0eca0e1a21036929dc2c2ec5976f4b8536c27a4aee6b5e4175af6c2e4e036cb73aee23c89ef776313a0846dd0513c3b1114f63c570e8dc5e7dc87923e10f96ee9df767843df35215578738984e676576391836f15df19dac7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha5f3b4ce927c7d99c325a0167582deafc2891a8328c08294bedb8d2b9e872dad6ecc11ce041372db12c4908e6a676f988bb7d30048596186af3fc1a7711b476d217a604d31aad6feb193dbf8af547cca55495ad768d3449799c15844e1e39d0bc5ffd9279e064f569d3657d72a297d670c5a22c1d405815b0aa9f9fbb02974cd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h66a038900dc18a7089eb2049456d48f6c2c9acb90538fe102035e11505a0eb4995b3525b3fae63906cee67747f867aebec4838f72cb581cf1d7f1c580cc3a3def0d97ec1464b6c1a226c64400443cfaf611b2fee62f5d42f0bceb5f919ef55d27066c0603b60b377b90b408bb7b12efa17412356f53d14332f0143a4f30a46af;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h38697d8137893dab4e7b74f6a987a510942fb157be15bd89a617a42b675c3ff03dbf9a3745b6e03f397eef70f8b49a685b7f038bfed413bfa08b5083be11539a6aa4cf00d2ddaca0131a57527423c34b53921b84fbc20941b4e90d9e649f6e78bbf83d5dda8a93bc1edc781b102b706da7d9dde0c607648bdd74b3c152a1df93;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed86a4728416fd264bda175e6482a268c19975e2d2ebe052af37543a5f35474ebd76c43e5b30027af7a07a5b47c55a4fea267819ec3a0b177524bb8d25d2231eae450f858a9758929cbb44641e9cbacee86061b3f810d8d2dfd8cc3a227d08083b9b31e66ce78ac1e9abc5f008e720e2d3576d8ea648836fe5f8074ee34d3f8c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h26deb68440af979590fd70371f50e9cc27f32f82e4ca34eb9512d1e5c99efd0e35540751573d45f6e04b3cd58642e81de6b613e857d74c4fc590663af66c21cbcb82a48aa4966bd70bb0ed21ddebbf2210f0b8b733c759cdb87c82c11ce39a715cef7ebc4fa577d83129de860d1a6e732109e8dae73435ea08255551fed818fb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbc787fbfb19b29d9e6916147181d321b1b629583141d791b1c1e80229d0290673245af5c56c866a830c4dce5b44e45df498ac5296befab1fc5825fa052110ceef62e1ad31ca9cddd8ae70668a6dbc12868a0cb0b466588337db548712c4944cac367986223ccdcba48433afd912688e452666547ca60a7ff6d07bd011d8f258a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf3cb06ab7beca10af5401bc494cd32a0e78eed11672089c9e11332c7cea134aa244f65cbf5deacc285059c62261b6b7387cb711e934fe93385c27be2e2444c625ff9b13f643bf5ceaa61ee834c2b9c3f21bf0bc407772179c23c06168ba2c2e906d1e73d38e46897998a1e65c1ff443277bdcfd997e48dba7e24d692127cc304;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdc5c145f0b1820e0367660533bbf5dd4e9ffa0f63208074773901cc4b3af80cfbed32a3392c0b474f07775916cafa84a72c8d7b040615685a7eafbca2edf29e57834a4b9bef6421ec51e073eb5c015e3fa1a0f66186903dcf08b92b30af0be6c7b0f1093fde532f25f08e664f162accd50f0fb306684aff971c261d2e0ef43bc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb127da153f897d0d6ad80d0ac1e63ee776b78cc8339e395c85cad17b5075d007bf6aa8266338f6432a74b6f7eca69a896258b011e508ffba958d8675d66b30e8edd7bedd1d34b644393b8f206bfd2c78cbb2ee60026de2e2c54bb515bf5af09bfcd1610afa3d878bf18b707a83d63f68a64791255d57a5c3401f05ccfa110e47;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba4e930c19640876bfa7dbf49522850526371011ac9d2e6ced3b1d4c8c861e1088f8f4e99058754522aaee9e4d271e5f3b187d4ebb090119a81b0d955d7d2de5fdab09216601b33a4a48ba7cd7f23f082e7672b4bf77929f483b4528a8aa177495f4154f1250f2e4f4a37fe87a376271245d645ac3873a8fbaa6cc3f5f5013d4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h91570dbac88b72c95698c80c6ec5df98508c589cafd3453b39180efaeee6f70ec4d827890c4a834c8e8eaa889eb01fecc5715cfc4bc96bfdc93f7f614d44609a0561a4d574b075a2418fb4b0999084798ea88145a87ff28762248989da58571cba2f134ffe88a9ff464428ab3598a7b16ca40b03a2a5e48deec1b21c72a5090b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha040bce5818df51ab0f7999fedc9f70e0456e3bc46b9861229fcaeef4addc812724d5e2ad35cfc36b17e13d3f6dd6c00e5cacd9882d37c53234c305c194e270853eadc43c8b709e6de3fa3cdf461bd80c9c9332733f59a635b51ae8f5e5ad8b5da1530dba7113ef68b99d8bc73a3c84127c5c6119c046f23d199d98d23a70abb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4e1787a053260c213d4fcf62161dfd7961b180cb5d3cdf3621f17c04d7de93fbc645b77f15909557d68144f68ccd21c199b9ee90ace129a31678bd13a3b3f8f50c39f626be5708394930bec808d8a21008d349dfd7066d458c63164735c8988983938dfe34abda9d5dfc8143b5898bac11952b7919bb350b916fc1d9295d2c0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab8b20dd8cedc79d34060c3a31e1b7381cf72e4f14a913966be07ccb46a6a1f0d742e148342589a912f32aae23653fb309e7c2e493290cfbd1adc2d0225f7138e10e6eca3293503805c596b3e141520a5fae51fac780e54b92cc7e68c47c2362db54fa45d932786dd76764be525b96e9da6a40c9c9c802070bf98424bc94cb9a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13a9672f1412c061908a5df0177970b0e32af1e21abdcd2aaf2cb81f3822a36214472b7eb36d65965e9c5ea65ce40407fa1d69e72e5f3df4f9c1aa370f73211643f53fbd1488ee576867562df1000e57390451976e90ea318e39a2726dcba28f96e3cba4e1de1e013bb32ffca49d746b84f381d61d3e8d943d4dd7a92548aee3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbe5f9a5bfc65148569696c792e6ef159fd9da3127cc9c8d75017386d9e53265d8d055ac82114ceb3a2ead736e36f9c23bc8eba84fdc308f0357c575ede57ce0eb752903f0ec201f44f433de0cb84333cf0c8f3fa088f00874a4e6bf6065ded117027bf23c31347939d26bc5235e72accd0e5c645f85942a4d57e71c357cea66;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h64172a97d90f2bc8b1ea7c4df97c3035b266a5e753f22a679fedf4da5344230cea5b382513f75b2956cbe9c8c8245ce28a5146b7923c3c5622a531c1c4dad1b323b8f79197de26a8189da026d2f5d27fbc960d6aabadafe6fe270be38cb2f72c04e77da2998aef4757c6327b74eb6aed0cfbc55db0876ba03d73d3005f25cb8f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf94244437b5e91e22b63784885d1dd19b334f9c144dc3e7d230c65e64e24a87887de13bd57f05930123ce7237d3fb046e1a1d5994d177394b90f9c0cf36fe108bf7cd930bc4d029304ad91cbb77f43fa8ca8645d3d0a50e1c3e621a6d032d550c6ea5e723c7f2d3d77fbc6488082be7db8b8e1db837a20b424e45cbf6d41f299;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37a1febba7cae45c36764e2d2562a83de4f19c48b068f0ee1ed1eaa500cf3e52b0e5214cb8a9c324119273fd7c891ac5e1c2d2a6a26de2f7cc0ce4eae7264e991fac6d4ffeb4e93ee19c39d29552c4c92b807ab222ea7ad2d987619efb1c9e60467e86d27ccc59d77fa6863e7bf902cb6bb83c1006570d4d085e22bdd18fae7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heebcbf21999376562f7e28c7dac335e6a9e5135cdbbe7f08cb7344c9844efac9d4a8a90caf649c407a7e7fd0f6d206624d7a453ab325e98407d5afac0e774d17702642dcdfc709d526e02cb103af30b6943e5f193e728bd0a584005cca2da54f5d32eaec31ba00065d054dc9668422864b2bc83283917fbc35707a965402e77a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h313ee8a952de935fe4dcdf91b97715b4f7624582525635fc4f3a81a7fc0fcb4d5fa591a2be2756ede904296ed7c532a1096c6027b44cabe4a38112386d20a8de68ac84b95f0f7dd798a4c6c0f1c5bc94e53f09db161ad25c70db39fabc2e29031d151fe79fd4f58e766bd4ea03955749dbc2a1f33d1167e08aba04578ae43150;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h164983c0531e421c2ce23acf8063afc8b124c98767471a51884f4b8c40303377503278a6a411e8b92878de4bf6406cd39904f0f4143d84ce0ed6621667720fced44306389ada047e4c5c8a916ec291f51a372832047c4e339ec64b8f10710ea8834964570bcb16881d4f60efa6355c8a4f1bd9f7a4439102e119b05dd45abeb9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haf6c0078d7538c406741fbf1cffa8d4f8a710ebc19ce655d2bd530dc9aa4fc60575283d28aaaa93bb098dcd0042e889687e4e8137c2f2765eb6aa320efb795958b7d87df98587baef5f619f4702e604429e1a8c2b5ba1458bd65d6a82a61eac266a700c1c2db052637993c9066175d2577fa068eccb5dfbfc7cfc0aacc72dc8f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h47702f1369cbabf5ef2bea17e960025b8bace95a81154724670d84c92eab3282dfdab4dad75382bc81a53b075e173738409c95fc580156f7bf2ab8c42c18fa181b2963dee561c59592e0f76059486078f1d83174724e7f260054d222440d43fb7facf8b0d29ffa73a21a86c9dacdd1758a1bbb850d4ad4166d943bdc754b23e9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc0a4fbf5f529826b608009e90ac4c9960056ccf3f12ca0efbce4cc44588b327e13b66588f7490736e3e42b408f1f4c6e96f3fb2735e47bbe069ff0358a3adf220604f92c98e36daae94e1176eb432d0d8d1fbfaae83d2474e54dffb38dff607b053ac4745b62b78d8f0884bba8c746394698b389e2bae707f178866b718270ae;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h70cb813666fb7030d8304fb48fe73a25cec6fecaf570e1127403c212e3e78122e0202a81a271af50432f20b6ae21e3f6ea280f5339ca732bb4af7e080561ad89cd1ac078c8503f0f14fa44297f27abda5114c3ea3c60094a1bcc450d48f22f17b94633b36cc3c8b03b809d149f97fb45331a76171e4efaf2335d7c0d0d5d3429;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13000ceeef035a30b2b23e19de20d72fc9c5bb2df8a9fb40085c5517948417a90ecbbfa14bcaa7fd6840d57b997bc04cba3541432700ddc0faa217731e01b5db8e2e670fd04cea7ed4a04250e83144a18e1c1f46bd1c137e3b8a05f7d7fef4996c0ab38bb52d85a422d799fdeca590541d2849ab0802b36358c512b92147beff;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c3fd7ba798cc7b87477755346cdbdcb2bb271e0ed01a32be2891d9a75f137d7942bc632d0cef983abb8486b08fed2a6d5659157a59b2f6947689d8de26952a30459d3827d94ed293f86a53518f7da757eb8f1383c33274b10aa23e032e61bb7d5fedfe9ebc4ab90c8348c3f109d041d9dd788634f06f2627ff3fdb522fb8621;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h60677b54539616c5cd56ad64aefa2e5aedb431fba60283449370c82eca88b6f539a8a21a7e2801090c959f2df1b9c5acfa968127b4c2f94728b3d511b4de766a096893785ecc29a03936420b1c6d428e69a58a1ed56f8a5e89504a404241f7dc2a98dc247bbf6a6162342824c7041cce5262c53566bf02a08259359ff6cf0d11;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9907f5c59a8d1d1cb0a07eeb431aa92f7bc02caf2d4cfb37f72f8d34314114ea069e4c41379b4df3a3ffbdcc090fe3b450ebeadfd37740f182cd0add89423fb3520d3ed61cde5ea3cbaafcbe015a38daf437565f30d8dd94f8c12a3800ca95ed47a7575ce310d6db8d17e53811bceb07bc9bc01b96e2325b05d566befddc06fd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9d9dd824c6dcb5ed29c6c868b0c7f9812b53215ef8eef32c4994eb18a2dc3009d8b8dbce8acb56865d3f5617a0995dd977889db1675054dddcd9462cca2047d4bc93fd8662e6234f5aec73bd6d2fe51687213d95bb38b5c73e923c7742fadc8abf4315bd8067a024a01912266a624818ba5525a7c203287d52280a3a808e88d0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc2c102a32388154b476b22e4b0b3a668f5e0ef2ddeffd1c9ba7cd6a397f5ef24e9f6975fbf12566fdb59e2e1ce22a117f2d8c15b67d379daf5a100879d96af9d9afae4aa9485b38ec16c1154bb8b9e1b696fcc123341dff8076c53054cba6e4dd0db95765f165114521608d005766b40bcf4b3e08d72f1c9783e7ee302510ea4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c8350e07de24079e8eed474bc8297a44b943b21deaf82ff2775d3f188ce17fd50be080140712d4a27ca4d6acaf99083b26f11d16512c5e1f3af5f032ed8f8440c517226adc1516ed41806731894f500728f2a458df4688f8df70a51c8c0628e0fb52edf648311f33544c96d3eb448b06cc061ef7846cde63e711dda969051c2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb45ccc9bfcb03042b236d74a8c6608dd46ffadae8a96c81ff52df100a4ee4559e0dcf401ae6781ccb77b2a3dd9dbd582a3c563089379088c49f2caac3b5977cb8de3892dcfa72b680321aa14c04859b66dcb3f096a33904e44bc16f3ad6c2b8480ce3c63af3df9604ceac4006c8b229d6cb6ad6e5c44935bf725db8952f56ae8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5616d821d527a6019acbe44f53b0a6d9840352afadf5bb5c6b7e405ece481258116e44d6300b59fdc593284aed69a66cb5eeeb67ec4c54ec6f8370768a14cc077c450581d55c3d95d6f756c8ca1facdb14711841eb4894ea875d29a7ce570e6b8ee82f900237889de75a095e8749d8136d05ac43789f57e0619d4b1829fe31be;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h128d138714c35f36fa1741c870401ef7eece5364e15e2adf947c894a71574b694a2ebffa660c21f1d0ad7198cd49c70965786212e4eb608a8c25dbb588153b325554afd3dd476eb68656fd0aedfcb783f3077b414bbb423438482a7c9577280bb58358a4a994fa2cba033daf179f6ba3f6cc2a57416291a71809846c397873ba;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haaca15020a45fa13a20fec34ce7907505671ff49c04f5194701b02a45aa3f684d9aebf0728581b3587d5b17b374852f62799a32163f6d1bd50ba6c04ee70541f1fa5ff2651080ae37209bc0fadd94c3910cdf75b588b38f8489ae90455c22246f8237f7868a86e55539a7c5e93f799c7eea2770faab7dab5106b088d701760d2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf3e68aae65d6c36bc2cacf2b9b4e532643bdb6b4e7849271a257a60627c44b2d8443d8488a95460daf6abdb52a56c7e96fc6447b0f24507ed547396576a7a9ec428b621e1c7c01d85dd75582d3a8e8c65a816942db266e405b70ee4785459389de25e56cb233ad44ad015ab85dfd98c72f5a68c604630b7163b2e62d60b00d0a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd1941b8d91377f36cd3a8baba7c90e07934389ac01e232a47b159928a19b1c258391665d2db1bf3b99e80f0de68b890c67f9ffbcb1fcb7ed8604c0fada5bbc41c2ff584e78da8f2873f482fd8797397094ca84afd8cc2f9e83b162035339b2c1424dc3951a7c155cae6c9f49c67011749b1f83a8ba14c5b1e1563baf14a85a4b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3301c2007cfce813b3ddbb6b75ba9fdec9f089c656d412a2fcd69f595f27d6c5c66a1a26fac50578f7105e2c611cd4555af527ebd32cb80ad352992519715b0b63616db7ce281b5db447fd9eec49368059baead4b091277e620b8e840d44484b3a7b437427673ac698756567cfc39bae4f8ae52c03f4aaa3271995849e71729;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h58c63bd1ca357850bfb58ee3fafde8642009865f46a926b8a97505705be8ca66c5107273c433c1a8cc9cc68d9e97d41dba32b70bc0cef64757d4b3d27a5abfbbb9d4d5d7cef5507c44dd55260bce4183c0ed0138133cf92dbe7db5833860ca94515a40cae6655a015961d792312f547918bdcd7b5d9bec3ee6915230ad9f4e8a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd4ef91b5818946afbe64af45d1da095558aecad68d11ffeafebfa94a9369cb0810dc0e7f6e9dd441d16f6686c79970c3942e2cd7455b66a9bd1a39796571a919db8cb2530764ad86d7750f1df2ffc313acf315359cf9913eab5b90945fb7cab64b2fdac30f8185d69e212dd3e4270ec6160468cd146ffe66357d8e40d0acb0f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h804ae4a95ca4a7db77be3af1fbf31d2ebe72606e31a64648293a6e2f6bcb850f6c25cfc62b9900ecb9c8482bc6dd5becbeb760b7ce60e5bfb1810c3417c3d92d71e56b3eb84f85c1de51de01e96c47b704dc227e63cf9f51a80cc7abe3eb6d15a22e9539ca878726d6e59535b75d19bfaec03e51310f263e376c3e10f34ac052;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73dcae24f71c70b4d8efa1d0364b05f3f418cfceb62751a17d5a618bdcdddc0e6b38ae8373ca29cd25ccba0d035e46641cf2b709e5faa0e9f9f62e8d4705a8c9cad47522f5447685f8797a65592ad44d6b06d4a3e1bc8a9d774027f7edd5d8bdeae7aa7ea2b5ed5a7fe778f0bee1348c397123e9525e818af30a2d8b46cfbfcf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8078065bc418cc3e66a9cca93ef3eeb2297fe4210a75616c71b507f2bb8567304f0f01d3d57244698f53f7f1f55b5691dbc7aab2267397d0045bc93163d92ada87080a71c476c0402428da8bf3cadc7ca850b8c86eb2701289b800e969ba1c80632fa1899ba76ff851da4be8f0a8bbb0b150aa21f603d39c2fc072d99b3f7321;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a3253b8515d94cb42ebb7019a277973a7e46c238c4c40ac7f88c2260bba43354375c4673024b8bb877e78632780c01ea58e2117b57c63e780321b70919e829cf34d60b8d75f1e9ed3466d4bf83d1f4b92f13e6c4b8d2f7ccde7ab0f3b9a81d9d066285e0b85331929ce5825a0ad4ba19c498846f9e26f0b101f6254b639851;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4a8149a813f74a79fe9ffda5e96342a197b331a49e9a0c07aad478f9ea2159e25e43adec4a686dd5146732063d062eda3d7b57c8701c02b1a49b44af05ba73062782eb19b4d0e92d41eeec1fec1e2b0c334ad401b3270fafc68d5d5f1f00dc41bac264c8065b19d7e157110105baab4aa318e5309d4686696aed6d142709a98b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2da908a5f79739b16e6919844fa708021f30200858be9813b416958674be98602dd07efa8ad97c997f7628170aa478249b8b1e09911216ec4b1728965bed9fbd2f5811e33c57972a8243fe4a8d687e63aae5bcf820a3c3644a9727b8df334e653c8a5ab536fdb2e62dcb1d404495b4bb0c527ae93cb73763ecef69bc1d19a5e8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9578f024eb50c5bde3c16d00755ae545b2886dc42174e6f86962ffd9dbb4ac20b7a03ee6519d52d8e1a9a02a140e6d0f6bb3e969468d083213504dae3a28e582cbf6dc19983aa4ef16053fddbb94742a9863f8935ed684f127b8af61afec006591819ca6bb34c2dd247328a63dd8c15214d42972d57af9a9d3abb492b6561b09;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97dc23cddccfb3ec6e99212757001191d8ecdf488811ca6a04fa87410300d2f29d5a1cc83322cc9f9ff511cef50746bff4d1d6c57ad5df4dd375701765ef18863c3db5615311592c31f1c218bfdf3f3c119e13860c1e2e0117237eb5da996e93caef5b6457af07b8bcc2de544b10697493e5b5253b4ff95f9800a83ab075c97;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1e53433ff080be6daf6f62c35c084812f92a4a34fee6ca0461b299db273e9be35d10d6111ebd693f4cf424bb65465233c42309a01a993137340d71cae78b23101cb64c3855939dfd6c6ce23d56d4b27726c976290c2a89158956bab55c7a4739f9d2b4cb80868e5d5fb563a112c12c607eceac240aec47220153a2db8a724ff3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdd1ada2431bff140488ee8ab2dd9afd5ddef8f0d672d78f85dd2846d961a1489430bc56855ae445e25289a5635da163e458afdfe5ed64d810deff3add1fc0e67cfced352845fb8ccfb8c7e639f71974cb16ff6765482b9f6212950d85d84e2a9b7c343f00b7fcfe24286edb292021e6fc7826b39fbeb546f3c33895b3643ddde;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc4bec0c7fb5ca070ef3928c0f76fb0ee4211f136302392056d329f5861fc5aceb018b1faa55f4b5abb30beaf3b3802f2769600127008ba03e8b4a14b25dd86789c5ec734c822581fdffed19d6f0a467cc6adf549d51a273f22d3407c7624a22f5838c52652cafe0f724dcd3097b5d39b169f94863db042fb04bbb30487e51c1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'headd36f8c0a73fff781767299cb74841a50d5560236021b1d8f749447684420b58adffcd187108a286aee21a7ec9687067a055acb2e0b9a58895ea489f33132b8a5d7d2b7406fe413351ae2e9920053331e6fa382425e5ea17bb7e2119d55fb48923ffa46a8701b0ea1a1ec82f55379ac824dd7c60942fffd04f2ce4b7dde3a1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha52111423c4e4f0def1b39441a1124de3abb80702c5029ed746f312c7687eb716fdc0cf47c6581186fa20ef0e75ebaddaa8e4fa4e0db4803a44327c50b74649404c2db2e4523f8c9e7b4a1d8027c0562918e68ac5f72d8f92f0c7cf7eac27e1ace6241ffdfa290c6eff96b7a70cf40293aaef388b21c1ad4ad6454505ed5115;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc26c7bf130a9d8cdfcf8b9b1c1c617bfe478a33ab46bdaf1df0966c2514dddac33ad48d7e4e02fc9ef948bd796e9665acb599f79a8a55414a0558fe0476387a59991190e57ef04fb7ffd7f39097503d617f4b5942c84115f7ce44a81850c8fd0db62e6b810ed7c860d84215f076642764bb4e0af41a635586dbe2c876fb5cbd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd5c557af042e2219579b7eb71ad74eba4d484bd1d804a0357ac9fb66cd5046289c1571bfb49770fe4855b85cabef6f4d27ef1c6dc70a4a98e1e3866d8394958aef896c07029f41b36a704ea80469a4c80f4373346b238fb53067be020f164743d4ff4eb9fbd47495cd16e1681b4b06b57883e857bd7d71415cb7cbff68cecd12;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7f8bf74bb5e2cb41926c5079369f83144c7675d4d025519152cc02a3141f3e592e629559f077f151129098552a55bd58391342195e812cea0bf4f6292c10a445cda52069170bec75895c460433f153511ecbc0f7170580b65a60c63eb0f0da39fbf43d089394f6a517e38d9b4fc9ac6b5230c75bffd351403b28e5806556c381;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd03d86a15566efa82e868c379e57696f366817e04852a035ae8731235ca4faa8b81c2430cbf97aa59412310e90333634f96f8f7f2c3a70a7e5c42ee823aacb1cb757b1aa9b0b6d352fabfaa9fa2b4a73171c1df79bd0df33b3f9944e6afd0e26da24b9d5216f62326dd1a364981bc93b7303ed3c3ab1af012a54f238e7841005;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5e7a116ec1ae91730184fade690b1b4361ebe401b0cde676b3707135fe13f9c47a1631032736166abc1c5378e354057f3ab42ad005a687286c178a49dd01eb731f78e986f2fb6d868c654aabd1332c1f0fc4693b3c32805015bb9850d8dfbfa3630c336cf89aa7b217aff7ce0e5d35b718491228612e86e926f49234459fc006;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9889293cf748bb424094e46221f9e30c4a2bf6d1761a32d416725674ae5f1fa87a13c59ce3072f72d9485efe51491a7bf07e603eeb0bc0c8d1a8550698dde3cf224ddb48f75e66965c97a773ab2d032f88856cb4feab2372d1cee9209cb98800bf74bcd4cf7093af3e9e9101977cc9b5a93c713edae97bee49d68e479bbe048f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb3d08128353d9303968f6b413ebc5f8d054db7120349f9e05447388eba8882dc553f295dfbd3eb06bd0a2c623768f7cc0b1dc7625425ad1e17ba9213bfbbd3c54af10decaab2af9c480d2bea63182fe8cb79725723d62a07691c87a9a2144cf6bb7cdb45d70da905a23c7898f5666a5d0e98f3265f553d1b5de9aa84d6566b3e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heef316dbd103aa079cf26c63fc1c8355f55472222c196d09d6bcf8551ab380e049e87211655f97d13b53d1bb05c70a3ab060f14ee15481ac4a9830fafe55e1a94e704b5f41815663531d14bd64eca74b3dff38ff47062ad1764189dc5f00f59ca5f177c8ae1cf5642f8358f4645a560b9be465ad88a302a473cdd8888e080a6c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd67342e9832ecacde06e024e0ca5be5c59f98193cce4427f93b0126cf77c0fd05bdd54ee2d6069d714bfc2c69c867579d12c452c22243f1ad10bcac887a6b5a4c92b853cd2ee9b2e2e177110d601cbdeb696dda0f4220473c9489cd130bf275391c6e2788618124185bd949dbe71e068cbcc89af11d56069b53f2f07193aea6d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h51958b3da4b556eadefb0f26c3f375afd041f00cd66a28df104055af62e23581a9194531507245f918a38d5f8fa00429cbea651918055a4ac2eb4772f8643c17bc7d9792a2c4f6ae8bbbb225ca717e8580f569fddb2f94b7b8c2e1d8cf711454ddfe3090b14c6911c408a195e29f85381bccbd7a0ba35cde66e1cf2b3065b0f4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b385f3efb1597aaea27f4ab55c277be1274ad157ad8d5f882b9aa198e23cf5482824356033620d85fdd5de7a5911ddf3f113d3bec7d9afdf4dcd27563dddce7c06202050e98063b19490b0de571115ed7859f90f15b9fdf5ea7e580828c38baeef78d4fa7bd7048f68e5422e7fd0d2949f245c25de4f4aae736ffc6b52edba5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h45f77b0db349f36fc364b27b08abd3f8cc500278f95e30328d92b5d1803ff67255ecbeb489762566a99ba8aa34f55f240c1f88b71687a5d4cf7953f95a2242dee7c8d5157f6e6e264f880b16da3cda45d9874c673517b99c470c19b25c0f1f836f53a23000f218ac19510579c6c62cb226fecad525d23859226bf4de5131763c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6f6de1bed1ad17f6e00b3bcbfc6975c39c86bb78bd3990e1d0872c36e07db19f52991e6e2d488498a6f2acc4e43738293a18aec9891f16b5dd7353100b2be93c3572239f0276c77480931684042cce3ad77b1e76a4e94db8b3d04996c56bea9d7c2d4fbb30449b3fd738fe15e4bac5754e9fbefe9d0d5c2942d851681db81b2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h325edcff951e1fddccb242ef1729859e4397774e21c843355076e934fc81c135b69d0177f117f120883406654d2fb87983b7f21f21e8fdd5aa20f845407df7e8fe6132d4740a8bebb667721c4b7d5170cd693e6cf30b1ad0f8cab2af4d3ddf2f82e1bbd709059ff2ac02b357fe6f394f26268409819afe596a1eb64a29791e0f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9d2837e58be410ca0b2c522b4b5c268021926836c93762d36159c61031f7c6dd00f9b3ff984112370ba030502ffcd1cbfb2896110117123dd3ae6fe725068918d6fedadf76138660b4cddf5599c2858543dc2353829fbae30bdd976a2f130c54283ca3839e955438338c6ee112a501af9845f237ad4b7276068d1b4551c0171f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb9cc468206eb9a8f6b4b654c35d9c63434c3b84bdd2b3d54e8cdb5db00d0357da45f1ef9738486860424afff4ec3a0eb5865a95168561b06e410a0a8fb149916a352f3838ad0e0655fa1a65f5f8b9eb1a0817179ec8aa88b9b85b0ae2b26a28a75410d1a3e43aed94a68096814b8622946810a0fdd7b806202e94260f1fbb281;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d9e917f6011ce2f7f029991cf89fab027bee9feaf58dcbd8775c8d9af0802e856472bd0a70286bcedd2c5261d6e6fa9dad0b3389b94f1d54b9068681cace6ede42d7d75bcb5aefc0e99bdf928a5b9c9ad1705a2005f3c0e9b03420b8971027b91fbe08ca834e2425e197cb9ba52eabe69d9480e79e535036bda15a5c9feb033;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he343ea6710fd85826b767b500ba3f89690da74f6491c2af7b8cfd9bb609fefd03f20e7ad6b93bb69d844a48f1c2728c153942fa2871159a487707391437df3c96d6e26fd8695353578efbb7a2716e6aef49e33dfb75d7ee54e42fa408637773c2b1f3ce3429974ecb9d1f01c3d5c3dc8470679b9856a15b4a7f149fbf5117ab;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h870fbd8090ad990872e3bbd5fbcc40e231d22526896d6f5950df0850da3a8df8de0cc183ae519a96149dc69310714c76145a365d6aa32078075519b2a5af08eca6fa16b16b31768f7ef62d9dd1b55012ebcd86e7c0cd26f170f6b183b92ee297093d440730d0a4651438fa253ae7755977cdb403d56de3094d8abbe7a908c25;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h370e9a4fd13b127a2a7773b94c2fe69f0720536d56afea71186d06274f6680854bfa7ab29f6d6596d0da05b61961977acc20b69db7f4263bf4b3853418e93d61a1e9f04ba80f13d63776e00a1c9221045d7288cd1e5c67b12c000f3e2c2e829d88b7e79556c42033fe5db80c6f0288af5c0e8574496cd8e71bd0a0f968b9a4a1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8585685cbfcdb1849c81fbbd159e7ff0ad321b3ae9dc1767f3a9af0f0cf3c920c93129bd998f65e5c9657bb49f01b89e99c91ba2f3480704bd79e3bd8995c23d7daeea34425120ae45230c32aaa9fdf8ac54f6a77d6135bda673a2df5d34b1c85c7258d706348dcfcbcb409015660ad9d4c8c3c1bf826e5b1c2968e145a70866;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he848d751d80464fe60cfdb0b33ebc792302a54e801e27799a33d53bdafe441519ad4815b90ec6f3a6e0a1c8fc8e723d4fbad85e6965c6f25cb1d7721cbb96730fb982f50f3eab4c32fd7aebceb59753f2455cb50bd4dbc082fbad8f269459657d76a9736d8986a4230e53f7308363fddddb0b0dadb51b6b853040ccea6faa227;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hff2a8bf231418d025723535b3d08d70b1bd50d7e6f5d8b688014317d00f9e997621c3fc1ec0170fda867ad8240b82787899566bbc91e9d5ffd6221ad7c4302de4e7d568bf2b184cce0b7b20e0c6cce4ce003e0901066b51b3792e1bb582c296419e6ce94aae0b8607dcee759940f58239ded47f23730091574a94180269839ec;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hde6f169e8d3c3b4b58591329bc37cb3b49f09fdf04463b8a1393f263b82b21cdd33bd826f099fb0b493658dd097ccddd5c5e9dd479c23c458dcd62faea193294f5f8327a8d58e7e5606cbd770ef8c98366cc7e1315adf9551d490420043de72c9c23a61458a5e5cd353a2d48dcb5aa84cadff1a4a626413637a953ace320537b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4b73d06f8b17a8a568522fe5bae02e8d0137512353e6d3d25d31478687f60e7c397088c1347c543b511dfd2287e3fae1afbecf48aef80d46ea1217cb4863ec86a3ad16703efe7b477c8c86abed9c5ce990b4610424978ca04067c456d55e90bc87a6c8cf97ec583a66a81442838ab9b95a7349126ee2f9c34060622d9fc0a4d2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h606e0ca699cf23eb5216575006509550548496c4975796fa066830074520356bb118d3304d2f7ff5c33afe3c88b82c095ac20ed16c4d142e810373dba01733d4f2da876036eac37951c1887224d263f38a3c8389267ff94425f5b5c440163b731ae05350c0407d39750b5c66d7ebc2054fed6ed90c32f046f1351653eb48417;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8ba10980efb9f045151ab44a4a2688e426dfbc18ebef8e70270a8a688bfbd55cddc81850f1bcf456f9cbd1a93017fdb5b8f75592b870d6328814458b5779426ddad8e78c43192ae29fb980d45eebab51c5b05bc8342b019887379e149a973201aed483f7671da1ae2ae6bc21078e0c0db2ebd191cd975d33ff50f67f3814b026;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h242808b43748c4bf80ed8d333a314f9f8d64145a7dfd688c858b56ae0dc761d2379171a2bf8e98a27d86d91dcdc5c628ae302541ab6293fbf29fb04421fedd1c2d69e495adc9897b662e7675e81ab8e186ab52233b78545f8ce895273d0dcd84e0b13484af72ec25748cf1cdf06ab53de3cb9dd9ae5f51d4b5373b73ac6c414b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfa954101cdb148ca9354d3f6290ab7b3684e8d0dbf68d407c3731ea401448a47a27a2a6fe7f82a802b9c8c42eca4645d0184501c951785cba9f3cc4796525a41438a0ef7df18d83f873d3a2d26bc954afa8a9272cc525d1c50f39e9fef108b93155c36f0b92cb856e1026b8561f0a8beae869bce25ac04d246e56ed8e4b40f86;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb6b73c107189cb622456f232716f39dcfc7656b8b22af2f708d679bdd64a5ea6d2b00b80fd4a54f8b1afad7b98d0c7ff1f8f472cf96ca530e5bf1bd996e1325b69562f5ec67f4103a6e877e9c42de4e9c361627d145747f4dbac521d6f8bbe3886c8798be8aa90ae404e6c5ccc4637e973a2bca1ceb73df7b2a451d7d80ba22;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5134e3dfbe0ae65c8326b34f3596c0f897e5ed994a4efc4c34259e46c4969df49d3015f4b515083ec656d6eb490990ef92b85c192e3fa9c4e20f034994b59f12bb751fb10b2606c871716e0e37083c8d1fc43218ed3ad89394ee4db1c73a0c00dc58938fc2e3e60b5cbcc11a0e969360f67a46131e9543b4a926b25f20f43393;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbceb0c06caf2d951bbcdd442f2add9ae2655f1ce990bf917c7291cf3134b3c183cbb0b33f1b4d3e477263375a938371c8ab4b76fd8af217d0d1711bdaf351ada39550ee0e66a2e1cc94e11e63fa34815b910d1fb4428a697eda99167190931b2cbf1716cc6112bb4be1dc82dd2398344d385b0efb174280155517730dc8284de;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he5ea47c64b9cc57c7a5c3d0e7aee0354f198a10119e303169d3a84e7161f5ca803a973867f8986dc51f2d4b71dc8bb91b71598d5e8943ddbefe3b497b010abc4c7d5ac92092b6efba8d8cbbd35ca55b1bc565a57f42bb1fde2842d0a46ab49a6720c87d64d562acd9558441591fe2b5e16c890dee4f146e13b42cb38b0bbb7ad;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2c0802ee43139c8863ebff0c291d83b03822820bfaafcc1f7e025da17d50df0b17496eecfe115cbdc8e1c499928dc0ef6f924f4e19349e2dc312987c37fd68fce5e1ec99a46aaa5572111a4962960744dcb29d66d88cfec079159f2f90e0c70b532b2f308e9aa9914601462ca7b26221849204ce49e56d3a1cc8d28a1dbbcdac;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc89afee09ff53dc07286860258a348a39ac6e9f34bb4d34a6b3c1ab83cf3effbafa712bec155d5dfaf4af5312bcff1a23c1aaef9493852a75af37c30d0c1ea1888be210b7a7793aaf3d5605896dc900e4b526d7c84fd23427e25411f9130920d1f09adb64ef073e33e3cbce233c2ee429fe76b3af92f865817d2ad3521ada0c3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97e5694832b49ce9def4382cbcd9c3c63197fa75eb1a9147755a6eb90b9c3244e6aee86f91ef0237963bec3276a83ac151769c7b5a9a47c3b363129ae53211a6498c31ab7606a927dd094f66ae9d2c67d953733618d9ab8f37f240a95d293ba8b7f5354a102fea19f77462f5b574ae36007ec7e9a5f0d0ecdb4648bb527b8d2b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hec3004b33072e4df2c5860dff11b6dcb35c51ca12309737148c2a27683e88be25ff6ec7ae747b7bddf1065cc0ee6a53a22284a1ac6f0ba50831946ad144677cbdfc61753b58bb11d7c01ae822d5f837bb1f5068546437f30490d53d43a904eb4590a1601f59005f93104422be8e867b0db92f814b8d99217716e9318b03edee;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4417a2d721aada3765ef9890edf665c58d9043f13570592cee700f9cd47aa3d607bdbc9a8e80a1ac1c9a2c28580a4d3a039e2c0a4ae9b2e5e08534b25b09907a9c34115e1306e9e33bf5240bc3d6729279da704833317f8e3bca140bc8f50db73c179036fa5050997218317e2e9ce0f0455215db17320061cbe95a521dc530fe;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfa9f58e262a97479b841a4309526aa22e6b8528c76d6b1fc395baa73b781c9c8f9ba99a7466db090324e0c87b7b935673983d9841d2413c32c0881d7cf37af5a0e2bc7f2c4218c4f70b853f3333d9754302d978355dee459345b2920d1ffc4ebe6f20418e6232ccccd1dc0861624f538dda42a35612ba3835c01a44668a8445d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h704656620075429f09f02e3bffe3db8b028c9ac0b9076a56fe3e234f274d32d24dca3e2482b9a381c06dc8c8d959467e03a8195f25c9ae4856f496138472a184752e555ab65f587cee7eda00dfa475a92fd60277850b6b1164ed946ed95fb3ec31802b6a766a87279849a6d6d44ba152e8ada7c6b4137811ad440cdbc7d4da7f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3acffbb0b8212b83571c5c331292fae5692f0eb4e732dcb1da83534543b325914053e2c4d6f56c7c05ecffa3bb572cb4ee9cad66e1ca17498bda5b9e5425db6f1ce5ce16616329bd44fc568cd3a1f5b3263f6164925ec3dd227c3a350803dbad19cc28c944004f3401335bfb4e75a0bb547962522b1bb3528f195dc256a5a596;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb35bea100b6b25b61394e6b3998ab3b66e8f529e1397d988154bcb577ffb91b983f60bcb9c1d934c95b2e6552fe766e9667d0d5bbbe4529d8b37f1bcdd1874174b3a862e21f5cad885f36171ee3af83a5f01b59ff45f5d50c825848010b8d8c2f929f5ec165be108166731a57a663df367289210d4bd1e97b5815ce637bc6e8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he522640e66a5dbc927b9a362d310949ffa91d196832013d7726d47069c92ff15469f736f85d316b070afc04599f49a8d043c18c6e277c4d1a609fbe274cc53f7a54c99d558fd6dc7fbf00d74515ca3cc1ef07bd95d7e2594a0b4473cdaac7414c5883be78119598d3304278d63d0139530bc52ea2d613f81544333b173df244d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h695c496d2d386fbe05a5e91ea3171a49f4f3de721fd70aa31263cece6cf5e21918eb4f03e42e2d1d891b2dc75cde29f6476819e334c5a68b01a44a3f69912e671a6a64e9b12d8dbf939baa9e7ae591f0e4e81fda4ac7ea5c74831db60d1de478af9272587e95429fe6d139ff824e0bf7cf756fe2ea0e37beec02a920b3d15070;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3f65b13344ab1c406720c45718be564550ae8d8d30384d96601c1de6dc6f25e3b0b8490eb7c7e1a56425569c232c187b9cc90dfc552ce858fa419838d89a2959ed105640591ebdbe1ac0900f96f582f40ccc2848fd377b96c7e9d39299520a7b5d48fbc25ce6a8f5e68d4c7251799d272f9697905d7e7e7f9d07aa81653d24d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h75a8eab753b850bf44f505dc7d8c3c51009c900e7bbd7e2b29d85c1763c2ab9665ac6af6ca44091947a3d25eb2e7343c88d8f1c72a9ee5694783be6228a1cd07ce8938ae0113345a36cd0bcc6c4401e4eacf9f75234a25fb5fa0e36ec7d630f07201fc9dd8b79bbccdff45c37f72886ac45380da33cab046549a8ae14b4d201d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb359cf916a5d6e52bbaf6540f440a236519f7ceedf64da1bf0b9d485957f9e6e719add374b858db12b8fb9aaf7ec337b7cc8afa8bb20d184c33877bed73c81cdac8f1dc3c6376081942088a5e8382d1a99e5235a63b0d281656e283b7e6845b44459c8c1a845aa87b89936695a9f320ec76c9dd8a7b9fb7827bfdcb5a4e0e420;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h79efb37ffa913365c847ea86967d31ee77526a501a1422f2d0045551382e95a5cfdf9f7fe26181c58faf005d3068ef924ccf9f65fab05ee9729dbf55315f3b469e3fd0aa6c9335f13b0cc2840f3caa91f4bc66d0fc0ff1fdbced2faff8a9907df36b0f263827c3073e548590d3b1d52e95d5051560007c836c87872c01a7fc1c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h494af60b9cfb30da625e38a2b8cf871eeabe296185a5149822da4813ea49158199ffeeeff9386d26f5a62a7e0e6b91d19cea0e92ad1d2f84885be3a1e03e7dd15737711eb15b3668d71f586d0d86b883ef00e3b04c7f12f802b64c74534d6a54b6f6c5952413b4683d3d9855580216ce8d2922da6a72ba6f515abdf7463e8173;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd04d659c2757f3bbce27c7cb5b9f6e8aa5f989889d0514f00bffdb0e58ed0a7c340535702bf3d915adc48642233241be2ef17b8517028e0d759e0e92c78e702bc60fa5c94ce3037a721f3666a562f0b55220e1b844708a619c3986967c0359b1c7c339f299cbef0525d7b721f4a4e166965c67118127567a8a69fd86bf74cc73;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc53d564f03ff68dc08fefb8722fe8d5095c9fc94ca5769c964abbfd43cf3c490cc4e78af8e29ca03923dd93a454de1160895048e1fdb15101dafc2c9dbda4710e98130daa9c3e42c28a1ffc226431671328f0daa4917d9b7f583e74126dd08ab4c8bd4e40c2a8db88c02ab5208616845228d78bff55dce364271f443601eb581;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8a5fc0d5ee1daf51d4a21aab9eccf69c9aa90f0399c6a8f1900015b31978a8da4023656cbc266af54f9b29e8422965abdd6a55a4e84ecdd6b9f785d433a85fbec4fc245a68a8696c62a0217221e3c14b39f5fd6f5d9ed84422fbbb7a627725b0c3d3903a8cd34771a58152213d95bc5ddf4305651a2c83e55ffb9904e6e3f1e1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he7a1287172d44143a8edefc865d910e584ea1b4b69e32a0623a51459372660487bb504ed790af1a282966b37eb196a857e797156cfc3d34ba463edc131b8f28fafdde582001cbb289aa6a882ebe179a0353fb0886be0f1613b10fc2045202bc8530c21b218292865212a99d7843ecc463ad364f7af52896f13ea45d46e910996;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hec24165f5077855831fa8a44b394d3f26c19f1a213e1acefd29957d5d50e67f520aab2efced361f09729c1d66218174c5c4bd813d444f0fd264399a0d69e5c17026d120af6d54c1ffc84a23e7eb27117be27fbf83675b5993c6afd63f4efa84d12173ebc16a23fbf79bb6a65e589d880be0e0e56f328c640096fba977322a312;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4fc245de7b3859dc658d30915121a558a798d203cb35319387e021fc4bf4db341f50c9720f57996245f62002850a7d5daf7d47838fab1ae1b0ffa3f25741eb93eb5ac302218a6c89bca2cded5d5495b659f8fbf7af2c2f3ce0d76b109d1f34ee66c43eba10b843bf7265eec953287ee4ccbbea6747aae1f1e7c1164b84c955c4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha7cdb14cf4d898f95c4af09fa3b235e62910380ee2e381147f2f3b5f94b0ea83ebd278f28a08a518c6911b276b946219edc2bab5b794c432c2a21e8cecee6051406afdd9c14ee1ac33d4a5829207c2d162a01a330f0593c84e466101ed099f0c1ea0d277c40a6aa943f22214b1b3492d3a86edcc42881c667ff1eecb274556f7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee718b6ad978958649d0c67b74554fe86f58cc822dd8b864da4b06d15353fc3434d6a1bdbf7ba7a9a66d7fcee6b247929c2271217ffbf9fc1f8de89f2f80f48547a8ea54d2784a6c7db53f2ddbdd2899e2783fddfcd789da1555feca9c945a69c0cb1a4bf9ef10bf67a8b349a0a96220b9eda863bea9964c663a2139bdcd099c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb27d59ed74274b4922bb707953c37f2486b7a366b13acf7a8df35cd43eba4d7c23293d6939ec3438fd6e8630e3074a37fcc9efd9750ecdfe4dda2b00a9f57a8029e0783572cd287d5b4ddde056f8d082247b281f76a40da9d9d5464d0cc21aedc02ca69a79c98642d4029f322de234287b31c04a02dcfc2ef04ca78499e0bd31;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9fcb00c1e662d18c2283bfba6ab8d5994fd91e1f5389a79d9916499a86e216c6dd868234f210cf7112d865472fbc9453e5b79527f4fd78eab64d3f4092b607b63d8929678005a11e9fb0019428169f19f6bc760e06ef1eac68e4541e73acd20f929d462b1521e8bbdf448bdff749c86de2f5ab716746a5319b1974c7e8340fb2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h51a7b40dcf11b55e4d8b1701f5be5b815ad17ab6f4af6aaf449472ccf8617fa994fb27906fdb1d3f0e93a2eefd24b6adef711ed8b818d56ece7fb793f67d6c388510b6e3d97b30e92f9ad2f53978b410aff852bb76cc55a0ef4f262740b43d703a9d796c3ce3ab2c5f153056969cb9daf33b7a08ea4aa02e786119245052d714;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf709c6a3a21cb164c265b06ce8f58a997421fff8ceda661f564f84cf05e9dcd6c3bfe8e687fa3878d6ed2ebb117662d875c30bde827c667bbfdbbf8f803b433c064102d0a6c82d247d5f5f118ece8c86a3c91d2469bc79c2dca8abfaca9623ff0dc58706c764fb26029ed5d571e9e74c582c64646eb6f1d3618403585ae57cc1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbaae3133cbd1e6cead12b5520789c9c1f25c9ed5d283c48e518c4abf4edd71e56179f3d6c07e47f5164dd4d39dc5c506fdc4413c159b331133c09252af949e82ab6def9a7b120b153195b41f19a26fd78edc59ef928ba875d98d6f7d081ff229a5c72da9ba6a6f3bfeed3c8b2de570b3b2868a856579c03029da4f59237d9f85;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha08a1dfb61380eb178e06c9cf36fe71247a544f44f77bf2360a3b13bc8a555bda6049bc668c54e9d72b71e0b1f9fd68528b786315d65368f1dde367ddfae2410a4640fc003cefcf1560b8d8a21971508eeae7f4affc79f7e610929998451eb82ba69ac2fd6efd7e6dfd89e03e3c0d3921644c964cccfceca876e3d7a408efdff;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf9880489a1e1c130b967c7419abdf4447c581d827c26edea5a2925c931ba73b2fcc8fb961a5b8bd3c8867c2a32a0fb8f37fde3af95b84aa4777f4509489ed3fe9da1186cc8a2dd6adab73f3000b03e628a4c074481b209d68aa4ddb82d058e40ec03ecedc81494fd102f7baff06651bdebd76456df6b73b449e57191d04e6b2c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha3d7781f325c92a5717c0cfe7c7fd8d22dd3d2c7da94f0f85f71cc5cf31c90ddca56be929e014cea0ba7e9a4ece371450356bc37b720654fac98b72c27eb3946555f72e3a0e65b006cce81368b9d2645b19cc35b67f6528299ced789202af9b74554791a9587b3efc590be68462d1552723d63bf07dba3bed94fa5adf79ae676;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h36b8c735d2f3bd46b77f26105d73f6c06609f1c4c61982b5e9aa4c05473545667c144cbcdd5c1356fceab5ad9235727b470561d34112a7350663b5a70d87ead92b65d7ba3e9cc595803c280b3dc1a0bfd3d82d146e2f24ef2f5dd38f82d7c5f2583a5ad25a7885f2cc67aad5b0301db6eefd4c22160a23abbc7c144ea6bdbbbb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h917c942f0de9ae29feb42c6f508b28c2f62bc9ccc282f03153cb8199baeb6e3f506548a16c0ad763bc16e4155a398a44e9a37de5e60a9f2a720a5eec2d7adb428c486be59e6ff22f899bd837060b674cb3832c18e12b243e85094578bf20d58d48925348c4e2acba5f863b72b5b4245c5c6caa81ec8f6922ff91b765310ef088;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha47b7464a0b6ca556a27fbc575d4138a7e507be42a7d06fbf493b0c634a71c4d4451da5689a05e7af5862a240da0d6ad6b2953a769722a34a2cf7801aa10c6cef8f4dbf83d68e9b995bfbe3c8d92752d701d9b5f1e748b7a3e833fdf82a44b1a888c3b453c9ee222e721de631c4507403734bea82bf3305e5a0a4fcabfb75345;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha5710d734e131b5c738e633d38244fa7089f728cc087201b887f0b7aa2de43e7b27c69b6fbfdae5d24638dae3597aa7c3ac4b97ff4722039412ad68649a8a162dbd8f2161de8ee1a6828f3356cfff53541d031e93a2ea1ef0859479ea762fe0270da08a3a12c4edf72d5cc9e5c3ea9ffd7fb6bf34523961243db293091f46017;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4e7502ecfa54f162fdedb3f4375cf2676b99fe6cf84abf4bc7b28630cb0ebcd32d099bbd801b3035208b572b96bedfc7536c49e54fa644955ca20685e0de53a6adbab9e97aa50760c161161849f472f9dbb31933e8fc9361e8f5d4ed81acfc1fca57bdbb812d2ada779a4a56d4881e8a17f1cc12c6f097d666f5e2a8b54b7c69;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5823973c930529dc30d6e512845848f712eeab08cad2dd8c8dd9acdafe44f207661d1e802cb2bc470a9a6e4039373121ffb74949851c6e970e6851264a227a2bcaf89db04afc78dbc24de479fef3af04bb1d2e78fc063c3e62128dbd3f3304e0d06763fce8c14e4d11602e3891f78bb2f8a41369c0d6d9cb7551cddf7e43791f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2edc35526c5c98fd2b72ceb274c0242dfe0646c3c3aaaf3d2a3676f7502af754d2197641a7e3f6e253b1e83348706b481be1f2976ed091b89ebf6c9adeb09694d885776732ab5affbd0b7b639baac2acba8164448aa0accee9b8c876cadc18de7feb87a9e094f1d1608e5aaab86db7b071acb622bea9b06b0f68f84033cd76bc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5a3f05d297d995b46006035ec69bd70bc14f7aa4ab2ad308ed7ac766a4cf99479619a55b84cf8d82b46f5b670de7601d733454071451b8ab3bf1221bcd570ac07823b06cac2f26dd4bbb14ad2dd559e095d2daaa8e54d806d392c49bf456e1161989373b11c57bf5ef313d72c53b34b15bf3489a2550ba53103cf1ecdda16de8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd32f7f89f44ceb88ff8b5a83b3225447a0945298265ff5b4901c374ae1fa0b1f3f487fb048fa62f0e05b95a497a3db18d928e638d6cc66f57c0a2de2593920ddd41ab3177b293a04fa8f9d96ecfaa695d72435aeff887883245a3aa29345e8035fc3110346e9be068dfbf1e8df521a3792001dc21237b3c5017f4f3e4b8f2167;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfe76182346de915bc1355f271c9d615f8c8ebda2c92775e753396eea0ba64d046860881c16624053c60e736595423992d9f81396c54588842ef1909b7594b9eccef2a71401cad1c13cbd11581f505c92bf6473eb675fcd03743221e19e63b4187713904ac023796df88bc905ac4af21dbd8e5ef2842fce97213ad5cc58de78fd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1e43eb8a4dd621e6a0a7113b8345ae8ef6b2c22a4b7ca9700fd7b2b3e616d4c47a7454ca57b889ddc99ff694c218a172237e1d21fd4c7ddddfe9dac3af4b969067fe75046e6eba6c60c6dd0eb67c83d01755c0fc088e9a3d860552ff92513f18af2d8a94508340baf8c2f5a8f3c77340fb792b43aa6340db7ac4a48802a98c5d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd5a4be71fbbe24620e3890e951378ac998e85a448959833ecf4bc64c27b969bf5dba11483410d39a52c0023b1435d116032ab3fae950d5372074a2674cee8fb9f563ef830ae3fb25c5915fb80992e6e763be69ee7de42a8b2f438eac24dc13095261734d1a19813642d6347106dc8c382b4a953a33150e2cfa666664ba95bdc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd87baa22c02ad8b7224efc8e0b026c1c13ac5779d53b4ee9fc57abda03c02dda9aeeddd2dbcf33737ee487f55193bec7013a376448552bcd99240537062a90618bc465224aaba0ef215162f310deb6701370557b2b66147ec03418ef344e210c18b2ed6373f5e768c9a44f0d109aa2b5d5cb3646ccbbd92d89ea2fc6ac721db1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd8cc1070b7338bcfb9e6d3b57c2b7eab2681dd6f395d1e5997eb126eff98b883b08db4921346cc963d67bac08f5074944ab0cf486fe497208ff188be2d3f2f00d5bb40226da2dc4d560ee34719f2c1f7d7c5d884914045176c2e7ed52bf2626ba6cad493f299ddbafbd27229c07904cc27a13e1add92c6bf700be53064e67683;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h924e9283292d589bcc351cd502dc85541367dec84526bff1bcf2c7e651d2c71bc6994e0cbf4a52723e657654db7ad41523b80e8c0d20113ff50288b2872d460a7163c9248a21af76da68f99538fb80d125c5096ee9dc939846984253e90c74a49e3a52693b7a7f4cf4d3108a4a241acce7951ef147612085d387d72cc7a47a33;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha02ad0f055d98044f7eccd70caab446459e55a9e18fd9e53b7cb5aa68dde721378aba5b2b30bd4fcadb219bf287554dfcb479bc706245357dbc38239632676e5ce71948513dbc387fb46829a1da5e79201ebdecb91b5ebc83b01814a5e8891cf5f0dc5c80986c19dee43a87b84f877c9d5daa6af507a8fa644f778a4ce605260;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc716ecf95968640b33e89ab63164ad9bd5e44f13abecc52f4ab601f86930ab2071791e147ec2bfa68f0f95adf487612686fbae95e188ac2b72f7ef961cad122182c7294352892f250c237df4418c06c2f53ab5fac5012ff8f6f30dc9490d2e87df20c981c60e16bff3c3f63d5df69dcdcad0d312f6e4031dccb0167bf0787b52;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf3b9e54c0d055f3eb57650c877f56f063f986d8bfa738210c4e8c514896a002de317b59d38cf386f328a9efda6d2366279f6b317b168ada85a3b52c57014d432e9171fc3203e8543b55503f4ea1bbfdc1c62085944a637c44865460992c9541ad64b3325d4b095277a79749694477bb201921041312c6666fe3194b6a8035c23;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbdd67354c6acc1472733d1d02e3c15f9a3380f56e3d7a1c99d64352d38da50f33227aabbc150046b4561610418b5ced2ace2ecaa5e0dab9132283d4c2a688bf7fa9fc0cbe88b672f8d1627b992cbbf12145d4695506b2eb2ef8d8ae698657656d56ebeca89962c0c5cccbb9e9412d87d52be76c25d5f6c3ec2601c1665d05377;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h43538a55297c0e8e35bc80064db02c50808bb526aa1344f3f310b4dc121dac28f0dc44b1ab43b42a9def8a42190d6e31c5ca1010915387932f9b1aabbf3640766eb376e7ee35aff183c1db3a086c54573c7d50f1bfd486b8739911d9d91270da59925a6cd30c666e3a1a428153980ed91eae7843a846d8203fe7b30308eb081d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h816e97f6e696e82c2e9bcf336bc38d88dac0520d9c55bb77a040e1c86844d8882903c59a257f7e83dfae71573745da3d5a51fbd8a218a0f2df936fe3a4164356206940ecca2985370015eb03a7a62fe586d80102cc53a436704de7b06faabaea941e921083b0595de6c0814b080bd17e36fead729295acdb3914bc11062db038;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haa65ee33815735eff85dd847ac4a6c052811b24986a42f4c82b5f08592d8b69d2ef075c73dd8a3b23504e9552ebb5a6241b4239e538d372a1a75b212271df59ebff0aa3b9cdd9255e4494957111c2ff4c647c2d642086ee285808fad4d4a999a5b2dbf53a421d2484894a0d3120c779bec5c306e85c6734315714cf13173e039;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc8ae3bfa8e10a9f0f4aedcdc30e58d49cdab19bc403111da0b079cc44ee6f1bc253bab59983260621d01b08ea156a8a7fba44d8e98c33cd6cdccf4aa662bb5e3c0cf49dd429c1c0724c5b1f87f8bf818d1d35d5ade907b645b88cefac2008d4c7260639ee3e660d47c6bf811d1e5b9a40058cd2d450fdad98ed4ab085468d53d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h82782a6dbf1beffb001f4a7629d71b7c4094e07d2a973197c82e72b230795e96b8ed69c90ca556ba330dfa526aef616baf2dc215be3c58cc414716f6c4fd3cbf9a56a5a7429cbe91b0e2f381236839a89c45aa36eb56c44277fca726dc07fead37fca8ae35bc286e57015fb0312e0997f9a85f8c17592e2148c92de28eea20d5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1ca875b9884f3cad41d56fc4d42f15fb08aaeb9051c707932b7d2f1855d6b17a4096726be6c190fe0caec0e9f6e6ed8cc2106b6d5b4dee3bfb8135425cfbc00819844b1b8dc8d93262c1fe687ef3dd6fadb8be77c6cde173e8cf59ed9ec2e087e2565b152e19b04dc84a59e9f628287a64d2eeb4781e54f127e31a9fbfe8767c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h292e835fbca7fe141a7d908bf5677c243a7aef33974d21e9bd36958d0da974337741cc3c345f2c6bc16804a593999e9002afe1dad87fda304e1d47548b92993086546b260a987df07a71c1cd34728292cd110b2f4cf81a14662513716c5b6a398250307a1b0b222bdcf918e6a941bcbe607135fe7460a86fc2fdcb46ab055dc7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hedb7da92e1d277ac079526f76a309b13dfc7bcc3283717e3511969f6ced8e2d8ee5df0427a4b4d1ee35fcbb17ee9977f9412137af20bed4fff724677ad9c1823504b3181d93b2b5334418e9d8c34c56e460d38ed152bec28bce7566ba3840614586858f990bb7f34225c7db56cd5235aca49859865de0ac0c960925188a82d7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha22bcebba2ecd6029fc1f05d1796f80e2f44f6d8a7702056c1b103a18833395c463b6f47a57d87758cfbfc9445fe756bbed5025f94bbbfee61a2c297899949d511c13d5caf2266c35f49de039fe8e2d4ce620296e6ff91888ca54bd4237fb80ee3d7765147f26805c71f365e362576867e143f5e60d1e460f144c363e403743;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h16c51219d557f45087d4ecdc12772cec11e78fe035d88cd427b4156ae8a372defa642609ce882ec96b143781cf2f4c159a35b0a685f110ccd709ee341c3a76f4852f4b16b0c3be7b4cc3fb0c225ec096b8a84ac3e7ab14365e09aced923be2be2ed826f58ad4bc4d8eb0a9fc8942e7f95b27a469aff0f697a62e39db5d324445;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h263d0235981d3d10d333b9a147ba259714d32198b874401c1d3360fad1ea0d463d259d92634feaf6628a457572a15b1f11e9c1e3323909c0738028f677eb01ac0ea9d83bab095d34e62b85815795bfaa2d04ec58f391336c2983457d7f7a7c20057b9d6838259b0038333bdbab11e5a091cd08c7a1eb28babb82134d6538a75d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had8e86b6d15007ae5df66d6334b44d1d991cd5fc0f255b76f159338c20ad3623be9c45773168e4f850d0933d10e583ef08d861e0ce4cca3dc9d431f3fa5630f4eb3673eb1b4df975410a2576014dbf4a47861ff884b17224b3b1f7fed964538e1d51e3ab3dfdaa156a51019bf4f74832282ba52a927478a3f4f61d3a5fa75d39;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd1bf031758c8bb4ff37dd484652833a1c557b70cb06b71e31575932dbbb5014414e85b95e600d1dab2108841f43c5ffc1a9b77940f41223d1108a645cbef6fab230c73b4f442c49e3d4a12968dc95eb795dd6babebba0355ab868118de64ee7d2068b1aa0f21be214eb4032b7979b7478233b7bf9282c0dba3d731535ab3e70b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h23472ff50a861a92bd8fa0fbee7114ceead457cf61e66fad14452c2cf0bfa00374c3c8654833b30a4733db83dd5d3cc0509c4c5205a2f05541fdc1e23fcdd544df584e4122b482c171e0b5fd109cb76ac17704b00e34d89b515d6efda99edaac71a0ee39727f9e016caa012e804c52f9640c54615b2e0a207b14a5aa9bcd4bbf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h554ac4cf7b894298a760eec896715bcef8861ffdd147012c891201147d7ad4762c9fb2cbec9efc321ddd404fa4d65eb564b987ada372c8bc234c796226707498aaef6c414fd3cb068a50c050ced3077d9acf2a34539af296e64275737ed4ccb39e42de18becfbaa4a99c9c4c618ee58b7e1f9acb39248544cbd3f1acafbb6339;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e43d7804301c0fb44bdb507e18d457b4264c0ee8084c9a0d4041f2226a5632d5f2d7605a3987ff5b305f5e3340af5b1c02bbbf76e9ac823b8f9d86d288ce70b572624442145b5926b034cf598f7562eb4eb0bd52cd20fe10a258bff3504c746b5f974cd4bf56979187508638f46f56171bdda2e9ead1c823f96c508f0f24d2b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5135c93eb29345bdb1f22f7f1ad77c2f654fd83cba4ad3d8d4be8a23f15a4e6486e8e870df9a929cc859b5b40bfe5a16d68c71cc802f6005273d231276c256a842579035eddfff9d4a6428417343caea438f0d18e8901aaa100e316adbea10e5adce44093f10f23581d7fc0729d2c9a795fb0984a390c50431bb880b1c03b5e8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h17633e48ef74210e711e8b0860bd995c95972f94278fd3086da900a926145a5f6bc484f53170a0d45d35975749a74e07647a6716a103453da51849ab4ce234916936cb820b7a320edbba79b8bbf800fc2c0fdf00f794a94b1b2edc6312fb599bdea282f155d4f4aeeb045557b1e8fbc52ce3e34852f8f13b9c6f5ea084c62b99;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hff3e179750b4389daf7ff356f4662c9ede8c89dd8ef7e9fdd03a39bbc4fddbff0efbd9ec69b1da6dc4c734ebbf0a8757262583b9a069f70dc7d2fa66b6104bdd8f037f85ee9ec196d8774558f93d1b94804420f6a302f829f61c0fc14e1457ba7adb9f31c0a9001fb71fd0af4721c8039f1cddaea52323e1c7f2bbe99bda672;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7be7a98d47c80b56263a27a326b26325beb34867800bead92bc31adf2d82f3f3a6c1e031d7604b493ad6f570feeb4bd2a80404367d2a1342104afffbf27349a84700022da043f59a62f3533c4d4d5142681a664b1e4b1d6f85066a80c4643102b208d8ddabfdc6d3391cf59238bb5a724553ac1bd4d19394edecade9b5ca12a4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7340329e6bc2aa79f837be5df4d484992d76b4cb39bf8023268520f1a1d72e687f712c7bb92a0ca44c557552d929068cc740a30065fb89b835627a6180f962823f4fa714982ffa005863dc4ff4df7285889278c51f0034abda32b3ecb14df8f3a3038badb93b9f1982e0120d12f43544f174c350b3f4d3e1041bb05153490021;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdec8d9f5ef85672c263fbeb1768879475e6dc4d2fc8666f55d67d93641e3cd516806580bc65a19c5a81f43fda4e2c5094f1b5630c3b094430742fcca99812441bdde43447a74046d537ae8e2542348c2593024ac56c1e5a154e6deb69be6a878a7db3b7d05a8dd914a5509cb26f7c9d40453c594cfa9e413104f5ed4069d3a5c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7991c2e723b18878363c88145295ece29f8f79caed99c9896518889d3a6c97277f6bc347aea4237b332817f77df0b671a0173c292d66a59a9afb731927c69382af73762e8f77fcf2a1c7cc139241ca0f19dd695bef3df5779d14920027fcaf093a23b04013b9f9d7674890dd4c345f69215a3f92eb48a97395e81184289f3580;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hca5c7cbe757d71d6d689850b7341d9cccf0006d9be971873520e31942fdc2854f5f5b8ef94d683974487d6e0b4340c15b24ec30ce26b0df9993530c071db6bb244bd3d36fb9893c2265fa09b1bd67b0c2128979f83f740e2996f51ffd3c5acccacdec47871cb708b4a0122154cf35460ab84ffb19f1360ca00472c60ac3d7d6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd59faf51fb5baff036e41543493b411a87b1eb81c68bfc75698c20638e6149e37360fd6fdae0bc48bc24d504000e41174723e6eb6d9158f0caf0a90424f5e2c880fee3d9f9a90c1f462501d9c624a373b826bac408829bf228d24076570e680c6a0f37db329bd38531e8a93fa99c9086b2646d33082af7187220e343cd3b099d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf204098b6a0faf0eb0672d7da9bb162ce08ad43ddc983e7801368265bf9d3112bd5b0815069057fad58af03dfba081df100d4086635b0cc1db80d00d96cbe13dd712f4e24c27d2b9714ad1e7536d997a0a981263443044c35438eea7f9380ddd2384f661045d92a9480be5a716bb1c37718757e4b82cbfcc67a17401e386c9f4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd81e44055a62067494678150cdae1b8ac3d7a1451f8976c50aa17b779815066bf99c1b58b5fa0e44c751f55218ff11dd7dc9860e63ef4ccb71ffce72f957f9b48bc3c7ecd515eb4ea4c14e034a4789770df7ad6190289142da413700fe4e4664f670174b7625eee037853c4925df79df7a893f0cb5343371588fa5d93fe79ae;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h78d9fbd31d0ca68dc0389bfd43075d2df86ca90a7d17009676e6a0e55240c48c3251dce0adad58f2f51072c223757727e925d6908bc34f929bb86a304d3926224771d1fe0ca65332272c5917ea26af267aea94cdb3cde52ddc29d513d217fa126694af3e3bbdd4d0393851ddc952731abe336bde1bd16f2db4a6efc3970fba98;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b709ba83d89c8775429ad7ae35c5a1e706987ec7fed8873be26f03bf77a6e5db76dfd5817810356a98da189ec75f6aaa3b0791c5f35d4b30393adc3917fc89e1e411cbd4160134ec07f588a7fe45d208a1dd67745a4ad5bf40321fd5e75aeb663c9d332546d622fc09cf1467416cccde24c9b787bdca6f061710357b9a99808;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd6f029b059258ea4cec6655daa863bc3c595ed7305b8f1f2f53978c90257a50b665800801e0156c6b1b3b8267ad01596001eb12d0701f1862f77e4526bc8a4fbb33a7fed1bb955b2162c4b65675423c61256dc33007b2b67e3eb5fac8715d08f05f95f8bd7bc3209147c93c5022277b0ad3ad6464dbe1a9aec90ff3d7dfcbe8f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h36e2b0b8bf27cadcc734adcce4ceb2e65b6433d03d205469a48891e01ff21f252ce27b823cde03e16874e083cda3573ab40c97ecd650cfd44d659c597caff377cede5c3bddfb6a47f877a9e6b93e45c2e82955cd8e25d5f499c97ce0c51df711d07b7aaa17644f67e7ff373a2ebd089a0b8d21d3dd4f1715af20f8f27d183a68;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h51aff3b935028a1f9fde1c038bd35cb23ddcd15aa45eb8daeb6297267c2e9f046029084fcc82cc443f2eaeba90fe00b41b7b3da460895b52cc9b1c7e5b2189bd79a771a699b20caf5aab6c2ebab3bf7051b9d37c9069271f8ea04c8c395969761b1f7226875d23554f0d0f7106b4a1c1ad1772ba4e4f5b7082708f010bc4a9c4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h11aa46f1a9d722ec1a771c6a2522fcfdf914b52ea52dfb0ae48283b92990862474aea68258f84305bbffedab20b1a93c7e6a5fd531ba065cd6e6e4e90df229aa60d5c162eff370b9ee6d74bddcf591eace221a71375347e7bbd44414598081bbbe78d66061abdad952bd97f4bac0eac02e1935d039160dc6c3b8905607eb869a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb82c05965df8ecfe1daf4e088ad28b5feca4eee11923650e1b10d517189dd4c91c43656030ec29b3c2f69ebaee1399da778af259c8b073ec2f2a3df0ae61087a465f703f1d2cba6113ede25c1a6eddf610ec17e67d6436c8624444810a412eb06ec8c76df7dd52436c7681351abd7018b79142ce65d083a5175a336544df35c1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha0c0df6e744de0fb7e5e8dbca1db6c8bb41b02b15c3a25e5d5a2d3fdbdf6b01671200f8649654cb891d6714e6a27bdd682c0cb6f88d132c59fe1b710abe21330a0763c9373b4f159f062915eaffbf9f4724eae70e025463bba3068db961ff5f78c7a4f193b4c2f0171f31af7edf6a99a7695d9a288fd5f1ef5bab4c0456a40b3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c2624c28ca512fd8dd2dbe672ea044ab8b2bb8808f5360342570382cbd8df93cb3c55da5202e6d82840f1aa32bdd92542a3b0d04e0250a88dff53c28ef3509ee63a6ccec55190613693bddc7396766416e8b1abc8af37068efb967a8b43f305ecf312f3243122e62b831a34c96f7740cf7e286a0465f07720b8c2def4f3c3bd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f0c1b728797455f8ff34257aa4c33068055b848fa5b3c6cac3ae0a933cbbe0972d62af0a28e755b8fafe2abf3946003908dd5173b90c77e82029021b2c9960ebbc59f39976652f15e3cb363b7f27b0148507f116f957c75ee7d8a0fe509dd08d04ec513207986831c147e9b41dc6b26dba53c47fcc411ce92e26613b90b1ec1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35766bc433e9f8d54dc0e91d6ef5ee46ac6872292341ed6df1f062d69e3962a7aa7e8aa0e53b3a3fdbdcb252b94d3f6b3a357791996201dfe0124181b2bd38147c1fd2a1cb655d953aa23006f1c25c91002b0cba0d66dfb75cbf11eee469c2d55f5bbc23741e3f2d23f62dc32bb6843a4a3f3579aba413d6ead050277eb68f87;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b53bfff2d705983bcb4d2aa932020590c49af1d3c11f68e0700f7b5e47845c33397d6326cfcb07b82ea265a84554f2305e43c93da1c4815cc86c20a1b32bae56d66f7f72c89a52816c9bd5099e6a361e6ccd57dee4ed7228bc230e8f1eb7a546f17892c07c812a21d6b29d3a189b232b0ddda540aced1bfd9d5f6ec710c7979;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2c4f32e833cd3c29df1fec96e8ffa4a821a7dc90c9b2d6d768884d9dfd54a7c45a2be652abd962b973478513fd94d3d99f0e27eb8fb138638cc3ed1e452bc2f80949d7ce7b7bdedfe0ab188611bd6a6ef8e61de79d04873cdb731f63dca4b06c46bdd22d3f27c59c29ebe349403019646b01ad0bad8f17f05fa22a7a8b603332;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h198a1472b0175bf94875dc7c091ba6e63322484133a270458052e1aa46beb773dfcfa4cdfdabae5a1e9dc0de5e328ebdc8036ccf585a1ab1e1d8d9f1d4a29432cb122efab9212db2394921043ac081541e69c2203dd4f0b29d60c20c49ab4cc465ceb1731399dbbd2160dbb22b888d4a212ba1de566bf7a9f9ae60d7fedeb3ef;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he6fa991aa71892dce498e74d5fac6ca3ff0e13c697877de57f7e444a006d356af0d402f7b6e115c0658bbe5f73298f7662f2819a340d9a14bb350403e29c008c52b57eeec2f1f17310e82a456c3e68f5a3f8de2db24e3d16a0440adf22d36cadeedb03307daa5bb1c878abf08e10ad676ff0e7597762ffad0c70d2e4e3bdd3f0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcbfbed030284b41dea23eeff18b12ba987309cc6d8fd1d32f37a03cda5ce3c1d0a97e865debd2a38e2b18fcaef0476c5c11addc51dd668f82a422d44deab85b69a2ac86f3af8bf384d62007187a18cc60ed032cd5df4537093c4ecd7348401ad6b47ea91207c14eb0bf0c3c9e75e301e4e1c6387b9cf2a44d4a665c354aa5f72;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ee91108450752ce28ee64888e88d0c4058b3149a45b0a2440adae7ad27be226b8d30eebddb54467566e5b2eeb53cb2f6fc9618c7678ed1df80bafe1e43f2a4aa781f12ce52219633a8a3c50cfd5dc6dfa6884880e7b459f131b649555bc58d2fee8bad1d24fa822aa9acc0b3b5657ba9a613c9ff115651c23137179aafb7513;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h962b0694eabb1a5252d8e6e49c675984c75b1363e8738f67fbe2eedb24043076d55c0657e78c2345f7c1b0c12f5325acd37a5c18e37e6e8c3ad13d91ecdf662c024c8d7801d6e1312f4a297ab3ac7275911ff756fbe3f5ca0a4c246f39b69fc37c00c309fe6cb95c57dc6400ce1a01f167963ad25b15fcaa7f40fba9468b1969;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d44a37d0060774969adf6c7d62476cbfff9656535fbccf3a1274010a9445627997cfcc6861b51591e99946e67445513bdb81fdfcaba75834956c18fa2a5c00433ceae82a2828f92d14736f0bcfa03966fb6ba55f49408a1155a06954ef72ced4c64f38134511805d8fcdc04da12f0884f7da6336ded80163df8c3826500d48d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h46a28abcab4ebd2522db0fbd9d2f48e843913037e6149f81f6ece1b4c1251c8587e4233d422b854aaa3c97d961d967fa0fa9f5592fc13064c88fc77ebee4c729d4eeecbd00f81394b6d21cf2a072d90a3068c26ec08ecb4a66a428c3a6f52e53f125a0f5bc10024252b01d70c9db998bb7de67fa042bd1e12b4c7959256a4ae7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4e0906a15e277ac8e642f672205987e595f936b2f07d4faccadcd4e36f568ab4a94235ec3fe48acd839368f32e5de6412f40729c50a6d16b6e8abc982de22153d538c9bf51e52ecc84e3ec4ffc8477fdc2592704986ae6e9a6846495df75e8e73896e1ced2e04dbb9ed2f0a93559dbd6f13ef36e0fb15e32cfc379836ca0451e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7941d6729ee68c7db84e007ea7365b2a7cc5e13b91a5da38b0bbc7ede5f38564c35f21f8842a33c66a209601af7db735d248f6d6083fce48573722ea0b02ad4acce5911ba111aa32ba3010ab1027e56b91a4c9fbb15acae9f6f7db778a1cf819e6f8ab00297bfa5cb49781c16b9a16c795d642533fd18d28d09420835308a141;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcb114df47368aaec693ebd97eb97f07e2482a7076fd7f0c76d74f6ed462090afcf4d94f30d33832fee4ddeca1ba52a45c906c29cd4649ec42263350430237a2d3379bf29a6e3e21b026813fb39448db0074bb0ebb83e0a0914cffabd6ffdd2da0cbe9df5ce9abd4143da8636cf17715f80cf26cd35db007df01ce3cdebe48eb2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97a85096fa7b92e577cf824c572f6cf15bc03f5ace8e0642b7b8285716cb68da94f4cea2cfe6b4728a185089d79c9f558225e72d658d92e13b0531a458dfdb70fe612a63dc997a34bf13bc735e14231b66ff7b4275dd379e21fb58ecb35e979f801c8a8faa7dd2b0293556b4ed841bc939a9afbf5a86ddd4376509dfd5deca2e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h23d8ec3a8e942f9b3359c913fba6a5fd95b3eda126eb22b4bc0ec9b4b42c82188ce8ddb7fb9f097cb3f656b649ca9575e5eb5c32ac906917a5f5e909ff35a3889bcbf1da474ef572cd3650d5a1f4b386ccd9bdcaa17f8b5d518e6bb12a02956633331686fe55de899df05702077aa10da62cc9b6df17560809d56fd2598b8469;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcecb6f1551a822a598fe64977dfd20c274f42cdb7d765c584d6a4b5a4ef133db35c22e88f5d080ad880147494eaae230ad079a6f0696ffc237ccdd7eb5c09dcd6f25c57d35d6c4605e1128a53e2b6de8d98073f66d1644c51ccf0c229f8a4e01f69387cb072302c40e22fd55720336bc38ceaf292a0331e556870e905aa2c1e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h62d726632884f8b2ea971a8b638d100b53dc3ca262e4ccd7261aeadfe707b0970a3f409d365bd80643b68bae7923e36a0df098a9c37db74e656ba28ee52eb4ba18874e0c90d091b3259a89ebb940270bbb2e84e2bcdacbe97c48fe84ee563954df343c5f3f8f2d8dd6cf09d37cf36fe20a12ea2fca2ff1d3a8bdfbd3693a2b6c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7a75e88004d75b9d422b83447f751fd0862d56737ba29d564f11f83d5f6e0bb1bda671b4e8ff64ee774b2feb0d02f28b1d621f4608e15a6cb7e1c1bb8ff08cb7366a8bfa558c1b18d9fb0720765cb2ed88fcdf2a4657e2cb6730a6b05bce8a998dfadce5d0d30704c7127295dfabfb24f7a29040a3c15aa232cc0f232c31806b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc04d20b737b4d7e52864730253201be935ac362863ae120f573b1fc1403cf9fdf6215d6c06be5dc1901769d4cb1919f0342eaa26b033be81b90b363885208c08dcf038eb0c498f2dd1d11f0ace284d9de1b9f78b2470c2e2b0791c89a227a995e6df5a8683f915bde6df63155b1dc7ff8a32e443d84060c13c3bceb9dc676294;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h60aa6d444dac07271d9cae842fef12439c1e7e6f7dd0d253f4b79f1c8b530f682ad98bfff20baa5c0ae2af7d4cf074debf125dd90bf70121e1646e94c8bbb6d5517cd01187e10328d8fa6b18d93df994b64466c8b15dae9088de26a1f4a8def7e473ea42831e492cba5943c9c6533ef180285edc9f450521f3f467e8ee96a666;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9ef7b65fd9abc62fb1532f6483900f95992ebe8fa04371f087cea89f6b353c3f889f83dca20ad85441e2235a00ec32acc12565aa59055eda01c5cdbed7277b159b46ca1ae20fb18ec302a37ce044dc92f3fe9c645bbad0d4546b15048c3c95aee7d9a2371017df6bf46d2400314b9beee982873fd01355672d5d22e0b7d904b2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3721a0bb10a9af373f80f68c31a49b4fc6846eaa8c8825d8ebab639cafde89726a66a3fe22ad6d949344a420c5e780461ebf7970d48a6352e4af90c448a4814e172c0edf89aaf1c56c7dba1f4145edef08f7aa463c7985c6b076844290b2662d8b0b9abe4a8c87d181b38fab129440fefa2bcecec8a959d93a8b254bb7a3391c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha2cb5ce63f4eafc87baae2a71837d297bb02f4c4251ab544bc66ccc97e7fe2644a19fd713eb897688031e7615d7feee893dcd616fa0363ddedd5e859a80a319ac4920401e5e7f171dbb2759c020127accf1fb4950da689aa6fac01bf235ed2aaf3eb6bd07a7a389af2caeb683f4642236dc65bdf280f823d13cedaeac92558e7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he735359942ea58acecad0db87d325a184c5f22c9172bfb0ee71f4f7d893349b92127a6cc1c51fae1f08c1093c9df3c7a3a7a7fc96863b97d63a17e201c8164e11d173259051af7f5f8160465d45e5a267efa871f5b7dd2531b42ba392a650519e68c0fb8b45d318ba93f02cda8f7b08b6a75b1acc0b70429d3e6dc7dc94d73b4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h24f1311af8dfb0c6a7a4c6655e049abf3371ba5b3c8e5e6e3b894901291d970ac8b3130dd159220f15a61dcf8605176728a0b0fc005d93b60b7ae2666b9118447832dcbd82ac40e056a227ec07fd6375e9a79663db0cc2f925e1dc45b90d8e0e8c8e98f4121657d84cefb99d8033c2fb47c59d64cfafa433c2e7d0a09cdcf99f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6408f7c48cc2a51871798e8ecccf39749a8ee978a5fc3141665aa3591b7d43307c5c60bcb4fb374ba59ce998fa7fd3b2612c51992da1972e68a1996840794c9334d01276e571d62b5d29aaaabf44beeb6820b746312d6b8eeb2b86c9baeefb0e6455afeadc740c09ffb31c1ae15df3f20f599a229d6f582da1f967412cfbdc2d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h26846bfe6f0e68c1eb306eade79be63f5a14e6f6e0042aaa61bf4de20bc5681d0c40110cca87e463e40dd225e37a15aa8f2f892886b71bd0a6f9bf46bd48622bfa5865a2923b2256bd42b2c219ca6ce1e981048c0820d73cdeafe2a69c1f7b1b583ba1f035c752ad6552a1d5f09e2c62ddfeedd56c954dcfcddd7520735e5149;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha299bf6348c7824fe5bb519e518fdd1e158d9f1db17f642f54166fd28f08125a3907bacce367cb9cb4184eac63ceabf17e6515d59bee8315ad7cd214e2d2590264e4ffef04eaccdd7540b3d2633c802dc11b3b598872b9643a38c03cd63a8c046d5e05cab0f7e8bf6331380eb5ee01d32b98322d9abef46f73d5f54ab40b57f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hedbde7cafcc50c8d130db98148c1c0680d09678934acf8fea45bda336a1597e111dc7882a055d0518678d3e0a22d8e6e0c595eb886f7fb9cfd1240c37f8041db20a5128f162f18d28f4c7e3f392761093cf2340146a4d5049df3d3c8b87ebee2c783ee08e85764dff98cd0b71c4da2699836307f9bf24a8d43b2fea588badd72;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h58756ca6de272f4760ff6dbe0cbefcf53953580f8f1b0bd73b69debc11f6b2e89501760af3e5b306141b938d5ce270c911cc02c7d075c039177d2450e8b72b7562e7e93838371b81db42a3471a51ba6c430d9f973ee2dabea548a10fcf307d4b8c217121d2d77d17f998863c9f954be0308e711a2c6b1f2d848a78f650d8ebae;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7c91c403702754cec2fea53288265c5c4605bb7b87585e466eda7e90bfa4fdf9e003e6e73fcb40594598732427608d0eb52390926a13d848e11383915b70979cfa275f8316e2c3fe790ab5a15be7d080eeece466ef4f8019ef9c50d1b21959fe2f49bccebab57391cc24e67b66f0e5cf8202da5eb4c4e9e581bd50d1db21d1fb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h43b44f7e6a1bddc23195e26c67bd8a0dbef7adcaef5ea1dc2a95cf2190aafed443fe95510556647f4b3fabea11c8ee888f8ba4354235b36df3cf2ca81103d0f23ef0ff1402b477b957a6b40e595a53312729cb9a2e89c8babb28ed1ee661238c496e1c0e58a1219fda6d140919a980c0251750a8b8feed1b5979677498eb94e0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h85a2ef050cdfd890af4273833072d7db14729a399ee3697c2cd170c3053065782d48e3f03d977e4bf6afec9754752d7fb1ed7b48f2e7e00e86b89788791ea15224fa394e46973587c82e747132b35397986e18bd1b8fb8baf0fbe9a2392a7f58790be1bf9b8eb3ddb85b1cb950171dbc24adb49bfe5610e1b358fc314df262b2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a191c8f88aee543d89601ff761da30f0411722c3577dbeccf17931e89f2740e492714777bb4ae3d8699929c7c987a69ae1cb55ed84359ecc883a38690d2fb9d1c9c8def6cd503f16c1e89346a1746b9875cf11f44571f9e23968b355149c344aac8a6f8d350b57e245a48bbdc45d4492b47b3f280d9a28433b4059cc58a6790;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8915c94866e2faa2662361e4ca60b3df300a4b54b9f5159f3c6ef1d9e1934d811cf19ef7204290d2fa008d76f9eac8275775ca0b2d095d670ff1f3ea71c7cb7eb28850d71a7c8dd8ebcae5f54fc6137a554c351064c91a55c81e4672ddd45028dd13444b3594cc729f1a2ad1ea8ee80ff9fca0f505d0709984d136d623d5747f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h143db104725fd9a42ecaea96b63c3cc177eaa575e6be72ffa5b112b3b0822fef3b2e7ac857533a53d0a963e631880f8fcb980ea3b48fe76779518adc9157bd8c54210340449aefb4cb38e39d5ddb7e26bb2c0240d45ded044bcabae078a6b8be55d1064c3700c54e2d04080f0d05e4ee9be037badb543d3a1b310b8368668412;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf7fb3d26729eb32a4e67d12293f2908b1e1d00b8c92e11cbfb5f027c125681fb9dc589d73611df4f377458f7eadb718e5d3d12b2f82f36aa618bc0fb3c64d5a20fd2a0b686fd4ff47ac8d630b3e3a936547506d1de594e35b1c4c0f038495210bcf84124441f24275ec2a47b19a2b3aff6da8946825e29bef6cb3779572b1cd7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha7cc67d212da8f7dcce77e5d0a400929810f4b35d7f8c59f620f7ee04a5f7a26dd98f4a52426633e658a98e77e2b79d93b0ed14f3777b2130275a4fcde3dcaec7c3c2b9ef645f61f2dd0f06f305f08675a321e051d433102154069d5ff6c3bbd0b3d7565f4d2a9cb485383242cc2e6234a5f7285ab370e47020aa991f146ba15;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he7485c98895828a6b5a662bcc9caa4dbb761ab9023282570fc9e5245845fe6ba2cd942d017384b3abd4ea514b69aa5adcf22f5cc6112236e32aceea6ec66f32386c5c69c9ad6fa82e0f127d1da0fecf9ab4dc7f446616043a306b9044aee65a03eefb752024abeb97988ada344de1038ddb7d0e8ff5914406ed622ce10de2575;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he1bbfdcc61ffcbd831fbd74fb5209dfdfcb9ab7b3ee26facedd614769db605c793e7ceef3917351e0a9a5a4ad170d6bc62c601333efa3cb24d14c071b52dbb4af9fd0bc651216a7bbc6f1b7513e8944d5972fedeb407242f4f21cf07c70fe03456b11bfd147a35724596078d7209791f2ab031da80fbbc33b2c2de650f061b31;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5cbed0a98d15941ee306d0019a3e1bcec002dc1041f3a2063b35839459e9d043e5516adf3c9fc62d7fa649b27c70add5bfc8be7001041239283bc364e3d29dbdf7890421d23df29ddc7ebb834a2765f57aa84b5e6c75e5fbc90f24ebef9da1fdc9e22c0d938ee0b739d9af3ff77922442eebe7ce149aeb3577db04fe0980af63;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3800d84dd3a528cedf77fb72b1085a41995720bb2e36e6072f889f548ebc589ee077a6bbbc3db2244a2e2a68d1b467c8b4a678727e23f52d356d30c2a6668f14715794d254c3c008f4f15e77a3fc46189eb382de03b664310b572a19ceaaad07bee47b010c2a8d752ae877d65b638b74ccc4ba605017ef79e3c83395ae7f1b19;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4128ed887af7863a55956605c8b984831873dd1682ec98e934469580bbd3dc6571e766cafbe2abcef6420679c4c5a6632dff69cec5dcd0df766a220f56a70116b0227c27498755f215975b8558bccd8504b5b6546699bb1b3ceb19e41a63879164e50136a011fc5368004a6628d9f527385051de10776c2dddc2317867c52662;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19d45c999dcbcd0bf99fd8e84488c93735d772e88e175923255b90d8a0f9f457fbaf7e3a35c62d4a8c700ac306d15c5eeb262c84d1641eb0fc25b2459a2dbe881e8ade4480b5776e82beca1a3672dbc103ba5e2d21754e8cb7af41ac7cb06f6c20009eefb101fb011df3f51df204f538684d1899d7be9a535ccbe34bd6b4ea80;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h32d2f335f387836e043e1687d09441aca5177a052f075cdefe13a73bc3773cff64da830dc7e4b3bb8f573424cd9916edc16bfff419fb66dcca6c95f2c720cd6f92a2fa08fb1e7ba4d929d7e23dd820787bc224495fef30c332e75b2fd7bb975e035675c0e2403e058212e41fe37ae42a62350bf6c4b6257b1783c7e2fe20b50d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf476f1ed3ef637cd138b1bcb0140db805ee3988a557b84382b2ead2300b06d62a857a3c4a082c24ad67b3226b214df422e3b86b742637f9cdd1c7101357c52eafbeaced54f6d04aca4534c36749e2fa73403f3230d51db35fe41fadc43a3a942b577963425906f6f4e4468d8e0b674e9339b943f3c10744cfdcefaf2568f3b43;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf3e9d5898c39591a39789b7955643cfa46325b10fe71e2b21f67b91a4493ffb1776447d53322b5079f96bcc4b20f64eda94cb7e300bcee10e33fe0dab246b8812cb7f3aac561ef7f29b0c3e887583885dde539680c21803b0dd829bf0277401cab5ea1eeb81333b85d35e544c4ce9df29e406c4b3ad3e714c35e61277efa3d99;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h400d8abf10ec74e4a1ec1fe68c280e12ae6c4fd0953970a3db2854ba8a79fb9025c7ed0ffc0aefb3298a863fab9c19ebaabb9f824e40e5ac9b8d5e407b5d28bfbab6a433b1aadc8fc121412c8d18a095c191f434d70024222739e43686deda3b7b09ab215fb731d4c99304d3e9123698b9be68922273872c15b66b19da7604a3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdaddb40b09e5c293e3ba99cd4926412a5e156c198bfbf6bf5970ae96dcb27aa1a6eca0e47e99f49d9b243a590c9111b5f9c7bf9a6439e91e28b0ac3eefa3acea591bf97d24bfe67720f4cb7486b9168652a97e53be7eae7af8088d96faf828ca7751a9ed2582e8655443c9fecc18d5e1ed8a443f44d8d5a14288624bf0081181;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he98890e4dab7b595702de863547c843df98b3c5533561d7ee5c7f264921bb85a1bd5a466ac916c7f6f606dd441d882537d340796b25ec0868bef3ea9c1b396160e2b4c63421762589a992cbd0811acf4d72e6b39d36ef443908f0ee9fea8866df8a14e005836f5afc73c55bcbf76dc3a4b50ac05000647e545a028887a1e979;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4a2b89eca58f4f55fa425977c07439a656b48760a14dbfc7454fc41d8ba45aff49c93d0ccf01a00e1b74584e5df05444a7336c23be005f65b5c0bb9d208d6efb7cabed25c9576127aed7bec87e5c796d9fc499a032d9f748159a835a950588f388ee50b3858027428b3618f54131421739cd7eb47dd26bcc05bfa104c9070426;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9a30c02e3929a903afed0e47f35b81b43f56b5892d88fbeaebbde950b2b6b8a9cf628f61051e5241e491944f72a18b53af44da6b1563c35698f6b81927895b6d3bbb4dca135d04c49f0167172321fd6148aa6fbac37473ced932915a71a91b76bc9aa05133baef90d51796f2f99d3b8374895e572b430d63fd9996e0330b2fbd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb05ff160d431c6cb4ab1bcc97f213104124a36b8b3633e58c807198c234387bcb332626548ad60438a612d4e8a2c073c01919c4b536d79294543e1b99b1f23c3180e2dc9bc4ec721cf93d57485b01e5b9269a80e0453d82559aead70ac2ec4d9d3bb10e5f75dd130e237e5dc8911e52fa756d93066b1a112a1d768d883e2aed6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1100e5c9ba8cd7ecd7b30a0048d86b091b038a1db65d20feb8606e8b767b9cebf0deeaae58e38ad083d5d03763587d1a40e128fecf120aadc4af680f2d0853b3ce13da3e3ed7e771782ae292d2152418ae541030638810b322955c9c89ad10160c501b58d63768762d8806198679972e2cefc78cd378df79f81ad35b89c58a17;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h95cc8bc9f07d1979346f2f392a7c2c28de6bd7e7dc3f08028f3d5c9b91014f352ce047be62fe74ccaea5625965ca5a8e30fdc25cbde2e6d29c84597e521c6ec4be86549b8687874d5b20ebe4dfa13f192c0b71a3c026c19b64210e25e196de6e1756884174263263f28559353b127e59db6c283f7f5b2976594388b4de685d5e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6d9a55002a7e6c885376246cbf7c24da30ec02fbe0a3dbb632b36df8e7569f357203c748a780f074649d579941d4da4e6ce0eca9a81b3e7d0d93b433b804ced0d7551a5c445160d9b3be808177a0ced752a64bbcbd36f47fa4d55ca94f28aa3fbb2cc2b4fc35fd6b7a7e0585f2a9645e1e0c9cdf4f263c4c7ce0d6dfc3c23b7c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h84d5392de2a070afe7878bd5c64f69f765754304975b5fd5485c877731174cb4f5e0553b6ea518eec9a69f29ab6d51f03daa943c493ebd5cfb2b21769c6d671f26a6a369d19849b7186ed219ede9b1639825c175c8d26f6e9b881ecc2cc033a4a97c7ee647c0886f588e17fcb945abc385af015499b76ee6056ffa1327baa660;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4343d5e1237b3e93c1f2e5908100f0438c3d71285b6cd6a27dd92c63129cbac964d666fb051c79afce4f85045cf0be6d3663cf4011bd7a8b2098318ab0d6f3dc1ad9acfc17e6e80cdf086ac37d5fda0f76839ae2d85844a600a15484786b24f7fed7377ec9872e0f5ac5436ba7f0192d4bce5927a202eb557cad0c82b30891b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h585b602d0044582971ad2e0444ce48ab3505b1f89918b24ab97632e20c00262efabdb23c691eb039751992742532af7a887fd880092646cfa8acff39591b1b740ec6cce6942b46bc239f98891f10c4742c04ca71a39bd3b8cdf1ca26947898a3ac2766adff7b4f9f2653588927b14ed8d0ded0ee7881a005a3a5299fa694d935;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h978713fb65bc1d546adb74ee9bca0411af6686946e024488866d0f057166d32ea3e0828d3316676b155d7f497a911dd791c964c14e5794693786491f3f059a0b1e643cfa152ff26741497b10229df290362f79371b9dd4ae2a3f9f6093e0badf4fbcee51db91a4b4525d361789e00a544f6a694f2891744e8f1ae4ed19c7f9b1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4aec8a123ef46b754c104045ea23b3ac554c2aa5d06b632d2852968e049b9f2c0c99dcefed32ff5dd80b4dad45992996dbf088b235c5f7bee8cbcf03d7feaf7092079f54a41336c3a0de141b57da631d1861f1b5d10fd12120cc971045a6fd6cc607a5d809bdf0b189fdc661c1b6d83d9e1ccc3f5cddfed9d8baa99a23309314;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9fcb66253473988a612a6a23a6811726752fd9ec5b77fc647b67c05c12fc5cd44e1cc444ca5646a0bb5cfe7807348b557316aa2a380e057d6c25fc34d12b101e993d41467f9dbd7675a3d8bacc9236fca36b2e30d25a739d890eba649839c3aba586d32a692ec5ab6a5872fbd7ef75809db29ba070db6b6e94e3261fd186c54;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h27436dea0e8571c91d00c1b6989384650d43d571d543eebc6f1cee62a7c88a7ba8b0133b87008c068cf35dbdec9b01336cad4dc3328a6cd137d21118cbc6200bd655128ae7d03fd84592c9e96c011a575e7b1974a81233937328cbb322bedaf73e0a7e71af0ed0d84f380ebe0ed7074ce446fe9fd0ca1191b8f027455534863c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hde165efcd7fa82f889dcb1f5a5d69611cc4ce415382b066426998650488c7b5c9db61bf799353fec84fc1903bdc86e6515bfa78ec4b019ada304b7bbae2399659dda9214757b65311872ed4ffcacdf04f8a3538d8f6d570691da581364db7d149a96daa990c46d434fc61f0ca1f0b4257a4368480a48154323af20d16dcca454;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h31562cc5f1f7e0d901f9fcf93b64967917a122c656de0a2dcd0dee8ed4b26f3b6b1434c1f6bf0de25d7c040a1f2418c4bc25b69004c357557a1d2d36f1a9a760fd8281d1f9d6b39163d9cb63dfdeb9abe4d2e8c2e3430f534ecef06f0975208df55660b9b2f9cb8220da715d37eab37fe38cd7cb97106a3c1f174e113d5f1096;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcfc747b2adae75ff646eb87eaa82449df8ad37466c85d98c22603cd0918eed6b5d746a9a3b66d4aa8c607f4372016404be341f408ae5281be33900320ae811fe41d735ca9b998db52460c6bb5e9e42dc6ee410996dde3dc0aa4fc75c5c611c839d50de683e63d265b517adfea79eecda23cc13bd54f6e0fb89e1784ec81ed512;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he3746cb25bfdb222383aab386e89ff55c87d59f84bbd297d7e9251d3ad5a85354b81148320bc0782a87aa25c311492b3576255403e6271117a9459701f60f3e567ca8c5d44ceba308e6132c95604d3ecab131330487fecd9c1f18edf1eebdef1d7eaff5e1fd757d5b6df2ffbe18762c834a9057147f92cb3fc54dc9ecd057a3c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd2371303395492a595504e95b102402742ff13d2e967c0ee16e2ab7312f1b38c868a81e6dbb880a4e8d21ff76ff020e2995e2da679491097215b1ede8f00035e300a34a3ae35d823af8f08cfc7e59aed59c7718d6bd8c62b2ca4bf7f45408472654a9c1e0a55b93ce30242b477e2f84401792a3aca9d93e1f924fbbb1218ef8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc52cde26de59951b501063675eda6b85b8cecdc672dd751e3aa333ec38e8f8efd7db2965beb70af88e57c682dfcfdc1b10693d87d1ada76043bc819a4fd41f8a0a6802ec519350f7a43d4e297df98106c0e29884c0c8baaf6db23768337ffcf8e80623837c65e3a9e4e464bc3d98aadb6796759e0044c272639adaec560a6ea4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5f67438a0d318e5393b0405b325b531a17938fabae04b193062c3288d836ad03e9bc80831a0fff9bc0dcd7591936f20d3b355747c616ea905a878805d1e9ab6c07da6c571bfbee35d59b0fd0ec30bf62b5239f934236f95a5a488c64b6114ead752568a2d52dfef274b920e671558921cbd0921a2ddd2e013e5d1090e5869c72;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc396d5b33e9147d3f00603025ae1e502b8446bbf832fbab17467e8388b8acb28ab54a003efaf289e9c2c534c588f3212a41923e734bbf0707d2ff0220e68770b2c0c4c0a9113040b75b3f53de1d47fe6e469350cb40daecfae2edf75e58d2e4ed6c7ed7434e6822d0aee981a3f8fe3062ac13126f9b8654799d0bb5960c4616a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h84984ad9b615904d905965224d20530a5d9e330227fc955cf1a9a40c6330218c2f51161eaeb19069ed905ac45f710cf0e1afc9726643eccdec255716a69b1fa4ef74f116e47299b1685e01afabae85536d71ce8e820469a110f7ef71ac8c0ce47a35ca8f3df718977417348e66ba9cb183700235f0840bc00ca7a8242b78eb0e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8b05fa62f1f0deafc256a4d040a6a13b9efb78859a24307047cc4481b48cdaf50092624e90d532fe0887f8319c1e2ca842b78394533c5dd2413d7cbea3f5e39f0d8fa90ecd4efd7607dce3cf4abc7fcebd0c50b5c27ca471083bb71bb0e2d8cfb5b13d4395ac1905be44799c2cce645d2adb7b6fc3809cc2d09fa1416342035c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h67c7a71bf7d4935c036fcfa7ff76454f7b7bcc7f57d33a6e9a3a4d054dc79d71854705f9965c49c0ad9ed2626c24e37cfd9b843e78a3386a2e18c84d557560f56f91c98e51ae4fdc0232bc8857971450af19655263b1539808c01def02a4eea819f756050cbde819278dd691a0ea162f7b0db234dd09e007f145b6f25624d92f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2402594a5e7f2a2947f9ab263f4d4b79a1e3628ef96e8c625503cf039d25293683c1519ee30d262e078590c449613e7b4f9e846bbf74fc004560ef72285188cb12992f1deafd1e99f6142c540e1c105b7022ed6330f3992ba21356ead3a0263e01df48996330597dbc335bd23cf5c2d132cb416e95616e23390941629f71debb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9189d0e532d41a605145834d0ffe8abeb45fe6948f4ad11ef635c316ff3e897248df8fdd6c8a102d6ce9c827187248eac11b97d21eadae6a3ad5647afb4cd24a559d89dcddf813e12c20385c5a2190b71835dc8761b559f158f22145489d113240dbea12dd7f47d0b92f5a116e62ab06b676786a88cdc9df5c2aa843b6ca8cf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h78e5d5d29da19d8ad56bfc9b289f976347208d8f3aca44b6d9cd321d1ac86fdac207d5c4bf5f7e5dd0647ee6abf35b5533ef3631eec6a43a2bd0c47af0c8f37bf3ec8531cb269a4ea57c1b6ea2d151e1451c9e607e9304fb800102533b6e12d0980a31cb0dbf0db98b99c4ec52d835a97dd73d4476a404890f3556f794dbde65;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h23dcdb8a0af9982b58402c72ab2afd29cb8f17b2f4aec4ee0813a5d189a70a40f9ea52f1e70edf1c3897f7b44725da9e899d2c5128420c9204965493cec5c29a0ac629ce50d0c52b341a092a3d70d21a8694885a37b40722c93130fe86684442f75d83c221fdc674df6642366b43c89774861bc8f0f18bcbe05160e0d0f73b3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1bcd809e98ffabf9efb8d18f18c61d557d6a7e93b471326cf90136924517ef01c5f4e44ce93baec1183aca6eb6eb649619b3e52815fdd2530c46867d2f0b45cbcc3c38b061512466d6ac7c8500cc9aa557dc33417ecb0752f0669cbd3303a3400cfab8e84c09e28a96bd63fc82398b5c7efa3bd9cd441a829b43bbbf0ad1ea0d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha7d8673cffa42776956d8fad572838cd60b8f6925470d69692fa13ae19b058e864f0b78d730e41ba43f4ade80fcdffcb17c763fc8939897e873f45a8c6f2c574e5b49d12b9105b03c388ff8d66c7160df5ba4a087f01295b822cf8a6ce801c999375c8c5e8eeda7dbbf9e3b4f25046462a4434db141fb4b102d2891cf9f61056;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7ddd464a28a4a98e3a03431ec6e4398e3d1157b05d86a7ea403e6e75bc053c65c889aad9a788fd19865138c17bb83b03e33b37f3996196e3d39db594a6f5e7351be70e1c6ea8156b0aed4e0d09ff7acaccff5b06aadf0ab03292d630151defc7478e16b52533f01492efef37037ce9d9896c1163a3e066c0339228c42ca893c5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb17cfe686fafd8e2f241dd529a35f7551eb30d0d7f0f76fbdc79af11ccc34534e7bd130ff24313389808a91a8151fca241af8d00533055d84574afa472a7d719bcc9e16e03a7eaab1d65ed2f4cdc81ede41ad1e5e4285acd864db20eae0712297f6796cc1fba14fe2bf47387f2e7c2ef9e223e51a8e692c6d9ce7e6a1f115d5b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7ef96a72ed06823983f7cf5169caf777542e5cb837b7dbdd9683905f4b64a0c6dc6b8f9e48452c9779719051dbfccbf083844d84fa8fc7c56c591e0218e33839e1b8addbf576257b71751a636d5e5dc72ad9506548d59160a97499bc8ddf9a950fb7417ffd07d5ff484c00d1fc7568e095462032c92c51e0ec1e7d3eb4359447;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h596bc1fd8e944b5859d2b4ceb6cf600fa3b418b675b51103cce46935d6131a63f45a8a91c2cd3798958dee38210bd70e814b6d1324954376320c55414a9d5cc625f7057a9b2706f81d4ac5b8161513c1cbe946790633fca005dbf8cdf49ce3482f53fe223e7dbbf3cad53695feb9dd07be9303e051532b2758cae612003a2b92;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h748fa9e8cac740718b552870baeab2fa317b67df5c44eba2500be3221f26c37ea8ab4687260e9f0c9d46f967ca44e6f58492038bd27e36c6ec3d3f989b85427681cf73aba5f81a646bc9aaa4346f1147f557c4059c1f9c94fec8f94f939991c91e5cede418870bd55a9d961c4c65aed93b7668fe63858ceb07c0ac0c32090a87;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6fb0fbd1386a7ed9ca310885d0d4305ba71fd2b00697fc644cbb4c285427a0ade91878c2761a8f1e49423bf851cd761c41ca6643e4e1c55523326eddc794ac17c7f81da0285dd7157f0383d892c83894dd436fd48913bb9a40229b4cbc34a36dabf31803a47dfa2aa070ab04bf4ddcea9ccb1c49c7051fbafb07084d0c6858de;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3094a28f29041c7c53266375f2c443cdcec8969384069ec6bb73918829adf96d31808b8f6aeeda1dac15a0071975353796ffc51d633d4011923f47130c4baee320274559bdf79a55f2a4afeb4f214eed3cdbe7ef4321e18a0c816bc4885548740f27448767561accfaf9b66d8b20803b1c7e23958056752f81bbed07b00bd972;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba061f0f7987518932b74e171fb1dd6b1a4b6c00d51eb84bccfd2525b0bc2b784f5f5c6fef4b13be42d404477f6d5c885a67f7b5e98af50c24c0fad4b7ddd76663d92d1bf034795b4d38d902264c855f43cce5d89ce087c352e8e308d8e53cdec91c689795a5202abd18a65dc266157a5af6b8efe45d3f90d069c3bfea80ad46;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf29e5cf3d4aff348b11e7cd8b5c6c7b704fb1ee5bc12cb4686c2f0e3daf515c34656804bfa4c637cb02daba18361554220c2be4074c5cf9db1928c447b2ca1b363fa310a2f7d64dea07e25f80c9f97799d5670803eca1ca60bab82633dcfe0b74e65c8b03c505c25f791568e9b7b7d1de2ba94b01285f5a01b1e840b166d37b3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h10bc6b97aef8714302416700becc277ed8a914bba8488617fc4738aa501b672bdd4496785defebff41ddc5b01bdcbd1152660d05f21bfce22e10ccaf5f1d87b406a8e5dd35ccbdcf8ffb1b55336ddb4d4fc8851afc037c28e2a4bac67e833c1111473ee6ebf73cae5617db97f362cb64a977eaae2d646c86d3f601c0ad9404fc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb4feb18002d8d8bae866956d2e13d29e88f665e885d6a672e9f919c991c57487b79f09e7536caf4b98005a10dc0517d3a7925b5c425321de413de67521bed74cc430e631bfa6a6e0fdaf8681d48ceabe79090753494879fecc5847ee7aaec61b8d99685d7376f70d14744d2714850dc5b717015d321db971e8f7aaf79d45787b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h36bdac7c857aac920edbaed068c7ff50cb8944fdc0f9822038278f9d6591a62382dc0636ce02bf71309acaf856dc1677c120743cc84f35958470136f6f11d78121bc11a5cc329887623de8f289bc0b36cafaff7fc02f7e4f0d168e593e99dce05ae423e22850fe4e6114d5f871b13660c32fcca05eded5b5b41c53e8ec8a094;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf5d1c5600f997b3056903dab8c7a15989087b50cd0958d29b184caeefcd9e5382ddb11a1489525911da01764c756473255067be24c8ed0eaffc1e0f1fbab9466f4c66bcde79fa63885776df7727f4c7aa2489241f7a44c4a73bca282b8e4cf4e1f869e3fc6fa91730b5d9ffc6ecbcece1fb5aaf15c22d78c6d3b3968d54f0b3a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc88c63cccfbca38bd5366a1a1d36a2e4841da4884dd109901531ff8bdfcc07d849d60b5330c8d0639dece7238a273f6a920e53f7a30075e918de5836e15e923fdf2539f04f73b4457e94e3f1d99c7d034122a9ee1e51190f94114bae26203eea4992547ffab1b02c840984c971591abaeb479682a80b377c81bfd60295fb8a34;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h106156b2625414a984c27b40fbd6c901304714f31612a30ea77c33922c9b1d7cf3b0e7d96346fe2a19262df4f66655cef53f532c0cd114e5767559370975d254c7d62bc0ba177f089f74bc97265106973a179878cf5cea7a5c9e7679b366616d8cd3da143d362eba5c9725575fa662af7023a1c4dc7727319ee2b6f3052e0fe3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3afe65c6f496700c94cf92f10104b135bf3cacfeaaeccdb0f3ddd54889816d0d0b5710fce0382a791cb6b1898cb87c4ec405719000359686c46f2ec45342d4ce30b89735faed993123aac4af1cbdc8cd7f0bd11b195e2bbb541ca41e21ecc7f5fc16bd54544e828f3ed0642f9d521abf26878fd03c417396245a66fe0721274a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6402f82e7fb5a9f5fe344d294d6021554d04ede5753dce8723e20a1c0dc2cd4e9e137be625a17d2dedd17bfde70f8cbb9926e3e984604ad5733001886094a51b882220b47e78e331d01c705f8c8d0a22eb8c3629fd5019f29d4c1d7600f3ad10759999ce7af75ee44dae656c157fd458e27bd8d6242b0fd5626d0aa427eae3c4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3ff906f15dd4b93cae5ecd640437d72c39ed52558ce661fa62068a109e2b05e71e56cce3ad1c0108505e189cb64c89fccaf001f2affa23bef1249c2d1479dd6453cdc92709ad04336e99172522336f93ef80b3500130a97a9cf10126c796f3982e9d09ee3b91573e778891192f9a8c12a1eeae67154dca52388907a4bcbe09a2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hefb1ac9d85b81b5eca3af4ebddaad4e48d4b8216ba96350db01b42210999b70b2685c52b772517268920918401ffe3cd110fc415c8a4e6865108d5e15ed0b42e7098f9dbf9d64e86743ea512bc2b86e2cae67bbc7c6ca05c4f00cd7293e47b8e3185d1e1fc6317418cd2e63424bc084b8237487550eefc7ea4341119ec60cded;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heae7c27676849fe9aa781dfa053798e08c17277c77078657f63cdea7b4021a1b0acd8f6ad4ae741b4899c7b414cc57df4b0e3f9c3ab923a116a69a85f582c4e888ade12f3c0887ece9f15df12a7f04512f1377f6a390c8e68ef6d84e733bc3d950add53bf5af54b05baef5e232dec059bb53be033c136d1f1e1eccc20ee6d190;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2263fca451fde479cc1ba9c5c017afcb5d8feb4aa896b01a2917940a66e6d4561ff71fe0378061f83aad14033f46fe5ce5a84f752e2fa320a46684e6d513a86be8f4c27eba1e3976eecac4a55bd50aa95e3d47b4e438a3b4e57b280c63c804b0b1d11a99c8da49e2838771a5742821bcf454381e783b79fc7bd2c65ef6dd88a9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4496eeb307f23784c750dbf550f4b610af92d77246c08d081dffa702539d464a90bb7a1952827498d2e51be63b65bff0756a3e0c8dfc5c818fb4ba3fcc3ec5d845d2431f8a626cc976a57c2df5999a513f9fecbd5de07a5dc09b4b1796d43f087fef469b3caa62cd6a8d18e44125f8e5c91921e5e3bf566715f61f2a966eea03;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h15fc2e21039b5857b391aaaa0be16046a96e980ffc44b9be21701bf314d94366e565c0d75e9619f1dff3fc3a40d52d724c9e6842a0ed3842a4a92f2a98d92853f1645c0ac56798bb83cafd1539a8dc4b3832fa73dce17f445e751aee5c642e32cec74bb43b8174b36ccf4226fdf3f75a4211c98b2e73a2853b71196fb42978cb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3ad40d6bc997ed522eb592ffda63ad4f1b592296d6561bfe174c461ecf8aaf99d7991d74b546de6322a74ac7acf9546fb8407375f643930d11c20782d7b07c40721670d45713ba4bdb58e8770657a050ac55c622ff937e7c2bf70a5dfc9b75e00c39ad43371eded378b1c2e18135cb85dcb1527636351bd3745f599c7e31c0a7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb06d4bfdfb88090fcccb044df0780bc895ba6c9f9349b1618ac96255ecb2123da9b785f82b4ea9919c2a37a2c8039fbd119c3f02483a920ab336894f41c775ecab808e625a8f00dba6da6b80f04ecd2a61b76e23684b839e6fd36e96e286aa172a5ac04b44c88c5292991f951a3665640041a6b71f3092e98470521f0113d6a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7605471281194b4a197122fcfad8b821802438c6e09989ae1476e775117650558fbfb0bb67eda3ee916d45597b54624f578e1efda9d7c7c23574fed9644b2a9dba85fdebf811863c8c39cdbf0ffde63ee235354341d91ca4114f8ebdb1616b16e38856fe8953d5ad4a440eca170a469bfaa8c1a4428e13a751e3fd08068919b4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5dcc2c362119f4bb2907f7064d92396230b71f83d66c0ec6ac71477e16d87a8f47126ba83ae84a33efaa9605c347099d4afe75436bfe996350e45ad48d40245f034d5e084dfecdafd77d92065ed4319604c1ed45bee1373403ed5e5653cbfaad1196f3f2e1b5f56de77f78c72e09e805a09ab8d8dda93f3fc13475659788ac51;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5773d2bf979dcc2c6b372d639a355d6a91e37896dcb3c1081f564447ffd627e29c9496cf78eb1818a21047d15f9ddcfeaac5a32880f86fade0a4e60b8a9d26b9f1317ee6b142af5e29e96da425f6207be4bb4c13d739303cb6983051c1949becaf03e1615ba31045b434861cd0a25546272064f6a4f2beb34451caa841759159;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h91ffcd34dbe929d33b0af652e9ffc4c71c940c9fef7293ff0a0bd900e23b98b006c79018ef00322f60036f3e41e692e13075890bd917ace3c5002886d3a7198fcf216f1def8e4e1c247dd29e93aa34ca5cf1cfea2a8a2a7652586ad89d248ce01945532eaec8b2ae593bb9ba2633f9001e33cb7bf3ec7c076de71c56ff36be9e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hafe9445577c273bdcf239da2d3480a8f6bb4ad42aad3e83efebf31939d930727bd949bee037564ab637aad0bda23036f3415301f1b5e1695103f18da217dd93fed44613d0f978436f74181d72642515904b27f82bbbac30bfb973e2bac02b470013ae62bd35631c113af00a569687ef7d1aea382a8fd36fad2e94b9a1a0b79b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6adb1f4b60f1aa9e75edf2c3e3f0f41a6ad3559eb73d536968acaa0c8d6c9176d58c71a4d40af4e32371c151fdeb32beb1a8e6cf7120b89164200c50ccaa14c7c142d5175a504706b4f11ea8c0bb7af7e8c86681a02bb594adc3ebb902e17270841b836158131f0d11a6f2946665632551b9059f498ff3e96fa3709f4f997585;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6dfc94bc884e3a370a192622fe37ccc41e2038fb658aeb66c9542122be537e892e57f14db9bb5081774350ab1f2c9803e39ca887d36f39da1212a9e5f3813b23e3b91686e8548774934c5048624ce79ee8eaeb373b2bc37ef7bd7e0d83bf7da95a008e10caf5637f7c4417ed5673a50b1b725df985c14455612936cd9ba276a7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h11de076a0f28014f3c6150ea5f149b11b57146430baa472518a90436e229bf96b62e8f9d06142f28cf8c6987475719520efcd3d8c5bc5a87398fc64774611ccb64230d6c0a768ab1202a17ca0f2e07b55346320fdb7469a9df1a14155adcee27a2cb802dfea4fcd84aec59ce64070123e4295862297d6c4555b63521d7a9079d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha7fefbff90de78319274922863f745b305b51bf9752ade5570d2e138344a2de6feb2204632ecf47f6d3b242320b423cdee79fbaba6a9f09321269dee5a5a19cec8788c7b378618add1cecd11ca5f30be5cfa28776a45e94e1e7fb44e1bf10f69ddede744ebc0d548af514a3b398976df21d896986a8d9c80f31e3774ccc447ea;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h312a0c34a4a086bf05aadcfb6c6c78ddac22620a068e6c25fd4b975ea73650faf3a711cdea617806c56971411bcc754dbfeec6f70642ce56ec602b7e523d60dbb7155604977cd9377449d0cb48cfb6d4a5681e6c5dd7d5247b8474f4d68ac9901e5339c8948192060f87627913bfcc677faa11d4682f39e806e52f855c2cd9c8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h34e7838b7e09e8d5a5c722296602e0c674a9143dba018c10e66f90cb115ea4a3d94cd3c4c8063d4f751c2201878f4fa57e3a49450c0cd2b304a071c207a22d725ba39eddd16d340190c1e1f21be8ea13f592c5a6a64578ac6973f9209899ff116d8cd1c246c8b5639ec6ccbcc0b0933d58655598ebdfc2ae9b7bc4e037353ccf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he56c7ca6018a3c90260fc2c4bd54da314c80ab7ac9969d23fa2d88daa592efe1d50d64b06a6498f7816f47f63a48f40b1b467199c2fadfa7351097c0fde28ccf4372737f43c3e83f9ecab5d48326bb2ed9f14ecb90ff2f5da9d112cb24541b55122ba525e222a6350ac249c5314eab12981a1fd9005048da9b45d55b2936257;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f7ead44a6a46e3e3fa39c7c8e5fbe6900d18384c6f5695d0367cb1a07a14c4b8284d386f4c5efefe5df2c0f29f29b6c9cb0e451b465857d039762aa6d7dbc8dfddd8be8e51c0bf791009c8ee4b301ac94a34c119ebcee692b77767c328cc4a946f2bc0851fece2d59891e505346dec939ce78d20f3b096eb484ab46bad6c967;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha3f18d71c5eb9e392bac02a034a4343a712a2fc1a1215964931509e8528e7f9e3aee267474d86e2ae29e1484a330ba94b7024ada211ee686b868e113e1553a9ec9be5a0c2751cfb4970b2c4de70a83a9826a422546fc8b9815d06e59292f76fc2282485a932bd02233a6c222618b626f7ec0e947ea978f2f644f0cc171a100d5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc7cc4ba4e772ef52dc0e1c866af353ab23096c961ed1a81146d0b714edd7890a0621a11d39578d1428e8e64b73b4f70230f73e16a86218fbc19e8de684afb3fefd677ca4a93c2a6d8a3b4eceec44144a1a3aad73b7c5826d9196778406ce1a4ad1cbcfb180eb289f852d728dce4643fe758e0cd943f82443400f76362b073605;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h33607d69c2119ecae6145bf9e43904290d022e3e61d512c3f3a57a2a91d0f85dc77473b38a1f3cb1c5bbfaacc6a647cff548b839348c274c57419fad950cb01b2c9552a6b259fcd898b2aa31f600fb405887607014fd81040357a465609a090a0342a846c1dcc298ff0c9beddd6ebabbfcebc7469fd76da333e5ff9e3adbecfe;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc2398d0ad322b11250805ffcfd9c530466021916aa8d2d19ada53b7ef1f735a80d6d8b5249f85e698e9c33271af1136e0a389dcbc9be86d1a189f9ca8e04ae54f66297df096cc4b4e6e1e7baba5de70ba5ec81c3fdbe30fcd8bd01e7d2f6267c0ffb83516f92ed41909ee055902834d4bfe270077b2f8532110ffa428c681c1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1f5e65e46b3c1ee53ffbe99b2b3d4177b7ddd1069e28a1f5a27a7979023e4aea0a1411242db71eaca3eba9eb8b031c28928f96ecc44cb92b92bf7a7886bf8511dfcfb6851ee0bd3f13d7ec53bff7dbbce51349dfa59050eb05e25863b65e71b273990905e193ca5b2c5fc97be5646c53cc5c0ab5c1547bf1b8de84756f22e249;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h234a39ed2c05d34f14117b632786970307fdbfb27cc6e02e7aabea8fa0717c19507db6ec0c9d99aed814dd8f7c06a2317e51bbbc25d6c792741e3fc675c58d2e59855039d24aa96cc9dfe875f40fb6c25ba77a8d49b0ac54dd50b60b2f91fda4d2e6008d4788f7f263a739a0da737cc166e23d722fcc089b435afa2327a57cff;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h170152b30f32d97dca0908cba112e9c12d18ebc6fd3bef4e1696f9ede742cfe46c39e5aa728ef2c71159907c9238f1b5e28d8396827ba6346d20551b5df372a7b09eb7745b3ec6db81bd1ba14109d19142a4ec901c7ad092374f7e3b2d37dea113905955d58fd1a08edb89514d919ff2843bc1c2bec1bb0e7a4959a9a6ceca7a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h22dc80d9e1a57a0d72ec473363eb4bd1d3527bf5b1efd9170b79b10e9a54e3d89209e8b7185e2ca0f03cfa64dee286eb2810aa28bd40b20825e159d0692d1fc743a5ae27e919c1b8aeee747a0c23a49d80fb90e738349fa72c9a155aafee830fa18412d121da4993ecc4e6769db9b719cf01230f1c236686a7534c75299d6706;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1ac06ad45e81033cb3cd0fb212767263fc029eb7b9c178f32a82822e64c34571c0c5bfe2fe62c11e54bab15e11c35c313c865c83d3151fd9ed1822dadf59f21b18a61011db0085c779cf857bb7b6c9aeb9fa4d04f68fb4763f68057be3698f8b4fb0b5161cd4e71ffb0a8ef910b33f6b076e6e1a7f7685a7b759b276845142c2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h28179113d8050e809b3f39f1db8bdc5061246fb9c39d9a818e9d69255182f2cb8288c7ea914f2adad8323dff32b10077cee194ec637b2b902189dd39e0b2d8309a04f5a4cd5c4fd9349ffd6bb790f957a99060cd3145bfd6ca26f8c5c170de683bf88b4cc6223e2a832c280b4d6683cb34dcf0b7330afdef4d3190e9b635fb96;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc0ff861e8fa73c83347077b57e1d321eed293df9248d55b35a1e04022976df6e058b8ab69ad1ec30db916404bb0d0f07f3dca723e8c2479d843270b9084125d699fb96185c8fb248d21064edda8c19baaff176c935b9a93085ac83bf3cb57b292b64deafc0dd5dc5fff4bb3723d506726f07426a677533577dfd4f5ae60324ee;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heff5cfabfb97dbcfef00814174faef16c1b5995dbbd45d9832497e20dc5787975aabd93ba5882fdacdc0fbfb68c63f561be7f2b946182799c1f4f149e60e488dfc190543e14e2bcfac89e0d25baf10cf5f9190b5d16c9dd75906e796dbbac3baf890ec4f93d0a4b62333da10dd0672b8355ac79bab40d4e3bbe022cf5312154d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4612688786a48c9fff7f4f6455c9ed8af96c26a8a49cd2df4544de6c6420a64ce4578998522f9932312de0c01cbac82aa81a4a1ccfbef26e8895661f9fdbc6c6cced2dd331872c578c3b0e601135bdcd6844796e5757642853ee22587fcedbbe0ec03e79340251241ae7cb83c89286dbf3c2f950263814c873ade6df77bc76b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h772fc5610a48266244370c21e8e7cf9367b8de05af087ced8ea0a90a3e86035969f9019b46ec1bf4cdbff650043c2edeb04600e1fe8825beecd6e5012d2704cdcddbbd149cff1fe190e27faac9abde1e780b44fc5e9032e4886ca1af9882e7233e6297cfc357abb6c30c976699e5b52e5d6d732f3b1c7b8bcb0ab3bc47edd967;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he3dab1c07d64cfc8847607d783fbf2f09a2c2c7c442c1a5e49de03a2ef60f367d3071bba0f312471aa35266c9911c84b181f7a5dcac4ea1aa97089d13e210fa419c8180cdb9ace8e32d42eaa2c5019f36bd5321429cc5d33dfa77088b62da21af0087b47d73ff75f5fd029e3a4587ea8d2b697b7740bf32a4e5554d88cfc66cf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h421461799f45eb84ff0049a062694e6083d18fabb279d59dfc41b909097a659b85204ce9607171252141c52da4e872988c0cde35628409d3ca6c16650e37c50941c3b7bad1f28f54024fa5ca40e5841f1bab4b0abd02e8285f3cb7a1b05da4a6326655c1f92a7bcf63c70b362e73f1b7c207e5fbf9daf4d6cdddb1fd1d60bd9b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2636d9e405138c7e073e3f11a14e7fe72343da552a22739430cc4675f00943f06e61987655e34c9e8767a77141685611c496c033c6e6a1f5de9e97f25bf1df2a10ada9f25c8eff59d25def84cffe2e9bc6f68372a3272a34ad066cead0043833e496bda0f5ae99018a869dfb9dd7c64cb18a7d7016f486db2d0c769fcbea3a51;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h67afa8385f9b1e0af60cef9b45024aed7a122a26788832f651013eab1a8a8fd2a952dec0ba4ebfe471c60945053e71920069d83b1b4755804fe38b083837ebd4abbd30f630e9d5e5683a1f83d3d7d0096619d774ca76a194f18e1f3171bfd05f9332ee8fd8223df41fa8c990c47452b12cff8a5729cda66d8b48ef951303cfec;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd8d854f302a0fd2f83d86b28e6e460b5bee1041abae7fd8792904cede10c892355b6e309c512a457604d90dc4d30091e6ee88ee390ecb9ba90b770d971787b280e4da957385f851815e41ccc6837d7e79b06c65ed8e7785e11a9a6e0741184febd92e90c209f3bcca0013784af89e3a54383bbc9062fe5569a3ff495e1606f0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdffd6cf9d415d8261e736d981354cacd2fe981efeb53ef2bac9b6b7354d42a6cc38659a80526a85b0ef174f08264b02d038557b4500e47f32c418475c9719ee76922691a45ee0dfcf6fb040f5223c74aaf75ce1b1f590556a27157cea4a58bd2b8703c63623e809cbf93834f4a7f94fa0cad0fd9a91506c4d9779ae224642f51;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1ee9371cd0d8e22acc04886abeb964e248ddac8a247767e069447cd7d66a481bab7baa16ea767e884bc59b385d9978b8a3245d876892297c814ae43464e6cf4904650e498d8907e460bafba763ec0fcbb5bbd3770aa7fc898b0ec978580829eee96fa08b8c7c0e0cee61cd90f15b8167c0bb7e19ba0520b6956d1428f99ac83f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8a9b5bf15851075c6d8e715b4601f2c79a59c333cf7e4c6322fb15edbe710135a65524d6ccf6f3f27e713317697a645ce0594f22d7c028842e0ac5b2627721f2b83eb22306cc117e248af3b07d094497f24aa0743a8835c6caa1a9f474339a7b497bf4908f5ee5e45ed77e3983b1cacc020a2f04d5000a36c3403e285a711a82;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h713d1a93565c6bcedd3e4fff9097c27ae7207181ea46f27f092f771d4b0f386b574b8ad4418065e43acc3a9d84f691319722565373cb16a44ba5ff6288ec1da19632c353e3020909dbdacbbcbee15e5ba4462ae9b3135a580dc96bb7d1f68fd58df0497a76dede1fb0d294ee9f470281bf40c9abf72ec95cf1b198b0b9ce1fd1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h863c835d585be9806f3374cef916c9fbb39dddcc25ffb6bb3afc981cff776b4bd26a1629762a6fc4625f8763b1de33eb68eabc7d98428b6382bd0604733dd1b06dcd256d70c919172a44252b5c766467925c76bf5b21fb88ee02f6345334f18117025259888b9fcfaf50bab5c4efdf59d72f4af4c8b753794974884637fc2199;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h996b00c78ff6a124380ec55ee9aca5c43bb7f287c4a17f3439e64eaea3038d5da3f6f0139c67f462f4c614c1231be516fa3c8bbb217bc8abbf5ae80986864c46bbef64c4d085a53a3e6f71888a5f5fdafff1f43501e2ad41155da3c56475157aad6f2a53f7be9ab5bedadfff66e0411faab18f60f161b0de00e5b7d125fe7f83;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha009679e8d6796c78e09a7430116fffbe691ba8ed91a6fe6523d4e0333ee5b7dc2ba2a7b9ed11dd43b492395f01e5ffad29017b7a79eb76f17bbcc4ea708854a6d12638c320cda04e38b77fc0af1ebeae8c61c715f658435b1610647b2bc18f5fc4c503ce95356a7d759a29863a6a3e3266996b5d73bc02668370be187dd2f31;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h25cd5176d243fea9bc2a9de66001932ddab4224ebea08861b6c64d678db788308ae13bc5782bbbd35ae8fca336d91c7f69184c5f2cf1655ee94593211872190703a26d839bcdee508d9ec5277fc050028742c78d704f1344eda2b829f637900d20439ae977ea42f9b6e81c756bb5a19d2cb65884273f25818979cad9438cab98;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf2fcfabf2033ec81e2253d034ca466ceed5d2bcd4290c4b6ad2e939245e21aa002a8021990843ff0f1720db4173fac2379b07d566a4e955d9d4f102d495382b05a5fd6d4124046ebf8e437073adec08062fa59ac0f5a4e19518d541bd992dd04b97151e0bf89825ff41e84dcf16e0959de4a52ff2214390193354f6a8eceedb0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d274ebf5166181e1d0901fbaa23cb378c214d05f58c1f4c4cea8cd5ab8dc774e39e8b6ace4b959762f8cab221a5de337f64e4fd8bc154d2d9c0c68d992b98cd0393c28edef2dc5e4d676c890d4cfbc97dc8b67c9e71739dc0a6eda7f05e7a037d69e0f6f2c2394ab22578f25dddb623b7b43cac96069dad586c56492b68704b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h31ba205582fb1999794a4179573bd6d48c71fa538592baf09b8ccbef13a85f4083f8e7ab79e7ec5cfc53894a36c5ca8a29b788b4203d3d3716f9fdf1ec1f2c70ee9031a89d70f8172593ecc1477b141ca0ca2461f3f0330cf65fe1b6b248188385c547ab241e10e75d535d8b63c24769f8f9e05bae0e173707dae66dc571e41a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha35411e1f038a158deeb57083960d1e213a14bf3805610b891646bd8acfe98bd050238a9b4a0b8abf7a5227027a062dc263d255c6171cbcf1c934e249e0b130c662d12f7c8f39473e63a9405d7b1171c2689f88c3ea5450da2ce534810772449d6d57a48bc9b1eeffbf5cd09b58043ce7f6937fc82742dcc7f9d3f511c8496d6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h906f9f275e70112ef8fb06ca08597498a9072ca9f8cd3aefe84831923af13e03ff478f0724dd66187870bcd4d402853b02e83491911eaed9b290b781f6821d51172d146a928df544a8d7872595aa152eb39f4cbd8e1799cdad4dd32c348dc4b7c9e8dee91504fe66e94dadb22f216c92bb8c7ca2f2b8f960319b86bcd6343d95;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb8b37245165557f25d099d72b479310c9747b4bf3bfcc92babe474408dfffd7895165f7d5e2f37d5e6f2764ad8ad02625b062c94f8163f326dba67f20fb62da58fb65627bc1e12dfd36923fb620537a42689f6966a151e491415ba8c10ec662a4b2b562db497b3895e42d9369a44e023d33f64d1b3a93c309ab717ed0fc890db;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h342620e5ceaa6f65ed0f2d4f22826bba28c8af15b6841709001415d76c9d7d6602c7044f12ef58175a64416b79d7a8f95ce69b8920f29d66cccac404f57218ff1fd519c28e643cfc2f505fe618cc38d31693a34850691ec571fb3b656b49e19dd8650af7e5e13fb0805ac54ca264236436d2468bb0668870923e20f0b7de0b14;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd5b2dd97b4c6b103d739ab8a13236db9946e6df679f12e32f09a5c70a080207f99a4854f741a62137d14c41be05e166c600fd4a9260abd7cb1e762feda50e98683ade2403d24f540e51d6daa55e7cdaec9a171dd932bfeb186c2fd932ef8f5e24ffddcfa7185886837925b9c2841ab82e86748f0346ecb64a88b554cc6fcdfc9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19d83158afb456af69bb8e6cf7049d35cf81ba74d94de407aa37687715b119c04a9018a3cca5782f35cdd42a82a01ce19c4cd62a1a64bbbd10827c0a226fdc2884b96f1ee231142f01a5d2fc5cfab8cf0b849312c08e7dbe24f90aa1a1c1baf4572010bbd8900f69b4405d31cddc308578e83e4bb0c24f06506dd71fd30db5dc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd2dfa207a4cfa555a92938504fde716f833c3fe1a1b5fa6f7ca185f60d73cc10a5f98becf1248cda1275bac6e3fb7177e7b9c368bef89a9dc2b0c2eb2ca6bd88cb351f020ca12a6cf555a2afd091a016ab1102984eb75771fc0f66a2f8360b87e16372c8ecc5d068d3ef7cbb8212282f518b45482fa49268048f87e1fc47dc30;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73faaa41609cb08eaca133cc2258db9c31fd02f703fe1ac058d6e4d10d34b1bc877113ceb2b6a6e3e72551681bb9422d6f750d787aa242b6364ed25e85fa9a3fa4bbe8ece4e8dbb24bf73f9cf4fdd1ce7e4f645115cb6beba7905c024497496bde18b5a4ffaeaca76d2b8e5486037c41667cbb55f4b29e90e19e773e1e954087;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4fc22c96091e0c4b72ce3aef06ea9673177b943d6c1f9f10003509d2ba52bc6f100389a78800119bfaaf61035c26adf4803e0f2fd424a0a7c37b34e2b011214692efcd05e20ec608ac5ce959c7d4de41e094d636b9613d76b9e60fd1f73868d2a424a512b04cc0bcebd1783eef54433d6bcbd154c8fbe6fbad55e28ae51de54a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbb001bcaddf998e6835d517e1a85c5bc48c34fc31c6a269097aa194390eafc2193299f0428a1d32095122c48512168412f690b458e7a1c6f785e13a13938c61e91b80172eed88a330c0adc01442b9f1da9b452d6cb1b93d725aad406de7790b2892fe7b0090f65b1e9e343ed4555aac79d8db540d84eae332392026b466d2a86;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h888501c23a6ba023d4174b2fe561371f520e347a7947613152d431a30cf50296f3ee8f18d48189ab472f16703ba3650136c1a2bb7bdf22858b7cfc701dffe300a235af165a9340a9c64dd0a2449e56f4e9f2c7528ccd178a3868d8ff758e16c3042f981777e12e038addc72ad9dafb05796b535df3999968e0b1ad083dfa889d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d4060347371bd915012dd32ded4a6b8186900f44203a06bed421d2fde5ebbf003e0a13d2e2dae6e1ea67e5fd09ccb43239e940646baa6d02082511aad70d25d5aecf377a374275478052aa15ff4accf5e5b923ce7acb62e8fe2ea7a44ee59e0bd50e5feee06e2680d83ae9036613b193811144e134e2b60df2b73fbbb208e35;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb91ae1bc1de478eb19625f43e3de13634b73f45836f3bbad2cdbb13659062a062ec93e220d0c0aff8ae35d4ed3c30755a9fbe91bb9bca5793a7e875c89ba5cb418c7b0d477fd315acbf5c0c8f5425834ef062d389666ab142feac3861343f9422e41fe4d90633781a794031bea556c4902aa2edbddfa17e6be4b0cec99054c3e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h11b768522e00168db11f1ac1eceb2bcc6125545cef527f832211fca88bf459b77e1b042cff3f75fb153d8b79532c4349fe78338234c2e3a41579559c8dd1b2dba2b338b6a8dddd21bb7b1323f33157ebc117c04c5f25e27f692608a8345db8fd0fbdc1fe6896be3379493ffa9ade743997f9ce5c8c21a3971193129da5cfbcbe;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc79c40ab832257871a29cccc0673baf7560c155477b0977ccac62bb268c369f051f80a2a41a344476f1a4900955ecbd4ad237267a828f064b52857120251cc90f0718a9e0e5937f40a1d55a6673b4711bddd14f24e3a89977de4c234a1da9a6f0c740ad36e2e6e1e4ba0e38e8a20499fc26f074b87a93244170bb07b936ce0ff;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h918aa93b94b696d64c9b051f4b8285a919d8c8e63bfced2b0c3ac153e2cb61474fed28231325e8ccc1da33a24449ac9ae45380c2efafc4c427cc9d630df202ac565b47a2bef52a75e882c599a12efa439f6a2b83a6cc7b7e04ba86b869d858efdebe5e9fb6d7738df7f667e7d1ad169e861ab8a7ae6bcd7ec9dea8bb4c1591cd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h747485a690a53e6c95fa9c7c846a990773bd50c38a3fd4409201c8e9ed15ec9d6a208e01184445961131fe3e48906b5b0baa7fba272b81988dd435da946fa41fa5f7bd432ea57e791cc2b0558062a66b1ac5f57c1a897b43e20bf10e5d2a98165a54184480351d8c26dc57f19044b16dc1258c05031d0bf836eca84abc715229;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc8f070183eb25d91efb92ee9e3604c11d5b60212beb18bacc95c2b76161970008de666d67ad5a6a78b243facc4b9c21a54a551277ccf1611f1e7a96b12557f617b29cd3c0cf42f4d398f2e6c0d8ccc0fbc56d58108139caa6cdde9f8064990de53f17cb0195c89108faf86726953c7c399184d456b5310d6a7284949923f9ea5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ef10c8def4af9b9e48f5f2d93a18787d12180b48f928a9ce421e780ec1863e0890f014ff420fe185e25730897a0606ff7643206755e6c086dbb863e6503dadaf02e1fc081e944121ad0d4564acef8af89e57fb00aca0ba90a96d8bd25230cefcf8f2f41bd9cceb6bc7cc873d55f82746da71538c5ee3f6f1c09417684af012d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfbf8aa482851c6dec04f133e6dd52f205cbe180a1d0f3bc2eea4ec391cebb4652a6d6222c5a781994b284d62eb9ab74480e20004d36272333dc5243aafb55f5c7ce03332dc7e5b9229f769206adb3e55c4d65e96393a55f3f031612e832a06d4c6b27979ad214274eabee29ce311c7c1a02611c8c781745c0187d5ecf7214e75;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h892eb3ac2f55edf1591ca563288abac7178305de60b1b3a22c51e8a66d3dff83bb1e5aa9bc209abaca9aea69645a828666fe0a526596093a964386af20782d89fb52824a14a8aca7e85a6004d2e1086b89f806c0b9941764d31cfd962664eecf901807a54f6c35dd41a3973592ec6c3ba8c09680139d2ecd2e644bc53ae6fae0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb3fbcc2f0c56e633abea12d9438392dc09d78e06ea4601ebc56efd380091c4188ab14ae41daa0f944278d5bdb6edad9349f9d7064e409ba6a039b78451868b41edaf308110b57542de8cfb477c3cf3a5ae70a143b68b5bec2b31ed79521c9b0d074a3922f6cc6162a61b9b4852930f6abe2d7c0c99e46ec90a3ad7541591f2c5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h20c079c057f8d9052ae4f1fb9d813f8ce9d3810c880d073bd8610ee91c57f556a19f8e1c023d08e2dfd1fb0956d4a8171983a466a0c831a07b91e4f88ce4662489477f441541320385ca8d135198f17281a98ffb3a5ea71c7318631b1275d1350cd7d86c05f2a302368d7db3bac8c1a55595a194d5ba5cc61713bd54d627d210;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haf791024757435de09321dadf0da404218320c349e4eae7166fdc5111602009e711e9f335dddab12a46839be8b9dab0ef6e9ac81abbfe20e78f4d920923b21168dcd33901ee790e5c49f0af9794e6f9aafc71be2d124f686d148adfe903ac48ec9441be2c7dc4ae43a2fd6ea9a1263a7bc7d1cbdf0ca4dbf103f7b860f62439f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h46bbf572464312db0fdd485d163247f036a493281ff73da5b1b55e864b11e40778d2c62dcab3253fb2182ff68fd06124e0bbf8834bd8e22fa8fd69494e2da1984ac5ebc12a440e31e7db8c016b46e235446e27c0cd4d04b68f7fb09e4361af44b21558e2d9bf8610a7740f4a43ea33409589577a71e0fa020320019766a25e0c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h533d674b95b1ec3bc768ae70ad808ac231ac2b77d15010fc0168533aebacb84d05885569ac0829c20d2a2604c21634957b0989d8d46dfd6a1754c0e7b7120b20890be54c8c56d322de30c57bf097c12380828e090ca830085a7f532ace572589925aa941853f099a5096c2af3350ff2dbd1e26c6eafebbfb67d3b2188a43577d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8fc71f054b8e0c9628e5bb03c60aef7f7bdbb066d9477613b8bb3f6a370efed55d078000a910dbcbfbbf70393eab89d77364dbeb57a9e6e7035969bd3df079e5f375e7757555866c5941136eedd782639e1c873c013aba7f477c6a4817872fc0e49e3a1bea9a6d30ba0265d64424b9a5b83853c53a1371d3be5c5be01740d957;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdcfaae986aee318685b6469535b7885784ffd588fa023bfb72827ed503535742014cc6cbce5dbf2ed158f5e86da11b4d6fb64e55fec12b9d1b8c21c653cb2a2c66b9a528cf9027a5e6fe89e8f6bf1d6dc1dc707b38e25ea528f1ccd91b82160bef8666638b5d987cc7d5d7bbd83d250ff2c92a10c2614f001b21635515745af7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h25a3f633e887035bad4e9c826286feb4ffbc90d7bb4845d08d0085f721b3c9be9be9d36e2194a008898d523e6a0bc1f1479e8684990650c280121e6464bcc4ec5fe93e6a90f2f8f23f359089134cd86182378a951dad8f63f4e820a2f5433df5ce797500fb4afeb494ae17ea34d950c94ef5780a73250abbb24e362c414abbbb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6211489319811a2a09379f3f65850ba7d4614fbd50f2f478f18a118e4a1c0e867429705fc36ce788ac55b2b1b85f6890f087f29896a0a1ba94ade13c8436f289de046853cc8b208f07659513059199dd2e86572418d75ae42ab474d619a8fb652b6c2d732b97aed180d6d5a96747deaab9f4154affcf83a73749743af4bce7c4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf54e6bfefe85dbf51657d7d2afab5077bbf343f40776379ce6e447a8157ee8bcbbae0b8a629509433ba23c2ab886b322a11eb150964a6f1c22910a97116fd961ff0e1f7330397da2808c8b4345faef872b8fd437c7b32d25f05e95bf4d76bb526750fefe55c19d2170d8aefb7cfd8d61513c63039eee026cbcef94ccc8556894;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h46060781298c12ed91f26fa014ce62a45dbf9c184befbaebd26662ef77dcfea7bccf190476ed8edaf20dc29bdb5864d92fe057225cadc68c58c2df136722fc5c03180d741df081fdbfdff430e3471c4255958b3a83f90808f83079483cebf64fb8fcc6d2f6a49996b6d74256b478194000d94edf38cfe529ab9cb9e650411b04;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8027bff412a0130843d7bba7edd78f02602539316dacbe27b0ed29030eaa0a96ba556e9ab0ee1ec40599f1e8e734666bacbc182191cdeb16fc059d3b00f5a9681f2f959bcc6bf5f108aab28525b4063a98e7361b05680a553a662cca1f930a1ffc906fd5b9c55561400dab9486a7e57d322502091a16727dcdffb21a5ee02b30;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hddf5a85e2cb510fc6332ddd6ef36df8e7bf95783c0c011883838ce0a341bef4191a470a9d580d83e18b363d81fbf84e85dd172e6b443ae178ce3fd468f082b8680126176775c5b07dc0e589d00bbcf0fffe6aa46b7019aacf8e84d2fe38d3992a76f87122593ad4d21256108a6ab06c88291076e7d0dbf1efaec3cc6540c6992;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8862dd08471cba29a461f7a586922b2be92c357dd2709a7e5b435392b5262fe600bdb8ffa8d35eaffe264ca44767abc0eb19cb4367bb823c5e18fb28f19b61b5198055bc12dcb52b0067f45a550e9c05577024ca97c92fc16d5eb60c7bebbfb5446411965fcee90562278dab8be1107bc2fa5a12308f96b844ffe83bf8feabb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd9f451a2f5a7d3d5ba7b87d778a0c805f67ec35f9083225a502d7efa2f9890a630f47781145dbd33d45203de74adf0fc036e3a5881b2aab677c0467cef96bb6515fcc7df3653ea7ab0c522b62c4bc4fad30bbc624bfde34c427036d9ea8810726ef5942c2381e1a08d842443d16fe0d766f2a7e4cbc015cb5fa8652bebb9b11;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc6e93eb1d9c23c67b7c26de5b3a3ff40371e622062d7a282df3f062897e01f92411013ae47e61f81a3b6f4e67beed98c2af70dfe94ceddd0da70cb4ded6a18e7875c814c3bbc62dce24d35329170f2aff52850d95b2c3f09e828e74ef384461ec087d44cb233dfc48a902f8c4bba0fa06db905de3729a34f1d098b3b8bb92fba;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h26876dac0ee45b323b2b7c98e15b15fa30cc7e2d03ae7655bfd5401aca1e91dfcb74d58c3fbf79f37ead5f8e43c4073ffa48d5cc98546757f135e86864924b071b1c06dc05863eef10fb37b1d949f76f26def318b1a0a17fcc681fdce910f71d89cf7914e3730af2fc0a7b1f14945b80d108956c8b1b0effbe00210a10289e96;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h447f4e8cd05f8e75f93d0847d5d78ab350b0ebb63cf7d8dc3fcb7c0a6e1ba44564f72eaf0dbc11324cbeea7de8434a7c191ab3e28ad3ad39e43ba60303759f38d7ab69f8374f1fae4ab94c2ccb84c6ea1608d9454a91a581702def047a3df011061dfc63c8a9b3ba6e023ac491bec9b6cb5c5b8eb1cf37da1fe49d9878357433;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3b15899ba9ab86b37e641e998ed9f73adb8cef830d111eb9d98a5d83f7c47e37d0475b3cd17e58e3913f85497edac0de67c9685e47ad6902ae311765d8ba243aa2a1bcc8e3a66fce6a9355a4417c152f5cf1bab7078ccd8d26bc458d1dbf088f8aff43ec63fc80242a3636d1d8f6b3944e7c6959f08f72524682986e79daa31;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h851f0fefbb0a8903a3d2d9294686f035a8b96bc11549acd0a43d55241c7e4949ee50c03006f07571ed63e98ab572207b2af3fdc275c786972672e3017460e3ba8888eb7f69a8485438421369462be565ecca424a5aca0404ce8b2f3e84e50c846d17aa9f2ac168b579f97a555aaa81a093db2bb2f3bdecc9971de2a96418e085;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h62162f25a631379234a04affa194174204f2ebca05b3e625b0abcb7a6cd10db6a122840fd02da53b3cd9c83c9040eac58abe5a151a7b61efc60472af0f763262156baa98621ea843d165aa56e31c9216d337ecd5f14eecab3c05ba4537b0399f2a2ff80c5862e73b39f725c4139fb6e0afe6a3629368d99a6a9cf376a6c6036a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13c534cfb257294dee5146d298788a3e057c193b17a00913ee308cad74c1450d08a6212f2808de452f2e63e675563e413d94b930abb9e9457da4eab53bb238d3e70dd4605081d016925d66070fa7e8af9398a5dcb23d100e152d0a5eb309aaa2712c955400e906113acad8543785ec0b3269c546f85d460f4ed47fb327ffe605;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb391cce5b076d70d7ebf096d90be36772a4763b358a44b3fdef2bf906e291fb8e7cb2d0f5e8d81d9c18e2713802e2791563cd6557d5817caced4b6f9faaa638fd1d6c9fe9d7e46a25b1af6a3eacb2d09bca7949039c83e39e49fa0f082ab8378fb795c8ee36ac58ac55c48c80ce221f589d6be03e7c8912ef068397bf9a2280a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf69d8554c60a545d0945ea821205b11da10074f02be1a1d865b7cebd5e6261a445d55c2d5815c35b2e1816afaa0d717fd73d0142a0d8aa9dbb00e6a1a3c350ddba7f0fa85f172c60aef4339f82781e573455b8714b22579efba271de37dc76c84f63b8f6e463a91818f2466ae4a03d24fd2a49b48d2f6e531961a69316aa88d8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h198091715f92b05cc748f9b4d75e299bdf1a2c1c3baa66984da4d407826b315a6989a718c09db1b6ee74586973bae17d8a83504e1c1f30c1cbea266b02d7ddc1a2ea15323523c9c72c14f65f7fb287efd18683e3eb542b2424e172d7d7825c25a62564dc68f01a3a09f9da7a946b43c1ded19e62596efb281b4c6007f8348fce;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h463ce6cb1613828a8ca9c616e124301f5c0a319799c4e590ede9fea1833b5e747b11ca474096d15202b9ecc7a0a13021e4142eb982226797a78400d28da503c5d03d34d167b8241e71e53af328203702c418e100ea61089637de960c25ebc4a6c3bf06602d7ba2fb505fb09bd43c4a90d9d8f685f25c15b76b0a74820d5a5d45;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he3eeec28eb786cdde14312c6bbcfc08af3c61bb58516502fa936e65011b5835af099fb881135eaed9a020c0af832d0413e09366d81d79f1de7c3740913fb062550f552ec61f56e7a3d3ea88c52ee42824e7891867dcdb93e27c34ab071401634a2dca6d50cb5133ca5fe0369ffb3332942113a77bbc183f4be6d3d2b24bc1ab6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h219a6169ad4f3d66c8f2d6896a7a6308782902aeedf4c56f0d30c014e38c3cefe9284a06dfa056f583784a53ebd0aad8422778ee9be7859d03c858c37854f96d822a02b7665f1808eef3ad6825442d9b0da54b99819f47a6752c6cd60fde9dcf1c29c06ea563dde3e8f0998792db5bf60d2d582c5c5433f96582f121866e2de;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4e74f2554e0e23461cd9abf7bb51b98b282de898aaaeef6acd6e0241a86e6f46fb9910e0e6f0ddbf3aaf605757625e1c14bd66bff6d338f866ed6694386a8fec1666767b1df04dfbd02a9ed03dfd5e0303ef7902899d690207480729e44444be5557776b4e407fdb10e0e95058ad3dd1aa5caa078643ae84ddb4f3751e2078f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a0fc1df1e19850b60b5609ff628083834185cdb3bdbd63ebc8cbc3499bd586ab123976f14229044850043337723c8b3ea7b89fe0da44686453a8b6bb79e47c4a8ad2d4a29938283f2d77d91de6c976147c563077db19eb7b4b33028733fb5a406aaece94a4a74e00efd13e6c2f00ed05b79d8d2a9aa939ee5024450aa9d78b2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h72c70505d983977a242a580d2c93cf2ff0fd88806679a7398205a8795175adba16d4826db7b8983c1bfa90c2b6b8b0c3db704dfbfead6a9455d05f633fca2b4bdb9cc430212ead2226b4cc3bcba35ad8d10cc87f49fb44b85ec1fee457ca29070382e94d51ac2b8055f89ef543f6d91e1d9c811b5d3c1467f21203f3facb24a7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9ee86798bbe9459f6ecdf3072c2902b40c643ec432db64ae4a6a179bc4041b95216320e88b4f07ebe42f902bf430bbe99f1ecb940160119c831f0e4e5fbf2dd4d04cd2cd48cd68f65cfc565bdc4aee8beff59711f2d357d4ab34948de247f4aaaa49b66c5da0174256b0ec9f43da0976afbf154650e4a681cf3ace9523a64461;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc1231f4a49f5da97999bcfd3a9726d088860581851072b00cce265ee4b9ee0ba296b8b448cbb015760d14edc7b4dbb5bc6deecb37368ce72a9cd34f8709a182f23ac191702636bdcc52e0929b8a787713680f93216bdda54aafddfdb6d819cacc293acc46af20099140bcfa945d74fe50327579e24f2b79fc9aa0bda3af607cb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9760bc6c7d2fbda5f2198d114e75ee53049ca5325322f8fae0a905bc2fad979c911025d69f9c9d346a3439961d51498696daf2005f60468b319671a18769a7b304933b16e40a09fb2c230743d879d558da6eb62b906f32f3b92ef7b14593aaeae132e43ebb98a901e4e2cdff82a9994b49fa4ff19bcc493f9247c309c462b9ea;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc4118b9d9b66b84cd615978fda102bd78b0ef4a11a21b97be6bf139044d7db1351b04849e79c299aa40ebf797cd2a05ca16cea009f1b95955d057f33f4c0c5236af40670d49076808d9dc3362f0b90b5c11e66a6ac880da52c4dd8601ae3536124d96da4abb9d0db9b699e2315156c0a84dfc9a0b857711332ea03637e35bd62;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha3cb740e7057b5a50739d89ee6d11c3be7feb33c1d32de5e100e43e3b19631823ec83124aad7b0de42e6a19e39e277a6119d34904639456f590c2a2f334c930935866d7b25c7d7fe6c8beae1996610a6ba4c2cac08d8fe18259d85b0421616902f852c201118243a42674abc30f18308afd70593d6ebedb666477e745ab2357d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d7e2d01aa9c95cceda52a507c20d848866af284ae7373520edb59dba1ce95188631a4cba97973b4367dccb55aca53d170bb602016dfe8401a3809fe89add316623d4d3714d1cae1eadc0bea285c44f24757ca878b30aa37296e5b240c967fb221796dd07705bd63fd646bd1813a2cd6027b6bcf551da2ee0b0e2bd79b889f82;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8431082d53a888021e84435b11efd2f932dacf006019add3bb7c6f4d59f698d048829bfca4a103eabcb2c15afd6c0af33827772212bdb298a68266f29500702db29a618a0b484154313433d8d2691f9b905c64be5414736897660bd69d24b7f3bc46e95c61caa17b01e39184b3f440bd75d32fc7d47603becf6d08c479f31e52;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc5e0235a60c70ea2e31706dd710a19acd597b1877801dd2b585a9a21cdac6a0a3e9de24ce35c67a34bde076fd8a6bf66cef9edbe0a2bffa371227f65d7ffd611152ec83102215594669afd91ce1477682e7578003dd8fef1ec71005f515cba537a077a567a6223056b13cb49ce2aa8748b97e134932b47ee5e3bcdaed9322ab7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6f169aa61e77a7303c55c5cb405f2330d8a9addf6b5fe015cc2a3c9675e0dd349a308ee73556ecb8df7fc6a006145e13f852d758ccb80af5e0996f960af7ca0d4fa9a3aaa7aae8f1215c24767e91c0fd161f503e149347256118c1933414875f82fde2ffbc1f2181147d9d0c55f8cd8ad09532fcfec218d151f2a3bb8857a5c7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdee8488d95b37c08299677484ccc884b9aed608afda581a52e6f1152f92175ae8cea18937e4fea7cfe56469f80e7b4e1641a284b3a3269e83346131dda9a6aa8ebdf98bd9a6a3e7c2f003cb4bc7c285027fbc6dd49e9093c3a52f28f9b6f34304099a932761d5acfc78d1a4c7a1b1e0455bb8e876298a495314f99ee5f184a22;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd966d612e48caecc8a7bd1fc551474874ecfab8bbbb1277613167edca3742ec024d8452ca3ce5e8fd4bf48ba4d366c0b5f52e8b249444640387e61a04396b0e7e5d02307305469a937db2be574be449c16b34f67d6a6ba2c3a700afbe7116e7f31ea2e0e3a65f394d390a78b92489d7b3ea6072b82bed9baca1915809f59f59;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf58d63fb402d5796c383aa9eb8e1840521899acc714588429109e962c9543fa60f325b919c164554722ba1d4adfaf1bb6747c0b2721d399c7b8557d59a71afb61812c6daf1980a85b1077de7de5605b6e428c70a18e33ae1ab21ed446a4fb5e9ec7b99913f06589728b608a1f185bb3c0c95b7a784e6dfc55507adca42f47574;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h40bba8f4faf23d89b9a5d3a817c016486d2c6634549445fdf4532cea087f3a8495c75e40b7bc7cc390fb201cb0d4fef4172d6e2441199d9c131eeeb9935102c863ce063c94860311a2cab8fb1bd8adf538ab0cd73ec8f3f635caebfeb91e7cedca60763b957e586d328a86426e216ecc12e5bed46860ac4bf3c52f82b2c97231;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h18f2283609bcf0c2fc1d35f0a216d32939075000637c93ab6bc54442c5073d34ee9baf947b7a743799b9e110aeafb7597b9e9d744b70258ce7a0a58cea1872c6ed276d52937a513fc3c4abfa89a0c5e88004228041fbd7be7a0899c2a9316bacaa5c1d0b754f7b28b8e58b06f02b2e94791e16a9eb558d5fc483e82a46ed7342;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd964789835fd2e557a2987fdf57ae186102913789fe2b4e90315cfae8cb07d9af1054ca1de160139077183584f4c87bda162c9ed3986e14e6ebec9011d538586187117330e56ca3fa9553493eb1bb9ddf0722d6655f415075e018dbe404749f5d1433fa2956b975cb05b4f420473475d8eeb1e5a78a05814a75bdf9467a6aa07;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha87c16638090b7cb447c6a6219fa162cc89c5e2535e2548dff378c49682ba78ce6a06b6fe163349cb11e832b54a37943154c051e2a05291753a87e04f574dafb756b99b5baa635a7ea915d454c67bd72a838dbb56483d09e71fd06a4f6ebad8fad33007622e218b6ce3fed2bcb9b364eb096cf2d80e00684e4921a42b1eb6941;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1f21704d8d8baa0511d594642f78e03d06cd53da3ecc2d5e9950274963047c69779f4ef8d27c8a1b473e1093051d3eff0715fea87616c7153f460c45d7ca15a5541260412325e18670ec4fd2c233af1b7b9efadb244a1f347adf9a9f11694e5d41ec9706bc7ebcb5a5f5fb7baafa62b8d83a9dc394156ea1d2fc6263bb798e32;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h75f92daa9932a539076af26aa98dc7ae3b9e2a8a46f3c200c2bb79115b74b405ff92e82e2674eec4aabe91633d1360c139668e943d78d9346a1fda6f8877b2adb3948a9c65ce4d84ccdc519101684d2c86d54da4d228f8dec76e28dc2bc3d89e0cdb47f316f0db60fa395d2da8b0ecd20337a342d837f7d80e0c9f53485f709a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5fa4d48eb0a86990c16aecd560ab5e2b57b3876d625a72f4c04fccd2902a2c5aaac6ac30827db6a0e3510ce7018d5704081d71a9ea47cc64aa07b9bcd7195b4f2065e043959b76e3f277ff845b78f09d5fb82d63be03366d35dff4d7992ad4f6fe7e9d963eb47eb6c6c006dd39d7a7bfe9491bca93eea4a3dea2ff42954deceb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcb8f670097188a9e5575cdc71d52ba0d7958cf81c99e684c8a6bf7db376fe0618c1eda019d5a81480095c677a72dc33733764924c63d1d03d03e10673958dc04277b3f6a5db1116e0d17ab0aaa8d49b5727af3c11983f32078ce71ae7b4e981817d05e36f420b3164653ca9f5c580e0b80ab00978683ab6645e94b53ced5a2fc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf7546b3705da946aa78afc8279cbd90c753de47343f3896979cc7f7ebff2625afdb5bb67e60f147e0c8c190c8caa8108915ccb0a21186d23cec38eebcc1619f39d41e83baaf9ae033c6098085806c7c1b8bae4afebb7370c403ebc53c3035cee0a35c1afaafe8895966f8d915f3646bf98f9a90ca53ac9b3634609298117153a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7303e486df2eb94734db04c805bd4e9b3d681d2a6eb6e842203f24828d1aeea032c55a157536c999a778be8d61edc4fcdc5a7f7123086b876930353941d494706e972b75029d3492bd58605a835cf97c24d8660c63764aa252d8b2e48be57547f385aabb02758f7741cf3454c35fbf687147790ef5a1b4eb9a83bae8000c365b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha5f73aa2089a8687a7b84e5a7a2b752985d3b2165c828ecd189f5a588d6b00ef37b6094b33194054c60bae88c632dbf2f554ec0ef6b328830ac8704dbb707a3a023cdf7a0fae23a8036bc5b380e1f7928ed698da24608e69cb43e84a1a5c826546d46c46aae42889dfb8c713de0e8d0aeacde2264f25f62c0da7fe7704f4e939;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he566b4a50239cb8ca3105446937b11c3cd054fe6400b50aaa6af439352b7edb6c72fbad549cf755019cb81c462ccd8dc00844cf2210933c6afab04882dae112d1a1256236aa04bb737499169157387ed3e0ba93081dfe2f8bab053f304a2404ef90c7cbf401f0104af33acfd66a6d33ff22f18a833f14cc3b7e001df7065c09e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13c3758cb8d541f135f16456b6fb5c86e005b9608dbcb34dc1b36b87549df0e9838ad9bc8db30dcae86291f0b1fed53bb96b9ea3ff0a338f1e5998de40bfa93a28934e7aad597dc5713ca43331a5210b7c006e7009a08de0b6b9af8c3b4ad097acb0c56ff4757798f394935c201a03ea1cc860a12cb4e300e3b7527d9d9a2169;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4660ca231927b3643fcd29aad7201b4b5fe89eecdb8f48fadfc7a8547bd530b8dc8428aa31fd50548aa272e807c8dc4266defa8d9eccd2cd9786e2c4a384e7d0078899934c4bbfbcc95b577d5250274b2db391fffe8cb32f9d16481de916a6886898e43deb1bac2505536b7387f9d2ecf11558f4efaaccf5747ce2c52473321d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h193f4e5d0eef3295d318ebb7ad0ca58ae0ce28d2319b9af0de1ec584568db7e0855051fe7dccf7246602287400a59cdf4e972fa0748c339a81b06499baa94a2121ebe847265b3dbb237f76d7be8361150bdfd3fc0ba1bbe5101b2adf4fbffef9f796b29732e60297bcd36c03b1944dcd461c602092cbfa4cba2c182494ece0af;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h747fe88aaaf07cf3f06485d139c917fdb059ef7eb269225341c063e3b474db2187031480080e3ccc2f2cc2a52e1aadf1efbd12a196c38b87587aa1cbfe66340a8506c1047a96325dca7c145bb908f0229714864773f65956c9f6104fe485795d0a037e8f9792de2ca5276e82efdd1d5caf85c71122686f7b173e31b8be933e40;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc7785896862c17ee1aa55d33d3066c775da737ff9c82059198214f525e39507c2ecc892b94f7e14b9f92718afd11a333e9b97f5c7cd17ffbf90795112b69e97eee29f3364e528eec6cbb3971ae01d59eb973c4ce7b25ad248846a6793a90f72e89f8c3cdcf6b5736934be18762257c11df4f134469ff845b3e5771b5c12c716b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he556e9c5c82e570a3ec4383b5ab18078bde7933ffd7acb8ec19f36ca2eb12c9d995c6e36fd4382c3b506988a6f913b4bedf6546a1cf0cf45839e3dd674e6e347ed9b8e81232337f61770eb039b96fdbd7fd7bb06c7258fd82aa337185a79781db1689465509d9b50ec4bf8a984c57e638d3fbc48e9fcf9fe25edc43463bc622f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97e86f8bc78691a0b242f9eb8189ad4a2e0caf2cd6a4154a932810a217f3d9d16ac98b0b9bac3975d16706f458d0e7d05c1007ec2ecd9f5526fc2a57030babef769a276fdfbf3c6cddca3a6b93d79cb80aa3621642826523a79b940d2cc1a7160b70af39af5ff73b9ee64a4e019efd7dea0c1f5bd9c16b722766c49d2cff8cea;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h376807054c215383e6521a46e7512ed055adf52163f81c0f2a403684051bfd604c981478cf06dedbdfe87e2e2171279ca9335a0af6e027febb29f79922fab89e5c693d017c86a9e78214db100df0221b1b791578fdb739327d470279832f2100effa634292cb1147799cfeb61105b649e0a85627deed2ef475171e8735328b6d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1cf995f75c99d104a1b65d81fc81d5d3a609fc1838310758e9ee65d70d4d316a41b18936517ad8d2692a4cfa8bdfb1e892e6f218017627d1bd9a79bb8d440e5ffdfc341f72f0ee866126294c8fa9d5142a6cff9dd1750a1231e829b1bb2b828f4662a8ecacde37b0bc68e865d63daedf52e5576f961f2b1eb94a390ac96e0eaa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9d828468ced0babecfe6b991beae2a09b5b3c516b42a2e4db0c1378c364841bc05c87d452ef8df59f0b478cfc1f7083f151fcf74f0ca0b82dccebd914f34dce1708fbb8e81ea7da89611524f453d8c7375fbd1b811e759542bcf82aa6962e515c7edee153c53a5faad34841dade683a5c0ce57a1c062d55311757c35c2ade5e6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b3a9173f299b21f7e6545673c87ef9a5432189cf4751550f509fa50137ffdebf01abfe1d8bf1dff87a613193592ab167a841f741fd95247056e0c824659864a903939bf9d360c0f9f47a8713043d5b5e299463befd4697f948d628f3511b4a0e48482a611ae410f21d372db42612683f4ed89ed7f182f7fd7ac454d1ab4d7b8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfca11f48547308836bd5ed7a2368a34f548ef64b88b22df160d283ed56ade799b310a719e099f43f2ba5a1ede2de1c60c0ca6bebef3d025fbf1bf52e1eb546295a1ff03787273697d9374450aa4f6cbff33f7589329646e9365c5111cc9d0b37d747fb10e6b228c701cb35e66a8d824175764977e819d056688a60a20dfe552b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6faa108edf3a5840d2ce0e10376fd006379ac4a9c3240c68f2bb71fdba8835953033e4f24637a53c39bbe1eddcc466700cd59bf79473aa003d6f038b2c49082dc3c6e3cebda3928ff52d8140c3a51cf1853b2d15780997b911c0987333dc2a16c09bbdc80b7f16b6f1e16a4f51682d2d817033d0ca4dfa76fddde2acc0de624e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d5bec96cc159ec3aeea4710b29789a8f220f3058bae1d92484022da0c49937e38e360173dfb17654bdb70d05e71425f026e729d7ac095133362e65504e0b97f6f4bf3f9d364f25e31f52ed903f1357e50a467a3430a672ddcccbf3fdff86c0da6e8ee98110e03f3668e8e5ca067f9f09d810baf271c3348e40e930046f56de8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4bd7dc1ae39f15b7b11fb614cef43473bd65d10ad51ac6f9bee4bfb6ce4ecc085f995c4e77a8048ee99d0380247a76dcb16f6ec0a65fa4c79be47f9ab41f4723ad42580dd282662de904530a4d549acca1130185d4d9a88c001376456e13a57d72bc478598a9dc4ce081a5e61279f39706bcb3c74ce41031640f839db2c9341f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h45ff379bc2d5dacc85bb30f4ef7a73075b867ac9f173a64a1ecf8b7968b29a9ad8961aeea08b699794bc34e0d37eec7c4d2b51aef3fe6aef43eeb1daca7f8fdfa661f54357fca15a5a42aea0e3391bf5da1b530546ee01b344d8018424ada3e2f3876e57593aa74adcb39972fed3b025ed1b5111a48382307aa5536984b142e7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hff7fe8ecc6fde917868e13eb7b0f9da121689d28d1d74894076bcb70b0a53892a833c38e67abef8d373dd90bbf5ef5624c90f36ca5de86d0f06930b62b3897d1ada8ac82f4ccb8772cd54b13bb493377e0b49078ba3926512d10c605865450461ac8096df278533fe886fcb1761fda8533daec2adf6329559e045eb26c316700;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3dc305e1042cbca2aad18e3b6643815abc8bacf4ed93e28dd71e66daa38f19ea02ac730b65a125fa79ffac6b6ac8e198fb595d516527ecf92df4386e9012132dbab8beb95076715fd9550acb9d9e703c5206ca8f90264b26b59b10161caef799a0227f22bc78d0d4496fad6c6e56d8d6df06bf85497b5b4913434aa261268ccf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6fda25fbb250a773592855912406210fe4fa3bda1720c3351c4470efed98449978c7e98bc0693cd4cd9b5ec555a5b048acffda8ebb4a395d99cd0286e17bad524effa65d209194529f7079dce7091a33ae05bbb8e0022d2c7b732463d2f38c8ba158ef441bbb07f4f9e8eca429c7de502c56cd80073e15dca09c5a204a7b6a51;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8795902d614de5dbe014d7062eabf8d892982933ef2bdcf3a272241bd7fbef3c7700bf51c451fccbe9df929abf48a7c5a6b40645446263bdb788dc64e0809519fdbcfed53de324bc54d21f8c60f65e106002f5b642c5973eff0c677f445dbdb1e2dda1b8afcc0bf1bca848fca3ebf66711c5f6d43353ebdddc60357e736b924f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf2542bd2e6d06e54cc276a540517463859301ea367bb22d84dc19c23484f8d24dad14f8969b35c07674027ff0a92bb0fa44e28c05002686947eb899e8b1aafd99e4c65f6a0a27d81a59bbd178fdbcd5f3c3692abc5c7cb5e89a983b8ff3a42efa406dcc6be9a5df95fa8113ab9409cf76cd127698891bc04508b2788ec326ec;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b1f76cd9314af0e1447ad41a3098ac8368d66fd3d03ae652aa51407f3a5b2c37a28027cb667a151119716100c8b2277aee534a427b440880dab808289cf99b2abd9612748130d6b9f48b9cd1ca67de9ecda44cce04325e9e80ea0848e2eef672470cb8d075263390ec7f53526997ff34703dc465ac0a4d6fdcc7e886a52f4d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbc0b4431425dc075edd406ec0e4181a18fb10676e317924e856760645b0fe89177afa8ee3a8cea8f262b96fe6898a02d140b006ac46efe00d9adeaa2ff8be76e9e912b39061d023fb1316689c77cbdabcc305226ad353316333ce9b26e0c3be96f80df308e137ed9a98b7e49fbdbd4879181bad44e988503d00a3061a024ca5f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haedef61535bf44f7f5a4371acef1d0b164f8ae360f53b3f8ee3643975877866b92223c728637b47da8a99a2b77a466641638377348e973d3dfe7a5a09ab5a54bc699ee13c1147dbad9028a98fd0342d31379815d01f8c22fed3ca821070fbfaf89c11aa78e8f67194688408604cca5fd2d04b9ee856de28bfc4dcb12d054857d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h455bc3f19d9867da901e8b99108f34e4225dbe645698e424971c41228329a809023e00923191d4c4d5f67533892ebcfc170c343dac10ebe0a51c9338dd504b2da53a56ecee3e4f07ee31e8286bc771b0ccf42456084fdb839ea17f2e596d286129c071234b67f1c4c97706b84d21bbacb83aa572ae0a428c1cc8e3d64bf27c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb8cc69982e2595d57a2a1578bbfc99278e261fce01357643abde115c9d860b27a1cb627cca5fc55884482512156ef669f2da8838a94673d44e382de7e5b76cbc0fe941ef5783aec212a346e1ccd9569016a47855abf3709a96228c986a6269a25c78f79a142b1f8890a7709204f820be49c8e5bb7072215e24074adc89f4c6c6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haccac437c8efee826dd7c79ee4391eb37c2d79cad1ce3266e4f4245c4b5df03cb9a3d73c7b39b4e6137470509263aa493d0e9feb9021d6cab6bf101efbff706bd421df366dde4ca6ea5ea6be57e3b97b3ef589511c39c5b137b2566cadd09236399e108b0a0e3addb57d534531efb665a3ecc470168be6968c59a6ac5c589e46;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb13e7341d19735c5653d68a616c90c0b0ea9ee56ce2f6948b28839c38363cf31e4e9e1e5337d9ede9f87d962f1938e2080669caf61941948be1ff9ab0432b3e4613b011a8fa10930f7bc5a0537fd73f1cec00de1225795a74fc00c25209bad87080724ad73a4488669991b9f78a84977b5c3f34023d82ebbdbccf6bace51856b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h23825925e29ee174920de8bb83eb7c97d8ffa251196285e69c5387314f1e99ed2c9ed7f890b1190018b4f6264a5fe53731bd4104bb8c8e39eb3f87f54e95abf977fe529a5c3ac136907594bcf45cb391df39defdbf22cb1ac4a6f52f8c3ecaad28a3fcab98328b48a1816848e76ce7afa9c1762609aa01c220c60b75394aaa88;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f80308fcf97597f35f7d4412bd9c53884c97dd6fbf10d0887accccad234bcb8de1b283e0b9847fff77f3902b7dac7ac62fd7921c74d7a13be1eea8929d9e766af4a9e6868353d46fd4069b980bdaf2d5ce2e5e2bbb296c23641c8d6c12773857e6a7efadbcc4cf25066b911deebc24c9920b9e4dfc947cf5f811ca0671a061;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed2830a2ec1cc3318f0c25a5253e66c98b56585982dd367bac241190549d6575b80eeee5c09cb9f62a38344198d5802b53d476d37c87f2ae080478dd2e25bb8e117d096dae99257bbcacd4139ac51e9faf6f6b8a7639277b2654df107ba5fabf5feaa3263d3618bbd748e2152a0442149861fb11f500b1959e047892ef789442;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7f07dd298d247d4680f3122d52908a89bae0e405322d9818f9b80c64c66c7136f3a40db0380d20f965a393436912093f706fe48dbe491a728595683f67e518ce6d3ab39a31673d38509e3d3b9bcdfe1139bd7be4f61220aacfbfc58bab8f7694117004285ba2df439d483d4dedcff0fa55bccbb6ff1548da998b05a4077892ac;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h813be1dc2f0a08312bb2545938115276f3c5748db1cbf44cc612b9268781c3219bfb41fe3f59ce6672ba5891e6ec1e9065be1647405b0da8c3ecfb1df72c6558a31ac0e3d4086148d875e9343cc9425b2a5901ffc99b1c9cbb9404a18d0ad7be7bf110f27ca8ddeb06e40e348d01a34d361e2efad723f74dba9f5ee84b356912;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2adec5bfaf4b760876650677cea1de74e9ce62ff52ca1dbc4df28bcf29716939fb0f03c091eefb33f41ce8572547375394d9f775878544975ec734b21ddbcc4873197ea0ed1ad793078c16e99efac25b3925888cf24337b94ed13011b3ca27abdca67e2d967bc934d2d60dddd6fe73fb29d3f6e47d55f06ffff1b7c6a135ba5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdd18ac57b6c410094381b0416b1c10a4c7cf72c7503e8d61524ef258e341a8fa8e59fde9d950900bb2c93dbca69e493d292730102b391d2c8617399d41e2c3fce9703ac442ba4a48189d58eed1942c7ce49a1c3e51e7fc1506ffe63b2de7f20e1c5be1156df9526c7aa5f7e734f27751289c6473415c8c4cd256a736aa870c3f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h99aaf7b2410a2bf04bf03fbc3259b1ccbefb9f18cdf0f6d39fa2c13acc7494076a0debf157a76bcd25e79459e3b6e70b102d3d424812729515be1168a6bd479327a7cd5d50c3452045b289a6473315f6b4f02ced3f7fa06e59857365486094b16786a791d5fc8d93ac9ba70917607b1e7bc7c5326632c8c49ca02c5397cae6c0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf0e7f7bb4af6b4901a01f31fe09ba054ed6e7d523f796ff633cdb9233998c9862e94e27a7ff4217d424d5f7294bc123e149b7c66d2b54c7d7fa11c6cfe503cd50af8bd1672741bd89bc90e625657d84a969ae2a14d21202926990188503493581a81b5ecc3cfbbc2704f3d5e1983fb22c4c0711d6d8bd6877ede88a74dc5d376;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9653482630a3c6b8b6b93478c9fc9cb8861e0d7bcb5ecf6e68662f2484a22124014314ff52d00ea6d20e555d7fca065c081a7b7c90deb5c6735f6b16a3dd3ab0f54d8e9010cb23c806d6607ec725430dd802cca5da3bec78ebd49d7366d4238b9e5730e34112469dec7673555bc87d3e78df7ef009a36f0dd9c7bd99ec820871;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9bc0e89c5c74049e4f61cbd13253460861ac98c094b201e531aa4c9428a3f98b2eebd55565246d862bb385c768f6808a0c9b9582be742801b3c6ef8b547475a678698d3bc44f361a10bf5b7e440ab9d042378bc6df053d36fed9a5f190646c3f5479d0ed5e96331fe2cdc4ea4f3d592db54bec0023b39df6269daa105af83bfc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he93a39cff6b771ed64e7a6bd0be5ef14166df98ed530a4caeca0fb681dde2be23ad4745333e07c439289025ce6239068d0cceb6911b3421b8930cc4d8c3e2dc4abc520045fda4c21cdeac87523e522ca44b3a3d8fd1ced72b862cf83ecf33110eeadaf61393d2b0f909b80ac469db4b3919f8231bdd265a81b599d8098a454a9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h572743e6b7378aae0b84d519d51f555fd1c01d0335052ec9d57409a81bad641ce9f87c33302c554c6d5ac43fa511b12702c6aabf250f2ee9f0f415cbec47b97a50046362eef04a66e352f922dae62a4c421db2fb5f02450429a949095d7d907bc8c425e06ff35962c5e5577d2ec807c8f457b1471ad87975720e7fd480a9cd66;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h91d160157b3ec74cce03bbed713cd904ebcba26eb092daf50f3ad8fb64d4317c8fe06f0049f4f03b5a0a3af1888ddbffd584eb5cf73844acf29d0bf46e01926ff44019bd7f085f6e51e6e02f541fcdebf9cbd2ec238eafaac1eaa9ea08ab02cb067bbcc1c29fd87fb6be5fdefcfa8f423d281400588f8bf20bdf1858c7ecb723;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha417eb9acd76344c229dbfc469f78eae4d166fd30c0d28b9b635ce18f2ff3f3e0aca9a0ed7ae9d717ee3981c1a35ce9ffda7d37162c252cc8cbb7270ad8f7762a136592c049d5dbd1ca8809863b7d69935a376cb9b3a1784ec68d7cb89fa5d8c3ca10f2cf339df33ef5b1f2148627346fed8ab6193dfd7ca0de136eb0e6f897e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb005ebe64cecdf8784282613cc03a2d9d281bab96d43d37d3755d0e7bc732b301a1a51975c1a8b9f8cb7341d2fc76e6a16ab83f3abf4c3416f8fa27a391a6d23c49cbbc15341795946751dd6093c88707bb1e8d2bc63a992e6ecf755010f0800f59bf2ce2bf75424ed4fe017de30687737af65b5dd61ff2cc1da4b05236b9cdd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha6defc02f7df648da4253ead37466a1b8cae82932111c0c1fdeb8fc0872e35f13305d465d88065fa89d120a404d0b293c11be905ef5920b9006457573af828f7c54a9f73821a02032898c54299e1c8c7bca13fe7040432751b3f6630387db0193acdee7d3575ab940e10141a310502fd23d034fce7ecb9941b69a2cb2dc00e4f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc4c86e073aa4485fd4210ade0a0f4051d7af2cedd6df9d94c62915155051cbe2ffff8c970abf8e947235f95a6d96473dd745f31c5d0f6d5afcb73825c572765b8272f6b5cb1053b0089b4f085f75453493f006f83ef6f6881bda39b0b46ae12c630ef8785c75c5681f1190fedae5e208a211942d3d0279dac9a7e92b8e5616ce;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19818aa082707a8b20cd23c1c49e748bbc50fa8a876a832ca6bfa8eacc76ebcf036ca2cdaed9fb8416e077240de0a270ec0dc294b0bbcc2751adde19947aebcf3945648620bf95626cfc49789db6de8bfa6629eed0b85bf01ed646b7f9582c54937e53d5da14d19b28e870f996e70b0b1b6b40d6dc8a54005d67174c8221d846;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6d5c5d2ea9d1cd1c7955cc731e2d44f66b4b33aa9a88ba8d5ad9749cb8b240d584ae93f29f36ce578a6924d96a3ca7e28adaab9a54cb641bcf48f9e5fe7531543001f232744f07011f12774f92b571fd2cb029174c28bb80ab5234d01b8d36ec6b25ee4cdbc2bcf7d47399dd6071ce34f45aa94188d5a3d6c1db4e349dd4d82f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3d38349bf6c6cb233b3f5be16d51b034ee8281e6d04aae420373667e6b5a520f04d0af2aa14e6d3a39a8486745e13e8443419e46c5202d53b480a1a9959a28a9308f517d9ab836de02fe0889a31fd8f6a09c3134858f523ba4a677539c2fb3a13eec637295cb6dd8b2a3f78be56377db5dfcb547ce5d361f27b8e79752adb54;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha09c24246b3a8bf94ed99997e4f6233d06fd1f0a23f22d63b65679c8fceed25fac293c0ff0816809a8497eadd219f87a4c6171ca76ac704416939bc52d15fbed105df9f737843c4a2105580966189c6ddfbf79fc1b021f9fb812aa246846246819a3155f6bca72d406a8dfa8d0987406f29ff3b0e7eb292fb61b9d301086471a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h233dfd9cdacb30e2c0939c7bac0b1a79d844ed4f848c050cf59cd420368dfc031b716e725b4790aa8e22a1f786dd55de7899ae564e8c9ef2b0789c3f121a517f708db1332053c601333f7a8f38a1390c1a98fa49a2a3f988a598665afe62d544994dfd1acf0791348cdd6e0d5c505acda4a7d4c27e087c53b99c33efdbcd02fc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5a72f8057e5f273ca9afbb7f5632104b3c8f21f41756216974032a3c37e17d2addb29576c251993def2a9154195ad641c97240c704bbbbea831a9f90650199bd8c4ea5f0d50fba43461c54cd1b3ead8f676c3d2093db2149a298835b6638bc4cc32c3ba52babcc82d78e8068356371beeb01f0992b986d20f5bb80d8321d9931;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8d779d5fc1f7962f64484716b0eef3f95424a2c88a73965339207988f73936b25a551877b50b0dd95a40201e511917b0b0bf99fdc8bf2b0b2a603a83c5457e33eb5939f60277f0cb71f8a5190d1e6b726783e8e90230c8a257f5c62c263be77df4d161e6d1878600165e29a5f4d235b5736dd4881d43713d6d5347f5a5d73c01;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h82628ddad105e19f85eadaa14b1af8245bf8c5be63aa27f627cc20500b8488c2bd330dd11ea2a303c5878b4fe2e5397cd657d4c4575fa10e1f7007809d28b65dbd3df3cdcc3ea56b3560c1f503386928dfece6289f6d1ca76cca8ee780a8cf4b89cadf66baf822153cf3268815505522f27194e1d4f3a6ad58f171d9ec10ad92;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d74a20b251e4d480273eac5320a312335ddac09ccb0eb83270c621d7f6ac9af13077bbc0144d349638b03fe5149e15b8a8e616dd15e048145249426833c04cf0579b91a0d52caa4b03c8186b755f59396b8005eee9e427875899c80395898cb8618381b7a76a27611dfd9a4dd33b5314a5ab546d302372b79e5f46bbb45100d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbbe205a9a19b96040f11b72782f5d61b4908fdd673c606338868d2f73b80531320d7f325947c5440e5665d483a826475c19e3971898b785b31bcde0a3d1ae3d85e2e64852042f11af79ec7226c85214e80ed267652106719d35bf020ed3de3c4f7ce7b8d25c492a412bc31ab8b091bca5c99c78424a6f5967607429783aec6a2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ed8e693663b0ea14b66c48f1e9c601d7c2977b64ada58f10ce32ec7e057559f78c1375c69583a43465b54391299ac92ffd9e283aa7b5f19c2f0f8f4ef10bd7d4fc268abf2a1b57a6f842813610f354aeb65f824be6f247a28d7a07a7c9aa61068745f22109a51ac711b8afb527d96d36732f485e8d19e691b58a43af346a44f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h46c9ce7adb3976429084f4962656f0f1a3ff52120c96f563be9389ffab535a60aaaa3eeeb49c8bacc7ef6409f3abcb4632544e90157fcdbfc90eaba40bbbbc10f7ed93bbd9cfbbea609f941d41a2b617789116d8f88f2f152abd27faecba7e4abd57bac33d38acd1a29c0969bd3cdc6ae7537d0a172ddc11b0f0da0c221db05f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had3fdf705c84807abc1789abf2525f3a13a2736a528b16b7c66d2a119ab37a87536f06f35daea7dc08402c79e2886a66cccb6533ec733df7bb6433394ff0e8dbdd4d26a829ef772b7ca83fe8af7ce2b213b1182a598d0967d9e09164b24b09421223f76e95a7a2904fbabf53b43b355feafd504a3926aa2de993d60db805b730;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9ae6fd6d0849c3c2e615ae1e7c28b6d8dcad00b2c219b1b079d4e2c635cb70f7323a130bc5f37dfe5f05f19a6025656581735d700c6bf165c17393405c37c1461e003458af49e5372780d28b87ac842d7da486feddb5129faba5a214d76ae62ac07113df165739320ff5b266892d96f808c3b2e4c1590c68dc147bfb9168d299;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h211ccf07afe2b63e96a6339282a2155535a757ec52e253dd807c8c9d71975d439885bb97e9b07e7492c991e68f22c69b4ee8834ea1f50d7efd81bb90e1f1bd4e83bfe9bb01a1cb2bc852fef547eed2df621078734b34aa4d7c399456099cbb9c298bc36ac7c8f083099a86d20a4af712bff05a56446a33515cf38dc1c9244b55;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha006b7604ca2701734010e456fbba9b26adf6558b6e7647185202f306d6f8772429aab5bcb8449a7b5b6c5c8234583e127a6be237078c857de045a3a7398c089bf512f6318b4a65e51630a1ea5880f70095724e0def0d1e01fe77f391536a01bb3b7a06f1cadade1ba433e72870107ecfb81cbca7d96927bd72a9183320c4c04;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6b4fe782df1f2a279e07c1975d195679dca48463802b5cd2d635282404720382537d956612b88cb391985ac179dde98a0f398bc0ce78422c6575e9461fee01bdfa55883fc16b923dc6531fe00160567d0470c73ce1ec33e56685bffd28bbc4a31365eb0a911ba401bba35124722dafe1556569959e57e4ec98f4f3d994bcce4b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha2aefba3f71cd67edb87b33a8a1fd8b2a772cc0625d59424117a2ceea6adaed05be2e9b4a1fa04cf08c67c6edab313b296bda8cc7a7799b219d3bc92304c0c19dfaf451c7211ac84910e19a016ee97c0ad2de6d285fbaf62523ea47baad1a659046836637a2ae8a25ebc35e577dab48999749446d56da19398b18f629803b06;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1ec14ae14a1b2184257758242248f8eac68017ea87d629a30c81c8f75db8f2458b58b695422097f5c8951fe5f84208036faa1046caf5a4fcacbe2e740615ca7d25a52d097c4db6f516198f52b54079c9a56d2e9769b469031b4bef722f6234d3ca2ca97bdd4bad064353fcac5406ebfd02bbc239b8de02676b96e3b32e9a963c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1e8d2c6b626983915fe4c153603bc4e612b887dfeff52e390bb737c7729508be3d6b739c3fc65348d48a0374586290cf8b6192c3a5dfdba8c24bcda904b160002c8f4dec694d0e3479e77fe2ddbab6287144c8137b7a48a8683716b92039911fb17e743cbb9aa6988f967e06337b1bff0b551954c40b8b20efd3f2b3d2d73d3a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h40fcfa61d9a8f099cc4074437328953d34f626fde11a498167c1d804f7805d6f275464f07f69bebaac929123e14e030abe472de427ff3fd6cc89cdcf47246f9a9d3104c4e03b6d1be76cd15ba5daa6d6689f6297e26fa4ed54a0b205529996435330801f9acdbc61288fad18dc6dab8138126970e6488bf25a145de5d4181ae7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94cf2570a3dc32b3fb6c3aed8cb1d64abe241bc8d6a6e41954162274cb6f73b914c618498a5618cd3693210d8f18d4e064aa9769cd8a0439efa54e49999ffbc1ae3bf8edaa3c16865dbcf40d0118b815d9989367e17ed5b4d306a00559c08977335ed2b9e230351ddd7f437115f2c9ed0f1533296ca53b5c9fbaac15a87a1b6a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h81be10a0502ed54a11e2521b6564467f44ad3e9949c323d6ef6df60462ddd92798cb20603e92559db51e9173592338ca71cf49fd10dbaaed282d44d26ede99f84a5dca9d39a0d8710cc3ae4347487d4a21c136d5fb8ae14193ba042f5465254d239f91fcd33e54929aee2c852f4865d7e1501df2be3c43e0c2d7de3e6ef26aaf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfc5eb32a82ed3d62c1a70107e7adb889e428062164f2ade6c9c92c718b2ae6c2fd5d5465fd30ceb6090de0633df18bca6e200a81925d195e4276406f503d8af28ed8b8beddd09e952d41ca7418144f5fddf7bec9fda24db1a6acb9d24a5b21f50f81d70d2115bcca620dbc2ec996b2da531249ea80f875fa8cdfaba47b92404d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6982bab76cff4825608d20fba78d8327c55f646c8329e19c93d4f07bb86781da68b338dffcceb9da929d45fc1cb2765f7008cb0d77f5c2c78c9163ae096b2a1a73ddf677284c0342b0183df663d37bfd13feea4ab4b8edc43c6c15ac6a7462be27cc5aa08ef89fdd33009d689047f02e1012f7c2ca01c5a229e935abafb3cf0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf91352511ffae0357426add1cf0910b3e50d99b04982809c4357321dc4b89d6bb6baa25870a0074c01ebf32a7c84eaf43e8879a5ff6fcd3e728170de49856ea7e2643aae0b5d3dc76c522583122e9827f4edd993ad5afccf6e52ecc0fe610b8e88e0e3f6bbed7796e5e97dbd9855df42ec4e008b39148098f52f2e5ec74568d0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf39757a2fdd97af9d24ea53fcf9d7e7ba9f48310a923e883ff30e68e024be3254e35e20e263386fcb4b7a12b9b61ff8ad3b09bfe818c864436fe381a31aada1d999f60881eb3b020d7e4db1752bbfcd3c856a92721dddd9c411831ef325b8d907d2fc55969e2e090c8e081b62dea348f63c2b1f69025426c6c1c9ff55691a0c8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h31157864a82972a71c80f54e5f044b3b8ed5ded96c0e4eaa56a4ccc72e2674c6d0d7c40b4eaaaf1749d1ad32c58b0f704aea8f23f7163474326fa20ba6b535d099e5846153037ee4c9a63d77a4b2a5cf4af67212f71f15ece76981dc0d5899e415cbe795dab3d23f25f825c8075c247bdd58ba2590f6d3f3cfc7708bb6929538;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf3d5056fb5954c718691f1e65819a6309fef4d47466539bed8b2a68eda98fcbc05f469107324177f1820e74c324b301214f1f39946b373552d32c78032186d9d2a5dc51aebda7ec25723dda9543fb400e7cb95236048866ab4bca939c3f72c3dbc1f8953d5ac1ac2c4bd7c2bab638deeff3044e0a2a83a8e517b6f96ce647c7d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h74ea6bf86e559aef70f829f404620f49de01036668eca944c6b0568beccb6eb8e1c69839ef9073431b97cc7a078fc69b3b10a6922b50e4ea4d977cb9690db0e628d8b5ea1ed4f5cb4c28fa629f03365dece58e032ef754c2e1425c84160aefadb6c108db0ac3625db47fca985e0aa5cb46c3688bd101ea02b79a508eb69c9367;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd81fc3e1f464820117019711a68110f4c6e32199d1c9f9d21dcf08af34f9d44ea78c8d582df1dbff7f6aedf7f9a9dea017ead549b02e451d0027ae8fedb74db29f1eb30978de1c044e16e00f73c597b52f5b0e823ac177de5fe818c5bf50fb72cb999addb165ef811ee0547cb2a222eaf6ed09222e15f4942d0ab05301a8a30e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd3ba91338fcdd0eafd5fee8fcf8d89fde6d6c29d07740fa9e61f0e35e15d3170a1755a99c932b355ba4070612d0b9ec3316100fab57e6e155b2a64c985b88ef5b842245e459d7067b87e136cb5a9cd69dfff1ab1008787922a5522e6a02ce0e806a70192b9dd595b65639db17e719b0c46054af6f9f99881baf710f6e691e5d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8de3c6d48ada950deb1243a79fc782c6253b2465a56478d001a827807323eabcd09e3380743ab9cb49de4dcd0a303ac1f9878bf8cbf8945a79b1dcfee063d5b4195a5967eef421778505112401bdc9742ac8cb3927ad27363cf115f33381954a3503df87a2f43b987a8d9f0ad3120e3b98ffbfa44303e21065a7c769ffa09a2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b54c7600b238825e929d8c3eaf27bb6261542fd548a9e00420786c45d6087c80bfecb67200ce9d56a89261849e48e4c3f7ca7e31cb527834aaf091aec6717f99019e853d3fdde4bf50d9d1e48159ed890b59ef5f3594e9577952d5c40afe27a56b71b1031d2ba9d98e31782b73630ee9802a3bfe731ee116aea451d5d6d3021;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5240b063aba35170064450a84e333cde20d477504375540e34c92b09168b6de00229cf3520f44a114c59c71e28a9db684bf0f054e65f706c7320500472e46c00b71e4ed667fb346d2a2803338493fb66c88c617a6db773168528b7125e16c11db12e0f630e7faeb8fe3f5b7b57aaa7a6c0f0bd1a4d46a39b6ac7f5a97c326e4e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8c65fae14832f8e5a3a0a9a529b0c3ea8b186937da3c533b131b57207c3fbe6a1ea560dde6649ad452e661eda6d492c1f77c607d8eba221966d41288a70c26d27d7d72619c2280ba7ef8a5c1623169242850935e353403ce44189e57fe0611a19fa85e2dc1a4642b7e1db18daca51efe41484b5fffae27b4f3efb429c6a47274;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he5bc49795197c235519bb98ca182fefa0b9bd09fe3c8261fc04f394eb8fa2129771e884bd6de8a2d6be63cb6813a3b68ff33dfa279ddde888f815659f77ee9e83f5822aa509677115212f7f52d440497b6284b8eb47427380834e7351f400a74451420114873b66ea90b98c980353159a21b056881fa6d02d9503b37a468b1ca;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h833c76e0bdd9a8652a343e5265170767bd80d732e8277d90cd7a83d672b3032ccd56a94ba7a2233ee0103d6994ad7163cd58cb4413f9198de190c48c0d48475ad8b1aa979cd0b24ab92aa7e222d1982b87650859201ebe76127fdf93df54c035ba5812796d9e596e6e0851a710d5ca30ccb1ca6dce7101f1734f723ab7d63106;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h236e8b9abf1a2dab3501782b3f8adfcc083d24970b7675d430373d7eff90d59c5c8d131446622ebe346215acc50d78019d86735be3ac7244b46843cda0b5ba7b86309646ffa58f1651c023a3511b33eeb7f181f8815f9d022d17021c1d23f12b8505c64bfefcc00dc44434f82eb982caa8f532bc269de332e5890fa3a8ff0aa7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2daeec8c5b4165705137323829c7db3f08609ecb961fad1e695d1436c4dde3f58b1db2efdbb701e34af1fc247fd2ec4c9b586e1aeba8f13148a2a5110a82df76d37be46ad94c7ae4a3207f939405157134ae326e5be82744f2b53318776f2608ed7964c0f3b4cfa62285e611116a87e3b018f19f74aa9c5633945e92baec41d6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e9f035c4f9c5a44df3db93c6b6ce57886adcd3c5873cafc2c60de3c0d1b48ab47c336a4cc36c5c3e0679343065da01c47271006deacb438acb110eb7afef412db3323e008744e5921abeda4fd7ef697601e860e79d2742209f64ec36bd34bb9b7590121f3df46670d57861b058e6d3395dd2bb9d446e4e7012406bed314d043;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc9299df3f66a9e2ca4ac4c5d158258ad1f222bfbb3fd0cb84a1a875171a1a9fde38782cb31f42e6c4e45409f645646f405f1368b1d8f03a56b5156de283615885ef5fd324eedbcc5d06dab63dbf92818863f1585bacc42f8fa0f6add78f55f7a4e5d399edd5c2a5910d1ed38e9b56ccd6f915d07aba40a00bcd50ca868cf98ad;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee27045b71122820dc8142391457ea6d34cf85dffe329c9c94bb6947c630e64bc45d232fb85ee0db3bd763399ddaab7d677de9559160df58fbe54b39ed7a5d97a04437c7de8e65f0d2a23d62f7dd4d0515be349c4deeb11b4cbb42fece17236c6b162984616c127143dc2131895c6f30db334719c9aafa88e77191f134dd9d0d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h21e515e6f6413ee9570ef693cf9fff28bc113f96aee6f5c6969899cde492f06da1595ae89955f37d8c90f3c9edbf0af5ae9a7d9320e258bd667821fcd677c8f503d747bb7840433eb28e3e4ec6d5623d1d3eebc39b4b273d83d93479e9a941b2fb663139c58cedbb3665b690b7ddf726c706fcbdb34f418510d29ee05a83a390;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf37bb21d5ba178f12aa6164b2bbead47d912d293f8674499563b6b5097dfa7272311043d835a281c7fb4daa403b340a51d41505763540b07a833b7cb3bf504ac7b89b3dc77d3cca3241e7d1ff04bd44d3ba2a9f2a266517b649b751512adeeed007f3207c3757625e10c2fcfe21526120a8f4a6bda5a657dc7ea31e9e0cda1bc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h70fbe98507c7a87c73041e7de67d11b4a4fbca113c7242e9a22d7cfbb89d1ed099456ae544348a98967d68a2027b0af70e5b81a7bba138448d5c708265a447a2a0d2d41504775ebcfeb66d26d97c4ee7380cb80c90ffb3b9087cbac6dff68f024b025f3bcfbc6da083f2a300a4ef96314a9897f7733263e044def439fb238866;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4239022ae5ab53acf03a90f9ecf8e74fbada858914f97c98a939d5e6f51627d886239edaaf4717b400203406b83413baa2766f4b2241dce5c5e18d9d6631fe53d1ece32591ad9585446e40d5963d59435b3efe37950acc8f0bbcabb1fd4221238c63060227527372eb36e27286db09df309518b8edae501f7ae4f7bf1fdac876;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h51514ab48e0af993799ab1a9be602efafcc667e34f2fe5c264bc8157408bc2cc9dd0105f80e5ede7020079eba77448bc2ed89487a371f17adc01ad2dd9d935d335022c8e7c06992029f0599af763d644ff19bdbde4747a92031a2df18ea1350cf86d17de6d84b900da7a4ba32d807cd536efc8e22c36677651f91e9bdf131c86;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf0c84b2a4e0ef74acb996087198e640017738c39de9d0ee4506c8bb8ee2dc0766d04ec9eab76c3e5fce75938481d317afecd39e6fb42ad83172edde0f5c42d2f260646e00f82bdc55e270b68a7d6a1e01a2fba87d237c4496568fbf72dc7c50419e93c36def8871e1b55c23b64245d3713679eb60cc90884e66691a772800ad7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf5be2ac9bea65b4162ae0a20a2eefd8f54f6ae53922fb15d12076906bc90ade026b4d05b76d5f1a3f9ed7520b840816d1ff34b9403daae2b29917a170ce27ee19459b45590005406bcaeda7b7d8bda6296f32d1a946ef0856ba6dbde85643a5bb3db007c744c59396fae1c9d0acd6b2f0da92e9cd459245e63a12e92ef8ad2f1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d385e22fad88b3480c0d3396b5f3ffda96f5c0b26f698ad8abfb3b32dc30080f4316c21e5b720fdb6ea8ea9f4282d1904c8033d244a7f317754417777af0ecb381bcfe26a0b589cf510fd480dadcd221b9f493b04523378b11ed1364c69cffcfb32fbd60925f5450cd7b71de5fd5b9aee9da2215b3d79ec45020d5dc6b6c676;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4b06e5b430509a41f3780fdae0d493b4bdd8d1afa09d90f25734c55b5f091f32b1fbda3b79164f304203adbb630db4eca260df2344d7e6002ade792151eca3b97422acc9933874338c1b6e25c6781524977f8bd74e02fa8d9bdad4ade5c64955aca821fc086576bb6f11de039ae4b75718cad4d3d19e069071fa782a33fef396;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2fe38c160e7f5da97833704f2afddb111043dff5b10547729f949d773cd477826d8bf110e20e1e35280bd4c7940d44d2643a2d8d8a6b91eafc379e34bd6038354fa0753a0ad8d45ab7e20657399f3a7e092a2ce777840a24182349fcb734a27660cff50db3e1e1a2cc5c09ec36e7c992e9c75079107c718aeecbe45ebf1aa9c2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2bb93221f97438dc16508ab6b81826dcc42beda33892873038953906346dfac1e41dfbe930241e691b390dbc72738abcab7567f464d082ff72b426c08af4a4c4e2aca7d0ff8d6d75c9ef46b98263fbf543f4a6d08c7b340f7f40fab6ecc137f453e74b198eb5fa4d55bc8a96d39ee609de4db1a0dd8c2925713173b7cb35a279;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haeecf8f4dc88a23781840f351bd78c5a69f1d98f1dcac7a795ae606af931407e2e26625e79058f4cc543e71530b8c9e5c84fd548ae68dc78da0b41ee67b31cfaa130aef0617a82e61bcdca6fe36657343b720df6a91ae67e436930c667b73037d37ad23d0341b8e13e2ec4cced08fd3b2a98c3bdf56fba4edf2533be64b4dea7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8ea4251a4c44bd90481d5dc594eb5eb0983b1f6baf8d26a528c74d1cd81f3e366f88858445ad3096b0130199851ea3e2a488e557f484b0a3068ba7d39e99423566773cd94ea2d18b83ba4c2527cfe3e924bcd86ad6cf412d83a868e33bfe0bebe51b563784ffc949384eb161990def9c8029c48ea154c29d83fa3f8ed913e7c1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hebe9ecb098ca1f9065cdb8e9a1203dec9015c571d9e411a84a8a488652a4b5175ca33176a381103c225024ef05292c7b900660564ead0ca92bad5ad323474af786b988b65aab20405df3a6ef52022cca90df4ebb6f65841e2c3149e77aeb1ca59bda3733ca19b34e783ffd686d6184d968d4b840e71ba37f376dfe7da2ad5907;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcb8c44178e6332cf28f64aec71dc81394d5c18fa01fe3b7af1bbc927e06a7b36bdf5945128b142b979e294df1ffc173cb998687ca8cc9d67aa5defb7735142175a3c4b3b815ea6abf3b2714fa57c314e8fcdff43c513e688e4121baf698ccaaa7caa8d19a229b0e1f13001c1f00c9c4172f47814974c1e064381f0b5d7a4c70;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdc0d386f2ef04b2a257e0986d615b34aa924f6bae51340edb12c40445a9a753c4eb1a7bbe11e3f515f43c24390800120687da17cf52281c3b9a1a5c0689ca678a82d1fe2e2c26130a22b1f36ce6683ab924aee09839fb3f091818a293e187bff2d11bd8fa917ca7783fe9bb064ae561a940cb497b67df67d6ae200544071c44b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h44611157609e65dfdf76525b29ff3217c0a1240e052299981e5c9cd3ae312e6f657247c74419f55c3faec627c25d7519f703a420f66d180891937aab4f8fd530e61ffe9a222c42bac7aef930dc8f81dd7a845866dc06a3525fe927ffc491d6452bfae4f0d340ff03e1e59bd9321dc2b26d0d196d45f409865bfaf9b4a12a137;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha689c997222d8bc929c7cb9cc158ecdc384256119f388cc71774ce98f3c04df977ec13a735a705d11dcd087ef462aa504bb7faca3bed0875a448e5e30b4c8d76a6d04ce0a820dfb2c763d0792fa0206916c3127cd9168a2ef619004467e0ef9c733aacf8220a49af209601c58436ece1f73e5eb603245174f44076b7eeff3f63;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb89f898c9db98d57eb2fa8d5703943f1c5b975e45ceff0f27c84838dcf04c533c029c4cfae2528c2e928f8120d040ece9c38ca3dc40756da055968be75a4d73c7c4d25f76ee8c622a8b0680be8c34278b790bc8ecd8e4f592f2b37721866a9846edbe247ea13fb54a9f2192e5200668f3f0ea5100f9a57a9876b183fa5f8963b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha0c7f66152a4951157595eb11686ab78c20e4c0c395d55d1249eec84c2b0f9b0742f61cd52f8df0ec0f66d08ba32fac50a7c0aee9f8c27a311a3bb533da51bef7675efa04bf8309573d008197b7f941f2b38fc2650d1548c50d5e6df69c196392efc6b7c3f688c363d0be0f65a301ba0032d9d282b7dfb47ebd402650b26b2d7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbb5a7ca1b33ef74e61f9eacc57183b54b18850b83fcc75244a3e0b92a1e5a1ea4098b6b43d53af3c56d6f4341b5249ff7b37be45677bf6003ccaefe8525fc817f948a5f6adc7842b6cf6430d70c361ff223e71dd421aed89499244de539273b2b62235fd2aa84cc2b9a882dbfdf049bfa774b91bd7bc6f5b63a2a4fa3dfe3d35;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc917cbe385e95fc8978c8bee401c8e91c4b72cf19a592e3482f435421306da69b00bdc3a7c2b219aab10cfa14b19d5afdf85ffd47e48f74bca29dbb92236e1aab2c5db030f0134ea2d610b255605ad22a766c19db08da3cd5daa095a440f024e95317f79496534c18a95c4e7882d53c2f1437ebe9d9d549a8ab21043cb9b8a3c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8328240cfc2dd177e0600f33818c81795c894b7f8bf9c515bbb4da86e1264f8ee5117a6cdcf319d798b551bda532ad26cb9ddfd43d50bff62c39b26015c60e319ee56eedffbcc1c844f03dc47e39624956d22c9c4dd2f3adb3a937e916f72742be343c615ee5059df59ee56f37e630d3b52fb2a32ffba13d9da73ba4dbf90f4d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h26c4ce18dbb01c7c20f5f039be6e0e9a283850915897f8e120510914220f4886b2328fc2cfd9fddd3a71b4172a2fc06b9c1ceb2f775388f8af3117f471713bf55183ae4f959b126d70418311b3de3700ba221d7b0fbadda10f78aea6deea9029a7c386f60af2229035c4eeadaa4d84aed7f69e73660cb71ab556314e9dcfb2b3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h47b29561807a0fe084340da71cb0b0ffbf43ad9f206d6a47314237a5cb719dc358fb7b26b8c162f01949a5f74b7678be1af3275919e9fbe81449b9aebc4ec291818cfc98f44521d60abaacc9e0b0d62185eac0c0588820cb5437f8af56d463c86a6ccc3a726c4e1136bae8f5c640c542354886d7138fbc321362a05ca7d377b2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc69751925540ccf904976f4e7828c8e762183a63fe92a5be2029e7d32824a66ace57205f7e1c4129ab4db781c389c8324ef5a365225bffbaa6452de5baea9713e7fe5755f02f5bd583145ff40eb2016b7ce026f032f6bb280ae7287b88fdab1bc79729ead0e03e24de574156f6a091c0166257e3593f9936b8721d1620fe647a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h898572ad0c3ac31afec1ff80258f74e146434d2c9b52f518938f106854921353771310d7baefb6924b007496bc56fda0923f6ce38e0cc98413d9cb51a751717a2966dc2837ac7fea63283d4f918453a25301dfd42a76e2134ccf51a8412da798488231e68a341b1684533e307d5eaa4aa13827f0afe04a756f666065229b6b15;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c76b79611c22f34d37bb674cd399ceb94355ffe69801efbcccbe42af1b7470ddba3504397725db06d6fa59d6ef5bdcbf5b1da22b22d99b8411c51543791e9193c42de1c6af19d2999064836179d25dc229b1289c3b725eae81fc2a51a69a6a2e3467e5aef47d0faa9bd400f7d2b56a9510a64cb8eb80f6e691339b447ee913f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd873c62ebe1a22f03c0f945d9b241324d2d2a4c203e8d7cdec8cc2502e428f8a61e190da29fc4088f3c26ecbf9c511675e7cd807cf576268b52d6b275e8ae7ddc16734b1e40c93b79fe8dfabbb74d856a0a40549d148abb8fa57b0ea6a2a1ba05cb44bf7056628f78d851c5709c81224beeac8617e2076360fff69f5d4573f2f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e87cec002f4692283747000b89f7fef996822f44204565c5ec63cb30bc79bbeff2e1bbd9a5f1c6173ab8bac86f8e86b761e0e131d0089cdf23604219d7a81023592da1afd3bf21a2e0cb83de18df96a8daffe96a09729b1eedd6ec31f977850a09c6873a0d4b30e77d3ee184dd939600efaf22573aa91332e4b0081db18d2c5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha11e0acfae35005401de9b896271d7485d0c4962867c35ac5e13e67be59382cce076d980e7b3430b7fe65f5d66d508f69e3ba8b1bbe9d923368eb9e4338cf020ee114693a4d5ecd70bf41390c5f080215d2f37edcb44e397c1d7a13773650688317042e788558677109911c56f60e2167efafc8a2ba3b498f85fed3a9f1a3830;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbfb0a556fe5e1be5af21b89f226a1a29bd09559db7981ee363c8fe2647047d25bba3ee9e6dcf7f624bdc4d4f64c6d4b628a0a49acc095acf00c6e8ab946fe6f092bade75d4c8f72020247d37d79c3ced601e7f61a48dbe3df8a1595ce714abde5e4c9b3c2f7a18683322292d046ac85c031cb03322472d4a134021fbb3cde261;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4417649434b538fbd1c0fc3f56bcf6066fb6334af2eddc6ed8303a438f46b0b7b7d25a225eb5297667a22dc42a70aa9ffa019b7c986a5df1e97e6a952484a1109a1fee4a831cb12d2a33128c0c980a552c4c26793544ae20cdc053755ef060bf2cb3605206bb46638ff196ee2cf04bd1f5b43826a78156f53d82517d2c81bbe6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6d1ceacd87bdb531edefb0d3271bf100a47f4c4535f5c29e9ffc997c7ab9976fb7783e95ce8d129451ca9306d5620d321f798f3fa7fa7915f185ac9459b8ebb43a033fc7944cfa356bef5c5a270c7d499381cf4522cf80c02fc91d5d80f4b8c023cc0ae4f3d6b645175ffdeaf541491d5a32cb64481c818abda173895aa13c17;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h463da04f5f667e7e84358c1296b3632da8d780521ea9d1035e14798d02835e411b30f28568b02d9625c062c82e9ff5eebbcdf809a18a51bd2999d0fb1b1e17aa675116bb142dc4864a9a0c1d47007494029d702dcd7a61a96eaac6e789feb5307096dd851ff3055caa0ce1a6f6f844753c2df9064982809e63f538353eb56b52;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h86faa639b2e87b55ab33f9d9a0fadb645c63a88b88ef7ccf24962bb8f50fe9b7308a6a4c80776c6ab7e63ac51f85dfa5802a9604385f00627804eb903838a430ea754e25360e955e8579a4129b22be05e07e81d272ae8b67d86c69974af1d633f981ddfde5524a647bf54f2429ec0f5f3d231d356a3206b32198c34df76b18d2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9c4a10508f22fabe2118dfe06a6572c5000e3d006a070bc3804967a865b988f10e9b233337dd71e6d6ad4f011d2efadcfa09b031a2d010b84862bc1d88ba4a45196f4fcb5c610b2cddc62dc8177bb97b8e9521f4e571bb9055b75eb597283c1a8a99b661bb25467b36de1d1aeeadc13a8cabe593b8c469f2c9bdf995eb15e155;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ef5dc1c2fd09eb98550cc36f57128f6078dcdde56092971af4f98a62b8031e065d87282f4a9aa67caf2d400e08f95ca4511054b4b7af134ba3bc237279dd3e2d5f9648296f5258df018fe58056adefb29bf695f0f500d3cd6e20e761f3557e6548c0e4415516da4369764c7acc5f9b18d6eb91d76e8d831a3dc6174a4b688d6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha74bbcd079cf0701f58222546c65394a1a6f968b9533c2994b4af2ab6f081ef5a1cc02e6fb38ee3c1c3c697e7cd9d213d60df852e631368d5fed799e2832264e1b6206a7ce037a886b167a6e5f2196134d5aa64dbc3c96d87cdf9cadfe75f4050a52e9e7f51b8d8db0e1dec39d23f81293a2ffa58c2c89b5381ec270d2c68598;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c092d6072ddee6ab47130ba2145ae0db43130af132cf446410c932e8bf567f2ee843113667fc6d519faef3c8d03e2d12bc9ad2f492448982c33bd428788d905841bb084c7a994967a2b5649751c9d47f3fc68389b288a55924727471a96f29cb96dcb8fcab3622b37bda2d99de0e211c1010eed786ee6dd6e331cfa70e6421d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h79da30490941100691163abebf9e1ab483484566a6cb7a1a5742016931e10ec5b544e2b2ac80edff525fe0d5ec4d6670045db5736a28d8ec1d51e56c26ac76c0ee99d7e3866d5841e61008247a5359a9c9fd0ab32dfe6282389933f6a985789b7d37c4afa30dfb2f33cd1c24cf5bb3b0a65db82332366605cc0b7ac53e049d22;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc57c88850aeeb49921f9afd790387c646e5d343b317b8df612f70ce9c5d1637dfb01f5ad00631a32279b1faca5d3a7a095e1ae4bb814c8b222a0e74668b54fa528f3b46cdb05afce1a1a5495809641c81fb68d5a7bdf84b68dfb90d692a7d6e6e04e37b9fb1cdc45b7765b7b040e3d09d84206ea7c8c682bc4b38a7f13a10e46;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb39b9482638fd9c405bd952a63b923c128cdf6ec6bb3d86e70f86a28c32bc2493c0be2f41c794d40eeab9db98ea929ef20e8df14805b66acf263c47cba61c4be1f03b1c89c9918c83edfe456644a592cea7e86045e8cee6b415107e06d320bdbcc84ec09cc1f04df709a7106f31c4fdba43f8deb025bd4069bd19fbdb4e5c740;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha869da5a034664debf4e3c216143f45ea84096e68253227fd3615bbd893b3bcc237b1d00c10969eea51a1537c1ca405e2d51d31e5797df663dfef9fcf64f0ccf9da3a416a8be296016729c7e827dffee9ef67e4de86849a45a8ff9b411dcaf7c69c2586bfa622e0cd0a4a383421fd1f509b598de6c0a9979ceccdf5e45135e82;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8bbd089db1e5996501ae4e5aeec1ae218850d97a11c9dc099d8b4259b70b467d784530d6b784625d06b8dd42f33c38290c6870cdd4fbc26635252ff83770c8f8ad7f50b2bfb690c08ffc408b491ae0ccc5549cfdeff4b89220f33ea6d0657b956fb826f22a2e8ba4bc557b1dd1e3917fbdd6ee6a0959eec00f2aa8eba041661f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcb50686ce4099cfa5a9f19e17202da05b4f4675ea5e5660ed12d2fe01daa1e9417c97b8dccc60d30c4a257ed0fe38bcdde82cb0eb3a5bc580f53f8dfba9eceff02b64cad7c38a4f8e039f350919ac682f911157707fa3e71d641a4a32cbbc84513e60fed81745e5d117e2b9692334edcba84e3868742247e5765343a4f36d72a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f424707e01d8e0169031723bfe94b1b7299b2f5681aae40ffa95f256e89a2b34ec67daef46b9b0c770ef952007cba713d7fe9498844535b6eac6d06330fc1e579b3f68d4ccb18674282748761861a438c379e6f54f44ebc5cc4f9ba3fe19416605ff37a162d1155d35890ac758a01719f7bb03d9ac4e2e9ed5a89a1331c6d95;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed5fa22062274839a51339939a9df72e5e5f7907567404c17e5ae1bc9d2e874569a2aecd573cd3545a110ade8c44732b7295fd7f76004918b47aa8830abda4101c1dd6b3843ba88ab7befc890451d94a43e538f5a5123c2c9d1033b8ad1bc2c44e029491c48e44cd6a7132bbdc11f385339bb7c299be643c8c2f7c489f668508;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h378f29f0855454c5909fe229eb94f2f66cdbd96618dd9a78c8ea5b0013ec42f3f523c8295b3e45d454adef3e13e0132f33ee10dbb834426b16326d2d7361a0e0a0b4ac2071d3e167e28736991164f2caae516c4e64e54aae23d7cc76ed6c45ec089f3cd4e0c34a07488239ebaccb98bb59e3433172d2bcd6b8e585ac86defb7e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb669eabf523b29382d16a04b882049036c1b752e01bf8012731cd82f536659f98495e3929898fcec6421b93008a296a5f893bef02a761c300126a9eddb15a8abbd8ce9f918fcd1ba7aeb4b3222d0351d9b2db034d189b437bf37b733824328f3ec3f02de17c9862a9bf21807e576eabef4cfa48b2f9683a8f7f57e0845c8fc41;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h785bd666fb2f2e026c758379adf53471238f3a648d08c2abb450fa6edca1fa220158938211010c33337b39c19ff97486895f9e9613449e3b85e168cf4b9eee601cc8253e3d0a130264fddcdf9731246d56faca518d9e4910140bfa1a0b5ed591252d23ff0f7e98fa15c004a09f6948a97f35a9b20652b28c670272d975186c4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f715158287e1de1ecab81059ca2b2fc16980e39603c7e300eda9906da87f7a9d29d83b5801e32ebdda01bdb01cf0370d60f4b96ff2c186deb16d52ca5a4c99cc4f0b0cbde46a11b3fce2265984b38dca9d7ff6be1c702e979f142ceb552bb5b9166a776423a976dc27f7b590942cd3bbe0f18deb960f22322e39c36bd7a5d29;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h127f5c83389af1b1d7147af062ada8b7141087aa10d0c55dcb38bdc60aa14e035e849e69292dfe0bab2b020b1dd81209b8ad1f61731c4cbb7bac865ac4bec71b773a2acb86b6fcb4ad40d37acb669b335fa36fbab168c6ed6599ce7d72e2fa788cb38d47d327d25c9e354aaa2928f9a4bef155ca80a8ea60c6bb1942324fb07c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd0bd6945662e6cd32d5a3a073e572cc27dcbd01b1b4cf891bb70452ff45489ebed3223df3525702a2bc179c6078bd8eb6d1fc88a1fc4f1868bd53d1a068a7ba610f354667a22a3455e80a5d3082a992984642dad2b04b56181482255b2d05adb935d72da01315ccbf5e09217897e97c3a559da190020f3c6ac12372d5c9cc60d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha233703905d7beadc8f23dfbbff542f3292e389d3d608e1917cbc4e879663ba7e2dcbb9d1bac687c6d125fb8b035483fdff57ad916909885b2cfd2fde191001bc5dab9ea896993a19bf322989868013c0bee02a88223b0d03721961b712419b139d4e65442a6089288ea54ad73f714e2941e67c224952184e716bce80c457b7d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he41fe4316d834229a3efd2087b0828b84e2a162baa534cfd486d9bb98adf39f2470657f2fb26aea146d7bdfcab1e57cd5e4aa9efce5e023a100ded5389afe911276ea28bbec27f5989eba7620247adc23eb00ba424ea8278ecf22b93c295be36fb5693df7535fe1e9eb2aa2e8452f9362ac3fdaf256776cdacb332b8d08d8041;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5716be0f6591c9cd8199801b5a1bead99ae98e94ea8634821b2a9979dfa4aa0c27908a71eaa573ea9ad5d9b51869f038057756f6a7b7867a739dcf14a82741fc58c173ea76a58b72b81c6d2bb4eb60be1c9cac565c6fa1ca1db61c989eb3a7e2dbd1246cf8a974f07372ccc1cf4c96cfd30d133400d82979e7a4764c50145ae4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h24709185da5737c470deb6ae84d59f5f79ddb4a6280515d349226d734787dd2fc54a41f2ec51456f97ab8bc1a95246eff412154c9ec55de91f19d29dd87f615064f1e83b70a8af6d3fad146fd207971d6504b316affb1aeb91a35721496e14d90cb98a27ee859be207f4f801b3907e22962dec16bcf4d5d17878ffa8f19b932b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb1f343554eb255de39043967b0e29fe23394e73f27b6a98803498bdae144afe0fce696dfd4d5e19d770d9c536549a5ba5079ec84a7ef82c361da4bfa8c099dbe4220371f2a3641122a2efc22a166ff8b569121e037de7a4f3699d5ddc9e81812c9586bb9fe96e456a97ad4b3deddbf8f910e727152fa7ec11582e52d254e3dc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hac2170ebbecad2a9269bbc5cbed3f8425f0240243d69a5486218233b035a63e9de2258745ea659f7877c274005fe74aa80198aaebb20e3453de37f2d3cce393f8209bedc6153fea66e05cf03d7d1fd70437329087d3ab06c453e5e937b0de504eb6be86d7e84b4c06cbefa7f22f1ef97817090b793cd724c15a58b56b1a61033;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h451be46f5a1d1023549c330a5ec3b7cffa4abf9c5a14e295001dd5011b47052dab80900b69ae5e09fcbee06f319e6b5ad9c44937e21a113ca73ef988ff7c5f05b6da373c992f253f5ae05f21c6919813a1cc30307176c699bb4c53d66d0e97e68252e7b1dbcb869ecfd2e75997969c47f3d47fc40fad64156b3a5897d65b8c37;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h149cb08ba5bef0974024d6fbdaf06f1801c6855efc99dcf74f62978b0c286a90530b2d43f5dd64e64be5ecfe0dec3ffdef4f489067e9823334515b04bd593e915461301cec5ac0c20b584f6bc003def7e5748c4289773d530a8b703b5bbbf6a8bf99244467454898fe4fea33d5f22a1747657a362e37314a861ea24fb211f4d9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc12233ab89464cef5947edad617154ac8e86c9ad9c94631aafe7fce60cac21f2f13d9c853ec3e470dec63c8130616c321b4b3667a244e6034ed034dc6c4c23f826c22bd3d6df73b6bc2d69e79612c60292a68f8b53be815b5cc95431afc11638f569302ed45c621505744d0a2c4682d55fd11b963b940c16f4a9b6cd5a479b8e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4dc12ff31fb3ea16f33ac7cf44191345842f71fbd5242dbc750d49862b41581f8e541fc35e62a1629b99888d00e548c36b9d16de9328cb4db144cb36a81c7ef08d6ad770a90989f1bf810594edd205a49b0b06a6a2120463b97fc5b03e0f241fcbc81b7cb9866e2462b7d6475b7c84e572b605d73a857a0a9dd35d8bfb14df8a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6d64d70d5b9635bdb1c5b8825e41c5dd6925c97fd193f739962ce651c96129a2eb3aa24464b01de856b2bf72b049e68fabc1d396a4d345a199eb0b097fa1bdb80b39768867cb3d1ea695e6cebbb537b7f6828e18e162f6d90cff75c2f00e310c077eb1342fe27daacbd2d5a7bdfff80d9dfa7dfd62635e18163bffe63dbcf1ce;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h678ed3273c32686124a4398363cec79deb62571159ad2e6fac21b0ac705f8f715e61245d5bbbffdea74185adeba0e7f7c0c1ca1a10d8e0645c1e01a2b6b80fd0486e986e517c190df1a320baf6b1e5612416f2cbbc092a9b45411896ee251a189f6776e77ece0e477519a1fc0c681163a785c911b674cf8cb46bec757bc26bfd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6d047d8f7df55ed1eebd20a7f04c0737f44271b2b9e89f6e339f4e6f92611a837e3841332ccfe85dded52ec669196e88b895cec4ec27940eed789b9df3a66b59fea37f256cb1f8e37f83a6e2e9ad40e0f91722325a9badcfe87f959eb7513dadca6496b8e7da497045be1645de924a32fe8d8bc18493f3c457dac10108a86365;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf0da3d1d4f24ed9cc3fe50596d021416cc3a18b3cda42bcfd8b25a4240a8d8df01caf293079355a1c05c75d20d2ec94d9238beccc60ef79bf44ca9a517a4e13596bbafd0355503de94c6704eca35fe03ffc0390bbdfde46a61b64b1be2f626ac3d930a4424afa5efd6d19471eac70939a71c74f1e1cacf66b234ca25fd365f36;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7de6d08fed6551ea4d354131eebc851bc8c8186f457d8de38e5601793e72ee5f1f4996b6ab707ba3ca3ed4bd1868967e734d3002444adc2fb1f3de7a612c141b270914605b7b29c6d677513bc08db630e3ec84d1a75deaed82989dd93d36a00c5f65666f2dc926d336055fe76d2ed0ab5fab6e1057ff2239e4738eea30a5606b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h740e1cc73d8cd178fc995afef466a5ae63e9e2666633843648ac4ea21aec42b52a740dae41b9246741a6aa191abeb28a56007a1528596ca770a29b590bacd9eea958b0a3047a9621bf684ae0a0611b20a5d5617ecd8734ee526d23f2412b3f827bca5e1f86b1423a6661e0e710cab7a07359ba500e1fb243f1ebc116b7802b66;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8a2418dc419542c0c031ff3025e39c1586252d893e7c044622e9a8faa245324f10113d3ac5cad3d479fe79e8b583d377ffb9f52c3d4a9ac23f90b96d2d55d1d581c80ba3c8c742cc1236512e9e22c62ae012b1af2d6b2635e34e3a205ce7060e52b5fcd567758009aad66a12b745e7d5f1c08a8bdf861634c5c7d5e2270e8fb0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd7b3060012dd67c585642425644bfda2fc3a0038a4e5fa3aa62044117c009b5abcd0c825ffadaa01947df8f83281b3e30b81e98d97edbdd7b8de1aab0490c42b34a6cc887c89933c7fc44cb53a4cf7a46168c2762e90172e949b57c6794afea5f4feb5cae537af9ca9a1dcd3df1a39823c2778e760b62cf648a9c446f82e030d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfddc5aad76dc775be294d07bedbaab00285518d25490b9b389fdb49c794ca17312708b8672704e09013f153af791afd5f2b323dbf87ed4c7cc6065fe03a7796251657f17ee855aa74af602647729a108359550db63910777962415cca00589dbb8202b20addd580fda091e030789a59942b7c891a6ae7a612a863a680b9c8801;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h913196a1fbc13e6598d1a2a75a67794d0c47e2637c07a00f8f2f897e5b92b0e3ae35348da9cdaa7da0337dfbd6456b3b54ed63f6ff3d200ccd72b1630372653fca6afafee3076ebc3c88c1bef1150f930ca1d2b97a7fb51d3c44030b0e886036dab40e9862e8e965d1977616f5bfdbc1f0e63df426694f4b1d701389c89e0ac8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h15ca1a4923af299fd951fbe169797e7b39c7c12d3789c24b2aef94a337ad875329c1f8249ec24526e8d7a1c04c101d137359d58c4f6b173e88e1a8261c8adb10a3280817c74ac88d8d5454e6e0ff208cb56449a036aaed40d5eb40a93befe0083ad400d0aebf32ce23e1f7492a7305ca2f8e1b8265c1660dca9d9c8a73cf1662;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f192d9f1bfb55d1a48d522ebd5512188c4717437402ae14ae43c7db84b6dc9ffb02514314236d888175692b319a3aeaa3d3ef34adc1ac84d38941d85d8f6859897c3895e2c8034d58e2299cf2f135c97bc459909d6fab6e17bb8be52bffcd5e96f0cb6222d33ccd7a8c6b3854e51667cd039276ae5ad49aaf7d0e75f2767b6a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc0baa51e8b40521b3eadadacba726a53747fcccd74522a127aeb2e873387cc506b47e4603332ced73d5c9a24278748879dddb66b5c112f13b5e1272b3ac68c11d69d78ed2502622ee9db40e5736c9b6d1d07aaf6f1dcb8288b1e87caca27e8c9268d7f54407486241ae8c951d52f716e7c319f6a52f45cbd1d35728300ba983b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha76c6cb922330064458d6b3a8c1a8c5663d997d351c48b9657a344fc82cea581588024a5fab73c9b8cdd1205e856085a546abebfa2b772c19a92ebbb8d6449cdf78c4d24dffe8fc1fb04c6fa12fc233792afa43037dfafa26a5af9c6a92489d1967e7ee4d839bf90c39d9948beb82c30aef384b55b595f787c28295af8322a43;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4c081839fb2f8006e894d8eb17af424da923d99d0adecfdd513375a0678caf3e73f0bce0b9ad84b0fe900e78932a2bf3352498d85d16972ccd43d348f712bd24fcc1cb1b5916cf14632180acc5e904b792f2ae50ca81535c8134fa74d69fed739fb42ad2550e9a3b13cfd660ed7358e7786d4ae0b48c04f83514a124f469b083;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hef4895ee676fbdd0dcce851e5cbfbc028799137b7ff13b88f53faa966c73ff307e64284a21e742fdb0858135622e1dae9ed3b3f3827a9899376207b231e44174ccacae58028959305878d74f97608d82f99ed71b9c1988e8926297793f26b5a14a08bd5f9a836c4a151e1c1f13aaf6d15a1bc1dc63cbd4c188b893594f852ec5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h135831d3a66eb87dc91cd182d916dbe894350c63f188e899e75c3a1bc2364beb289aadaa02d9250531a9df447124ed8a7ee7bfdf6cb67001262852fd7ee43996003ce52a48dca49aa7dc4f90d4c365276ee9e18542357c08a3e95714be48a97540db948b450567c4c8c0e316bd62e578df88ca4c15e59f482af54172fd055987;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6a3d9ab66725ff7e46fcc601f14b4f8c2d6a8f826c6f09a750b120fc4f5d90f678fe6b67b9f62fc9ae2057ad7fbad6b90bb8e4d151508118304af8c4ea104ccac10f5066489312520b45199d37fb1cf4c4127c7db8073e9465dce1b918eb99f401d3a271e69b56f6805d8d6ea3c045f1a2eefa130e99780ad5dfea18df1c3657;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd43b12780e715dcb9a2a21596b9eda24a8a4f581831164a534270f40abb702b4568e78d296c5b50739beed9ddbd703945b6f4930cc8acc140954acc64c17a3c978cc60aa982b8a06f6d259e9e41b19fbda590a253f4bbfbd07b12e63969eeeda29f87626229bffbece2ffee80167c30a53af5917d8ee2440fc4190ac21d05315;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h283d82614261929f96dba122f0365c7e6cff25bbaf82ad5d2cbc63167b06873f806e549c3bcc4ad89282e289d2e8d4ca83bc973b46bcdc488ef5a552e9109a1c46cf08d445cb540d1b91d9b27aac4845450acdf99daae8fdc94507de4a37e352207de6e5cfbb7cd7f74eb3d3427070baeb4c6ed63a195ed68c4b061c33e2ac28;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfa0cd47ed45702efd53adb6700b1d5ee3f45714ea7d14c0150821216fdbd6f6f366f19c1b35f34e022df27d04b6d186c67b18e5c7b66eff6ffaecf2911847b600a8a9a6f5b888e65dad0e8723126e54ab42095293c55c584e33b00f97717ffb61174b26c7470a1b99bdadf53a18ec8bf1689706f3a9035b38ace442ab6af7de2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha4e145233daa2e53e255b80dd8b6151f18814c10edb7943e595fd7f6431b5f0b450589f884ec295007fd65502b494393793286a7ac1b0272f2bc61cd73a93d8afc361dbe548f7270e77bf04219f92d52864c50c707a172e26ea37e48cbf96d8a0c6b8f6fc144ce38fc176ee712a9a2745cd5f7785d438f643ae446adf38a7700;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h50fa3a29d4f5e4c70a6325ae65509b6cae911d89917f0f525b4b6af6c9fedaf39a3e10f9ad2e432ad660ca4487954b9852b4589668720f63f0c4d0ae5ae5fd25da62608a3a5420aba2551ccc4f34d253c5be54647346c0810c04ba1dc76aa049f0038a0c5c059a28c342f37ed3c2408738354733df56ac75eabb244fcd3e8c65;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6589d8df0e25b47eef81d1b042fd7e80abaf13e9ac5569457d9647372718531a85874405fd2ea57c01e87bef57939e43ea82ec6ff877ee767e6f2089e903353f2ad52e817c496c0fde65476b00968629f594ccae10c0017024cc75fec45c4b4a13e083b3bf35de49006ad25010c78b3743d569a9094eeb16a47cd9122cd06a74;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h900fda50860620f5ec3f8d8be81a85355c72d271b253bef0df751db7c7da699fe5e1f0af382d92bbbfe0cc68a99ae1179af77b9371ba27563495ec887bee9607b1f7c566d9c0fd80007840f8f9a3f061f54cb7b6f04bac641d17d465a10e88e23f617e15922248670c4bc9a171c2aeaebef2ee6a98efa59079016e36941386d8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4ae91c7e72036c1153042967b1cf1add5e10b25f7b24795a76f20a5ab6a7ff327020e85ef28ddb3fb94a2bacac730b96b252de0ed24a9c35bfef9af5267210aa58c0aaaf4530fb89c99f63b27250c4dc010a148aea266870d78a76c4321fd66a1b154dcb5f2aab31c34b0e5592e82ee5fa5c30602f8f3ca8d8a45c7074e804de;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8ff65f3ffdcb674c5f88e6d27d7cd20d54a052620276ca0800f7b2a5f1f9a15c9e95bd223dea1a42aee44b226c3dbdad467ca7ae1e217b0d26824edb6c9e1a86fd2a7df936deb5f5a746e40b856367fd296a8e9dea710c4a24793d3cf27ee3eef8cbf2068dbce7881fb0ffac62aa50531a8edbf0a3bb6b3223eef395a61075a7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc298e30841790d30e04348af502f910eec144f3988829add147013662e3c1f6d10fb287f043a85854dafb9af33ada0b6b9cc5a3e644c06fe8e92dd2239ea11a94e205e1a6bb38c13112e4cce1f324241da015409fbfe59c2ad6e89e3c8c3b32bb5a61e7abfecee6fd02d0e6733b07eb28524f3c958ef1900f2bd83eff35c98f4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc0bd91d8c1a1e78f916b5b86f535ebfaf7624ec2520a699d3af7180de34f1a9f86bf19ff832ecb842d9172ace6660c30483c1d9c2bd1a44154bd8a435e48e187b17e53dce4014b33ba62be3198c4f1b65a6970507920f5865df2f73e18142da4b74f2d044e8d9c25659e922f1799dcaefa1ece4cacaeced4f385d0ba5fc9bc41;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha28f3e6130976131f5196687c2125ea762f8f0a8924fe34488f1087d8035b43b0e7417a504b079bc285a127fe030a60ab022d6ff5d4fb8ee430fa6bf65b9b5a6f5d5b532ef0811bf4286c72bbfac1be352efb7779f17541b9a32f322f6812517d27834cbdbeb095eba99da9bd61bad09f3cc5841986ed21fe631bd9c11e95da5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5bc8bc6511a4f3160455f21ee0bee725d32924330d44998c0700f7d115850c86a78624f2b1945d3cf2fcbd3e0790922ef43e9a8e53b774a91b0b61494b49b8b94efbcd69f78b52ff8f1c95966e3b6966e43a5c507d460df832e66d20f9f5d7004614742a6cc6b366f45ab8df37b5d900bbed86ec2c2549c6a0506166104b7cdf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h443df8b895c29eb2b95dad232f5c32ab5b8d75a788378862185c23aab61f011c7f19412a44c85e6433ac8c8b49ff47ae48d005c1fc1385bf60e3b9aae181747d64ee2c0d791e541e8f1fd31df9397b0b844ff31635f75a3e0cc80418fec7c6852e90ae1968f8641e55c8096e0e30dee500be1ca7053ea2fc9c6e31cb498ace01;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hca469ac94cec329092e20cc07845b39bd5ea1bd54624a933759157537a24d4b0389601a23afc4ae5cd60862585f2c25dbb1312d2a6d11305cf5e313696b42d137443cc1e00e7664fad6db5a7902a743e8c615a05e15a87e2e3acd27d3e80c53176dd1ac12e4a0bead232fd79a53a215ce3b07a497d417e5900c38e960821d673;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h25ad7588db047edf7f93c792f6303218bc6ef230de11072aa4085dc8dfe96a80a768da3aad58e9fa3409aaf657c540fa83db85e58cb0b9e489ae2fca4b5b95289c823ac033832788f354333f2d460baebc5fe2544079f6d29edbe9cfd7d7c6b9e44ac6ec0540727c25017d7e3b8e4e4400663ca36a96dfff6f62067cab2fdeab;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9258507ce29d66fbe15d10c8b93f90d41134bf30177ea9ccd1fdba1f47a6a6aad2793348710638823a7f58110f0dc09786a59209b956a20cfafad12fb2d880d61248350a07ae5eb6052018685619ed3676299a5af4b2fb12266595f849f0dba3d7bc5c7bf1f428527c6420f0441bd2eceba002e3d4eaaa6a67097d94d6a6ad4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha11a03ea11e1a951f199120cb244a4f4be8a94e599617006abbff651e965fe639a094a14680aa99c77c70fb516bae6ff654a7bf747ff5afecb4e70d93e9b7c9ec9506d4a9bf8c9508fad7aa16c86c7917e4ca2fdf7b912740c50088587a98a1d2c6bc25df104781d1340d8890e4f1778d749e11afca0004a943381519cace2be;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfe76d640ee72e872cdbeff2dc535751c311427aa4c297b0538f3cf6307326ef0e88229e702c85d10ba0d0e98d79adbc4ce860505fee8431c3df64beab98b3d6b86cadaf166ecb634aa161ff9beedee2923d6745871fdaf442f969f5fa1433a51669d8a55fa322858de83594770f2f046b61fb5aac784b02991610e41af812bce;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3ad4f6b21adce4dd532378905f7e2fee7e293f6905865cc569e108beb31658f36dbc44cee04c780b1a809b867b0487dde261dda0a2439bac8c55a83478ad553a0605b374799105672621b146007386fe75fd9dd4566493271c87f3b2ee46694065d0fd06d670a1f6981f1b323a484a19c0d832a4877765b49c223185057c991c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5afda9d79a0289c973d46bb8fb680afc8e36060c9acee3900db657469a792770913f12025a397d73807a5c3a63123ca6076cde880d4cc77f2cba0763cee750aeb2c5b589c1ec11e2ef89b4440a8db809c043382e114ba42d5ede17c9f69fbede00b0cd1f4784364d4d4ab8ee835ef7ba5059a16e0bc5bf23755adc0143dfa05c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h59e72716ec1f6927f31791cdc4f71fe2d33271c809aa898018b800ad4c878495c689fb6e570420fd404abc85aa12292575a0a2ab2774a20b43efe382df5e4f4cc01be751c6d7e02aaa6caeafde5da2cbd55e4ae3aa63ed48f2b9bbe87b58d862b5a230e0a2401e2c9a1ffb081111fb611d42fb7d09d565b229bed4210b160ee0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h12c715f7cbf5a26156740a07584421009add9fe12a520a4ce1f46d7a7a0fa09e85a49ebac78401c099c06d2e4d0474075d9f66e99091e023daecc369d59d3769cb1917e206aadc2e9f839072b2ca0707fa603f7061ae652a10338b5170cf899ce016238775697a3cf6c608cec2097e34efe6d31c2039aa7875b1b466a3313780;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6969d6e74d1e30b78f8f864a8788331b9795bc156a948e76d801e74afc5435e589385df75a67827878af182689f5ad1b477c44f375a848058a0470a117c3a0558ed4c3aa345288c67893f2df0c7b92ad2426cd9defb5a78d2e68a39a23360f17f26198b1eab884c440c9eae7c59db8b863249a8d26ab0d3ddd1a90ef6e1da2d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf1c91c5c8e6a02fc32fe2edf2fd1124437d44f622855acf3a9b6a39748d05e2150788206c54cde273543d47f4f257640673dd2f390a15942d6cce297e3b0f1088cb12aa67f36c97fcd0d5be3912ee2aff3e89d5d0303c9a202232e807a8c43091f043b5ddd5e32e1cde5ba0a4c9da87c89d7e8cbb36ebfb897c24fe0c927e4ff;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd30b1ef27502576e21a8f84584b62f962c7cd65e14d9491c7f9f593211744fb2597bd052dfd18103dc6e6f4ecc7d6f6a6ccb1bd89262fa2daeaee595cec879fa227f9bf249cb4d08ac9047e88f0fa15b52e0313402fb8523cba88561522ef5544853d0120e01976d54cc2da8d2e3c4ef8b4f039a8568eaacd8d82893ebed65b8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd5d76bcfe3451d8056287a11126fa9c146a75b1b742dca072960ccfad2776e26b700a088ce5846cb6505cc3b4451b3072199ae45f547ebe55ccde223f09c7c8bfe6d651beea548613d4f0a65777abe673756856695e4d845c4e743ffbeebff456b1c0e2e30dc68096548757b48737d990cf0198faeb0f30d7281fcd33d76b620;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h32b7dcecb2aa88cfdddccb652dad746bd243d41b786347cb2bb2ea89acdbec564d02ef2fb69df05973a1c1def5e63d0899eb87e6bddf8f0fffe4166c6486deef7c17792992ed50a4ddb44125db1390cf06eda0f4d4992c07037edbdf84d1b6cd23893c523c8a21e8d00f8eefc5a9402d64425500afb1b88e1222e4debe2e5263;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7193bbe520c9fd2aecc687902bfb413f7a9dbc1d4283e67220388f440d08e8e887007430b6b12654811ede71172279bc73086817517453ef8ed2a9bb2e4f8b218a5849a9c279affc2429bfadc690ba2436705acb1259b6ada9d3ab5fc5ee4812d2c90ce2ad9cc025c83f7b0dc22e3935405069e2c2c623a0b45ce65622200f13;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d591c5c13577eae5182e9b278124e72cb8bebec0efe010a8dcb060f4b0d7943f8142637dcaaea7781e43147b6328e40c599c3013bec4651eeabd9c2f3109466f6de55b409476aba840be374382a9aed1029de165ce0e535fbd09591ad667d3543b011c0cabc226c8bda98c61587bd2b9a2a383a57b8de4fd7edb445277d74ac;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcdeb4820dbcf8c1a530b4e8ff98d22ab8310d79dff03fc7639c25abed6a7ab2679dbeeb1c6c8e3e6049006047f3d887e253ec439bddc111d0b2f898ab226fd6004431ee6551928d011090592e20a3510f59d7bba7147fa70831af2f0d6fe659bf622694c3fefe833e1aa698b6ec4473837851df21f7dfe28eba30ed932e16e8c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h137cd78a9d48f3f23a91260b00b2a61f5b7c25622c65344856c3d836637c81560c871bb954200aa992877bc8a9790385fbda15c9f75b56cf973a8b24b0392bd2238f8463e31b0d368a8c34c81330aaca906c225987c150e9f1e876f1cb8382189bd697c9f781a1ee21310b07374ce18863c66a68fd52cab2a31885020d2874eb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h70437d6544d209c81dda632e6f0a78969017957019ea68367e052411626b399f5e63f4a87c28476ff3a4d6628ea7ba93de9b97091e27ca7c925efbbd05b1d08378b9c31dd7551a8c4ac639fc311b9cb85595cf87bf9bcb213fedae18a35f363226511530b0978b9726128b00d9432b025be4968d28a5a6a4c4b87f07e5e2c0a9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6a70f46309faaa5097c8a944760d81121e18e0a2ea59c818ab5924937d2bbc95e3cbb00e91d40d4134fdcdff0199565b148dc5ee7cbb77f1dc6bb91cd21f0041cbcde60ff7366b5496d2cfaab5bfa67018bb351889ce087f808c1423880f0fceeb44a4abf4509d05f0a5170b4c78f309609233d5df1a62f721ad9ab617883e1b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf232f2419cf1ff2f0cae17f173b76b2a942315ad1177ff8b1656fe4decb6fbeb0e627f8bc93ab6428c4be1f998cd937f14049762a48a959503fa43be71e1142142324b7f489a23e78de0d61a3091e3870ba76cba7452fccacf34f9f083812522ab93a5cd572cb7b5ba019b2d5a93be88f0f4156636d76579d00249a19c5dcba5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5bd328767427bbb4aabd229a939ed71f10a395f7c0447e75461502f8be3dcc91c186e08cb4982ef85644f11ad55376ea96f2a4979a035f9654f0af9ee97f9d704c7e49984702127b9bf17344eb631b8b734cee9fd87b0cde834f33cf05c5745151493f676ef58ec23163f9558045400d880693e53fbd993c8a6920d18bca0c39;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4781cca97037259367900f8d7439abf175ebad704d4d0e7ebbf056deba9e0691c8ce93de8d26b9c87b0037abe08c6444a7071fc3c687816c254dfe0fc3ebd22bf076eee558977d2afaeed2d0f47a532af2e2613ca60d949a10ce39152753048f8e272489d6a922cc35e0b04fcb3021b1e12eb726755e5105115449b3cdc20ff;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f627467ff0e2893044771e9186329eab3d91b17466cef8fe42ffb17d3dbd58fb7a2154457c5d13bfcf54f7c1ca687b193560408f80929893f525362b2fb404df8b0b01bb709266dad9b9f8d03410d20293a8f74f8b00dd8193b3751dfb56fc60ef091c7da56e1cc4a7f3b9fdb6008cb4dff1def18334b686223511140c9fbe2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd336f6191365103b9706c37505d0bebf695a04cbfa32daa8d924b87f3476486f331f4b959b196a87581e0ec0a8b7999b6ebea275b4af61696940a723ead75c2619ef7eb491b8be05a64b6653fdb62dd0111c38b8280f44447124a83cf3821e4e13b50a348d5acd692eaba38d9dcd577868befb0ef1ed4f782be70aea1a9ced2d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc16b523e1ac60d618ec9207061efaba345bec100e089bad80980a27f2d536aff8b53f590a6eaa6a8d95990a6909e24769040c276f67eb04316e6b7497fbfd602afc1dfe6c3a46f312a5fdc750973f481af6471e28d4f8dbd6c3c8ce6d96cf8b4c6e69f12c6c573add2bcae6982308a33156fc8c448200e8e5c582ca3ac572ad8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4b0e3a31e2fa99b8a71b095a242f403a7f36cabc295e8f8bbe71982a7dd113dc6288bcd55e4a58ab11e44aa8ab1dff71f1e824f891f649acffeb0561de3748a2c603c0b226524f7478f4f1e86ce3dc2e57ed5a132f5cb175938645bb40411a360a2d18aec857891c12d97f03f426c1888298b030f923c60b978c2eeb9a5c4ee;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73aa8de7db86a6961aa06e6d913040fcc912c4874e6062fd49be79eff0779f6558aa82d5e88e041dd3b7e5f2588e88ce3481e7509f6d1d30edbce46f2fb342334737a582e2113e7a05b45d8de61da477815da245630dd3744cb4970cc39bc24703f23af47639534a5eee36e8bdf2d3dd50b44e8b07e533a37d1db36726650201;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8e04f1b96a35798ff166be80b2c1bd6b32116d774ffc501b0d4879c37eb705e4d87879b17821394f555738b75c7723a43379e1a28337ffe9b0ddcc200cb97619d964033e8a02ec975dbfa2ed14291528738a535d2450ae0ef5637508c59d6f240986ba1c5de97cc8a977e2f9bf0890964c21c8e56260d76016347d95acde0cc8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h36de72a26516792b43680b5a88390149d12d6b37323e2eb96bf6b879660cffe5e8d6b55e16673e72d7278ff8eb91e39c6cc49c4b6f31547058ab4b4c91bac5b2511c1dec2e644927ff5a14459cbd4bf7e39e8707dc60647e8162d6df2da4a7df41e740d86bce5d0dee202810b1671720950914152db0cdf85003585f94f85b12;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h66dfcf3861d7cec06b2eda56f87a12052b0e563409cf7633eb46a171162805905833907cc00e6740ca8aa0ea7bdb4c4ca5b0d5420999292adda846b9c2a4fb10820d1364427e44870361f8cd803ad8e68a051497003a30556bd3f7bb19dabb30a7d57e163a112690489dcb7e9c9743b62b7e42cca9310e9827e99da2e8951cad;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ad751d061a5dc826cc175c929b3e2e7411961119fb4596f53527da9eceb40c220a1f8c9cd172d838d728568ffbaa10dac18ab29df1d5386343d0c119eaf4dfd8a9c6b63b22a757c612f5cb590c834206d148a521aef800c01a042921dac7d11a497e5732db4a91883d620fb02ba79c5bafd391630122b09097e596de27d8f94;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h292a13778a6fdf2113f77d74c3a53c2cdcbe32a0188b9eab9619ace6d18b13f46ae273ce118d46424a2aa4619f351b34ac826120014e9bd0c6eca6b38d105b5191d9c4f5b67c1eb7640d0c69d8e49399b57564c07b7441ecba39c5b8eb8d4bf01a59c4e36b8e1ff5faa0abcb86309c44eec6ec5fde42cacb0e426fb153f1e0b3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6b92a9e1e8b5f53b25c2fc96ca0e0e084f91b774f5d4b468fba97a0b6b2a08e1aa5d6099e4ce37798dec5cd558699afcdf5984f0b3aca94df3f026d41d83e4df9429094384fdc1766b71bd9d4c277209fb2267f4d706788742642a39123bd3d7fd74075670c09dd8b60ce8caa34211437fd93de8bb96191d5320191152e69eaa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1389ba148f236cdeebcf9e5772b7f93b6cb8b00eb7dd8452447647c23368b3cd380e2989e874f102053e3bc0c187f23ab8cc9dab56b353504f0f6a21bc5cf82815cca363a8581719aebc76980eba3f60ae6988b8028678f85a42dfefdeae29b3dc5d9e8528b99faa00e457c44f827e654b4e0b03a6b9d904a6d091f70017a3af;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h62ca80b48b1ae8d52b162a4dbfa8d406d50b2e66a7b4f6abaebd5370b68353834c036d3c84b9deac9e54c08f2de5a07e512981a65f18cc14bbdff5c24834c31b3165ce75c3152fbd66b9fe9ab7641c98cfb8a26f779215ac0fe6e87752ecfdc8888d17cbd14746a09a7b74c8b08d55827bed01707f4fa2fed27cbfb63ba2f397;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4c3fea423fb3ef701cf3165980afad94c70bfd3aa7cf1ec4613d2c168c2ee38f9217bd50fb1b791000f5594c61a15181d3086aefbb84e5ee5e24a895c22a201829001d94befce4c29438d2420c156a8e47152209ee5a023f63350d4cf3634420e10cb6adb87c3286e952acfc9927af7872afab5ab0c29a86809381a0b5e15fb6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h90ca0e45eec287fbe838673bc9a983e6a5789f719eba2fdb5db4abffe16d0d92cd6c85ebbcba30f10624086961c2f9bae2531febe91b8b1db8be5e30dc16fcd556ce8bc64d16fc77a836affbef36f17f6ef6426dbc7e26bb5405126e4e2c2f4f9c38c11176950ea920dd978cadc3b815f5f3370398f88ba4541b31c437366853;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b260edda0d1f7912502ce0dd75a273c6862e2fd854716d0972df2fa2b2075a092231185bfb7e3868baacdd65ef7ac6f41ca88d995b288b64fa92f498d13edf23c9e9b12f6bd0c759ed9398329054fb19657359abe6468ae7555ffae2118e5238fbf040c39c1ffa2d3d5b20378882567539cb73084576a7027c6a12072a4133a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h454ae5c6ab0a116a4b4d8d35d55b824f974a520de4baebcafecac6c1cd3d793de350ae09c9446ea7e0216da07c17d7089bc97757f2992b8fbed95ab8fd57b6725472faaa45f513ff51f00a49651411653881970f819fe79514c6d45d0d65aba598c12a1a4524ffaf109da16f164d362910a2987b8fc472579fbf171ac20776f7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbbde456cb84c47dbb86c2f417f058abc00bbaa7853087762b769f1bf61fba5177ca09be1e5b934a9abf8d548e90ed2b76099417735f9baf486112adca32378dc83ecc4a531f983ce5b43adfa66f08b796d1b8a1043161a9cf6ff2943ed6ce6187693ab6c77e65baec7263ae739d531e59c88c1a45db4de757fca61ffd7a58bb0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6b4f0506459f1b95f211191b4e081957e66a300d96aa26ea5d6b294eae65bd4cc92787a77c8e0d83d0ac8561171165c0a926a930c85f7f1bf300f36f8495fec94dfb0628f1007ffc3dd023c3f282422b6ad376d52e9d0fd2668cb58f4d8a8801a7c07bdd8249963594f5f306bfcfcd75845c429f8ecf9e0f51a9e4c1581b2ce;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h314f3f6ab92ce623ed317e45f3261db8877a9df15436bfa23bdab2a60962765e33952c5d0eb1951007c8daac918bac6556fca5896ea27bb94ab6efdf2efa46b834a9520b59f8860c5a4aa87b1a10e331890f7cb9bf2c418717fbbe28ea3b2d81f6d392de01ba499f44a9ef9ffb65f6b4f789cc1d26cc5e1abbc0c115d712dde0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4b8d753a57d17396988c28ed426726ffe5cc8064bf6155b9b8e954d1ec8488ce24db6f32f78c046d507491880bb6df4ea151d9de265aca213be0b9142801a30736d33aae765313d4fd0e1fde6c30bf207466cff0b1e6280e98998689cdbe53afaf5dba784c43158f546905787cea6af6d0200f9f04ac9fbc2deac7d0daae24c8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd0a1ccbfcc566cb10b481a114aa6e7dce57b3139c37c0d3e8084e214c23f5232be2c7b3624b08a56d258f99c3e433180edf02e51acdd4147007d17f4a1e938e7ad66381ed5aeaf695d3f3f0380d6ca34be2ec2ae5b6c87c2619dd4871cf253d4cea037fe7c42630421bcdd0cc9d2d9723ec543091e2e1e9ae05fcad05c42cdeb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13b72da3efad3e9c2a12e23ad4d5a3a6b182b95ee49c2069637cccefbf7c932626e3996d3177f688d8223b899762179530a9409ba30d67f55690b46678ae0342712a5430c01ce07a51cc7582616dab2e28f29ef33c5c96eaf2b14a051b286cc95440b8981fa822243bedf5f965aaebe3e69a009359470fffe3f54490fe6976f4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc0b3936be2223d08e5044ce24bdebf1626f652a226f2a37d7b26593be5ed2b5b364676a7c23b44acf04ccc8079005b30d29d785a82da990030c681c2ab343cfd291c8a660b0f6d048afcd623e0a2b668bb5709cac90315d87ab824766e4361e1bb7b2d12b6fa8c1f5d19b9cbd8b19c49d9899aab8aedbe163a97fffc39bce673;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce231854bc33af5655735d65f1d1531a4ff9cac20abc315d93c86677bccce5e379faf155f605f11a52e00d7cc0e111eaa65a8751706df552e765f36ea0634722a62b041238c34446324b424de7c979334220e75fbb6a8fcdbcd1a72b2edf4c9bcb3e04e0c048ebdf11c5e2c9fe2d31ae10d5e9e26172eb6c4ae9cf1ca4f9e64e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6cad43697a2d697660947c65aee1bcede1b3f2a546e450a7503dd2c09e6d315757c7482a9c647c7507910db69d9f923ff96317cb4cc62faa792ba85e927194f01f0714c2dcfd9510c9caccb5e272292f10102457563ed2d6f7cfe32f06d769274de5b1815dc9e467ca5b4407c3b0e725d2bd6a6772f817f1ea489a79544b916d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfbb7dce12f80c471ed1e6b40a0b5f769bbeeca52a14f98cb40ffe0dc7737b48c42a4c1755f581a959f57812b674eee1afcf177eb4682c50bfa3d157c576cf97a1a3f6641d273cf809214a51f16a3349f83bb7200cdb35e1f430f35ec92f4f675977d58f7875a83ed1745d9f5b1e2855d5ee30afacf7e2b54776dbc71718985f9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf61d90a2777ad185f690c74764a0535288968fbbc116eec5199b75ab48713cf8466a79cd89abeaaa9a76aa7aea9ac2a028ae3ee5f2be54d46e022ffd96a9753171e7b538df8cca7910114560a6dffed8b659f94516fa2661266db06803672ef05d79a4f0602c2c3da17a8ba0a8847dbd80660dd4483d4ceb5f8f46214fb6cc1b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hecb4cfacd36c2b7322a21a4da767bf30146d3318e2b5230cbd7d6ecb4e19bf841e874c7e874c5b9a702cc247ddb47de345d7c53f438ad57f9538e0885ff6eae897fe6260ff85837b0116f824ec90753170883790aab5e1602afd26146a1f2916dc334f24370a09fa4d4215981129e23b8d6d3f7791a3ac87733b7129ee1418bc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbae9d6538efef744cb1554f1df16605b0ea4fe5af8c6f53322caae679b7afabdc23226b10e11a730e326d40ef21ec5f62723b981faf2bd56f9793ebc7f1f9cb2520befafcfdbd57b08601448667fe26c64afc331479338787f815d487a0cca63f966be7bf5a4c60f762dc0a9a7848e7b789408b40fadc015946616f0dd76cfcd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3be527ba600281aad64241bb90affe233a6a4fd575923d0cf874bd6fe383f10e7ee95ea51f1accd07c57dfe1f642477a416000afd426a956ed3010587228688a3d9dde28b19d530119415718f5f5a01ba7dd9282e9d60a63b0d34f598019db121e257da4442b6a865dc01b31488effcb28c857ba3ea7a207b6445f6701e0c448;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfffa510411e1078518d924f73b49a774b6a1bcf868a407ebd228040fd28af765a6a1a3c7d749c42a180d30ac87ab9113cf5fc7d1c571fbffbf50ab43ef6c0bb78bbbc6e09d65a2147eca0a42c94bdb4c2c9b43df532ea687f0fd3dd210099c9c9e68c9883f85c0f460c141b84a25b2280a244cf228193da6cb0f7d6251592a43;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc9d0369c07166b89e2086455366ce0c9e4de6e64361b6ff4a35e4331e7af37797fd8c66a5f58b81abcc478ce2a7ff9a716ae0a84b7092cab19a5e35cd3d9ad1cd1063598bded7e8a6314b73553920aaf1115b3de721ed16c2cc772845f78eb9356f13b8681ef57dd55f30db3055577cba0ab6d3c75a806623e2828384dbf3f5a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h83ce613125d4d9e3eb4483c4d8b280a800d68df6f1c85f0054ef011e1a7b5fb046877154ae3da5ad48223eed4413993e37ce6bd5b1d43a507ecb5ab5328a8b6b7fcdc1cde8d75dcd8ddc39ac2d818f0dfd22797c5238c169d31b7dd8a51350de47d13da1a639229790e34ffcf03cbcde0f6a731e3cc6398efc3de16208ef49d3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h87172d45b8bfc125b43016c35cd9c3dd75cd0196fd02ad9d4d01681859104a8af5dc0e85896757ef23ec11a45b642f2ef9b796d44d7d5d537167f772deaba485d2d90a88ef2e5d5776b3fa3d645bc61f0624e524b24e2bfa89d390860d975b4239e6a5e15ecb291c8bb163ceb03e9c56dbf9a1ab9de0d11189164148102a4cd9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h36b5babe6880faeb2c4f0eebaefe1ad3eb767a76bd21505c77104bcf3be26a1a7cb67e0fca22a2a69e335659608c6babecfc800db83391acca4eb5879a21d2ced237f473bbaba8385b08e3dcd4a65556af59c69107928655a87715f61cbf0b19531e5e1284fad38d2e2467c36303a65478c3896180e2c77e18ce60330246d6dd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfe5e1b27e7d38311d8fa2eb0df71f06893e0eb15c433a15429b56fd5b4e6502af7e42a078c1eb7fd371089b44470ae8ea6d84f5002041994f4c7b41507175213fe9ed0cccca4ab6eb5744141a06ab05d558c495f8c424422740edd6190bc2dfbf63fae1c60c93216cda67da27cfa9f45b9abad8804441e993ee9b2b4cabab3a0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h57fd0272e9c6a596bda25e199d67cd796e14ed814f3b2f27fe593019b2dce8ea2ed71d55ffd2a3d808bd726ff5652278b9b56decd360d4f75c55d318256a5160771571b0959068f47274509daa1b287c96bd66b6661283bc0331e8be90aad272d602db1fd2af287b473cb7e38831c818c1ff60144c81b3f027c8cb7902482eed;
        #1
        $finish();
    end
endmodule
