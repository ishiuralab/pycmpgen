module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [15:0] src17;
    reg [14:0] src18;
    reg [13:0] src19;
    reg [12:0] src20;
    reg [11:0] src21;
    reg [10:0] src22;
    reg [9:0] src23;
    reg [8:0] src24;
    reg [7:0] src25;
    reg [6:0] src26;
    reg [5:0] src27;
    reg [4:0] src28;
    reg [3:0] src29;
    reg [2:0] src30;
    reg [1:0] src31;
    reg [0:0] src32;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [33:0] srcsum;
    wire [33:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3])<<29) + ((src30[0] + src30[1] + src30[2])<<30) + ((src31[0] + src31[1])<<31) + ((src32[0])<<32);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2e2e9b2e82688b72f90cc09efb67a631b4376c18c8584123430fcf921f3b41307d11c0e1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h172817cd90be2bbb365e3b00137183f4245ef669f26e61fdfede1292b98043d6791303d2b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hff176e8a7417d0aa79e426bfa1c0327ddd6f5aa91f4c2294e24c1085836182e348d04357;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h32b4626b7f75bffd20ec13cd78cc10f52f03ee42f9a1eaafbe89d7fa45e77ed5340fb031;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc71b38b18fb4955544000ee5ca3d83bcb234220910831bbd03a19836dddd8563484dee7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b613447d7dd2d168580b06da44f007688788b1bfcc27a02a5bea795454af5b351a95295f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18a393153725c6599c56c6e1ef1b1c5eab29218e88f8937c1cf9ede6717752a3ef14f9b42;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5db85605a31e53a47efad8064b6c7cd07a60721f717ef6866c2bbebd819271f6033ddc58;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15709124ab6231c5ee35e3ada221a760ad3b631bf7a373eab062c5615e5da7a5915622661;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hda713fc1ccff75142e4240c1051c06c492a6ae33fa9a77792e1cd5683e87e5b15aee90d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h44001690d5b50ae9d97ee15ca5adcb73bb87d1791d4009707ab293a542413259d284f07c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4ac3946b3d359decb150a57a7e8667cfaf32524f8e03e28e5d3e323207fb7b7742263127;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h145d2debc173ab892c7fe331b9e2424864e3043da8195c4bde6d07a08a5642ea4b0d8f187;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hadf8d6e37cf6d73f3fc48db8d22e90023ef95cd55a28365587912437b432b22014f1b4b1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h129c72208cf5fc83f0bb4747a290e7bc1fa031f8e444bebfb003becc39e48d5f4c2ce085a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h47f9f99b92ae82819ef9d0b84cc0563bc64930878e9b043ebb420c613d9771ee2b41821b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a976afc344a87883beee0a0ca4d8df7ed70c4ed42ec0ad1a6633236baee5fd93728714a1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12ede1667e2d0c7bd95d0add683bb0224c6ae2ea45e06c245c958d6c3a14817a2d482d3b5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15cb040776011a716786ff5ac6d7065938451f4a30cab96aba64f44faa7dc837f2aec9cda;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3550a8b27492e3a075ae48ca4ddeb39f07fc23f61c7228695fd6d9ea5eb287e9835cf829;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b7cc7da0c6ed08414705e55a4073f65f1e95ff74ba7d5db59aa979756d0cdca777d045fd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h58e717a5b6f3fae130e96574d8e9589f3f8f06d058488e77bba1e0d11ca30e3435337e6a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3e068168b3cbb3be6616feb93216efa771a2efcf88cb39a16a9fc2b535c594b5bc726fb9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7b3fda90ed85d15c363718c8a313c31c82f211313d1cc6f85081fa11c49be176484dd631;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18f217c07995ac1c89f15aedab4207fab108de21ef1688d07cec3cd7a7909c696bf8068fd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h45a66e10a936729a4b052a889678278487fb4946291b20e30433a43d0a63c1172e6b2fcf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd473fa21e5166ab0613b6f30c9c20e3f240332de933a29a887ff33d5af98fd98d357f905;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1012f8f00fe521d6a5d45446980741915326d67401128d648685e3580196b1258de4a167b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17f515c283389195b630ef6d8318e756b714386fdea2dec08de414aede250b0bc16011b9d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16c7bfddc353b464e95c6fdeb0be0f070ec4df162cc82c8611644390c7259fdfb71980857;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1639b732b275ce8ff5f2f0f2b597aff8b0a2484f1c491d06821d8dbac4b6513288660b3c1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h144790a2dba23428d3fdc2dcad18f3194b6dcc53d1e220bc9a354c437d64cc3b65f3c20c5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc1b1b7ead3420adb63695fd2cd77252f077c5177e4194198c6f8af7c07da0d8e81428be1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d61719dc60f8f734a45648c29a8a502d823a35e1f5b8ffdfd8e826bfb541567d301f310c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1702f29b03b0c194eb1edaf2ea775cd6f9f9096ca32952cab4c7899017173ae634183fe4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f63ef5b711489fabdeb7217c5e4af3edfe1a2f06f8207b9d4b08c0c95b105d3f42eff8f3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfa34f6fe0e2bc5b8ec8c876b57966d25ac52510d2c954c836ce17d56a4ada2e2167537c9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b5e0a46b0fc88014607957052c0fb97f27cb24924da3ee3e0ad901d635e3eff1c0d13907;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8abc3b05e961d6dcf771414cb881a116f2b027127c3c0bcf5c7412b13e2ae4842e95392d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1671a12bd3464db25b6b68023abee35fc4c4006b55955276b9d1a286ac32b28c4b7218f03;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h994eb9e3db87e2067f2fa0ccd2571d1985f6cb9f38f3f73adb82b898c5077203e7691c1b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h155e48b7a61fcd662117930be7d141067b781b3aeca7cfe1cd6f39d9e7bcf46ecce2ad22b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha2dab70144f760f86fce6d3350a5c0d3283d04f2071ff5f64dfbd944f927de38c06321dc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2551ecd2646abbca7e17156584eff7767dac887eb2afd64ab06d36511c82e899a7bf2d5a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h884d61a7d15943c5fe92a467aa8668a5003b4cd9230c5c453ff945f228780a77632f8bcd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha016c6116a4cbff9a9422c77a538501c0dc8aea62302546720b4ebddd264aada4526ab90;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd882f36065de7c37ab6396d4d06b4ecb754ea55a43ffa987baadcd2b0f0f14c4032a8928;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1090e405091e1555cda741c70a27760c37d84c1ebea2a7ec12fb116d6734fc2b11c628127;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dac6e6df9effb3681e1767928ef28a79362711a7e62ae0fb2c8e9c4a8bd3099927e5a7f6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h166d9dacb313080ad1d21133a27e180fcb578a11fc67ead0ad17ee57716e16c5714f66d89;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5c54d36eb6b44c4f4ab9143328a18cf0903005db61a7cadab76d9679333b81720fd448dd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha2fd074c39bc5abca14bc08933cc15e934bab2e5c4363c2e0398c1f804b035fd81178909;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e552814423e10ee3cdc6420abd2b7609bed892753e2fc6b9d79507ff69d57a1daffccd96;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h155d6d05f07c09fa50999632b2901e3bba53832360c99c2c3b9c7afdfefa39c543b34c6d2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2b6b4f40fe523dabd36119a2de71a19b3e0eba4fa03803ceb0294fea9c314c28efce080e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h131d73e6a94fa8816b63f1d3bb56fc9a4ac34cf64206db6bfbc03d079240e4418b8193f98;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10cbeb1fcb364a196db3786692f8b2e71a2bfd5bfb4c9171dcfa9881c3cbd35a56d0fb5e2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hee39a86bf4a97bf2b9c0bf3d23f45de32864e1a2f1830cf0e963d33c20c90232160e9872;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfd0e2528e8aec56c5d44d38f094a091edd7bb8b975f5aac382949f28ac98541cace09b91;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf083eece04f32a4b6d365a2f2ed2a31f6e41763f6acc62ccd527415861b879fc4e283dc3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19f03a81b3d8130f75d3bbcbc48cd4d97ad7d1273c469f62267b5bec826144c07b683fd18;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13248c0bcaa7a19ff1a4c84bd95c941f323565248c64b7879770dfc672c76404f1e3d3d0e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b72289c0ce9ab4ceb888b3acd635823d526270f59d3349726e632a2d04df805042fed540;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1735a0902c9476d9af6b7967b4dc848881c399c4a8a8aeeef7524d9d5177654b3dbec77bc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10445ad6ea7f7240a9c259f81e02336748ddbf778eab92883d273a089696baf4bcfa8c8bb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb825bbe845b4808873ae4d69b4103f2cb122b3036d2709970aeceeb43c7033aadce0b1bc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11481ba73b6c5b9b8eb264098e65c5e5550a9a8cad5d943667ebec5886793d8533a75aaec;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6d4f268b1a8a5496b099a538b9683b9be39643830443c2ced66cf504943a5a5e03a83244;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfa01cd512e8ec24b01d6d4c0ede043a4a83d617f6b6eeedc7cce2cdf47b82ad5aff53fb6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he3e865b1530f9ca15b1425b6eac604e2770f5e31ef35e50b0426de0923f5613780c50459;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16d0a0d2a1bb2aa431029bf1830ea35d79286704b7147e75986547d0a1a6e54d5dcea74da;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h185dd00fa370e9fa3a8dc961f9e9b791fa1437cd4caa720e7996831f4218ec64b25d45c12;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf8e2dc5abb906ff897780cc69b60064e791b47cb1746b246b17ad8e6aacd7d64b3cb8d58;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10ada240f36663aff4f977970cf1bda1b69abd0d305ca60634957eaacc00f9f8089fea097;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf9114bdc7450e064752e56080b0230150c9ec85fd49a0807885732220787a734991571f5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hea64d5f519d88c965bf2358b1d1eb40074ab4a5ec68e741bf939b837d6d64545149c1de8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he80c1953cdd4a54b8b184916d87ea1460116b034eedf11b6eb529a244173ddf73917255;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h621034037b434f2692cc98f57705ce4d5cb4bf6b2f60a0d98607e3082a41c00142e813c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11412bc6d226d609d915801a6e7494aad4e221f371c59652627fa3ebc1d6e7dd732fdfe25;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e0c427dacfd8700e177e3fb4e3aad54723c6c97abf47efc129a7843ab97f57ff2acf81;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h106b7ec6653acfc2e0288a246888169fd083b54fb951d380db5a8176e788bd2d36c353bfa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb4c6377208ea9bb6364ad58dd3514c908573a71684a342b465674e919149395ded90789a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a3299c3dcbc144cce0dfcc308e8ca846d3dfe52507f7f19b24ebfc6ca596b6b6e2e5fd18;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h131f3153b4231bd3275c8165eb93118650cdda39bff0f962719222dbdbf3377edad511c8e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1035d61fca8ba63bb4526a9e751b2c1a955ff7da9bf8d8831a45a6887fe25dcdbeee2e11;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16e777d8dd0b8787db0010050f4110fafee8131a6aca83917ab789cb066d7d04c80cd60f2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10057c447930e6ebea49ffe31c6c35d207a19d62b0a1c19f6c540e50394f2b405287a6379;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h56320f73cf90ff76dc48c437b2a0647e6ee3c286088b9096bf13a714511a9eaffa1a5fb7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6711202a5aaf8b9d8c1119579262fddab37ce34ee6e34f1e2201d610e3a5e6792071b23f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8994a48a394ab3787c76eb61598279e73bb3ce8fb1a74125d4014028ab53f6ca19a81781;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12b7721d37c4faf6e9d404f7521ad5f01e6ab3290eec07e7b379c82882669abe8d9796745;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aa918fb5ba3e6f5e087f765ef14a731bd311bf63a2ccde0851a776fa042e3ca0efb3ace3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha9dfa16c9b38a6a732a47d4ae8e3cf8032c33ad287c4a8cd3c18cdf327a1da0e295c383e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a6efa3b6aa6bdf7b17aac53c56f80c2a39a71aa494f5c467a6b7a3ddd18afb59d8a2fe3c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he1f66b6bd1904400cfbf274c2981f18524ceacd0919552d7f040ac7d18db5ff4272532f1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3de3023a836d1fbf7dc71e730e2fcca37c39df8599c415745cd32a462396b0b527f9e419;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h54ea6dfbd8a7a53f5b06709ecdefff7e076fcadaa70a518697c3df73789df21ce0ec1d7d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hedae6a125ffe1ca64ab0fa92d7ce9fca48846052387a18a538b0f295ee8ae53b6aeb0250;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19454bf388329282313a3061281a0072ef1c4515fc7aeec384d76feaed047b9cfe36e72ab;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d88abad765931cc79d8a33cef646b758f06984e770b132bf95e76b7119ef62040ef448ec;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb400df719e034dc34c662ed83656b9b1f0452c303188c541cf1b36d1b65b67252fd63f44;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1906de9dcef5fad0ce1af177371c5424542c072eec52f066541421fb4772dc9c59113d70;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18df77695604bcfdf4a35ec60b1190390fe2d0c400293d2e3b9f08dfc267568b08c00c8d3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f9921442509910aa49b2fa3ff096498116c28c777d975ee0aae45f4a0bf5ac9b488b4628;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha97c3b4e262cda777031dbc430dc2b40fba205f4507dddf3d2eb9419a3b13cfe45fcb77d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fbab4e423a817661750ea49dfe089234ea71ffd83563d1a72f4fc9d9916ec1ec5863c665;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h94210e7b688dfab2304a2a7a39f0489296859270cf483ac6283d24c41369a92fdc2380b9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h130ddf81be67d2dbc309f911621851f064cd4bec5f26244b36880c5bf36a1bd71bfdd4f6f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hec76a5b785573de717dfa852b8c4055f537a9c88bc5794a7f0086a20d7b1fce3e81b6bab;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14812c7d7b393c86239e68fc380e6b80bd2ba1086a9c74ff458b5aa1a43113558c7c7c0eb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fbe57fca1ef171572f9cb5a3a01b6c8207fd43dc6c05c333f16928e0acff3454745985f7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bf72c7804e83bc19e6440499dc4776d8054933b57699966a9c50ed55adbbef3ed0217cf3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h36f80fdc808b92253f440d23a3ae006c1a62c996c73bed870b7663e45dd5a43140cd5746;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h237f07efedd40b8032ded762f808fb803db6c2e34fecd960954a569d3801ac6b7370b7a7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ad7259f88bcacc57080e8a36d0ef8dee1086a1bb07cf22f3a04b351414d7649611104ba1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18aa6b4d5ffa3b3749f2e513ce4d5663873cf5a59c24327d217e1489ed72ff4574d72566;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h183356eb2343c51b0be8641c16b67ef62b10eb6cd9b80552ef44d0f405fceeb68741cbba7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ee3f6dea6a5466270dfb9026a2ad405ba0fef7c8e2226709329b3cc1de97c96325a7bb09;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12ce76aae40b82d2e151e570885d09cac1e64bba9ec73b62648fec784a4db52f22b73ca6f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17599208b3f38a9d19ef7b7b480098dd2e8e65e71a12d1105e4df92397f8d71545b25701;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16881b64acc40cf9bc15091a8fbbcbe2f7411edb8cc10034b8d2f1a0a1b31e068e363fc59;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h175a28cbcb58bb95b8e52ea47bbdd8e808413cea2cc892b2cf722a3743acbf7f9f5792d60;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h51d2483e389155f396c3de3a5ec3b76dfa903ae6182767e1257d0e18d0cd781424c94eea;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18193578b83c2f95ebaf98a67704a3564ac348dc5e0445991973e8f0c4b87d15784087e4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha702a0770767cfc0d35ee282b4f7becab5c39e5d7beb5d269ec5eed81964148a61d52155;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h58119ddbac525f3e96232af09be587d59e2761a72866b4fed6d0d22cce3fa322dca76fd1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b2e5af8264d9edc0bf5d5db210dfe6ebe1483dbaf7eff60900f7774d7f286ea1d2dff00e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9f000b942f8c05098999519c97922bf7daa08ff2be35993c612b4318a0d8a08c6539eaa4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17345cf41be405b93cf985b2faceaf0808a462d09f4387f264a567803beeb9f111f0e9e1d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h345e1b96e695eae5d6eb6386f13e15411147530d5ced3173dfff0b16920f504ff735d664;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h92bf4faf4d0bdfc40500e5b5b164783fe4bee1189685f36770778f4b7cf3e776d59aac19;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18b6c9db55f63641021c2c3f6391ece7a1001e01b5b0c3796661a97a34fca81b5bc04e257;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17aea13a9f9a3fa36a8499c9df03bb7a89c01663e59d2d10e78893df9df3e6ab34b3240ee;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb40d785d3ce8cfb4a3c54e9440581b29830c620d4440d1508f817a619211c2e269663456;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1867ff7612ff1165260392048ed428c982dd03f1ee8f9a2fa31d05ce8b0d742266477a5b6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15533491dad3bcac2f9d76de64529619f233b00bcce83cc14ca42c7ed0466426a95efb052;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8d9e230f83758d735fee8a6a577081a6360e83e6bc4c09ffb20e8594df6dea0d9a6784ae;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1577cb006d4e38149c73c85c8b4a4e771e47ff04136225065c927020d6c9ccd3832a537af;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hefbb122c72a11a598d4b083f740d6c8eeed2f9e2c4454ea7d74d26474cd9e3f93a060777;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h97187706d47865e56ce58b78afe8366e52bfc3935250930e2bf9cb379fa4c7dd48fbec30;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfd72cd0b5597ebef7e070f5dabd44a156dd1a1c4ba0deccfe4d54109f01de16b87130c03;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfa7071dc5666f07ab0b1881ada493878d8aa1deb119354bd42e5e952d8daa8b0d9076606;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h697fc41caf9d3506f05c9fc37a40f1053302a40e944e0f713248d9c2a186a1da482e81a3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b8a0ed39f20cc31760c924fd5879f4c0e6a0bb20e9dbb73b27fbc4451fb9381f5656fc3d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b26ec0a2583c44dcabd02eabd462c74d73ff148d6b833823e1aaa2a18acc0efdab2b6889;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15d671cf914fefc28839cee580c81bfd54540e99be3e197c2dd0e822fa3557d1abdb9b97;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'heece26afb3ada8db3f2d3ad826f1a2b83763ee781b176ee95d58a374a2a24b42356c00a5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha515044d2e9aa7ec5d947197747a89707ab85b071cc002a5cc256d1c89a818bfb26411e3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11cd3390327e872b91baf569373a35793e5f6cb40d31efd6027f052c1e29943dba42cc914;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hea5cb9f745a783a09c849c6582c9a49982905cd894caa04666e45472574c98f6691263d6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a51e259bf3655c1ae615a02131c74d20305d5d08f37e57d6020910ba4fbb186d6652c284;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3043681d8d01ac31e0fab0b9ecc14d5089dc15fd6cb5c9de28b349b197f3335d1b0fc7d1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hef1356dc6a780fcc96567ba3049e62ba9f1865eb3ed297d14f0b99331957e0c2417463b8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h180c38edece7a6abd87cf5a21da40426dc7ac6cf23ecddc134732fbe8b5830b56c0b88e0b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2d7fc91dc4a2c5974cb5e728fa246201717032b0d3099a0ed099eaa1eeac6e131b4546ba;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3371295fb2193770169ae8ec380e7f515e2b164f6095dc696468ddb51b136e805b50f24e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfa409914ecf04c36f1c0a329cca67562a704776c8d5df4e92cccef6c788440cb5b58c7f9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c3b251b83dc6d97364c65ac79f1216b81b003f649066453640b6a703de6d7966393ea198;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc423ea460e0c0556e00b6d2698a4e1021380c902651ccf0afa1a0376b45dde388d3cbacd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfc3854d14ba22aa168c9047ba39a5fb3db6ba13c1d956662e1d51dffca562f218b4dbed0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1526a131b0bc473fefe9a60d885405f4eee160c4a1fb036301479260fe0db18e3270588af;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14866df6a7c43bb09be77c87e1b207af0b1f9e7c7bdbe96e538cc750d1db8e39e785002eb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f236336ecd30701488308757a4efd53c3f29aa38291678218f39e0fb80e2b4ea37c6a78a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1283d0952db78138ef3099cc5fd3ce2140a5d6e2159d4c533695aa7a7770c73e1785d46c1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18777db5200906024b9ed61275063b8b92cad8b5b9f1cc3c7ab08c30ce75cdba05551054c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he92873e18f85bef1373c6ce779567405f7a659c368f65d73eafe89202ebb0a65ecc30c89;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1894ffbb47d7e603d4e2e9285f6518c783ecc74fe760e2b60188691605dd5a03609921dc3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eb930da11d9790bd08227a3008dfdb44a15855d368bbc8d6a5a1bee03922616c960ef5c5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f31e736760f9a8ee0041825a6ca3665faee615e5fbbe3eb152b792a44f8054878a945968;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd8ac3845fa11c6a88c98cec105ee4f3159a87164afeecd39bca82fc210ebd0fdb99343cb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16cfdb14a736318c780d2be6314f52a010f223260e074a28433900ed0669aa413ddb3190a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc7f56181ffab0677a8fa4f604652775383fe2d6d86e6d503fd34a5406fd21f5ef5bc00b4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h188a994d8ff99725d2016ba4efe7b72709c7f1d51a6ee902cdb17197c50fc9ea1cf8a4533;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b09985b72b2fe31c844b531967be2bf63cb2ae7fbb62ec455a9979b5a3355dff4d716e63;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h22083ea701d3ffe219a77b1b9753407cd80497bb9450d6e4286629c74de4990b07fb52d1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h133e50fa89ce47eb4b77a05248177d1d45d3b18acd01fc9adc9670b669ba99d3f0244be5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9672abea221d743249845640e9d431a10a1d4bbaab1311e7632cedaa5db8708f341b6953;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e86f638d60c01a7af201a7a75221c8f82fe2f2fb888603cd92a67053a4fb5c03591707d1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3e3966cc8d8196e0f2584311e9095cb2aeed99f283f73c0ecf91b344dab6b4305142fa9b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c3751e5d9acce2115a7c85d21a30049393f0ff12a78c71ff30afd5858b1475b9692a831d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d519bf4668130ed3e3c03b424f5056f8559312eaef56faae67d5fae292c0db1c9b7a322a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf8c876053f974e9fbbe86d20d21404acc7bd93d24c96192d623142acb5ee67cded258cc6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17905e87f12033c91bcdc1ed009cdd27beb8f1bb39f893750ac21af3d6c28c7d92661d1ce;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7e21ffca6174ee1d5ad0e3a06d630c174da28ad4b6a7096f57bbd2a776c8582715ab866d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1659f68c2b0505a88a105039c68674a2d4f14723d77102e6de9b5193515f0f4f8e16ac6e2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c5d69ee0a7268fa0fa8fc13b6cb1f7990c23e06ef8a1f22b329b3ee44a45c3f0e47fb1fb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h534c266c4af60d9328b24a5782f01682f34c03d587a156b7f3de1c2f05a7009afb4c3375;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1220dc9a37a9b5ebcb7f2bcedafc557d1f6ff3a0de0e1a7060938b1f71c8fad7ce560ee42;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2d8900f0d976b2fe8a03202a0131566c258620ca23cbe9321364a203fac0fb4a1a0775da;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ae0464335cf54c8e41a76a53b70e89c5a1f6f28a3d260b7f1cbb41756f9ac6ebc1eed03e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16205a8a843c82039add210dfcb082b9fbbc6004080174c3dc381a6f92ee0a0634db89a73;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb6cbd8940c256ccd2abd0f6c48536507d6618fd3eaf61544b9b1e1be61ba0cb0c2119ed4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1599a5aad19ebba7ea7c0242a257f9650921cd218a7fa802ed3eb2985885a8bd871bd81e2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15058746da317302fb1997cdaaebfb98ff1825a6f57b8090654b8d3d11021f549e3057c7a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf5f467dbba6567fa05906164e7aace1258b9daac5de1b22be4afc3df79feda6405a46730;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha220d1f228acb69a78c873f63269f763264bc6998fe86154dd5007a22c67fbc972493143;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a8d6aaff7390103d4f07d2273d5ab0fb630ef302210ce0f173db5497cc8b81a3fc8cc72c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15bf1464c9e80aa0bf4898e76dbce6e274b649d288e0c8d8119e51d4c8c413510ef0bb0a7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hba5dac241ffd4abe2ff13a4844d090ec3c674c5af1a0d5d201690f3552bc5fc9dfa17e21;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf3e5df55400b986b3ba7fe525db865bf1da6b260575efe8d803cc02d51a970c04f939775;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h134d908f6a569298d7e498f9994c2b986d01afb7e23244430986064b60af690e6fbdeb4f6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e68d2bffc6ca5327d18471f28e238a4043d52e7e8118ed3c34537231daa5ccf4471284d1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18ecabf08417d9fbab8f4d100bb16a6a9c58df87298ffde174beef11cd559295723325ba0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10f8e4228738f704eeea98f8b8aaf8a4cb4805d9349c43a5c232d37d9f1980f4ab7491574;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19a7627fc172516c878937669a9421f5df77b2a665fd4715edee2272e0dc9b02cac25f6bb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdb941a5a147787278384b736cb525c58887bf61a2f49982ab96311dffee954f2ac740da0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1327eb7254c7cfd49109246bf3ff44760fb4010ce8fe804a553bf35f5070c097c54522503;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2fb52f90ba614e5f6d31602396beff3b27148321d1807de76c0068f2cd78d43c8d60e263;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h44db47b2f97f1b3fd9f7d50b0bdee22024a5e5e4a8f9cf6a2b4f83e30959995e8461eec;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he035426115a0fbc474e149a60dcb1b355cde245b154f0674af4a99d29facb5855abbc591;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hde055b96592596889ff0998522d19bb06170422913288f1df3ae5578bf852c3eaec765f9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h199e38fc8cd54ec082132ffeb11a93ece42b3045138252f1901e0ffac0286f4b221f25d1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha614e47556e9be9a40a9ac62d03c2b369bb7b75fe972d90030409388fe67ab11cb89fdd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1df1607ff65298e8e05a12b8bcddca130b3396b524f41557fa4486ec28e13a47d761f4091;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7dea91a666c4eb4daf75c724908ec576935e18de6929a341b88a72cd468c5e4045b085b5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10ddbd458c79a47dc37c3931860a0ec6c637c46d0705062075ddb74068fff8286c30eca47;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h175c1563b184fba503751c7962741a3698202be2342997e9a7cf0189600a1ac8791d031e8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcb8a9ab8f5627526e315a51f4abbc2f7a54eda9b54b03655c5ad516adcf2f86b5e0caf04;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cbbe8bf4e4cd4593654f1461ba5857e0663dcd7412757edfe582230467d7eb9588818fe7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eac88002e6eafee6c03185a037016058d19832d4e45088a46e0930cef5575be33bb31129;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10fe071c078d720b119b2379849bae2da6145b9c8132b38a99fc5e761fc31e4c67ade0a8b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d9e6d7c672f0aa1bf435a44ebb43e4079855d191e35f091a9a1cdf8010baf9a3ae752b14;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19b0846abdc910a2e214113911cebf759a26b87cf9a8364c4e71dd59c2f75b601e3094b4a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9149c8995d4bcb44e5fcf40bb2552fd8d006b0a0501d010d06cb72bc55ff98ed70377eac;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb48cdaf6be965a5743a350bd1756b866d320b2e2bb3c295b7dcbcec429dd273752981ef7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f3b5e248af9eb31266e354d9edd65fe30b20c45601f14be85c7c471eed2e4dd5f12fcc4a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h140d64efb6e7da00a9153bd3900cd01f948394a44d6d01b52c8ba7fd2f5a9c7628132b28c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9525263d57b8b6d1482acd4497f6bbc16d5bfc544d0ab4f7b9e7658a6e7f92f95cad037d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d4b3858ed97aa18d05b877ab49fa911a5af0f7b8de688badc69784561a9a7136972dddee;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h154f651cf20ad4b193eb39a70aa5371f90b403e522711168dae08ca051df331e1b91dcb0f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8342e47d1f71480ccd3c88c0c089eaaf1195704a83fdcab7f904c1aca8dbb0aaa11f78b4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d4866694683e8efb4be83b5d6e5d1b62c175d49f4b6993189c20bb8c603afd640baa4203;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3b7f7d750698817eacb970093ab383e3d9688423fefecb15f48816d832a42e56a37fdf01;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15a23efb9f1c816990b0042c179b111e1d4f58a27e34663bf8896ac6fd511a0026f242e7f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h42f24a0e5d78cf1b0d67bd3176872035ba5cd0afc0562566b907426729dbdd3ed4adfde4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c8e625781e08d7d0e9299a4d9f8cf8e241a8ffdf8ab173a4a3e8a6a8effe9e1a7cb3fcaa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19da8b23e2676d274091c854f77753b314f7caf156f063777710e19ce1e9c53ec0459ea55;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d09104f0ced411703ced771860e63b21b1ccf7caa25d8a9d570c19308f4447f86d066089;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6dcfa201ce3bc067388a1a6c020baebe9100f5b0d61a5c966ce8e1636670a535b62712f7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h116a66b8c78ffabe1bee9ef0073c5f66913d746acb85040c3b7ff4d40d21c1adcb618893f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h37b769a0c868403c4ee71cb40ee3562d7e8f8626e22b7666d61671a8c1fec891e2a8bc0e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c7441b8a9605189793800d293a9ba89236177a95d2d35cde6a514cbf32c59acc4fd9e215;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fc8ea08567c29b6f3c044c83158428340464c92a8ee7431ed3437a63abb55822eff257eb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h342c41629e137d2e1089352cd18435f62c676cbf18391ee1eb97703dc704958e1c1b9784;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9a15ddd2fd45b455604e454a2bf5e6880119e98ce4b6a7e52d7efd16566b4db6c134b212;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h190497b8519dd3d8ec700230607f81e9e23a47a01cf8795653676f66a5686f6e7bb59f9e3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c945faf2ead055f144bece538171690437183eb220b136535f1e2bc8af92ae3f4d4702ff;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ad0ad0a1892b474cd23e6b15319a95c166efea33a14df58b7707802b9d9517e6aacc0154;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h64710320c273f39d2f5dc8e46c1611a7af6fcc7118251cb03d6c0ffc7155ae0018bcc92d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1521c04ff0fcf0958926dd79e9bcf3690112b33931f96078f1a8692e580a7acf3bcf8c4d9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13fdb34a83b1029b070646a05f8898e49d8b624c4b489adbf5b316d47c23b86c7bfd04892;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aab1d1bdbadeb451cb1c28d9a7719564922bae17c75542c8594a62fb1979183056116033;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14c7eb9f6d962f504a182d0c1ad848bc3397e84007411d1ee1437a444ff6daf4a5e105c96;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he0d1bfec0ac551ca6769be00982753ab6b26f634d20230660f3ec2d274a6bce1b4f820cb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a6e213a19add22283f07e94a9ce0de49fe4863fd1e8f5ef17c26535e2927457a532b3f56;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdf8b0d3c98f4e424607619cfc00af97db0e4a43b37101f2efdaeaa130ec134ce340d303;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h160831ba0aadbed11b66f53f7059a2827f37461d2f46e8f802eafaad319dbcbcd55ea4399;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1df4c0111cbf62b9cccdbfa1e584b2cc1826ebd96ea1dc69eaadefa5c77621447a8f9dffd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5158251f4138f1b0d54cddfc5a7c64d6d3ace0d934947f58b46bfb8a401d335ced21e2b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf0d76bf951e2b32da80686757734bbd0a5b472170b774e0ec7e7846124553b7f0ea0e5f9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4f3de70eaa4f50e6f4fe2f700d44e6b948e728bbccc72dc76f098c39a6114092b17ce117;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17774ed15fd22b2affa3c8533f4906fbef20ba532c8c241d60dd180e98d9b1ba3170b588a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bbbafd7ba9cfbb0fe4ecc07b49b7ff4f222ceed156108c5877e92a286de1183e9dc02cce;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14301f9389f248c172ee5c7ad89ada37650fc46602c2183a3ec548bac9e3588887bb3a791;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h551cc6b5ebb366c422ae1050352b96a0a0a1a0330f3459c80ed145c82249a5ef8ae30070;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc795f96756aae01bf8e4306b2f56a0d8982e7b4e252f7da559f1e6087a4beb712777b54;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h73ef6a87fd37524fe64fb9b843d764d2a6a047d4fe1a2ce57477bf5d79a35275723fc849;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6dd75913c54fb23e3ea5dbeeeb95adbb3c2466d58e90e1321e8bb889c3b793b890e96550;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ab2b8ad261728659190c4f205e347fd5bcca7a8728226b502a28a2d176a296ac133e0805;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h448afbd7292d9b31adf4107f098fd2de18f26ad8e15bb3d652809031a532289fca41d99c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10233698c567bd3949e20aa09c9b7dcfa7b7790c3685a5a5c3b4afd119be2e4f71bd16f29;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h676953666c6b3e3bcd7f30b864e74ec7546288f107da338e909778136613298c2be5fa86;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1734d62b2d4daf23de01e31c54de68276b398f4ea6874d3a0fa204118702fd029002aaf42;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'heb31a65e2eebd9565000e7e7b06102cf34811079a1ee2ddc7103e8c5a7d3ae161268d813;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eec15f3db7af08eddbf7a07da00c5eae08b0366533c1265ccabf2561627b6c57a6019376;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7a09c3de3f57fbe38d844676371b0593de82ae05f9dcaea8498d6a5305aebaca768629cb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb6e8e155837004313db23d3d07ed79f7fa640742264d365114ad986a2c4719ef4fc2846e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h78490c8eef0f208a0b63253e15bb4cd555326e63a41d487bc03a369f99fba20993d2f62b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1db9fd531f2c883b00bf5ed9eebf943abab1802142c5638178ae476e5d23796fe7459ed8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9ebe6316d28e9a4dd05ab378e32e483f3f770379a2cbff3bd14417800a210f51b4f51523;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d794f212e559e4389d14ba6abf95e4edcc5a8e8f62784843c6719f4bc0a2c2573d9965cc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12f870c79a92f6d107e0e8c45e26e7f3ed24706b6fecb5454fd45667917fb8c46aea4ec35;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb18cd5fdf0d18248b8fb184e5a1474757259079ace518f0999e7a29ff168b58f45dfae9a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc60a6ef7eee7b267d7674cf1e701f9f7a1e97b7e4f7a57e02e6481146bfa6f5ece48f18b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13d371fa102f483de63cdb486831b6095b94ba0a2b720f9615e90514ba90ed6471808af90;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h58f5394b2031b0b22e0a9115172792556f2ac7415002f071477adc9fb82607f0d184baa7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10a273506fb985102ea2cb751267a8e7f8b09e402925d9b484850fecc10e88daa1f963f8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbc7e88b6d7623b168dfe6eed3db1fa249743e7642d12217f69910c6669fd236ceb13439f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18e6e3e0125f51721e21072192f20122c6489e9ef9ba3b27eb9db40819a1f8fa33533d961;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19d1c05be25a09c2e660aabc74716950fe591c16ef8785d237a289e4e9b1b0d38bc81fd0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4222e9748d2bbcca727fe78970f54a6240de0f077786a5ca28228dd5f0c9e435d5fc0baa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16485c7c37644c7d9c7f44bd0b295cd2b2a9290586cca46bea43ea95c0597045ec4d6c8f0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13722721c7d74319fdae1da952e5a4068e32ee64e6e67b542b6937c0e14079829b6036886;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14e8f356d03b2a85bb08d3c3abd42b7731cc0ce2db5b99a858f6701e6da3dd6ed6820a165;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10aa7d4b94984030599f5a02cc1c027e50fd44cc0f8c7c809f2a524a45be9e13be7f28e66;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13fe51b4818429ccf2a70a5a62427a6664a1d9cab27f7b21601f14d6d04c3971721da0356;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14e6d4b9bd791cc5bf7e7e2963711ed62ab9906067ded4dc022dc964c7a7ebfd08405855a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h129afd666ca5e91f786ae6d7960841ec4250ef8e80d33fcf36103f263bca959e8614fe3b3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ce84bd471b6f1079182097342f9450241b7248d5b22980b6f85dcb2548066dc611e8ba7c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5f319e586f4ccbc2b595238cae6540d1197c8007b587a2032598610aa695f8a1cdf99124;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h59a1fb332406b3d2630fb4cbc043d2781fb678d6d017d3763e071312f888a19b4d74348d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h89ee91b79359d2cf11c1a21fb68ebd06b607d308f2b2ffc5c06726351b375685825d1e0f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ff13c1ecfc9cae037012d87cf4323ff2741a39f76b598fc49b13873b718ff87aff8beadb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19351b5b2507b9c7b7b04d88ac9da606c77e0be5fdf329a83dd84e281e885ad379e0dcce2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d7c5d90146308c1ffbad58a9808d67183e7f65584011bded990abc22301501ed0f5bdddf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h74110698fe417a5596fee3d62249443c99c4172677a96668e40ee7154054b31fd89dff7d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7cf243e507c5f8d6adf27387590cfafd51e1234a7efe0cfeb32ea4b59a5fd1b1ad6e2b87;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a8c905fad08fdc223564cab05826158bd9bacc9d0f14da09eac4ff08f17871b0c97a041b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hce090a1a3fe9ca5cbbfed8070bb49d4e38fd496742e4a5ff0947ec071c18c327a9efd58b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11d9d967a25c24d30f3569571c9396173ea55dcd06cd46742cc9b0eca93e282b99bd9e1eb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hebdf10c424d68661b84a25f75afeae428bba521b5f83656e9eb064140a1e3ac850a7e160;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hff11ca33324c54d78c367407937f40b6b6707602bd917779278da5bb49e5a8ad1be1097d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1413fc243e20eefff2ca5611c9f910aa9aaaa2aaca1f3e080268fae03fc2222d0f3434bcb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h112deb58f944cdcbad6fbb4496465d15e1d11523dc02cb58fd26cc5a9b673dacbabf624eb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha3f38f9faee770a7bb99456b3a123d19ad0c12ed134680c5af2619e0c44fe181edd0fbed;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb90785f9ff5852b6412e1a7e3368a70b22d02a9a4e5ee595fa7557a46962eb05fd01f629;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfd805f2b04ac1de0e36a8a74d7a2b88940351ce7f544dbffb7c2eec66242b86cca5e6ea1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f9d8f019820be11c6293a649de76f8afbdff6778ffef49cd3e2cc19412b4696d0bd67cc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13e7c9e337dba837eb1066c4a32c93f870377ef4e902a5a9b82831deecab0a1f15e50cea2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5eccd58258e4230306b5f69200813e7616108cd8344f9381377da88c8d1450a66d76794e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h177bf406d3642c1167ac1220538d2151a90bca8ce1e7f3f7117aec2b54fb0f2aadae4691c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdbdb0eea7e2fc0e88ce206f0b7e0db9a18f6b7c19c5d69f3030de215ddc1ce9fe32bc825;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h752a0a855fb6d228019d7fccf161b39b4b852dc531cc44bfd9965b51377c80507fd33251;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d353e3a1ec8013775d631a6043b4c848217a72042103d43dd4869ed846e70d0cbccf3f66;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h179ad0511a3bd60215167b1a6f6216b10c16ab528432d2d39b06cf907abce4a6e579ff17f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hac4034884f48ca09f3610d3456748642c235f4d1531acc19e2b6bf3e67a0469b2923ee95;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h179e7ad20242077602d503479604b6bbe3a86e2c97c55588267e3608756c74452984fe15a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h26132a6c0f025925a4dcff47a31f9a272758b51ae35ab558502f8424853e17a3e752b881;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1578604859c86af904ecb97256ae2d008fae5b3cdbc149ed13d2aa8d61e3bfc41750d2fce;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h71ccbc202ee4ca3eadda51f0e793f9871a5c707641ed255776a4f8d4a5efe6741212e9b1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c88809fe292f31ba4beff2101f3db10fe2fcde8ac5f41e484863e7edb6b2461bfa178a7f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1217ad2560f0d7118e598f92e9976a677fb8bae91a9e449447e28dce9ffc4c7c6195146c9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7a06b936c605180672896e4904f8ddfdb292ea61ae43039f4c3f78bd4e3f9cee4ca33129;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15a5a5d611183678ac102b8f00c96e0e7eba4e0a6d12564937de877aca9a534ec9e1ea098;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d8c1ee26898bb7a990b4c94163881479c6fd8b9bc2f76af4e2c0a2d0bff5dca4909cbcf0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1265cfb8914a72999763b2cf9b6275d18e31ad949b5536ddc6aebc0830fbff32d7852c4f1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e8d51aaebfee47d751e0d7ab7b69834804cfeed850c9a5cb1021940ca092318e1cd13e50;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc1672e8c0829d03e9891e9eff6c3b6f5beef4401f8158fc53e3cb908779ac9bbeee1db5b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12e3165169a3922558351d8edb904f1c064514464250af063d450dd0957ee37164c4bac3c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h172e522b46923d7e63f607d86c9eecb1ccaee870ed46a48307b31e0fdab41b69672f13bc0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he4a6bf03d2c487226bb9ccc39c638451adfb3d68ab8b95a462b234bcda44e406cb2eef0a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha14a362f2ed1b8741a23fa0cd1918319efe3be974a049aa7972ed86873cfdf86467daa3a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h176fb6ffdc891efbf1afb2744b79e1a4a12a87a81678f61aaa352322f10b160beb02887d2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2d37d212ccfdb5e399f8cc49353ab9df4da21b5f31fd137aa4fef12466562eddf8d1602b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6142708679b258c82d4f75a4fb93ede2001b204c7d68d4e0e6ae39ef9ad62036cf613a3e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha3089e3c001967b41ff063de5c2f39f3be982dc6b7bc44259dca810e112264f2e039e1df;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b5d9acf82cbd36156983b59710adae09931900af3623e3972a2b1bf3b061995694b4cef7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h615976240c7ffa0519d82cd0a82c21582ce2af587612b3b302aaf9a20903934b6da111dc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7b96d34c6bfc3cdd2d868b681fd1b551e13736d9a0fa8315fcc137a35fb41a1cb4d59e4d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h134a988e0df5e7a09f4097a442d0fd3644d78350e36d455aefbd942af2751263c714b0262;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16ece1fabc73f58233bea727b9cf6c3cf9831e36a9683dc0b54851b48b8522ba384e17975;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cb80a15919e72c55eb9c4bc5c61a27ac71bb596d672d5963b7afd561c9c8136e295cdeb2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6a86017c3a6f140c05e7ebbe369f6d7c6e7faa72893bb34a3922292e593979fff529c78b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9152f201fb0f8c5894512142069eccce64f9ba9aff7f460cc1cbc94cfdc14a5aa9db2bee;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb58b88500081b0bbeac86f6965a8ac7a4204da84e09fa23a22c54593b6d2a2d573039b96;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c5dca097718834a05d97050138c683c41d2e873ffb778c7d19e5efe8b2ccb46e02b74fe1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6ea2c4a2bf1c1b0b868bcb6e20dd037d721413c27f6767b17feacf182e820721531821fa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cc0aad59daceca38f687f74c33121312391d807327d2f7ac96a49b26523156d571b21be7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12d4d2ef901fc477c16227a651bcab4860f387459cb6d14e65f59b1685d29fc8f4ebdefb5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c035f1bc4ae3c10e30721b0992a3179a04a5d7725a537437dddef863b84eb2f258e77c88;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11e20e6fe24d9481745c1bcdeb767a3b7110baa242a33f144f03b06be3a6a07f3e187196;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a4d58837c3626da71c2df356a361cb7d08cf085dcb552e0169e3510559dafca9723f113a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h53614eba38a0e3fda2ecc34d3d108c2104d93e41f8cfb68743f4d032f22be715aac94f5d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ce969ed6e17a972b1bd715e28a8b352862e5048f2f526116ca36aae1aea6b08b665aa914;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h101742d508d42a52905895335d535110d4e8ae99b9faf2e35f3768318a73b470e95bb3dbb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e0750b74e9578c044ff3e709197512cc8f4156b97d7059aae17c64f218b736deacd7b94f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha0f14d2d7d6988cceaeb6a6a7b53a7ac36ceea19cc5c067991895b00a5c04ab3f27a1cdb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc8213ce2bad5b6f22f3a452c5ed0180f609943495f320c4e6cf377fadd2700897a1a0f2e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eae37942796b061dc594e2ae117f70af3ca59d8683979e393d7d20b0fa0caa43e52e18b1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16004f24eb04cd9a6a8998fc6e6eb4fa7c20f37f41236e476a154d3ad19ac2e823edd5877;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ac4bb36046bd56c2f5912745d7d048f74c8c7352fbb26093e284370b09a6c7c8596b2042;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f73674831cc2299d065f3464760a299539570ad63e28518b9b8c278379958ec57a159158;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1968b898e6d1a2cef642fdbc28997925b5bc1ac998f7203047a08bc47bc254b3821a3991c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7776293f9b22ccdc625de198117dd6cff5234967a2e05ad6e945628edfccf37397883619;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14cf8c521c37a7a0454adf14d5bc88770382d4cff6064bfd015c08ac30b5e1787165c203b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9c2ad170dad25269e50f36821ddcd97890a715a4bdbee9590b51fea9f4ab7d37f404c28c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h219293d2cc71a1d09d49d49b7e156f433de0e6f27e2effdec68849b21875e776fafcf71e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4f5dcd130cedc49e26cc70c99ddb06fd6e09c90c8af486155f2ec584fb359f1a629cbc7e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h147086fc89ebe0ee6d4c082e6a02cba728b193eed736d06a34d53a2535511885177709224;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc0d99147fdeaf9bfa84d68dc2720e337a4f29e4847a58ff17b521596963583a1bf4ca4d3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h158a4e9b1fa447cb4a24483bf5c925639b310cdde1d9cf4f3508cdd876f87e1a188d35ce5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h57ddd1539a717388793c83547ea496508dd636dd4dad7a0fa31096a286a47bf7960029b7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fd6114248e5f635f88b39b97110b494baf6ad75aac436a40c4a73b9d0b74ce101b43704f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1279b3e383d5930ed0d57dd1881174930c0a9eee9655af202ece795d86c2dd813a17b5fa9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d361a389b6d115228a96c5d10bf8a418ee0c09b08ceb7ab25fdb6a6eb67757ad3144c1ab;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2121d23c4de5b8506fbb4d459a913b97443d01fad57e135aa9b398eeffa27fc2dfb403ae;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h105687beff65031389acad78eb23bb2e901c0107ea6c41d9d7df8c8c3352f270e85ab8e89;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1583a68615bec1ef4700655c093afc9b01edfc0aba396fb3d171a2279becc2ff3defc605b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h141c393cba40f613d14b63bb7af1d18d5cd4e69f153b285600cf51f01065f423aad956faf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18485dec28fd5ae16028843b5ab1a32adc09ebe43b263b57299861b3f111141c2136c66cd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfd9b99b23aef10866c04a07577e3ee1de10fc661b16d6e3feb34bdf0dc174e367222510;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d87e2cc8321d554f3ae317e8ec18997cdb001776e5d847b1cd2dfee127ffeb81e14ab81b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf27cc24906d74d57cc622b04b8dc9a000f67384577b33c1cea4dc89002b43eb37b8db1cc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfadc37bc9ce8cddfd52cef3762323ffc64a7c794a4357185baaa03c20752505409fc18dd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7756ca2725ef7f32a28ccf927731143ad8f220c4387e0ebc2cd8e53b87e485697a119767;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1827ffa747535d500fac76b45b3edef831297c2e0c836041dd21a3c83cc7f44e3fe34265f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hde451a45ce72ce1be42f24e5a9150aee2920481310cb029cc801edf825182207481a2bdb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb3b185015e2a262fafca59065e648456f33b4d972b67b6c9ac58aefe3b07abf549baec97;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16a943754861089700550cedb71888684ceeb6b833fb1f64be45ecab159575d6af3aadbe8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e9c5fbfcd276210bf857b65b030a700fcbdbbd999feb22584eb20b3dd962db3d9a030aeb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6610074331c4ac932750c3306246bc3c7fb8d36922ae36c519bf7eb80a78fab348a7fcd9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5ba22ea133eba56f8262821231030bf8d4d02154255eb7a15548c91d6cfcb22bc4995cbb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19ab78c0ccd716f1296cdfa7f460ea22a988b39062447b27ade0034a50355e73dfd427610;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2dd423a8968b4e8daa60f790837862e45e15797d295c157a3026449a7b838ca884015d3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11e385583a81de5f7b05a4753565ddb8c385a8d9471990582f86f7605ae0e54f8ac1fe824;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15b18f38b36cdc3638a49a774a0ea675a55752ca996649fd94e8c068f7a7cf23ed16ed2bc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf8fa80685b6d5fd18cb96e385548588dfdee8147f4c0e8ddad9288cc22b93ca754cfb0d3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ce150d3f7f4838adf829bc55e75d02341f3daa4f0fa9f5cb16b118dc0c390f9ad707f7cb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19fab307f2f8f2ded3dc6b244b57c69f37478a4ce22ae56cfce7d54f5a8d23cd0ab2464be;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18e32737dec4d86ae407dc2ee2375a882c8c71fee241280a742a397b4e9f5421fd2983567;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he4f1edbb03a09667862783bab43aaef94499caeafa84406b06f39f22c40f1d0bd51172c3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hacc573294b795afb8e53e736f19d44a99dc1992c556673a23578a2e07a15f5ea37224030;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13b0e4ce989c33aed0aae0cd0fdf211c632c575005f5fdde9705f9a4001829513f3dff9e9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6c74c7f1e6d5e7d61b6e7e701e004aa8a0aab80d9b0ba997c2a9d13cf944675aa6420f0b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6af638836a6f2a6d317727f3496eda8715271dbef5e13fb4a739b5dc4d61976308500891;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9f73fb0dea1b6f917fc2de53b4cb14692debbad25c92e333477207a1b9e4a165633cef29;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b0c78d3431b01357f0f511b27ae99cd073313d2b951ebac7ec0f5dddfe73ece3cbd6042d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4e7836c5c2f7fcb2659e401d6ec1868dee3f51f3aa8d7294d734b18a108b93d6308fa380;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19f4dedc4ec58ff8f181f24dca5dfbdb53a896d06d82a963253616427b4ed332747d832b2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12bca7ae61a56ed9bc04c96f18892c26d619c940418ee19df311c3807666d97bdf3441323;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf0fbeda3dddd25e593f1ec38b9d1ae6a68bf571e14250d44dcf7e756cf5f768c99eaf8d6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b7850ff0bd57ea59d596d358d98696bda9361b38465572086d613a3d248ffcf7b4eea7cc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18ea96c353ababf634a29aff0de6dddd87d8a5bdef60994db146907067870501ed8843b9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1db9037337e36db3b167b2f72077a2ee4b8ebd41f962014834ffbf2654546a4942610726a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf4b83017e4cee276606b625352699fc70fba5f8dbbd7724ba69cd0ce6b3235a183ee63fd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8c8da6635c94490e6b80b8a3e371f2e32717730a83f97751177108e0ca9312b43cb3d0cb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h38607db5fbe70a83a60a5238f685a13a6ab0e63d7500cc49995fe4c3439a800d0a79f12c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c538ab09d5e59c80b48f99f7807696baf36195378dabe6f7de2ff279f4daa2ff4d3c9e1e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h537a7e319abc50fe7cb7f9389033207f93c19fe869930ef04cf774b16ac9be3f16c32696;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h869bb72c6eefb27a265e061fe8f1e7a8d2ad529ae62129731ae8983235802d49ad516e64;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha221e12c02f825a8e18f865dee218d0bdd4fe85462afd3e527ef8be304fba5163fe156e8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h192ecabeb6ae7a62ea363a9c8c920ceb5b460adeaaac07099556e6a8f9fdfebb09b6a8c86;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h90aac5aa1eaba36a244a51e56c16a74949945d2785407f1c25680e6597a0f3a92252a815;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2a093086998028dbd7a5b64621a3f9cbecba6dcef413a6dc223aaf3a8e1a59cb2dceff90;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9dfcd43dbc12bf1219260456d1545c80c934ab2d91ff8d2b95e03c24a9c3e189f07a072f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bff0418a5be88561dc835423779cc28869c5e4150a6d2e40aaad259b8ab4277766918d96;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf5efb40dfed461fd916d64d8efc36e0d7bcb34d405edab21035b56598e33052c279a4d30;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h143fbea4ef80e537d22a42d088829a255d18585bc45d85f94d13d24d8507e242b8b46ba00;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2666a52e911fc943095882112c1a291e3a4a3cbd8f71ecac4bac5c671436d34a7db89cbd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h613d0d2933a50c26b2e493625bf98b48c6c63b028ffc76aec1a27963a03fc060270a18e1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1605eb7ccb57ef3d8491a96019b368506b2ad71eed87b4b7c2a9d6b6225da61c1c53bb5fd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h182b5391709b108017ece90135586f900aa1cf867afdb9d43a1644e06aab95f3c749d9b34;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h33cbf48436c9fa6410432d39893c16090726f675f8f1807321c30a70a814bd3a641a81d3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hceb8add0e72c6d36230a0aac7faab6e6b9f5c4f12ca7e6a248ec36873acb7f2e7194f1a6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hab7e9ec6062caca37defe043c11fb32c700a25e761add0ae1733c8dcf56d3224990664d1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a892daa927d2bcb34fa63c2cb02ee60cfaa341c8df666ac4f8885744123737b318f08071;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11c52708e7751031223c0d7f111a78dcfa78795fb83dd5c0d6602f7fb5858b5c0dbcd9a62;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h327f9a168fe8f36a3051bd67dee5470e5931b82b4c0e95fac6f85ff003fbf69fb19d2129;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hed01132ab4bd5e09b60441a9f22db2debcc900856f1ae70cdad4a61b9cc1f96c2e1aec6c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4f49d90700b49567d957631571bde5eff3ade8ad3e1fdaefa0f05a6f3eb272d39815ded8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h186dd9b3734090bd795889b1408a0b31e7edd0ae9cc10c391f97bd97920d3ac6b5c77eaba;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19125dce065d3c28f1483df4d78e1c57de7297f6920b1d71f1c49f0a79148a1e5924b9686;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e513e1d44ca22728c648bcace194c4f138f05450e25cdff7415693fd73b96e9ae266c001;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1081e5665744f5e983fa472c62e0ef4b99c99ad3050615201bd8f60f7570df0a6be9b5691;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1769134dd9b51475aa7b865408fef64670d8c787171f9f48cbaaffa2acd76d167cbf6ac3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h193109a84b52af835fc0cf2f86ea8735f645fdeb72d12498be8d7e2dcaaad20562d3c0aa0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h176d9a1e4bc4a63581f4b92ed0d7792c7642a6b1cee6a1cdeec76232b0ee92d003cdd7418;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8304cdebc5ecfd868a244347956a73f59d665b1bdc25ff4b7f528275b8a96d05e8329a79;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cc20e843a4bad8c41c056d6fb6b06698119d739b9968314951f0d44a3264c9fea6d94472;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h136572197af89205d40e42d849c3045e67175dd095b55913d05e23507696c79e1d078b6cd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6749a883f51b4d30e62913dc352c0dc69f46cc199daba2cd7c29f7d53b337f14b135f2fa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cb1561d7acf72ef38968d10c86384f4b0b5cdd5203027e95cca664042e48c7e58b864e10;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12898fc87c7ebc1c52e9181ad6dff2142db28fb689892de42806e828ee9c1a3ce29d597e7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h61ba5e194bdd7b71e77a90827c8e82101aaeb829b11e3fd49ffcfff1e1c5adda80b4d771;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1894b3542c3faa9fac69fe51da76b40137efdd040f65f0132c3517c6273078fb82026f436;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fbd9c0c6af33056d37b459b24ec3e04b44557eccbf088895bf8396bd0c778337c6c1b479;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15e9254b808b70d5033d92b3b37db5b362b973b5c1528370c564c0f095185faa6e9181271;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf957d977a9e66a38bb6e54f996dce8ffe8a4f0f3595afc9f54015c327e591243386b0655;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f032918589ad0e5191582545521f2b3b6cba252326a7ae7a28277ededa6b620ab7263b82;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3aec74c062bc058f44f27d75b2b8be48b4a94691ed8cd75f5310a720a91dc173546b9d44;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14c6467b12665f8188c7d44d4c59ae0fa28e697c8255fd7c1fc77b4f563425baea9d43a83;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1216e0370164dea41684441b62e2ff5b4b4fb80a0d6947448e0c331b1f9d1aff59a1f107d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13aec5ec0ff948675db5210b2c5d68821d193a44aada98b5ee983041e59cc00c4efde5948;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h50487536eb3459f8348b6442f6ffdb0afdb6b184d28c9beed5388074ad20b219c4cf708d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6a2f8a831b8334805b38d57cc49551f58c8889d46a60b1aaf9fdd1c61ffa73c3da08ea8c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha78f32012300e5b04a86115fb649ce082df807a01f0c2dbce4ecebf32875d97a4a9c27fd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3f1ba80675febb32708db2f49f3378c9bd0906cc51707bd9f71b745bae4fb2f59676d447;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h55d8edf0ad832196d3ddf021f58ef9ec2003a2039dcdadf8d9212ff52059ae980b517ae3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19acd63511ae3793c1852384caceebfc8b23ca5ae531a992fb43bb445524d4dabf1207a7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h717b924935348440bec16a9d61be554665059827bfc91093f6cad043b10f805f445dafa9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1015eac8f4a898849a8bc00cc35f9898f39909477927957ff88846dc737ebe814877f29e3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c91135f2f2890bb565d076e6452862795333f78194eb84fe9852c76ebec61a51f5ee7d16;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1372ca8e19868232e0c7ca93f8bc13deee4b0dc4f722fe276268bb38136750116a731a2ec;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h183e829f2176b81ed786dea5ee8a01dacf06d5894e744faaa02456137cff7034df0e13f26;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13c298ce9d269c6351fbbe3a03dff5f72c3f34d50b79c350790614cf692cf4d4c562c8d76;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d0ebed722ba9976af2f7777a8de947f82dde578ae63bc00afb6aff0752d222f80a061c27;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he1c9eef98f20a7a4d2435075ed801e54146b58d3b3f29e0a52e45742b1137f29b683a67;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1080ec2f53e98da31adb80c09e3d39a693f5c3c7b7e76ba7a59431081deef4a7d08f048d6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h139b8a374c0eb5e29d3e742995d78f3e6d30c1e9e65d73d42a39b56d3c746669d1d16528d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17070b02e6e8851daa2560a655a9dd69db2dd1abe43f91d78238ddb3fe09515abd591afbe;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h73496cd80f253aecd49b57182ca174cc63f4ab5cfbddad60ced1a9dcc123197c89fc19bd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8c5fdd11684a0035173e0a2e15ca87ed45d8cb25a3a866d985d7f4e210e38e3fe49bede;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1997fb28612828059abb350da2003a50d1f679a4ad10baa8ea9aae229e4ea9607425ed3e6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h288cfa070b42d5948f7bee82298431d12ec8a169e6268bd425069bccceb4a82f6dc7a164;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f334efef2627024535a0de0de040faea8d4866d0b88a4886ae4552153f0571e0f8b9e6a9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1859fc6407d4d66bf5a125d1ee415cfbe24d42c06f8e8bbbca11b5387e7f0a66203a6d420;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he18efaec768806abff3fd84dac49f9440c8e744d949016821cb267cac82e0a4a2441fde;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8d936fba3b1209e33959dbd35892b62118504c777f46eb2e88d9b66689c9170dcdaae279;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9468d8cc865fbf5c73fd3d6dc2caa425927d5049c9825755480fb57b6699aff6d11885cf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7edced41d7ab4c76dcbf4c4aab081f8f6abea2ebdb62c010af7620d69c954f891ef13be3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h122ef43f2ae71ded3b57d611ae20f036de588bbc1911126c27e0e4b1ab1abd283c81485eb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d3615648328eb61d571b9ca0e28a8c28ab524e38f3ff2c7527eb19ec9de6868cad60d506;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd0e5c255cd86312b5f9ac9004a76dba82107c95b88d91c000406e5cd443e2f37737e6320;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5a8b8f677d4220c1573f276aa9728e7f4a2b793c4a9554891f1f188e7ae967fe3a77086;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h206372d5eefa39df905bf53d3e752b7599af4d614f0f2ea48f870268a00e04be0edb3c04;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf189b9d260f68cd2713e4ddaf701f07defd12f7ee8b90e35c4f656496ad04f23984239ec;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9cfc5ac1e2cba0d18f25fb0d374cad67d976f349d015611c661be843c945b980ef9fd22c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h91eb73ca4df9177eace395c7390a06033cdb451a465305a529fcb4371ce54e7d9b303a44;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16d57b811c69f249ec468b1d34d6cdec412f27b178bf44ef16d99baedf67f6503fa140bb6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15ec7b82eabbd8ef5713193e299e01e56d700030aec149a36cf6c0c86b08fb3903b68400;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf6c0a403afa632d8e8a78bddad2a90895ac9185426b1918c0b2e7e98c3439b282b9cbcd1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5edc3f56e9df38de5c410b46690a71dbc965466168ed58384206e8e244aacd01b437ae0c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15e03a4b64cbdb0cbd61930a304a7235a546afe445cd54269c0408f70aa50aadf979a5188;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e2ded0f11c1c953641e1ba9a6f50a19537106cccc21e64d27cb64d81259474d41659a2e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c068f44e7f0d9c6e670530a55ffc9d983329c31d7f48dc799fc6f23aafe1110e586a864e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h43c71631d28d21fed3ce205b99a1e382be54847a765f2cc584015a118d86e1ffff4204ea;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h111459164f45188ff66cdd7cfac0bc1e18ba6c097f2fe459b3891bb725cdfafd858d03cb8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h26128fa237842561bb268b8cc3f58de2acf5ccda4497e990c83e5d77fede1ec475dde6f3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6a0b83b6cb31e459f996e3435a9b64e8f3aec4a5f916db6cd4ecbbd7d9a42926095e7bb2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2a5ea7642715cb69c65e795076ff9144ff70c0082127e8d1470ec2bf5e38a138a6b146af;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11b38de9ac6d4f4d05611a97f204dcb83c858e30f7d5bccfefa539ce4461214aefd6292b0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h43eb8345199897353fe3abe8f82fca1bd7c54386fa520c461cf5aed6dc88fd6df27d9d25;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b2367ccc55a6abd8900c083edcf1c00cf7919aa0c71077aa3613ab20d510b72b43db4c62;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h101fb36b016b19e18c7eb09f3199fda6a1e6bc466aca63bf0e7f9ebc032b0d64e87e636f8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h422fc2e6a2e44b9f448ada6fd00b4801620bd163c36d5812d3ac07510832241c160da26e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h37f194cd31d52db09329c62ee0b7f7184abc767d4da3e30ccee19606d6885128b4e8da49;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h218d4edd5c7c5f97ec934b3d9944a3e79888ff4f0a3022bb75dd58f29e49e998491949d2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ecf7114de53ef9c7f44b6ff4ef4f88205e8f79308dde67be942d4da64fc4f12202a7f2ea;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15985ec3b97f1c621fd9c14a7f7bae38d2f5c203b299bcf7de81fad8d30c2bf35e239058c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9a901ca85ce9fb1cccb75b7c0f67dc56cfaf3264737232aa1d0a5319845c53152aba9d72;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10f315789f11328c6454f031b1d7151fe06bbe779ab2aa99ff0876505476267db147d7aa6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ced26249f238cc254f3267fc840ff5233446bd0402060c9b38d96cf31bbf839b46765765;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1215ed302fd6447afeb1e7045666beda450b3b24c9d62206caa23c31a7b0c68c893b611a8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17a13ea71b8a9469c4c10aaadc268e573106a748a309d205a1a2d147464a0b6afd49f9e43;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17a1b6b3f96c50e64fd8fded387bc5a6da12656a69154d9e909860262594bc5b574ef67f7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c1abcf5f3242a2c7d9d239689552226fa37ba9510068b444d1deaf36ce603f115ff3d415;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha5a7c7ebdd188c51a7de250a37e2129db3c767e2cbae30925dad898a761f2cf553187310;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'heffecfdd27235f5ae9743d859c070b6482e0dc7a1e65497dd63dff6d34c72c2accc202ef;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he665754fe748d7bd4826ca3a1e1ad828342f7e8e3dff58c5786fdbdbad9d2f7ba060dfa7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4f7b13e69c40b6529eeb01523d37e7fc219a50a319f1333ff2ce1647fb694ff612bbbc07;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h189e050dc2de9c9e2dae316088a74534e941725b7bd64934a89cb78bd8f769a791f4ef61c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h58d0f69ca4c454570b83696d256d85e17ef359a26aa6dac15dbb69dbcb28c9cda7ac03a5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13410d0bd8e6b95fca7421722c429cb84432e74c55bdcfef35786c4a88ec50aa1b2a04c2e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13b3545d5deac7c0cc13339ad9ea910e023812271e2b9654e044697040b024d1273b16873;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he18403531d58287f689028c37a54cafef11cb2a6984a3c1d82260aab5c60c1f4a322ec7a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f77fbd624cc1d483d42eb1d2fc99b0d11bede327bc0b819cbe3f73240191bcbbb13fc467;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc8755d52c7188bf029c0706448c7c5fffc379f10a7f522f0918f45e37068794186e22d78;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdd7b2874c907f592c001cd820f7bf1fdeffbb9e874548cada75b9e389c82611754dacc4e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12f505e47a5cbba7d2e6e61c7bcdd2dea08f74027094d5a15fa4d953674720f4a9e012683;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14188a3ddb60bb1ffa2f18e1b8092c489e14825b9fdb676883a2d1932504881a9f1703f15;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7bcf7dea2b6624b5fbeee4930e84081578003e6606d88def048b8d2d70beaa1d5883ad23;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c6090699c4c2adcd653d6c8ea0df742dedb6e9f6a3cead7c3f97e444b7d6e45a3dbb3537;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hec833e2f0b03ae75a384b90a816b2e668955fcc66d240afeed4d9442d8965119122507a1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf01677c46d49f97649751cd17365b661c31c54ec410abf48e2fe28b33a5a2c5ca8131edb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he95e9e7285824a79c9ed2ca23ea6573effab3cebd62ed6dc03a080f38a1d39ebc9274d15;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4408da5e57dcd8305d50c1691ca94c33fd28143100796f608bc8ce35d8c6ef097a79c1e7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f0a244a12f27beb91c1aed4624e8fe89a36ff2d72d6e35f520f1cb48acd40341baddf8a6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e31a73ef392cc54a85e9fa02710bda927cef6c584a32aab2074e1eeb9dcb508dc1f01e4e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h49f7e1633b017f0773596e2ec7ae743d57fc77ecf1c437c001a8f5382ff107cd9da300a6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h893ee81f8bd663fa7dd9a0b5270b9b297bb0b6219f62677fbedbd9b86e2d5ad92ec34f3f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hda11a8d50903f4ad783b9d1606388c01eadb6119e371b65c597c327272879cf4f06dfbf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17241f40b15e6d93f084dbabb4f0505b3491ca3910079c50a6e2b495720c05aadff377347;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17789f69b134af5bb9ad76e201f26a018ed47a29577f5876c235f2166cf6b1ba0ce13981c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h178259ec884b43e4d4f60b80093728778754642e6d146186b296c54586d210470f18c6d5e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1412f5ddce4f859af0adcd6f55940badca22b1461d1fe9ccc4359fdf7019cb58cbc8aaa8b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h67d7136914a47f7c854b2370fa5d772f77823bfd3a0b932ced4fdd885a6ee06af54325f8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9dba63c59c1951b15f6b1a47896cec7d7e3395598b4440f5b4185f446a3866171e25062b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h810bc227f1fadd1789d9203c0255069d5c61d10e111776acd5e2f84c41b1646a0ebd62ff;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb8b1caeab5d99208e3cd581ea7999040b8bdba865ca3d9821344327ac53c2d330fa3c18;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3f963640820027e3a9b311bf4fcc05ef9c981f4f5c703721e505b267602d44055e1c4cf4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h971aeb59e4906e862f57cfd7acb4ef033e985a4d1df311525c6321147ee94ffa3a140cd1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h183dc1a0ffe7b1fac85d3e0899217743c3172df3cbfc5b84b4ec3ab5ea03e4b3e4dc26e02;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hea55c21e67cbb5cf692eedf5e838e98856a00316ce628760e7a1bf458f6c07e8ac7e7bcc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd28bc40a7a25cedd7470e76880b818cdf7288b6c773a17f9da621b1648d0e2aded531cc0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8e97adffc0714f1123787674e255ecddadfcd099382d46b0287e7953a6c34752a5913406;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h852b0426e8d7a89247bc420ff79b6411add7d2fcb33610ae6ae963a7b1b6ad305f2afe6b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16e74e4eea2a3019024ade279b44149c6fac3178c35eeb0d69e2eed3507753a773e95b5d2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6cfade783a5eca522a799f584d60da5933d0f6a445fed8c479621eed6f5ed3a4717b980;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f7a29b240369bd62f2288e7475ae827a3dd583f1e42ceea5d0543fb4d838d4c9012d40b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19f13c9a5c08471764f97dad3926257733f352eadf7cb0a99ae40eff4e76c734b41400bac;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha9e48ade3ce3ff3ced06066b120ce44c69e3bac0c255a6f7c7db6bc29feba2b8cf962360;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h185cbe9e389c6a9c07808c5e2d15d8b23c180abf9d63ab74c922b450f844dfc319888ec2e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h109943aff84552af251cb19af5a023a4bc0bb5896ddecca537263e4496603c9ce6885d905;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5cfc542413cee9ce8798db092e99756eb68d7f84c5d931bbbdb7d0bc6bf39adb1fcb1fea;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d8ddb8891a713bc295a303030c1a5127524319b51d986ff708cbbfe1eebe17031c5aeb08;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h465318dd2622b18aa03d637ada5aa89cf71def64863c1fa5acca842ea06f14a1668cfe65;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h21bc97d5c01f1ea1a6153c050f2b5f5eaa4593356785583f4a8a905c0ef958343bcaa3b7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a47120e826c4ba1d79275c3d3af4e3e01417475bbd70539cf6f9393dc7da6af93c276ae9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10df989c39408c2bce03c8ed7bf3927b02fca0f7eacc2d7f70ef4176d1b22f391c602ff4f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb397cf9a7326a15afaa536a8afdfe5308dab86765736987f8e0d799a6db304fea2ba0d2a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cf008713a1c9b3fe5b72b13a04d6a776be75a6a3d5a1b14615a5b5b05119d789e020bccb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e72094f42aab5f2f03f62d251bcde5c87d64dc2b54b8339d93e091766197519036621d42;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h170e8433a7e32c049ba9c07eb2f522a24c4cfca217f5885f0032435370ed8a43e12d62f90;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1073d1651768ffd99f0b80dd5f534b9f9fb97cc45afb2a0f4696edb44c1d75836ad784f08;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf8dbf484203e003a9aa22018d7a5e1ca729130378dd03c60c68e2feda3204161e36eec97;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h96fb25468ecc33482bc382c8a936e3d08aded64cbc08f26e6cffdf8bc01cbddebf666557;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f1d396ab251245acd54548ca5297319393e3df06f6703a03b9e0f8b5ef8d763baf322d35;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13e10b6486408a45d101f5299de99d5fa8fced6229ed53030e3b223e7e7af1ed9942fa90;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e1195dfdfb9c110d357d9b9013145326e44ad39021069ef3172ec981664bca3fcdb7b732;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha3bca881f63468d1333cf342df8deba1c0962e3fadeaa8d4e2e7195989735d0e8a6522b1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha8ab1f130f4ae984670a25f8ba0db3017fa7c2fd46c15e512e2461028ca1579c780faea8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h601a62845064ccaa1b71a31e35bb18319c582b1ad658357d2332fe0b92a354e3c59ac62c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1283a56fe3a08e7e8f07099a7adfe995dc87f59b1499c8767a374179a2abf0d38ec958f14;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5572f0532c67615f1d1b7d98349ab332bc969997d473815924f466ffc9adc62f1b168652;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1baa208597f8a1fb50ab27fe4a2ab204562297df0bdf2b035809f96f2710cf2a96aa33dae;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h230df5d8ee64c8410279d9a4af16f85a9adaea381ebb0655c5cb8c6a207981e813adece;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10490e7cea044ef28ceb2e19e994c18c596e665cc5d555b55511a904741e1af06ad17fb51;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h174709cb58f036bbce018d05732e13b90d002bf1589d2536f2902367f544d648bddc9288f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h81d1dee0dc00b85b62e9ca6638552f661868c61f4595ec94498d14470a83046dc3837f44;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h64a383703fc82c146b5202d08970b16d2036291a7844c570959c3e03f833edbcac5a5be;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17aca4fa563e64063748287c0ce40c7fd0031446764d3da738d118e0078e2dcc71dd87cbb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fc9eb0327f21d0c8adc0a3678f1b4b805ec4bb4af4476a0e5daebef598c7c135702816e6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h93786ccc104b51b2d32200fc8ad84abaf73282eb31e17e90d23fb69609f631e76f27d00d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8d6701ba4bc826caeb2ae26087d93110cee31fdafecf4f57f07b9d32299e1b1d2ae3c872;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cd24e4cbd303d03d7ef02bb29039bc10188b0a564b13dde9d657e743a7accf6438fd691a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15d18726aadd6edce07608a3f2eae462e08d6fa6e4c40a9e0439ddb98c615b522f0bd8d71;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17c4a6edfb021fb977e6c12bb07b0e843f99a2011e614f11bcf1509875c0040ccb8e1a6e0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14bf7bcfa9149e696e2254c482dc9dab3d4b1cbfeb4323b83527ea095f33ef46b50ec806b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h124b805cbef87ff07335f9f331e0dde0f7f3babfbb3d15ba4728506f0d9571dbe8ac60a1d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'had0e5c80e589fc09ffd221a65a8e62c4c41d8e16a2c2a928687c507490347b3440aef713;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8025355138fb88c1c8e9241e4e7384450fbe1f0b88c1022ec86b30ffea2a8ab0b98ce771;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19047fceb3e772999df2c7f5b9afb127baa186f393650d62240232b89126e7f74979da760;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8d211aa28d073aeadee35be1d32744ab1166b4d15f6c0f7d2b9e4b26e8a1243a2e081218;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5b6336149976fe0ad8f5c3b86cde03eff49c1e3f4e37f60dd96cda7f2e2f845bebbdb0ca;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h26ae8430f7f904cf1c336ffe7578db5687653fc04ae74f999ad503267502135381832821;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1947876d6b881e272c35db3e9380721cceecd00ebdc68059daa502527319593c5bb29b552;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h130c0d1d7f9c75155aeaca3a5045301a5c347cd6f47905b6a9789daa6e7e6ef45b0f45e46;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfca1ddaa08cb91643d7cb2b82b0211ae10278e3a6d593d53cf218cf47acc2351604eb026;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'headf95846d853ad3cc2504221681108df5f339b3a1cc7fa3ec3929bb6d56f8468a565483;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11065a42a2fbacc04732a2bb8e1b0f48f53d1af1bdbeb38ac8f7799eb88e62d9a9a21a235;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h65d3d4a102f573974068b6cdf3429773da39221dca1cfe1e73db4fb1c75deace7012023b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he78f4599e7cc9c5984d62bde933c811c38d6ce0eb49adb9a377595de7a769f26c34c164a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h724e045c61b6213d1c991a3a44914323bf3673a74dced55fbb15d5d05c2a12d67acdd93e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19e73cb1c20df7cb8997b434663a73ca1d6e020936f5525616bcadcd1c1a718ce73b4598;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3006294a99690656afd4ee28b29f8443e95fcbfaf4386ee39800ae3a60a673e9688f6171;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha834d4d06e43f20e1a330daddfc3c88de4abf9a72365b6dffa8c40794f9d877d75b70c3b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a1b89e33d12770b1e4cd9e3c156c51c2ce7f7737a1f0eaa6eb6fb5b5c6f6562d823f14a3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fd550d05dc6b752c7823f2433cfb3fa1fd6f46a034b5bcef17a5ab6980fe6aece289c3b0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h161e31516e985157eff2201450c341f77447d60252f7cd7d990b95ad47d193b00df49a2d2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15169845f21922adf1b16f1528a0790dbf0683e645f95b222404699a9697f41644ea87c19;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dda3fc24a235a76311a479d4f56e6695dcb531ef7380b0f73f3f9b2ff6d5b039c1cee5ab;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he7ce253aa5a66db40b495ad0afbd2ddcfa671c10b9dbc49fab6950ddfe50e03e8cbda377;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7710b260be653bf019d09e06e3aba1d433955d65653aa414c709d1912a275afa8432da63;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he9a9edbbe19476c0a4c47c8933535f3df72367135177140f89b72a83b98379692a4176b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc06983a187e1ccd0bf08c3b9c2e57d232ae04ae409ee9f2c7444c93616da9692fa8022b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b309610bdc8447c572ea17d6e8f6db774f1e8a057df54894695897e5b9751897ca25837;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h125aaed7176ab492b604a3a890294361f9eb116bae816a15a9e097a54f880e1d9a099bb55;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4277ebb3a9dc871e294fcdf73eb6f5416377193722c0db67d2e911c64c87a0a1f22083f0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h134b383f5f2f8e3ad3276b22850eb524db3bb4f7912900e8bad938996d4b3f5941649f5e6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14bd9dbe2800231039456cab745187762f3ca878477d93252b9c22980ba353860fbd690b7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h44b14c9f1c95967fd1ab116fb0144f155bdf3bae897e3369689a34f8f6f4ed664893b697;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1515743f332ae0eb240673af14e766540e78f150b58a9adbb5738fda10660c5c316d0f391;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h169944924e1222cae3a7f721a3f06953d8e9b9eccefc759a56286412949879a9edc4b43f8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16d9f7e88cfd2f355eb8f3cc0648e1f8ffa4c8245f499d1fca954aa3d240e64982210f6e4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5dd7a1c6723af5fb9cb4dc456572d67ef078ab010f392dbcc097ad5143d85eff3acef5eb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h476022db56d223f7c74c9cd4b263c8b29d4b4a69a317111bcaa2a66a215f33b9c8349887;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h61356291bf88baa8be4cdda91a8293bc2800bf8ad22c9e53a083fabac9fb17f9fedf8a15;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bf1237a75177032b196d75d751ecbb799e7bd4cf8fc8a8a50e6acf2d725a996a3ebea226;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b2239fe7264e3f65f59cfe81b88ed9673c53a6a43722b0a000a2cb8e50263eb58b91ead7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'heba90a21eb856cc584659160c1b82e765c79f19d60b9c89ad9570be5d195e00df687b5e1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h592647f43ad25ae2368f7705b4aca348f46ed7975e2a7bc0ccf4a4905fd8b7b293e9edd8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd22ef2a1036f1b2393d4002923e0574c39fbbc162a13b7fd45a1a0641fb5cf311c6596d7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4bdb937882bd7310c811cd1f613cc545d54c750bf325ce8a61b92a3d4e91c2248df4fc77;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16357f2d700ae2cc208d12ef51ac36c79464adc20e96a849a0226bef347e51f39fc727914;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h104ef67b29ed30e3b12e9acd7a32adcfb4ad5937f1af21404ae5b738551e79f25a38640b2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19c1b912f32a44f2fb350094357667b337be8f6dc3025f6670c657c89b718e5a7a43568b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h791c428d660ea0ea28bea050632f099b14edffbadd0d2f13a98b685685aece59140f98d5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdd55fa6fb1ff61cb4793eaf8603cf298d303f1d69de5fb61a23607f46f70df3878620e8f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h391bb3e0673d8ad9b096bd6b10e04fd62ebd5aaaac15450045a9324dd9295951a1ae6da9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11e5202e50583595803d213b4e9dc9e5e1bac49d3ae20005bb4c7d7ccf0ba2a582da1037a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha7af2d06f74c219ef583ccddacb6ca3e678170978dbf195f883eceb5817e7b75a33e882b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h283ac1d18afdf8687c684a32e54a2b7ba56646cbaa54e517ba9f5c8cc8225246b9939427;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd1a7ce6be4fe856e3dd4f3f5cfe596a1c6b1be9cf2687c1a2d040ee76db0e520320c3eb6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hae2833e5a81887047eb301ce7537a540cf5f22c49fd546e493c0161a2832cf482e4347e1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he908d1a045c880345f163f00d62549a97edd775d767286821501d09208f7c81c2ed00e5f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13ad044a6195e93473124b1d8e48484c3b61ae2fcd046fc4cb9e6926c239a722141145e1b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13f99fe06508ea5eaf9c6f8dbaffadc38663fd9254b6266a0613810f06ca41ecb0f6b5db2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1afb21712956f8fa807f496ed094ec00da60628a1599fc0883028a40994fd725f0c90b321;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbf2c5b87a6950c58702eb57ed8110a60155f297d11c3927ea41846a024bcb670a7000bc9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h102d90a5eb5d32b6168e3ef1b34b4081dde222ec3e1417b4373ea60a36c9f576a7ed60d2b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h160fc561a3e40890fc992df417ba8c7e7222a7814f26500d0fe1c8cda1e3155f7a5bfbf6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f1d7ec7db9cb4351c914d0394eac9ff28b98269afb2af8a98368537066f30013e75cb3be;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e48dd7cdc21358e9028a8b30ebb82e591a0a51f09b0100b6e062fb448c8379cea200aff0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7d79f50b650a7b7cab8e0006e1dc84863987603d030dd5ef86d7ec12f739dbbc76597a91;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12e4bd8d45c7ae3283f0ed501275cd4b425e26d1a6f10485c031862b4f8dcc2146f8adedb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h104ab9e9ebbf0d54aba31330635ab8e2267aad1ce4704982de73cff862058a019f79ddb21;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbdfd3d34e529ea5abf2d1c7056e1820e08b3ec1b9feed2ed690bea26a181c9e12289d11f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h732b18c5c1e5abb1fa495ce1a5cca88949318b9fca4624a3d304a9a80a0f1e5169044b9b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h178ce9c4646df754191f11510405b184c6e8c76c5584b58b23b7077bf4cf280b08fac240;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h86028691fd0063890a87654df56e82d1b21b905429bb394c45b18f891fe96d4f8f01d19a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h174ef9e3f16b35a8862428c02b24747e8a8657918c98ecb44214c5e6b181ebe0bc0629714;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h71fd02542b9fd3c219590957159852f5a46a29da6b885074580c075b936a5c0fa5c5a566;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h136b446ce717c621aa2170bb91f1b0dcad66f8665516258fabd1d34dfaa24e3c2fdce6494;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10ef4ccd60703942b8c20ac7e3f294985e3bcb4811b5e9759cbde20ec800dc96edc99075f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7b071f559e9619ff73d650b216de71131c1c3faa96be976609586ddad03fb6d6174e4a80;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1615129c7c7222901cf39fcb29ec69f0bf5c39234fd4d3d5329f5b802d0f7e277fe21eba6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e90552feba41eba60212143534b1bf822b2222337b9984449779bba1a569db454bed3a08;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c17d5c47206c7edf6fb5c385b58a039e27c37e76932c2ac83789a869956309282909876a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cca21d41d1839a5ba4db37e99850e1be4602e49d707261340d7a0856b0a12d434a70fdcf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8c1a985898e1942cb31f9f0c364aaf79e3fe6e2df335836c8ff2953e3e626a6336d0643;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1089abf001397abac3e0bd67bfce29a43bf9c31901dd7ea759d518848bd6d08bf3599d46b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h365f5416730f16d4988a59c18df7e4e5637b665dfd71462f6ba2341c3950b7eacbff0958;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9e24e0b7bb8f7d509b989154ea919a95f5e35f32f3d5d2e7b2caffa3623ffd2934a1bf15;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h149caa42965c9c8e31adb4336851a641b5ba2e15261b425b87f312ae78d635cb48cef5ac7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h360b270bd458ac46988c604860ce839573d6af626dc0382ef477ccde068c8eac5fb653e5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1037b7790dce3eabdad72ef178854cf93d05bebbf4339fd6bf88ca297eede149400a9f519;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a8155c3a25b0c34d70afe03eb1847e9a5e00a82b90af12c47670308ec0360a440937833c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d6863060df387233597473819d3c1c923c81cba788feb5c5f649d8705714126e7aac188c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11920fecafb960f68b9bf359bbe6333e6e1b8dba174fca5859f2195f16879675ce75eabd1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12a3d68672ccafa7fc663c411bc938d9932dc92c5c12478556cd5e75e76f21e794b225d40;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he09076e183e8d7151e616646eb64c9770d6cdb9e972509b61b73e029636ee7d699679cd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h872626e52632ed456440b7c0d089c2049e3b3eb5a83b9ecb6a17749e83d2f61109f09e2d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h151dddaaebbf35e986f77129bf646d1e2840d4b5d2e007a44e96c860607cc123cde35f2f9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9ce1991d3e2643170234bdb4de322ff085e7ba4549624e42d9b778a5b33f850ec877e7a4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha97aa674d0d578c12b1bafb58be3127e92bd9f69cfc09b2051335ca1cd834d0178350ddb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h187366877beea23b60ff7e620ba00eb37481342e99c43260a907ecbb07a7fd77d39626fee;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f77492e10a25194e72fd912dd30ab2f9693b73c6df06c68cf575813f8e30b12c6647f684;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fddea48de4fd5217b0c2eab723fa193218ea01cba1e2cf17d3e51644f1b7b8affaa3a2d3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11cfd681a3ae11d22b57f3a27254f9f2fa033450962bea83376912d9b279974959f190f71;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11d5186058d0a5e17d278231793b9e724f65822da282eaff2a3b14646460024f1f717d2e6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6ba6213f9ded6c3c213a130caca56be2be495f5ad2de4186e195f8f2b02e473321a868a1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h95fef65945fe2227c669de25387766a49d0d0e11cb73899bab6f3fff2f4b9826b297ac1b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h301a5cf74915ec990e20edcd828663cff2920e95422b1684e801719160f022b2476bc59c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4548648e4abc326996b23206986cdde2ab5da3406f43ed8900b877ef88b63d5b836e0314;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13e8eab5ab51b7e8ef39e4cd8aa22c2d9b5bc1f54d4cd055480c1848b5df6d721a66b2555;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12ab1d01c16d0a45d690681576d6214fd644680c936ed2ee8083ccaf4043270f671812685;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6880f5751d4b5114ea6b921a6d16f074db729f62d4dc23e8f5b7134f3cba6f40ac51f4ea;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h168947ce02cce645b0e3b901e6049432bc170aad816b43af1b4c72a9a75a4e12bae401c33;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9e72cc59f89c0aa647b8dfffd092b0631c087093ea635db82dff2d25fab1301d26462793;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b7849ade397ce22518603678f72e930f1f0a9ad519bb0fb0c6796629ddd50e10ae2ca5bb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7428857d5089313606e54e630b2aab19c2d2f1cb6b035a5f8fc11e1263c367bd40c6f1c3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdb98073de75827177ff277bb25c99fd088613c7c7ea8263556a7a0547587dd5a44a95901;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2d9990f5c899c09b0454db6d71cffb217133d678785584795ddfd0ba463a00838116a3cc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2d814cf00a24b1c714bf6b87f25615e1640a9c9dbe28d9108d984a9afca42b6fefa8de89;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17e8b94ebc54a9edec3a6e604680001494a2f612f3860e2e8dc174364ed3c95cab2ac959e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h171b374d16ea580c966437eecf1f639d77825902a62094bc21baddb29ba18247ef9f00921;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14636761bbd22cb1985be47d757ba9d53f5e15aaa1796aad6ca605363d501e317612e9c7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h196b39f03481db7b7564ca464ec52a08161d37e9c28b9de36511d6d8a4e9cbf00beb1754b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc6c482416b3687bcb6c3c0f4df906d714f3d20ff1b266ae497ab1c32feb9452e91202ff5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2312c13b039df518d4b5f6b22cfeb663feca4490bdd3ee458adcaef453fac8fd69f28cef;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aad713342245bc0947c4047a6d95e86b8af377732c12a24387b50d469214fc575c8d4fb0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13c15ad22c61311eabd4c5be6467f302db7e76526d1be9b21b7d60cc36b9fd05537065acd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dfbe660392e92db4b18444c472a4483de36d9bc7544be5e323cb9af760d2a2dd4c9c8417;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfd8f6f80e9ea7239e54d0a9b613eab99d4f5867d41e8ee8df3492f25ed73a61e18c74f48;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f4089a240a4b437fc73f674698029613a2cfd874159f981cc95e32986e1ab6e765b4ba9e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc6fa47a024285e29c4d7d5888cf7313c0a6ad2248dbd10c8db754a42e8cb4a69a7cfdd1a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h740ffe9deed558612b14cbf112a2cc8469a0d263af4ac41723730b4494496353d2c1f239;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f76024942d87f2bc7c34939f86bd537aad2d08765f67a233f57a0bfdc9d694f1a2dcdde2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17118af7d80f5bb031f858601a23ecbb9f601157cfc56c0daf02c6db6c1599a534001c180;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h181a22bdc085e9e7977d498d50d52160e49f59f224a7eb7f25aa61b5b8600411612ece85f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f2d8e9f726ffd9a9f1f6f47e8b2309e660463dfc2bfc3a698f6030620800627122d9bd8a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ca20974946954ab6463823974c46c0770db45c6518b7a7bb7940b4b4c3b80814df14255c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10bf99ad1aadde2829f53b13c26f070d0c71a3ec3c3832b2118edd3450cad906676942a57;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12b826357994adc3a92dcae8e948509551a835f8a8719c2fc065284118a56ed5f08d988ed;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17d9e01b9d7a09b26bdf9d51879016b326136a10836fce8a07b2262b1f000701612896982;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ee12492aa3516ab81629a89b767632c7dd7d373d74cd302e4449a2c8320d6f126a93db73;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h159fa8d2b397518662b9c276c06cbf87ea6fa4425314a0a8f84885856212e27114424d18d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dbac076dd127b49b616a934ce5ddac07cf25ccf9e07921182280d648b6ecc149dcfb3365;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fc394d1bed362b698482c2cce07f0d3cfd023e6cde9373e78d2775e06b04a43a1c2d96dd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haacd975e3f9b30ee4bbf723a1a75de654a94c3d49873295f676b09f4705d7f49f817111e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf2ae7e2b9a6f66136ef1fb6003ebee9e7dd76c6728fc5199e5fffae7790ab99adca1970a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c98cbc8f6738aac07129c3f9e5bf4e219226d0d6b62c30f573c42c12b6bee9de74998d9e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ed60b57cc9f9c2a8bc616c83c0cf2efcdf9f3ded48f1c2a7b9099e328f8ec638586cb809;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h376a2b7d2dd085662a2f3025eeee181fe2f518acbcf2e20be8374e2c479902e610e0e3e2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h50e659526f9d886daafa8e33ff5a7ad8f8825c3218e21578cb99f79abc7f0c4778d1ecff;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h145ba0da61c244befe566998667cd107c23ce5280355abee1e91e0ebb73932393eeab105d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14617676aaaf32b8411d7b3d87f485c48e37038499de03bf3df4de92dd25dfc2976b52f38;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f4c26364a6698803d111232bf3ccc9e3f3e16700203f29cb17874e67e83a41b3841cc00c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16d2c47f2053395f58d87f60ea8b461a7eb66f99afa9e2855f8000df9582f93c6161940f9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h55688bc80f423ad8c6f4c192771be17c456ebbef9b970aeaecdf1739447b8935f2f3d1d9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4d82c00a26e9374c4076659931521dfd3a747b2ebc860f3ef63f28503940f4f5dfe89bb2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a88e8d7d465b1a825aa2203f7d253a653f349ca2b1ebfe4cc8336022ecb75f41b9d2aec2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10fb87ffa6050b9c91960bd06a8324abf96db55049a5a6b426d652a0ac0658d3fbd9460df;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ee50dfe75962de3777788af083b8bbb13e31ad97cbc49b0b7b85f9c9fb807286ff76d023;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha87c515270ea88bcc31bad6abeae99a826a2307c999d982ed7eaebc71d9b7e45375c20cb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e82ae40e88bf15aa702742ee4fb908fd76dee9f8ff367069a1ef0c75be1390ad3dcd694;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d202051cf05892c487d01b01d2e9b1b53f501a4ea085884f2b2970443957841199a91807;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hee222d6df93070a11a012d7a65fb6c8bee98715bbade0267cc3f840ac5060d6d910d771;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb4b4f22cf8d57d51cec75ded0eebaf9ea0ecb7e66f1e919f7162dd208bdf703063213906;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haf3f20a631020365e1d8b03f198356656bb6dc7d0d363b78998be2d36e7b53b82ab4fd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c83174b1b943052c3e26e6f180e6d4b3eccf32e1260caec4ef58daeabe3ca5caba3c700c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13d2b59c599f4a3a231720e2e99ce5a563e4021e7cf7bb44385ce0008d5138a8e6a60f092;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f2a6025a855c4688669886ac68bf00504c879e30dca1b17ae7105cc06e4b6bc8360986ab;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h57dd017ee338515627c234a823d2c54ddec557596955a776dadcc67777ee3ecff780bb6b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1188213915e14c7eca30498384b35f59ab62e4175cbfad9a6ea3b1746d24811964d5baf2b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h47220022ea4056a659e272b8cb0ec76f490b601e751276aa9ded75f0fa34300ed0785064;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17e7ef7add3e332ff5d11a884519232a842614c7e8011c804dc873ed1a09372678f30c4eb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b74dff3911bf28e1420062020d6b88a229ffb7943c6d5ad8872bd7108b97a0b400fbf0fb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1800f1fc3ecf89051d8d55cf9957334950aecb6774d874cf4eb047807411af437ace22ba2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bf4d55e49e0a5b078138c58711a2cba3b35aa46f7ea34aa945416cee28b66c1d91d5a07;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b6e7ee0d200e04e873c51215a1be01fb18e547449a799abb0f555b5d4f4e77a49deb067a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c190dee3bb29079e471c327b3fed7b51b4adb5ed015ce0f7770d38573098a4b1da1218f6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h114a499a82052909c9dd912511e0a6464875c0a65de5d570dafbe6b301bf085da5d7c8199;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4213447bf1536fab8dc2a118032fa86a7014936d68a77ccf53ec2385859b92eb483ed259;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc7cfdf0ee493e2c10d3aefb98a61954eba7045464869eda3a5bb939674c9a2015a13969f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h128af6757d74539dffb51db9908c79f1dd43d6304b27844a7fe23e611d8786f2f8de36bad;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf6f51e4952565531615c503ca71ba8b9959fff3c22d85c585df61a47dd1d7022309ca74c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2942f6bf2374f8b54ca9d3de75bce3572d6a795a2fc7e771f5fa5284d98190bf16639037;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18052a0d53dc8028245da69e28d24887ef31c45bab6652c2d000adfa259baac743d21cd20;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h126e4844382cd4109f040bdf6fa6646e8861f4fbed5ff96626b3c9d1dc61ca93411daf45b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14cdea2b5f279df0cca717587a80affab487ddbfe9b1b870a273e55776af1ca57ab7858e5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d2ae187aac963fdb1c16282066ec36eb654a9838952e6acb905d8f21b2c00a917cb3658d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15fd5a814549fd11964b751009ba335c5dbf6d966a182e291a7de59d5f95744755678fada;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13bef7e5254ed62ee628d0f02634072e80f3f20d78c648ab04b2fdf94ac4f6c410cdb7f99;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc71d8e784afd10a0a4f2b7f9c2763273a770979bbcb047cdda67039f48cf3bf958a7266c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e9ab276fead093080e006de328045f2423231ac7b0148eeb85d6c640892504394e5f5bf7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb5f61f5d27a87c548d093a43afb20b9e689537ed4258c0cc23a75e5b3fbe1928940b2827;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb522a9723a37e142c48a51188ed35b642909c82916b098433913b73be1ed10bf59de3fe;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h138117254fbe4a8603079f250b1d1780c0a1e3c605b93b996773e16869fb861cb667f39cf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h436475d14650c952c7bed5ec42d005ae45f58cffb2d7d86f2664320b76eb539a93d1abd7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4cbd449af4caa3d6095158dc7246f8736f71bd777ff5c00d657a6308e732f9ebf9d955d5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9caf687754e11a47b9694df7389e5f71f38172402f2f68557bfa835c847fcd3f98bcd476;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h182aafa1a8f3eaaa7fb827b98a3bd9b55363a4ba7a532330a8899ffdf03491dfdfcab064;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b34cec32dd5dd528146a6a14eb569c3ecccfa8949a310bca2685598042789d213480cf15;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha3bd2d94859795027a5d5e7c88e161a0e2c34286dab3fc18a7c1e384c92608af5dd62fc0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a7ac891c578dc09af5c10dfe4c0464f2957955a32501615099972277fa2e15660d068ea7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h167825a9b2f3612e4cc3f504a355321c434f54d44bd214d5b8066cdb9da1df23dfa876dd1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h31479564585a849bf79d47ebb4762e36de8339919dbb9d1bc8f30b147132ff235d2645db;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'had7fe524f2fe5f77ee50a3ca3e8ca49e7c8850bb630f18282a5106b3f252542334fcd6b8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d1f37d7ce2568b2abe7683d674540612e32aeab787bb76a99769cf8e3e9ad15e4600ea87;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17c839dc4cba7d59927a16bda7a0389948e37942dc26b713e542f2eb484de81a6891a0297;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha9d44c2fa742192bcb0e3ba24ad4dfaa83d96847a806c565ce454467c7dd5a1dcd69fd6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc77ab961e0c11b3d4ed79b539800269c6c035f5165861cdb97eef896591008bc7f3639d7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11c8386b2dd4559a4c75b6d119599b8968ddb665180d80b2ff75c7d15a50311fe0aa8cdeb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bcb4e2e73cb60fe887e5641d5adb116afd6271640b97d3faf740b1952b8ae67630a9be32;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h153d008e399660685129d3bf8986ce9ca5e451e8449523bb5d39199db5bc45fba076d2715;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c7cd6c9839a359de88824209d937c0d9f0df346e8b46a8d1ef7dbabc0c9e23f351845a30;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h122dcfbda14f0c5646aa607fedd5baebaf93fd3cb1e806d6730aa1eb794220bf2019a0636;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12f7789207aeda2f8a1b9155e504fddd46ac3da018095a2699b06bba305d9f90ae0c6394c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h196d3e76b80bd933e8327763543b01a42f9ab0e8f1a9b7e8bc78bbdd4ca56f73fbe445275;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16f7e82f79e83013d3b59c3a24c6fa0a54553e70db71e04b39fb102b1abe3f54799f227d4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7c75a9d3d729172021c4e89110a68e5d8250aad6376f9e3ee4c50a8aeec68d6f77e8fb4b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h78f2af18e5d123ab6df0806e677fceebdddb42662a19f09351b138afbd6d11dc5d3909db;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b82eca4c40c42d838ab76d62d3a6f1b425c0a312f6751a701c32c7cb9daf4d3ba263eb1d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19b1eed2b1b26c13c2abcdbbfcad65271c278423e60e52b5dbdce851bea299b9ba01a78aa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he4c02f217046c6a4b9676ec6fe4b836850c12e6eb0ee5051f904b3425e3658eaea9365b9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1246a0cf0da963ed9710090f2a3179c109fb81e342d148769de9dd9f9426c6dfd01a8be3a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aff71c9fc9944a74b01b34966f4c1d9da8aa1a65ee3caad1c2e3ac249bb306786a156b12;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10b66264aa8d19f189277fc6976ac747962e659136438ec6b47d72ea86d7be7347bbf5974;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h239db8b22abeb6d9d736e95442e3d841cfd4d5f1255e783e5f2348811c10dfec3cc7911f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbee618720568b38a96c60df9c3fb81838a96b8e3215c72725aea60a2032f9ff2af654cf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h182f53bd897bf10b27572fa19656da1e8cd9ad1c0448d57a87a09ea48f3b9e3d6bd6f47ed;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf23eab3a91ffa7367e4b77fdac625816f205969ce9bf83658535567c8a95c8b979ffbd87;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1901f7d477c0e673e57ca4a420a11b320b4986b7a46c1a8ef4bf6fce012911534e79dc84e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he8e6e48fbab54d9c713d05533d9dd36241232c61ac92c1e840c09a5d260802ebf56dd229;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10d14f83ac59294e5f777f5e411379b3e910ea76d8f6cec9e27615a0dfd879d5c2fcba240;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbab0be96f77b5fa4864c36465c756f59d5b491db39d3ca042037c74368a2b5a08a01ae5d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d40668f3b442e07f66aa64326870d936b263d169bde09ef9f6247b6f2cbc70c5df84f733;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1faf4e22135a2eefb8be4db987d29026e1f3eb200a9f5cb774d312270ae5a21e7a9784a0e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6e06cb2dcce6170b71241075a8d8dff5de7b15a1155c5374ea418b15c2d89eeef5e9bf54;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb0dd29a12cf45afcc4018ba6aa7cc9d840c94b5d2f2227c9099a767195d2ab6f582e2ea9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h408fd693af00e78b0ccefb85c470d4153acb2a171d8adfd800c7d6f017a2d92cbf87f0b0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc72573eb7494bcc52a5b101eed9e425c9c041e9bedfcc301a11d391d361027bd2edc0b2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14b90f17e010c3a00e7ecac1eaa4b65a191f75c932a4cdedd5485f94ffc3ef0a2d09b6cd6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15ae46c32001dbcbd86e357e41773fe64b7730090f84f6e5320d3e4ca9b28b227c9533df3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2b4417f582790e2be22dfd6915b1d9c5d8b9a7f1b63be460b07a78993497d7d1665585b1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d1267aa9b544fb41f5aac2ee4c0e2991a3617243f7b9528e0c458c050ec9ce825cfb50ed;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d5f0a62f04c2537eb31e58742dbc04a02622e5173ad0e16009abb0acd099c5fedf83e40;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dcd80b041e6f1a66e809e252a23d4c0bab578b43a6778cf37c04547f15cba1dbe660c176;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14eeb758a3c246b581f7b312de9c8ecdefc510b00ba94119379c2008726657f8e0f64a97;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f8644fd67d1fca4b4df6254f235cd1379ff8667ecd4df484946091d08848fabbcde318e2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16a9ae0087599566d30f840e6bf46bccc9cda6ffc5a57bb670314943932a7f02343f86953;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9b92cf86da034c512c314dc3748036a8bfd182e99eba4326d0e70b120ffb8a73a9bc41a7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cff8c9883b6a2dabb15655250ec59cfc42f4eeaed7f55fe8d4394005d4bb87e4c91638ca;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1228353d992193b3b054eb22808c71c50e2b943278cd71cd24e7676b3987175232fc1f7e9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha3b7ec43cbfd0f2a580f25dec2b4dcfe5e2c81b6e0618ed8d17e3c6e34e1e96ee48b9d96;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5f38e3d257cbc2e3cedf5a040060ef8c5fe30646afa5a9248a16d06563c463232ae7cde5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cdd412bb5631237a2c5211b9116651184c27c53a5bb4bd2177989418fdce7f6a2467c39d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb3eb9b146cb0f7f5da5c948d4f9b43d426afd5eea03445328deab403fd8464ccc1bb2bdb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18c0de5113cb42826357f88b87a4922f429d1796633767edcfcbcc5a0ef429ed2b29b1fc6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f8baddda77e8fa896dfc510d285a811b15473a3b6fcf22e09407cdf6dd29ef6fc2c5f0be;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbf31a72352a06e30d4575239be4b43a4e9a2b1ade64320010b088b2b553bfe81083b35ef;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8a7fb91c2f8c58ce69ed4a405e8b6d65dc1cb05db9872bad1b22637e9ace68069d598a4c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12ce906596f4b6ea44feb6aa479e1592a924fd09a7e06d1c256ca6e105b47b0f6e473dfca;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h104225a07c85b6d5af96ae476912d2c1e2fb82d599a494f0e3a82d2660b0aafd2186a18;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5934bd06fa7c745995e5a78f2564d25b3c884422a6c056ffbd54709e47d93e3cc2f3aeaa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13807b4e8ab472b0779a0b10a767ab8de96b26de511b98bd41e2794780133bb869dd9afcb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3a713366a57db4a8fe1197d286e928120988601c6f6e1f9c6e20d6fed9687580bf018e7d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c2b7a72d4c9c477815e3ddf5ad4855b6c129dc20908a34c8821e6c77b1fa8ec1088e0431;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc78a16af362d715b04181fc94654fcd1ea6fc1905317be1d54b7926f1d769bbaf1e82285;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h152760936edaf221a5cd20b7632ab676470c32f1bbd1c0a815eac42d15852bd61aae7d87a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16d82aae88a04798de8861fc2dbae7486f020f01426ba5a53f81d3a9518c7099c09255a5b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he1baa4eebc63f49fd3553488ba8535be2f9b2b8457183e65d9c4d57b1a2a98157c05108d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h150bc1f8bbab96489d0db8338e5202b0952e3425d18a9f3b3a8b02c4fe0bbd664bde4c322;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf45591c8bb9a5192f7351cbe3501add1279af9e1b2e7728380d6d1eebf8ed7d79789e0d1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ef236ef1fd28cdfce097862460b93e6d80e07e8268bba5621233490ec0112d421024b222;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h60f5fd46bde3903631fd6843c94558c5f4c7c5392acb1212b4a3b1eca1c24a79e1dedb18;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c6b787bf99e312a942ff6acc6c3f2c06aab9df4142552edad6c2c21ae70e5f648b3ea748;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a0ebeb6802ab57ccb2545151fd8b883e8cc40639940d5007b17b3111cd69fff5441e9f4f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1301e42de0edf438d34db10dd8980eee855be2b946f81b8edef1cd20d3af1ca9d41aa2f2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f33cf5df9f0daf519b233cd017b2371ae467984275ee64e34876252a3636acdb7ababae6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h113472388bf259a34828786cef471dedb49aa3aab54ab534f5d2361b21b0ce414faa80cbb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h66328ec7493a34687e13cd67112f369000d24e5f6cfcbd3a83fbf99ee642107b95e05f29;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e8d2c981ed9b05d4294014c223c59a185c4f7633615ae69eed2a767db2618d8a570c5386;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf308851d5fd87ebf1c4a6191cf14a8e4defcf91418d03294e138a6d2d8a9da82466ca040;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1de3571c5d07d829f57cd9bfeeb0ea968bf888dceffb052d6ea0f6d8cfeccc37e226a00b3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfd120d50a85b321c539c21e69b04cd9313360052844079fcd86a98f938ffdd709b0b346b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1786be486d94ca0c58fdf2ace7e10366a7ec85826bd806e3713a41b8ee5a481e8c8dbccd5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e287ad316dbcddcdb2d189ccc82a41f1ea52aa46ef3f7c3056611296fcb67d86d20c0a66;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h261fd13bb8d89d535c2adcd3c8e258c7bf35c9d4658f0eb0e2e6df09867a19c062e43032;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8e0a17b3655e0ad36c4875c9086aadf73b2189896ea2370a79d246ec5921d3eaeb6c7aa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13ab3560d6521ac4fa1e2360ed885c8476995bd95a958124462df1ed6df4fb15f484a01ab;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2fb211e33d9777cbd3b677f0bd5788148d7f6c71667b791aaf9e27211b5605d32398c373;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e039ec7aa42be905990a24ed024b99f198421618e897881ac55cfb4fc40ba73354c0a1b9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1175c2e934fc927d1e7d1b7cc3e86862a029eb216cdc1f0e4de24451a034e128c9cac8263;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a8230a0c484acf3d26e2128f80f8170f5fc054fc89217337302e296f0eee0c6b195259e9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h124e49c0902d1f384197dd4de292685a180136f70b7528f2590d749ca6b8bbd04d5cee1b7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1da6c0f494b036fc1dec6ad90cbbd7ba721e4c9a1933c6ace919899fdc78ac0d3561283dc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5adf4f24a4e5c7cd706a570f9fa33b869c9d7f6ea71023c9aa51f9f965cb385af6bdfed5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc5a82fe2cdc63a3521721a8eb2ed6bb49710573a39f56256bae5152773a2a1be090ddd79;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d506df187155507597c3d78e1c19af9e7d17e9969af28b4d8375b6069b0e2f492fe24ff;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ca8a15637a1740917b5b64523714e15ade69761edcd48bc807d323daac3ab62c6d53b1ed;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15e6ba0d373c4d1bc498d3198b6cf35c0bce5b550a8d67d0c14f9a99ec0139ef2645bc70b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf0906773893e787f194a425f7d79f727af1dcf56c8fc7e2c536b1db7db30ea3b14ce26ed;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15750b8d99a8855258e60523058ed94ecb006791f94da94b3e976fc341b781cc2360f93ee;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hffad2390bc1e47ffd40064052d92cfb37ec88dc603b8cd320359b810ea270564fd06d6df;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he7d26a6e0cea612eb77b694bbeeb1ce7d5f643dec47b53f4a6ee0245ad7995281f0429e3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4c304558110974ebeb5fa4be3e8102cdfd6b282b4e676aa84d75447d0b7724497e98d1f6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbc0b7b4d612803b87a2d67782541a5490d49f4c498119fd6089c78fe2da78ee63506e727;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haf7db7e87fbeed402391d5b84990880f2d0532d9c095b4765fabcdcc0f49e1fdee5d829e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dd112856e16e2de140bdca7fe77d51af4a81d4d3617ee3cf07db0b43e963c8f839fa49c3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2ab1187cfe89b6d9f4f8c50000be3725d6ffd33e02b38b43c42629ffea11d03f7b47682e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h24e75732e6ac3acbfacc75bead3514c3c6846854931135affdc321d79555ba4585f5f3f6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hffa8cf28e3d248499f7b184ca63a777be22c5b920a2f3a6a3a6957621a6e2b1d52f320ac;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3bf900d5c5b9fd3be6f08a09c09ea6a2866bad8398db68aad2b8677968b812318c07cd7f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h180986b7ba9dd137ed8d62a1f7f3e61346dd40ab68ba0a53e5e8a2f440411543451f95323;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2552e856812106985866241a456133cc15bd0fc03641b93e7dc3f8b9e68ba778b5123993;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13068fd7f4f74efe0ffebb4a8e359b0ce1be3096536fc796acfcdd2b3044ee1837da8d6f2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfdaa860be82b1e10973ab2f039f34ae4c61b5a34a82a50c6df361eb1f6279744550d1afc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h87eff75df1aae7080cc9ab26a07d97577ed529b294ae33874192f8d19f57e8614d8a1224;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18df5569a874d5319f29039b59fdfa0e956dd80134cdb8bf6dd5a106886276847619f4fef;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hed00a7ab71c4be4f3da8d19da0e24fb18fbcde8bd7a3b7696a4524908829f8c181207757;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2aa126d9904183eb485bde6b875322da8d86c5788df03bd7ed5d10ecb5a638a284749282;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf557ea3bd10e33a3a40f9f094868e4ba74adffc575d4746680790b9d52f348708486fe87;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfe549f7182f4ddc56402d3e9e74d6b2692b004a12ee227180b997b4aa395589ee2e8355a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h29fc2bf85f011415a4da6bc098f296eed91f972e277a6ade315260009d45ad75c6da400c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12120a72bd843c3789af616eaf3cf5dad5969be32dbfc17474c495d3042b3f6ee9e6e2e3d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h108e32bcae6f1c32eba0e1712a2eb6298c6e9e8cfcf93c0a2d58defa171fe207d45c1ea4f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1418be41813d382c8e14e14d0f2d5aa62afe19215c9da285a663c96b0d2df15ac935f082f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1442a45f17f0dbe437788250fe856c40cedf246ec6653d5efcd8995946698ff4f07861ef7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1103da96f5cf6c1512343ed7a0691c823388db6531abab450b9d0d3d2dff5b4580f0b1107;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5d46ee744de0463ff1305d45e3171918361f6d02c2f72492d5095129f93471d44e02997d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16ce8a3ea4c1d328d758a174886ac3addf0886683ce21f53dfb5874a32358ac436de1eb6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc7427aa6a6cb971599584c7363fa15726595b1b915ef9c62f56666d67549176f5ef9c72f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hff9ae633a2f084f3f4167fe82e7d84b71f101ee0b226deb05dfb24c0be1c6a7d7023cb49;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1955a19dea687f4e8d496c15a7d86f792cd7e898f9c736253b5227496288162bbd3ce38d0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc00e495004b58a44ec86afac5b870795ec5493b12e7a7dcf4a6fb05dd2fcc0c800bac4d5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ce87e6e08972c0e18dfae6f88b1de484353b657591e5d6b0cec35bad0d9cf4cd3f9118e3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf9560330205b783d8283335ee12bfae472e9563bf223dc6cb6f4f1456773bed7ee3a161;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf004fd9ba995a0a3ee72c312218b4eea2975b4762b1a4fc0f519a20111b78fcd37974078;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a456a93fbc92201bf50991b458279218e0212725507d7aa78c98aa04bd4236a7f0c21ee9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a5cd1da73f013ee2c15506a2d2f83001a3c0a5ee31b7a4fb2c52dfc879863bb90e715135;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h189bf3820c65e6774c8ce70900462f812162c70cdeba06b4b7466bfdf03348f0f1036598;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc7f3fdb75bca32f68c5403941ee22f18ed4a14cf569a8fbfbb39a7b43c11553feee67c46;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eabb174c7734f6d6063103014782d928d0d90cf9b02011c2ca4c8ecf6c39d0380311c3c5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1737628a62fec0d8e46430607ef1372a57d2c964ace4cc7202432bd53a1c0d471979c89a1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c40ac9eff76878aa97cc26d5b39a75151cfd7c0c88a7ee0df2769d52ec5477deac3c4f4b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb4ee5659e23e9178809222221028677e7728b7c3f9cece6e519ee53d5f4af17a6c3b7c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b0a3282cd7acc2b51883d570d85cf992c3b6d87cd0246015b6e8ee1516dc509f29e43b09;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13cdf45863cbd8e24750deb919bfb6c3243654f780482e723c4bff9517d4363a852aab1d4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ecb90d656e4436bdb2b7f440909889bd71a9c3b910e931817d2dd20c6d35321ac7bbd6b3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfd2dd7f0ea65898dd1ea584cb4cefc4df1e87d5526b584d153172bb87136e792b4e40fff;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h131a345ef60078f5bbc365b5d251a1ba9b21db849f255e42413eefef399e5b14152b44dab;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10a5b67597fd3f5dbbce0fcff271f657812da476dc0e9b3025c15a6312b9d26c8699a3179;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h877042f061f9adb7cc66e524377677d2638861ad88fb29b4d74da3f64727c08e8b55d2cb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d396707f899db78be5e61af802b39be98ea0f12b900eaaee66589cecb52f702476c19429;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12cbefc855a2a15c6da548e997a1f36c22c50f0fb3a9cbf9b33c911a3d280d48529b44c8a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcbebc89b536ed1d664abc4e1a4f11beb9cb86fdeac2bc68b361c080b8cfd909162dddb27;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h157a02e2d6c9e37e3a1d22e538fd5da273d0a19cec52f0d0050be3ea33a8420ca0bef828c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd6ec4e70586588ad785cc01640ddb9c23bddbe3cb80780135001f9769c69c13282220f0c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h133e742bd4d9fb3367e5cf7de146bd7a8a2d39989e34244c3ffe47dc7b93a0f5e4a6f17b4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14acaded72ef885323869271d47893c89bbb3ed4a507cbf79df1b7ff4b4ec3442122ed2f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2882c9f9fa939a08ee7a494c83e611d53f773246a32ddd3ce77f6c4cd0264ce1d83b322c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fe51cd69a76203272b0a4b3b7ead201de5f0a516c5107d56a57a97e86cdf63ea50c3bc1a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hde280d5463f0268a91bbcbf7cb8ba2c16b8bacce5e15535f9adbb70f688c733f3e8b8c28;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4f91ef71491752fff3303859d0b9b9c91cf6c584057bf1fa294a9d084a8a46f7fee4bc6b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hebeafe8743d9def556ca8d52e20442c820bf92a93964ad1347a061d7b6250672d0f8855a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb2b2eb417353fbd50edcf625e057f3c76bd65609d6435044f3bb6c907a3e5bd29ebf5d9b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he75c5298714594328bcce29b1937b63ac4f90474cc378d24c466eb9c620d70c0b2f4e829;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h118f6e9ddd7145d32607187d58a382da537d5c52b8f99cc9a8b92db457cb663abcf0e1af9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf1b82664d1e32e5103125788329bcc69856f8b0381c23cae47dd31d40d6ba8dc8a86a54;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c8773c43386b71ab2496b856d3bcfc9848193407723d646ecc2dc20e3e5e66e513121e8c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14ae6e832f4481c1cb542f8592d0511c3bb75ac2b2b22a9be3835b7202038abf304ca7257;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14a298ea7b4055d1f056415c5f90826f67bb261c5997144a2b9464ed2e715e93da3545dd1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7593ad41f5753045ea5fae0737945e42a749de0a20af20ef563e9972410e3ef72dc2a078;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8671fb1701dc37047c74792a0f5da1442d2bc4c5390e0027e9b520a59f0c460c349e57d6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h86c45fce6d455e73abb9453752ea822f499ee9032d1be32acab73872ff177cce243e13c0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hec202320cedef070629e7fbf9cc243c3ecfcbe9e33191766608c0e7a6f29761d2b2cf62e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h29b17fe43ff37ee8a174435bde0bc05166f503342ffcf27eac6e1ed42093ffa03c581079;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h23d8ae2588eb34ae604b1493053d239a1b43bd9d67a4930f09f25927a5b3e63a7246d59e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf3953fa53f613889c23990c7486d4fb9fe6c46ad46701e953d2dd98d733b69564c6c736c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1118a201b0282048c4faa5dd7ccd8afb7ce9e8be334ba42145a7a2b58000d85cba13a9fb4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cd7404069a538afd44f4a60ed044250803ba4df0ac9f409218f1042132c6963704c3fbe2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcdce3072a12a74cb5c14302f6aabc41b9c6fb447f828b994d5625a033891d720ba493f1f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h168d8f50f5fb064f6920dff1d8732942209dfbc8d08dc2668ba68b51924bfbae07c8c0d1d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7946a0c39bff7277f90a226033d5feee7fde62aa3ac56b99ba9dd38d1807430aba4767df;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1706f0a42e63b615fed30c37a011a0b323833f0776214cceae17c0c8270c535fc5b8f6ad1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd257e1fe852d99d92a5fc2c0ff0c4bd6ce92d8f8cc464e9a31317b8835127af84bdde6a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c7f3ca9353c578106692aa1546d5b603de9f70631fe13fb00f566dc521f762e9a19494ae;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h129701882af96d5e0d8b1c0d060a4a540b36f801f1d46dbbadb25d82b791619f3213f12a8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h105b9d5b13238651018665d9d3c2f36a83ede27745e88ddb5999fedac8a1a8aef7a6b5c67;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h134800f49aa3faf6ec6087d40899533df20dbd8d1ba0a1116f499990c251be13544355039;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h101e9eeb923446324e0468dcbed283b6d88ec3da45b4953a10689ee829c43a2cf8557e0bc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h967b082f84f8a1de2d1cafe8cbdb338961fd6187cc6271308b592927221bae95d3a1ef3c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7f4a155dd89a4af77f8e2dbaa889a67ccbe21764f49abd77ec96c3f10211457a51de8211;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15d520427fbe00b5beb102ef8d1f78f66a00ec6d578a4cc92acb4e9490a230fe77a48a555;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c4d5f342a7b468dae8385ff0cd490b52d6d00691eae41061ff44ce746269044ff59fc01a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7c584c19c1db990831194f8a24b3781956d80c1031509b28314ee989b54f460933b99ffe;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9470bbf529539815bfd0b4f35be743bb961274a1d3f90abbcdc16ac2ac7ad5e936243aa2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11be40b84a63af2d2fbbd1974a94447fc624f711d7713b371505c474b135f695025529075;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9a99f2c6fac5c3ffa21a4f464b76e5108eb093b124366ac54a86c23d53fa77a3f2670eb8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h158343f8a5b551f9562f0d69ab8a75a96b47519a4fd4828353ad7d9b91acc818a2826430;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e9b94996b685f5c4c21dcb480c23e0d0b559d992efac272b5a37d6c0b85d0ad5b77e0542;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2b2b510b37f82a8764684f771c01f4504237a3ecda6e91d3c4ceee584196509fd63381af;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h124637fef51fe7854c7e40696c8d2afe91a3afd82f391b26e17c3e6f8febe2da2a1fdefe;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11c91921f3508ffc2727bdba4f93abcf36f520d7c41b62a96b54da23bcedeeb5a11b89aa1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18a8c02af70169f817cea872cbe6524dd97467f24a05b2dfd76e0a6fc1043caa9cce0948;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd37eea62bd3d48d268c1a24e6de8dafd50fee5f7199362fe5d3d3892bf0bd2ebae6cacd3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11f0fccca3526c11b3613dd3544ceb8baea55e5b37de8bfe3dabac3690893e1b2630f9ede;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cc84281b1c508df5202f6feafece413fdb9e5a289e8be9927f3e8053ae2f42ca652e173c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h107a0d21e8884d1284b3673cfb2478f58c8a1e5a0aca4c01a634269d0040e5dc4402b6b39;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b37d4b3ed5441d8034486c083642d5430875db5ba45dabc2a6b7eb2f2689335840436d60;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11c6afc1bd1f6905951d1d04edafffbda7f5e457dba6e62c78fa0f8ca25b26bf38453134e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ddc085d0447e5a3a91e4d5e3516f20ed41ccf1d6547936ea7738b4de49c50fe543f314aa;
        #1
        $finish();
    end
endmodule
