module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37);
    reg [63:0] src0;
    reg [63:0] src1;
    reg [63:0] src2;
    reg [63:0] src3;
    reg [63:0] src4;
    reg [63:0] src5;
    reg [63:0] src6;
    reg [63:0] src7;
    reg [63:0] src8;
    reg [63:0] src9;
    reg [63:0] src10;
    reg [63:0] src11;
    reg [63:0] src12;
    reg [63:0] src13;
    reg [63:0] src14;
    reg [63:0] src15;
    reg [63:0] src16;
    reg [63:0] src17;
    reg [63:0] src18;
    reg [63:0] src19;
    reg [63:0] src20;
    reg [63:0] src21;
    reg [63:0] src22;
    reg [63:0] src23;
    reg [63:0] src24;
    reg [63:0] src25;
    reg [63:0] src26;
    reg [63:0] src27;
    reg [63:0] src28;
    reg [63:0] src29;
    reg [63:0] src30;
    reg [63:0] src31;
    compressor_CLA64_32 compressor_CLA64_32(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37));
    initial begin
        src0 <= 64'h0;
        src1 <= 64'h0;
        src2 <= 64'h0;
        src3 <= 64'h0;
        src4 <= 64'h0;
        src5 <= 64'h0;
        src6 <= 64'h0;
        src7 <= 64'h0;
        src8 <= 64'h0;
        src9 <= 64'h0;
        src10 <= 64'h0;
        src11 <= 64'h0;
        src12 <= 64'h0;
        src13 <= 64'h0;
        src14 <= 64'h0;
        src15 <= 64'h0;
        src16 <= 64'h0;
        src17 <= 64'h0;
        src18 <= 64'h0;
        src19 <= 64'h0;
        src20 <= 64'h0;
        src21 <= 64'h0;
        src22 <= 64'h0;
        src23 <= 64'h0;
        src24 <= 64'h0;
        src25 <= 64'h0;
        src26 <= 64'h0;
        src27 <= 64'h0;
        src28 <= 64'h0;
        src29 <= 64'h0;
        src30 <= 64'h0;
        src31 <= 64'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
    end
endmodule
module compressor_CLA64_32(
    input [63:0]src0,
    input [63:0]src1,
    input [63:0]src2,
    input [63:0]src3,
    input [63:0]src4,
    input [63:0]src5,
    input [63:0]src6,
    input [63:0]src7,
    input [63:0]src8,
    input [63:0]src9,
    input [63:0]src10,
    input [63:0]src11,
    input [63:0]src12,
    input [63:0]src13,
    input [63:0]src14,
    input [63:0]src15,
    input [63:0]src16,
    input [63:0]src17,
    input [63:0]src18,
    input [63:0]src19,
    input [63:0]src20,
    input [63:0]src21,
    input [63:0]src22,
    input [63:0]src23,
    input [63:0]src24,
    input [63:0]src25,
    input [63:0]src26,
    input [63:0]src27,
    input [63:0]src28,
    input [63:0]src29,
    input [63:0]src30,
    input [63:0]src31,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [0:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [0:0] comp_out12;
    wire [0:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [0:0] comp_out36;
    wire [0:0] comp_out37;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], 1'h0, 1'h0, comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], 1'h0, comp_out1[1], comp_out0[1]}),
        .dst({dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [63:0] src0,
      input wire [63:0] src1,
      input wire [63:0] src2,
      input wire [63:0] src3,
      input wire [63:0] src4,
      input wire [63:0] src5,
      input wire [63:0] src6,
      input wire [63:0] src7,
      input wire [63:0] src8,
      input wire [63:0] src9,
      input wire [63:0] src10,
      input wire [63:0] src11,
      input wire [63:0] src12,
      input wire [63:0] src13,
      input wire [63:0] src14,
      input wire [63:0] src15,
      input wire [63:0] src16,
      input wire [63:0] src17,
      input wire [63:0] src18,
      input wire [63:0] src19,
      input wire [63:0] src20,
      input wire [63:0] src21,
      input wire [63:0] src22,
      input wire [63:0] src23,
      input wire [63:0] src24,
      input wire [63:0] src25,
      input wire [63:0] src26,
      input wire [63:0] src27,
      input wire [63:0] src28,
      input wire [63:0] src29,
      input wire [63:0] src30,
      input wire [63:0] src31,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [0:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [0:0] dst12,
      output wire [0:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [0:0] dst36,
      output wire [0:0] dst37);

   wire [63:0] stage0_0;
   wire [63:0] stage0_1;
   wire [63:0] stage0_2;
   wire [63:0] stage0_3;
   wire [63:0] stage0_4;
   wire [63:0] stage0_5;
   wire [63:0] stage0_6;
   wire [63:0] stage0_7;
   wire [63:0] stage0_8;
   wire [63:0] stage0_9;
   wire [63:0] stage0_10;
   wire [63:0] stage0_11;
   wire [63:0] stage0_12;
   wire [63:0] stage0_13;
   wire [63:0] stage0_14;
   wire [63:0] stage0_15;
   wire [63:0] stage0_16;
   wire [63:0] stage0_17;
   wire [63:0] stage0_18;
   wire [63:0] stage0_19;
   wire [63:0] stage0_20;
   wire [63:0] stage0_21;
   wire [63:0] stage0_22;
   wire [63:0] stage0_23;
   wire [63:0] stage0_24;
   wire [63:0] stage0_25;
   wire [63:0] stage0_26;
   wire [63:0] stage0_27;
   wire [63:0] stage0_28;
   wire [63:0] stage0_29;
   wire [63:0] stage0_30;
   wire [63:0] stage0_31;
   wire [23:0] stage1_0;
   wire [19:0] stage1_1;
   wire [23:0] stage1_2;
   wire [31:0] stage1_3;
   wire [34:0] stage1_4;
   wire [34:0] stage1_5;
   wire [27:0] stage1_6;
   wire [23:0] stage1_7;
   wire [34:0] stage1_8;
   wire [27:0] stage1_9;
   wire [28:0] stage1_10;
   wire [28:0] stage1_11;
   wire [43:0] stage1_12;
   wire [22:0] stage1_13;
   wire [44:0] stage1_14;
   wire [31:0] stage1_15;
   wire [20:0] stage1_16;
   wire [34:0] stage1_17;
   wire [42:0] stage1_18;
   wire [19:0] stage1_19;
   wire [37:0] stage1_20;
   wire [27:0] stage1_21;
   wire [19:0] stage1_22;
   wire [47:0] stage1_23;
   wire [43:0] stage1_24;
   wire [23:0] stage1_25;
   wire [27:0] stage1_26;
   wire [21:0] stage1_27;
   wire [27:0] stage1_28;
   wire [37:0] stage1_29;
   wire [29:0] stage1_30;
   wire [27:0] stage1_31;
   wire [17:0] stage1_32;
   wire [8:0] stage1_33;
   wire [18:0] stage2_0;
   wire [5:0] stage2_1;
   wire [21:0] stage2_2;
   wire [17:0] stage2_3;
   wire [18:0] stage2_4;
   wire [26:0] stage2_5;
   wire [10:0] stage2_6;
   wire [8:0] stage2_7;
   wire [16:0] stage2_8;
   wire [15:0] stage2_9;
   wire [8:0] stage2_10;
   wire [11:0] stage2_11;
   wire [16:0] stage2_12;
   wire [17:0] stage2_13;
   wire [12:0] stage2_14;
   wire [23:0] stage2_15;
   wire [13:0] stage2_16;
   wire [13:0] stage2_17;
   wire [20:0] stage2_18;
   wire [15:0] stage2_19;
   wire [23:0] stage2_20;
   wire [12:0] stage2_21;
   wire [17:0] stage2_22;
   wire [16:0] stage2_23;
   wire [23:0] stage2_24;
   wire [17:0] stage2_25;
   wire [11:0] stage2_26;
   wire [16:0] stage2_27;
   wire [17:0] stage2_28;
   wire [17:0] stage2_29;
   wire [11:0] stage2_30;
   wire [21:0] stage2_31;
   wire [7:0] stage2_32;
   wire [7:0] stage2_33;
   wire [3:0] stage2_34;
   wire [0:0] stage2_35;
   wire [6:0] stage3_0;
   wire [5:0] stage3_1;
   wire [6:0] stage3_2;
   wire [6:0] stage3_3;
   wire [11:0] stage3_4;
   wire [5:0] stage3_5;
   wire [7:0] stage3_6;
   wire [10:0] stage3_7;
   wire [3:0] stage3_8;
   wire [7:0] stage3_9;
   wire [5:0] stage3_10;
   wire [3:0] stage3_11;
   wire [6:0] stage3_12;
   wire [8:0] stage3_13;
   wire [7:0] stage3_14;
   wire [6:0] stage3_15;
   wire [5:0] stage3_16;
   wire [7:0] stage3_17;
   wire [7:0] stage3_18;
   wire [12:0] stage3_19;
   wire [4:0] stage3_20;
   wire [8:0] stage3_21;
   wire [10:0] stage3_22;
   wire [6:0] stage3_23;
   wire [6:0] stage3_24;
   wire [8:0] stage3_25;
   wire [7:0] stage3_26;
   wire [4:0] stage3_27;
   wire [6:0] stage3_28;
   wire [8:0] stage3_29;
   wire [5:0] stage3_30;
   wire [8:0] stage3_31;
   wire [12:0] stage3_32;
   wire [6:0] stage3_33;
   wire [1:0] stage3_34;
   wire [0:0] stage3_35;
   wire [0:0] stage3_36;
   wire [0:0] stage3_37;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [2:0] stage4_2;
   wire [2:0] stage4_3;
   wire [4:0] stage4_4;
   wire [3:0] stage4_5;
   wire [2:0] stage4_6;
   wire [5:0] stage4_7;
   wire [4:0] stage4_8;
   wire [2:0] stage4_9;
   wire [1:0] stage4_10;
   wire [2:0] stage4_11;
   wire [1:0] stage4_12;
   wire [5:0] stage4_13;
   wire [3:0] stage4_14;
   wire [2:0] stage4_15;
   wire [1:0] stage4_16;
   wire [4:0] stage4_17;
   wire [5:0] stage4_18;
   wire [2:0] stage4_19;
   wire [3:0] stage4_20;
   wire [4:0] stage4_21;
   wire [2:0] stage4_22;
   wire [3:0] stage4_23;
   wire [5:0] stage4_24;
   wire [3:0] stage4_25;
   wire [4:0] stage4_26;
   wire [2:0] stage4_27;
   wire [1:0] stage4_28;
   wire [4:0] stage4_29;
   wire [3:0] stage4_30;
   wire [3:0] stage4_31;
   wire [3:0] stage4_32;
   wire [3:0] stage4_33;
   wire [4:0] stage4_34;
   wire [1:0] stage4_35;
   wire [0:0] stage4_36;
   wire [0:0] stage4_37;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [0:0] stage5_2;
   wire [1:0] stage5_3;
   wire [1:0] stage5_4;
   wire [1:0] stage5_5;
   wire [1:0] stage5_6;
   wire [1:0] stage5_7;
   wire [1:0] stage5_8;
   wire [1:0] stage5_9;
   wire [1:0] stage5_10;
   wire [1:0] stage5_11;
   wire [0:0] stage5_12;
   wire [0:0] stage5_13;
   wire [1:0] stage5_14;
   wire [1:0] stage5_15;
   wire [1:0] stage5_16;
   wire [1:0] stage5_17;
   wire [1:0] stage5_18;
   wire [1:0] stage5_19;
   wire [1:0] stage5_20;
   wire [1:0] stage5_21;
   wire [1:0] stage5_22;
   wire [1:0] stage5_23;
   wire [1:0] stage5_24;
   wire [1:0] stage5_25;
   wire [1:0] stage5_26;
   wire [1:0] stage5_27;
   wire [1:0] stage5_28;
   wire [1:0] stage5_29;
   wire [1:0] stage5_30;
   wire [1:0] stage5_31;
   wire [1:0] stage5_32;
   wire [1:0] stage5_33;
   wire [1:0] stage5_34;
   wire [1:0] stage5_35;
   wire [0:0] stage5_36;
   wire [0:0] stage5_37;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign dst0 = stage5_0;
   assign dst1 = stage5_1;
   assign dst2 = stage5_2;
   assign dst3 = stage5_3;
   assign dst4 = stage5_4;
   assign dst5 = stage5_5;
   assign dst6 = stage5_6;
   assign dst7 = stage5_7;
   assign dst8 = stage5_8;
   assign dst9 = stage5_9;
   assign dst10 = stage5_10;
   assign dst11 = stage5_11;
   assign dst12 = stage5_12;
   assign dst13 = stage5_13;
   assign dst14 = stage5_14;
   assign dst15 = stage5_15;
   assign dst16 = stage5_16;
   assign dst17 = stage5_17;
   assign dst18 = stage5_18;
   assign dst19 = stage5_19;
   assign dst20 = stage5_20;
   assign dst21 = stage5_21;
   assign dst22 = stage5_22;
   assign dst23 = stage5_23;
   assign dst24 = stage5_24;
   assign dst25 = stage5_25;
   assign dst26 = stage5_26;
   assign dst27 = stage5_27;
   assign dst28 = stage5_28;
   assign dst29 = stage5_29;
   assign dst30 = stage5_30;
   assign dst31 = stage5_31;
   assign dst32 = stage5_32;
   assign dst33 = stage5_33;
   assign dst34 = stage5_34;
   assign dst35 = stage5_35;
   assign dst36 = stage5_36;
   assign dst37 = stage5_37;

   gpc1163_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2]},
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[0]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc1163_5 gpc1 (
      {stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[1]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc1163_5 gpc2 (
      {stage0_0[6], stage0_0[7], stage0_0[8]},
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[2]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc1163_5 gpc3 (
      {stage0_0[9], stage0_0[10], stage0_0[11]},
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[3]},
      {stage0_3[3]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc1163_5 gpc4 (
      {stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_2[4]},
      {stage0_3[4]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_2[5], stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26]},
      {stage0_2[11], stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32]},
      {stage0_2[17], stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[33], stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38]},
      {stage0_2[23], stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_2[29], stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc606_5 gpc10 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49], stage0_0[50]},
      {stage0_2[35], stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc606_5 gpc11 (
      {stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_3[5], stage0_3[6], stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10]},
      {stage1_5[0],stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11]}
   );
   gpc606_5 gpc12 (
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_3[11], stage0_3[12], stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16]},
      {stage1_5[1],stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12]}
   );
   gpc606_5 gpc13 (
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_3[17], stage0_3[18], stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22]},
      {stage1_5[2],stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13]}
   );
   gpc606_5 gpc14 (
      {stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26], stage0_3[27], stage0_3[28]},
      {stage1_5[3],stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14]}
   );
   gpc606_5 gpc15 (
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59]},
      {stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32], stage0_3[33], stage0_3[34]},
      {stage1_5[4],stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15]}
   );
   gpc606_5 gpc16 (
      {stage0_2[41], stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[5],stage1_4[16],stage1_3[16],stage1_2[16]}
   );
   gpc606_5 gpc17 (
      {stage0_2[47], stage0_2[48], stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[6],stage1_4[17],stage1_3[17],stage1_2[17]}
   );
   gpc606_5 gpc18 (
      {stage0_2[53], stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[7],stage1_4[18],stage1_3[18],stage1_2[18]}
   );
   gpc615_5 gpc19 (
      {stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39]},
      {stage0_4[18]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[3],stage1_5[8],stage1_4[19],stage1_3[19]}
   );
   gpc615_5 gpc20 (
      {stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44]},
      {stage0_4[19]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[4],stage1_5[9],stage1_4[20],stage1_3[20]}
   );
   gpc615_5 gpc21 (
      {stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49]},
      {stage0_4[20]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[5],stage1_5[10],stage1_4[21],stage1_3[21]}
   );
   gpc615_5 gpc22 (
      {stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54]},
      {stage0_4[21]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[6],stage1_5[11],stage1_4[22],stage1_3[22]}
   );
   gpc606_5 gpc23 (
      {stage0_4[22], stage0_4[23], stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[4],stage1_6[7],stage1_5[12],stage1_4[23]}
   );
   gpc606_5 gpc24 (
      {stage0_4[28], stage0_4[29], stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[5],stage1_6[8],stage1_5[13],stage1_4[24]}
   );
   gpc606_5 gpc25 (
      {stage0_4[34], stage0_4[35], stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[6],stage1_6[9],stage1_5[14],stage1_4[25]}
   );
   gpc606_5 gpc26 (
      {stage0_4[40], stage0_4[41], stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[7],stage1_6[10],stage1_5[15],stage1_4[26]}
   );
   gpc606_5 gpc27 (
      {stage0_4[46], stage0_4[47], stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[8],stage1_6[11],stage1_5[16],stage1_4[27]}
   );
   gpc606_5 gpc28 (
      {stage0_4[52], stage0_4[53], stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[9],stage1_6[12],stage1_5[17],stage1_4[28]}
   );
   gpc606_5 gpc29 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[6],stage1_7[10],stage1_6[13],stage1_5[18]}
   );
   gpc606_5 gpc30 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[7],stage1_7[11],stage1_6[14],stage1_5[19]}
   );
   gpc606_5 gpc31 (
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[8],stage1_7[12],stage1_6[15],stage1_5[20]}
   );
   gpc615_5 gpc32 (
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46]},
      {stage0_6[36]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[9],stage1_7[13],stage1_6[16],stage1_5[21]}
   );
   gpc615_5 gpc33 (
      {stage0_5[47], stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51]},
      {stage0_6[37]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[10],stage1_7[14],stage1_6[17],stage1_5[22]}
   );
   gpc615_5 gpc34 (
      {stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41], stage0_6[42]},
      {stage0_7[30]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[5],stage1_8[11],stage1_7[15],stage1_6[18]}
   );
   gpc615_5 gpc35 (
      {stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage0_7[31]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[6],stage1_8[12],stage1_7[16],stage1_6[19]}
   );
   gpc615_5 gpc36 (
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52]},
      {stage0_7[32]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[7],stage1_8[13],stage1_7[17],stage1_6[20]}
   );
   gpc615_5 gpc37 (
      {stage0_6[53], stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57]},
      {stage0_7[33]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[8],stage1_8[14],stage1_7[18],stage1_6[21]}
   );
   gpc606_5 gpc38 (
      {stage0_7[34], stage0_7[35], stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[4],stage1_9[9],stage1_8[15],stage1_7[19]}
   );
   gpc606_5 gpc39 (
      {stage0_7[40], stage0_7[41], stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[5],stage1_9[10],stage1_8[16],stage1_7[20]}
   );
   gpc606_5 gpc40 (
      {stage0_7[46], stage0_7[47], stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[6],stage1_9[11],stage1_8[17],stage1_7[21]}
   );
   gpc606_5 gpc41 (
      {stage0_7[52], stage0_7[53], stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[7],stage1_9[12],stage1_8[18],stage1_7[22]}
   );
   gpc606_5 gpc42 (
      {stage0_7[58], stage0_7[59], stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[8],stage1_9[13],stage1_8[19],stage1_7[23]}
   );
   gpc606_5 gpc43 (
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[5],stage1_10[9],stage1_9[14],stage1_8[20]}
   );
   gpc606_5 gpc44 (
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[6],stage1_10[10],stage1_9[15],stage1_8[21]}
   );
   gpc606_5 gpc45 (
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[7],stage1_10[11],stage1_9[16],stage1_8[22]}
   );
   gpc606_5 gpc46 (
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[8],stage1_10[12],stage1_9[17],stage1_8[23]}
   );
   gpc606_5 gpc47 (
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[9],stage1_10[13],stage1_9[18],stage1_8[24]}
   );
   gpc606_5 gpc48 (
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[5],stage1_11[10],stage1_10[14],stage1_9[19]}
   );
   gpc606_5 gpc49 (
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[6],stage1_11[11],stage1_10[15],stage1_9[20]}
   );
   gpc606_5 gpc50 (
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[7],stage1_11[12],stage1_10[16],stage1_9[21]}
   );
   gpc606_5 gpc51 (
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[8],stage1_11[13],stage1_10[17],stage1_9[22]}
   );
   gpc606_5 gpc52 (
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[9],stage1_11[14],stage1_10[18],stage1_9[23]}
   );
   gpc615_5 gpc53 (
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34]},
      {stage0_11[30]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[5],stage1_12[10],stage1_11[15],stage1_10[19]}
   );
   gpc615_5 gpc54 (
      {stage0_10[35], stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39]},
      {stage0_11[31]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[6],stage1_12[11],stage1_11[16],stage1_10[20]}
   );
   gpc615_5 gpc55 (
      {stage0_10[40], stage0_10[41], stage0_10[42], stage0_10[43], stage0_10[44]},
      {stage0_11[32]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[7],stage1_12[12],stage1_11[17],stage1_10[21]}
   );
   gpc615_5 gpc56 (
      {stage0_10[45], stage0_10[46], stage0_10[47], stage0_10[48], stage0_10[49]},
      {stage0_11[33]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[8],stage1_12[13],stage1_11[18],stage1_10[22]}
   );
   gpc615_5 gpc57 (
      {stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53], stage0_10[54]},
      {stage0_11[34]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[9],stage1_12[14],stage1_11[19],stage1_10[23]}
   );
   gpc615_5 gpc58 (
      {stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage0_11[35]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[10],stage1_12[15],stage1_11[20],stage1_10[24]}
   );
   gpc615_5 gpc59 (
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40]},
      {stage0_12[36]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[6],stage1_13[11],stage1_12[16],stage1_11[21]}
   );
   gpc615_5 gpc60 (
      {stage0_11[41], stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45]},
      {stage0_12[37]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[7],stage1_13[12],stage1_12[17],stage1_11[22]}
   );
   gpc615_5 gpc61 (
      {stage0_11[46], stage0_11[47], stage0_11[48], stage0_11[49], stage0_11[50]},
      {stage0_12[38]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[8],stage1_13[13],stage1_12[18],stage1_11[23]}
   );
   gpc615_5 gpc62 (
      {stage0_11[51], stage0_11[52], stage0_11[53], stage0_11[54], stage0_11[55]},
      {stage0_12[39]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[9],stage1_13[14],stage1_12[19],stage1_11[24]}
   );
   gpc615_5 gpc63 (
      {stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59], stage0_11[60]},
      {stage0_12[40]},
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage1_15[4],stage1_14[10],stage1_13[15],stage1_12[20],stage1_11[25]}
   );
   gpc615_5 gpc64 (
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34]},
      {stage0_14[0]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[0],stage1_15[5],stage1_14[11],stage1_13[16]}
   );
   gpc615_5 gpc65 (
      {stage0_13[35], stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39]},
      {stage0_14[1]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[1],stage1_15[6],stage1_14[12],stage1_13[17]}
   );
   gpc615_5 gpc66 (
      {stage0_13[40], stage0_13[41], stage0_13[42], stage0_13[43], stage0_13[44]},
      {stage0_14[2]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[2],stage1_15[7],stage1_14[13],stage1_13[18]}
   );
   gpc615_5 gpc67 (
      {stage0_13[45], stage0_13[46], stage0_13[47], stage0_13[48], stage0_13[49]},
      {stage0_14[3]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[3],stage1_15[8],stage1_14[14],stage1_13[19]}
   );
   gpc615_5 gpc68 (
      {stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53], stage0_13[54]},
      {stage0_14[4]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[4],stage1_15[9],stage1_14[15],stage1_13[20]}
   );
   gpc615_5 gpc69 (
      {stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage0_14[5]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[5],stage1_15[10],stage1_14[16],stage1_13[21]}
   );
   gpc615_5 gpc70 (
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], 1'b0},
      {stage0_14[6]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[6],stage1_15[11],stage1_14[17],stage1_13[22]}
   );
   gpc606_5 gpc71 (
      {stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11], stage0_14[12]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[7],stage1_16[7],stage1_15[12],stage1_14[18]}
   );
   gpc606_5 gpc72 (
      {stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17], stage0_14[18]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[8],stage1_16[8],stage1_15[13],stage1_14[19]}
   );
   gpc606_5 gpc73 (
      {stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23], stage0_14[24]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[9],stage1_16[9],stage1_15[14],stage1_14[20]}
   );
   gpc606_5 gpc74 (
      {stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29], stage0_14[30]},
      {stage0_16[18], stage0_16[19], stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23]},
      {stage1_18[3],stage1_17[10],stage1_16[10],stage1_15[15],stage1_14[21]}
   );
   gpc606_5 gpc75 (
      {stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35], stage0_14[36]},
      {stage0_16[24], stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29]},
      {stage1_18[4],stage1_17[11],stage1_16[11],stage1_15[16],stage1_14[22]}
   );
   gpc606_5 gpc76 (
      {stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41], stage0_14[42]},
      {stage0_16[30], stage0_16[31], stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35]},
      {stage1_18[5],stage1_17[12],stage1_16[12],stage1_15[17],stage1_14[23]}
   );
   gpc615_5 gpc77 (
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46]},
      {stage0_16[36]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[6],stage1_17[13],stage1_16[13],stage1_15[18]}
   );
   gpc615_5 gpc78 (
      {stage0_15[47], stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51]},
      {stage0_16[37]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[7],stage1_17[14],stage1_16[14],stage1_15[19]}
   );
   gpc606_5 gpc79 (
      {stage0_16[38], stage0_16[39], stage0_16[40], stage0_16[41], stage0_16[42], stage0_16[43]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[2],stage1_18[8],stage1_17[15],stage1_16[15]}
   );
   gpc606_5 gpc80 (
      {stage0_16[44], stage0_16[45], stage0_16[46], stage0_16[47], stage0_16[48], stage0_16[49]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[3],stage1_18[9],stage1_17[16],stage1_16[16]}
   );
   gpc606_5 gpc81 (
      {stage0_16[50], stage0_16[51], stage0_16[52], stage0_16[53], stage0_16[54], stage0_16[55]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[4],stage1_18[10],stage1_17[17],stage1_16[17]}
   );
   gpc606_5 gpc82 (
      {stage0_16[56], stage0_16[57], stage0_16[58], stage0_16[59], stage0_16[60], stage0_16[61]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[5],stage1_18[11],stage1_17[18],stage1_16[18]}
   );
   gpc1163_5 gpc83 (
      {stage0_17[12], stage0_17[13], stage0_17[14]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage0_19[0]},
      {stage0_20[0]},
      {stage1_21[0],stage1_20[4],stage1_19[6],stage1_18[12],stage1_17[19]}
   );
   gpc1163_5 gpc84 (
      {stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage0_19[1]},
      {stage0_20[1]},
      {stage1_21[1],stage1_20[5],stage1_19[7],stage1_18[13],stage1_17[20]}
   );
   gpc1163_5 gpc85 (
      {stage0_17[18], stage0_17[19], stage0_17[20]},
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage0_19[2]},
      {stage0_20[2]},
      {stage1_21[2],stage1_20[6],stage1_19[8],stage1_18[14],stage1_17[21]}
   );
   gpc606_5 gpc86 (
      {stage0_17[21], stage0_17[22], stage0_17[23], stage0_17[24], stage0_17[25], stage0_17[26]},
      {stage0_19[3], stage0_19[4], stage0_19[5], stage0_19[6], stage0_19[7], stage0_19[8]},
      {stage1_21[3],stage1_20[7],stage1_19[9],stage1_18[15],stage1_17[22]}
   );
   gpc606_5 gpc87 (
      {stage0_17[27], stage0_17[28], stage0_17[29], stage0_17[30], stage0_17[31], stage0_17[32]},
      {stage0_19[9], stage0_19[10], stage0_19[11], stage0_19[12], stage0_19[13], stage0_19[14]},
      {stage1_21[4],stage1_20[8],stage1_19[10],stage1_18[16],stage1_17[23]}
   );
   gpc606_5 gpc88 (
      {stage0_17[33], stage0_17[34], stage0_17[35], stage0_17[36], stage0_17[37], stage0_17[38]},
      {stage0_19[15], stage0_19[16], stage0_19[17], stage0_19[18], stage0_19[19], stage0_19[20]},
      {stage1_21[5],stage1_20[9],stage1_19[11],stage1_18[17],stage1_17[24]}
   );
   gpc606_5 gpc89 (
      {stage0_17[39], stage0_17[40], stage0_17[41], stage0_17[42], stage0_17[43], stage0_17[44]},
      {stage0_19[21], stage0_19[22], stage0_19[23], stage0_19[24], stage0_19[25], stage0_19[26]},
      {stage1_21[6],stage1_20[10],stage1_19[12],stage1_18[18],stage1_17[25]}
   );
   gpc606_5 gpc90 (
      {stage0_17[45], stage0_17[46], stage0_17[47], stage0_17[48], stage0_17[49], stage0_17[50]},
      {stage0_19[27], stage0_19[28], stage0_19[29], stage0_19[30], stage0_19[31], stage0_19[32]},
      {stage1_21[7],stage1_20[11],stage1_19[13],stage1_18[19],stage1_17[26]}
   );
   gpc606_5 gpc91 (
      {stage0_17[51], stage0_17[52], stage0_17[53], stage0_17[54], stage0_17[55], stage0_17[56]},
      {stage0_19[33], stage0_19[34], stage0_19[35], stage0_19[36], stage0_19[37], stage0_19[38]},
      {stage1_21[8],stage1_20[12],stage1_19[14],stage1_18[20],stage1_17[27]}
   );
   gpc615_5 gpc92 (
      {stage0_19[39], stage0_19[40], stage0_19[41], stage0_19[42], stage0_19[43]},
      {stage0_20[3]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[0],stage1_21[9],stage1_20[13],stage1_19[15]}
   );
   gpc615_5 gpc93 (
      {stage0_19[44], stage0_19[45], stage0_19[46], stage0_19[47], stage0_19[48]},
      {stage0_20[4]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[1],stage1_21[10],stage1_20[14],stage1_19[16]}
   );
   gpc615_5 gpc94 (
      {stage0_19[49], stage0_19[50], stage0_19[51], stage0_19[52], stage0_19[53]},
      {stage0_20[5]},
      {stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17]},
      {stage1_23[2],stage1_22[2],stage1_21[11],stage1_20[15],stage1_19[17]}
   );
   gpc615_5 gpc95 (
      {stage0_19[54], stage0_19[55], stage0_19[56], stage0_19[57], stage0_19[58]},
      {stage0_20[6]},
      {stage0_21[18], stage0_21[19], stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23]},
      {stage1_23[3],stage1_22[3],stage1_21[12],stage1_20[16],stage1_19[18]}
   );
   gpc615_5 gpc96 (
      {stage0_19[59], stage0_19[60], stage0_19[61], stage0_19[62], stage0_19[63]},
      {stage0_20[7]},
      {stage0_21[24], stage0_21[25], stage0_21[26], stage0_21[27], stage0_21[28], stage0_21[29]},
      {stage1_23[4],stage1_22[4],stage1_21[13],stage1_20[17],stage1_19[19]}
   );
   gpc615_5 gpc97 (
      {stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11], stage0_20[12]},
      {stage0_21[30]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[5],stage1_22[5],stage1_21[14],stage1_20[18]}
   );
   gpc615_5 gpc98 (
      {stage0_20[13], stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17]},
      {stage0_21[31]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[6],stage1_22[6],stage1_21[15],stage1_20[19]}
   );
   gpc615_5 gpc99 (
      {stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22]},
      {stage0_21[32]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[7],stage1_22[7],stage1_21[16],stage1_20[20]}
   );
   gpc615_5 gpc100 (
      {stage0_20[23], stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27]},
      {stage0_21[33]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[8],stage1_22[8],stage1_21[17],stage1_20[21]}
   );
   gpc615_5 gpc101 (
      {stage0_20[28], stage0_20[29], stage0_20[30], stage0_20[31], stage0_20[32]},
      {stage0_21[34]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[9],stage1_22[9],stage1_21[18],stage1_20[22]}
   );
   gpc615_5 gpc102 (
      {stage0_20[33], stage0_20[34], stage0_20[35], stage0_20[36], stage0_20[37]},
      {stage0_21[35]},
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage1_24[5],stage1_23[10],stage1_22[10],stage1_21[19],stage1_20[23]}
   );
   gpc615_5 gpc103 (
      {stage0_20[38], stage0_20[39], stage0_20[40], stage0_20[41], stage0_20[42]},
      {stage0_21[36]},
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage1_24[6],stage1_23[11],stage1_22[11],stage1_21[20],stage1_20[24]}
   );
   gpc615_5 gpc104 (
      {stage0_20[43], stage0_20[44], stage0_20[45], stage0_20[46], stage0_20[47]},
      {stage0_21[37]},
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47]},
      {stage1_24[7],stage1_23[12],stage1_22[12],stage1_21[21],stage1_20[25]}
   );
   gpc615_5 gpc105 (
      {stage0_20[48], stage0_20[49], stage0_20[50], stage0_20[51], stage0_20[52]},
      {stage0_21[38]},
      {stage0_22[48], stage0_22[49], stage0_22[50], stage0_22[51], stage0_22[52], stage0_22[53]},
      {stage1_24[8],stage1_23[13],stage1_22[13],stage1_21[22],stage1_20[26]}
   );
   gpc615_5 gpc106 (
      {stage0_21[39], stage0_21[40], stage0_21[41], stage0_21[42], stage0_21[43]},
      {stage0_22[54]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[9],stage1_23[14],stage1_22[14],stage1_21[23]}
   );
   gpc615_5 gpc107 (
      {stage0_21[44], stage0_21[45], stage0_21[46], stage0_21[47], stage0_21[48]},
      {stage0_22[55]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[10],stage1_23[15],stage1_22[15],stage1_21[24]}
   );
   gpc615_5 gpc108 (
      {stage0_21[49], stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53]},
      {stage0_22[56]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[11],stage1_23[16],stage1_22[16],stage1_21[25]}
   );
   gpc615_5 gpc109 (
      {stage0_21[54], stage0_21[55], stage0_21[56], stage0_21[57], stage0_21[58]},
      {stage0_22[57]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[12],stage1_23[17],stage1_22[17],stage1_21[26]}
   );
   gpc615_5 gpc110 (
      {stage0_21[59], stage0_21[60], stage0_21[61], stage0_21[62], stage0_21[63]},
      {stage0_22[58]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[13],stage1_23[18],stage1_22[18],stage1_21[27]}
   );
   gpc615_5 gpc111 (
      {stage0_22[59], stage0_22[60], stage0_22[61], stage0_22[62], stage0_22[63]},
      {stage0_23[30]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[5],stage1_24[14],stage1_23[19],stage1_22[19]}
   );
   gpc606_5 gpc112 (
      {stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34], stage0_23[35], stage0_23[36]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[1],stage1_25[6],stage1_24[15],stage1_23[20]}
   );
   gpc2135_5 gpc113 (
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10]},
      {stage0_25[6], stage0_25[7], stage0_25[8]},
      {stage0_26[0]},
      {stage0_27[0], stage0_27[1]},
      {stage1_28[0],stage1_27[1],stage1_26[2],stage1_25[7],stage1_24[16]}
   );
   gpc606_5 gpc114 (
      {stage0_24[11], stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16]},
      {stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5], stage0_26[6]},
      {stage1_28[1],stage1_27[2],stage1_26[3],stage1_25[8],stage1_24[17]}
   );
   gpc606_5 gpc115 (
      {stage0_24[17], stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22]},
      {stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11], stage0_26[12]},
      {stage1_28[2],stage1_27[3],stage1_26[4],stage1_25[9],stage1_24[18]}
   );
   gpc615_5 gpc116 (
      {stage0_24[23], stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27]},
      {stage0_25[9]},
      {stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17], stage0_26[18]},
      {stage1_28[3],stage1_27[4],stage1_26[5],stage1_25[10],stage1_24[19]}
   );
   gpc615_5 gpc117 (
      {stage0_24[28], stage0_24[29], stage0_24[30], stage0_24[31], stage0_24[32]},
      {stage0_25[10]},
      {stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23], stage0_26[24]},
      {stage1_28[4],stage1_27[5],stage1_26[6],stage1_25[11],stage1_24[20]}
   );
   gpc615_5 gpc118 (
      {stage0_24[33], stage0_24[34], stage0_24[35], stage0_24[36], stage0_24[37]},
      {stage0_25[11]},
      {stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29], stage0_26[30]},
      {stage1_28[5],stage1_27[6],stage1_26[7],stage1_25[12],stage1_24[21]}
   );
   gpc615_5 gpc119 (
      {stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41], stage0_24[42]},
      {stage0_25[12]},
      {stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35], stage0_26[36]},
      {stage1_28[6],stage1_27[7],stage1_26[8],stage1_25[13],stage1_24[22]}
   );
   gpc606_5 gpc120 (
      {stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17], stage0_25[18]},
      {stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5], stage0_27[6], stage0_27[7]},
      {stage1_29[0],stage1_28[7],stage1_27[8],stage1_26[9],stage1_25[14]}
   );
   gpc606_5 gpc121 (
      {stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23], stage0_25[24]},
      {stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11], stage0_27[12], stage0_27[13]},
      {stage1_29[1],stage1_28[8],stage1_27[9],stage1_26[10],stage1_25[15]}
   );
   gpc615_5 gpc122 (
      {stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage0_26[37]},
      {stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17], stage0_27[18], stage0_27[19]},
      {stage1_29[2],stage1_28[9],stage1_27[10],stage1_26[11],stage1_25[16]}
   );
   gpc615_5 gpc123 (
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34]},
      {stage0_26[38]},
      {stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23], stage0_27[24], stage0_27[25]},
      {stage1_29[3],stage1_28[10],stage1_27[11],stage1_26[12],stage1_25[17]}
   );
   gpc615_5 gpc124 (
      {stage0_25[35], stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39]},
      {stage0_26[39]},
      {stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29], stage0_27[30], stage0_27[31]},
      {stage1_29[4],stage1_28[11],stage1_27[12],stage1_26[13],stage1_25[18]}
   );
   gpc615_5 gpc125 (
      {stage0_25[40], stage0_25[41], stage0_25[42], stage0_25[43], stage0_25[44]},
      {stage0_26[40]},
      {stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35], stage0_27[36], stage0_27[37]},
      {stage1_29[5],stage1_28[12],stage1_27[13],stage1_26[14],stage1_25[19]}
   );
   gpc615_5 gpc126 (
      {stage0_25[45], stage0_25[46], stage0_25[47], stage0_25[48], stage0_25[49]},
      {stage0_26[41]},
      {stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41], stage0_27[42], stage0_27[43]},
      {stage1_29[6],stage1_28[13],stage1_27[14],stage1_26[15],stage1_25[20]}
   );
   gpc615_5 gpc127 (
      {stage0_25[50], stage0_25[51], stage0_25[52], stage0_25[53], stage0_25[54]},
      {stage0_26[42]},
      {stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47], stage0_27[48], stage0_27[49]},
      {stage1_29[7],stage1_28[14],stage1_27[15],stage1_26[16],stage1_25[21]}
   );
   gpc615_5 gpc128 (
      {stage0_25[55], stage0_25[56], stage0_25[57], stage0_25[58], stage0_25[59]},
      {stage0_26[43]},
      {stage0_27[50], stage0_27[51], stage0_27[52], stage0_27[53], stage0_27[54], stage0_27[55]},
      {stage1_29[8],stage1_28[15],stage1_27[16],stage1_26[17],stage1_25[22]}
   );
   gpc615_5 gpc129 (
      {stage0_25[60], stage0_25[61], stage0_25[62], stage0_25[63], 1'b0},
      {stage0_26[44]},
      {stage0_27[56], stage0_27[57], stage0_27[58], stage0_27[59], stage0_27[60], stage0_27[61]},
      {stage1_29[9],stage1_28[16],stage1_27[17],stage1_26[18],stage1_25[23]}
   );
   gpc606_5 gpc130 (
      {stage0_26[45], stage0_26[46], stage0_26[47], stage0_26[48], stage0_26[49], stage0_26[50]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[10],stage1_28[17],stage1_27[18],stage1_26[19]}
   );
   gpc606_5 gpc131 (
      {stage0_26[51], stage0_26[52], stage0_26[53], stage0_26[54], stage0_26[55], stage0_26[56]},
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage1_30[1],stage1_29[11],stage1_28[18],stage1_27[19],stage1_26[20]}
   );
   gpc606_5 gpc132 (
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[0],stage1_30[2],stage1_29[12],stage1_28[19]}
   );
   gpc606_5 gpc133 (
      {stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[1],stage1_30[3],stage1_29[13],stage1_28[20]}
   );
   gpc606_5 gpc134 (
      {stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[2],stage1_30[4],stage1_29[14],stage1_28[21]}
   );
   gpc606_5 gpc135 (
      {stage0_28[30], stage0_28[31], stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[3],stage1_30[5],stage1_29[15],stage1_28[22]}
   );
   gpc606_5 gpc136 (
      {stage0_28[36], stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41]},
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage1_32[4],stage1_31[4],stage1_30[6],stage1_29[16],stage1_28[23]}
   );
   gpc606_5 gpc137 (
      {stage0_28[42], stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47]},
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage1_32[5],stage1_31[5],stage1_30[7],stage1_29[17],stage1_28[24]}
   );
   gpc606_5 gpc138 (
      {stage0_28[48], stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53]},
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage1_32[6],stage1_31[6],stage1_30[8],stage1_29[18],stage1_28[25]}
   );
   gpc615_5 gpc139 (
      {stage0_28[54], stage0_28[55], stage0_28[56], stage0_28[57], stage0_28[58]},
      {stage0_29[0]},
      {stage0_30[42], stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47]},
      {stage1_32[7],stage1_31[7],stage1_30[9],stage1_29[19],stage1_28[26]}
   );
   gpc615_5 gpc140 (
      {stage0_28[59], stage0_28[60], stage0_28[61], stage0_28[62], stage0_28[63]},
      {stage0_29[1]},
      {stage0_30[48], stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53]},
      {stage1_32[8],stage1_31[8],stage1_30[10],stage1_29[20],stage1_28[27]}
   );
   gpc606_5 gpc141 (
      {stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5], stage0_29[6], stage0_29[7]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[9],stage1_31[9],stage1_30[11],stage1_29[21]}
   );
   gpc606_5 gpc142 (
      {stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11], stage0_29[12], stage0_29[13]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[10],stage1_31[10],stage1_30[12],stage1_29[22]}
   );
   gpc606_5 gpc143 (
      {stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17], stage0_29[18], stage0_29[19]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[11],stage1_31[11],stage1_30[13],stage1_29[23]}
   );
   gpc606_5 gpc144 (
      {stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23], stage0_29[24], stage0_29[25]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[12],stage1_31[12],stage1_30[14],stage1_29[24]}
   );
   gpc606_5 gpc145 (
      {stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29], stage0_29[30], stage0_29[31]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[13],stage1_31[13],stage1_30[15],stage1_29[25]}
   );
   gpc606_5 gpc146 (
      {stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35], stage0_29[36], stage0_29[37]},
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage1_33[5],stage1_32[14],stage1_31[14],stage1_30[16],stage1_29[26]}
   );
   gpc606_5 gpc147 (
      {stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41], stage0_29[42], stage0_29[43]},
      {stage0_31[36], stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41]},
      {stage1_33[6],stage1_32[15],stage1_31[15],stage1_30[17],stage1_29[27]}
   );
   gpc606_5 gpc148 (
      {stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47], stage0_29[48], stage0_29[49]},
      {stage0_31[42], stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47]},
      {stage1_33[7],stage1_32[16],stage1_31[16],stage1_30[18],stage1_29[28]}
   );
   gpc606_5 gpc149 (
      {stage0_29[50], stage0_29[51], stage0_29[52], stage0_29[53], stage0_29[54], stage0_29[55]},
      {stage0_31[48], stage0_31[49], stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53]},
      {stage1_33[8],stage1_32[17],stage1_31[17],stage1_30[19],stage1_29[29]}
   );
   gpc1_1 gpc150 (
      {stage0_0[51]},
      {stage1_0[11]}
   );
   gpc1_1 gpc151 (
      {stage0_0[52]},
      {stage1_0[12]}
   );
   gpc1_1 gpc152 (
      {stage0_0[53]},
      {stage1_0[13]}
   );
   gpc1_1 gpc153 (
      {stage0_0[54]},
      {stage1_0[14]}
   );
   gpc1_1 gpc154 (
      {stage0_0[55]},
      {stage1_0[15]}
   );
   gpc1_1 gpc155 (
      {stage0_0[56]},
      {stage1_0[16]}
   );
   gpc1_1 gpc156 (
      {stage0_0[57]},
      {stage1_0[17]}
   );
   gpc1_1 gpc157 (
      {stage0_0[58]},
      {stage1_0[18]}
   );
   gpc1_1 gpc158 (
      {stage0_0[59]},
      {stage1_0[19]}
   );
   gpc1_1 gpc159 (
      {stage0_0[60]},
      {stage1_0[20]}
   );
   gpc1_1 gpc160 (
      {stage0_0[61]},
      {stage1_0[21]}
   );
   gpc1_1 gpc161 (
      {stage0_0[62]},
      {stage1_0[22]}
   );
   gpc1_1 gpc162 (
      {stage0_0[63]},
      {stage1_0[23]}
   );
   gpc1_1 gpc163 (
      {stage0_1[60]},
      {stage1_1[16]}
   );
   gpc1_1 gpc164 (
      {stage0_1[61]},
      {stage1_1[17]}
   );
   gpc1_1 gpc165 (
      {stage0_1[62]},
      {stage1_1[18]}
   );
   gpc1_1 gpc166 (
      {stage0_1[63]},
      {stage1_1[19]}
   );
   gpc1_1 gpc167 (
      {stage0_2[59]},
      {stage1_2[19]}
   );
   gpc1_1 gpc168 (
      {stage0_2[60]},
      {stage1_2[20]}
   );
   gpc1_1 gpc169 (
      {stage0_2[61]},
      {stage1_2[21]}
   );
   gpc1_1 gpc170 (
      {stage0_2[62]},
      {stage1_2[22]}
   );
   gpc1_1 gpc171 (
      {stage0_2[63]},
      {stage1_2[23]}
   );
   gpc1_1 gpc172 (
      {stage0_3[55]},
      {stage1_3[23]}
   );
   gpc1_1 gpc173 (
      {stage0_3[56]},
      {stage1_3[24]}
   );
   gpc1_1 gpc174 (
      {stage0_3[57]},
      {stage1_3[25]}
   );
   gpc1_1 gpc175 (
      {stage0_3[58]},
      {stage1_3[26]}
   );
   gpc1_1 gpc176 (
      {stage0_3[59]},
      {stage1_3[27]}
   );
   gpc1_1 gpc177 (
      {stage0_3[60]},
      {stage1_3[28]}
   );
   gpc1_1 gpc178 (
      {stage0_3[61]},
      {stage1_3[29]}
   );
   gpc1_1 gpc179 (
      {stage0_3[62]},
      {stage1_3[30]}
   );
   gpc1_1 gpc180 (
      {stage0_3[63]},
      {stage1_3[31]}
   );
   gpc1_1 gpc181 (
      {stage0_4[58]},
      {stage1_4[29]}
   );
   gpc1_1 gpc182 (
      {stage0_4[59]},
      {stage1_4[30]}
   );
   gpc1_1 gpc183 (
      {stage0_4[60]},
      {stage1_4[31]}
   );
   gpc1_1 gpc184 (
      {stage0_4[61]},
      {stage1_4[32]}
   );
   gpc1_1 gpc185 (
      {stage0_4[62]},
      {stage1_4[33]}
   );
   gpc1_1 gpc186 (
      {stage0_4[63]},
      {stage1_4[34]}
   );
   gpc1_1 gpc187 (
      {stage0_5[52]},
      {stage1_5[23]}
   );
   gpc1_1 gpc188 (
      {stage0_5[53]},
      {stage1_5[24]}
   );
   gpc1_1 gpc189 (
      {stage0_5[54]},
      {stage1_5[25]}
   );
   gpc1_1 gpc190 (
      {stage0_5[55]},
      {stage1_5[26]}
   );
   gpc1_1 gpc191 (
      {stage0_5[56]},
      {stage1_5[27]}
   );
   gpc1_1 gpc192 (
      {stage0_5[57]},
      {stage1_5[28]}
   );
   gpc1_1 gpc193 (
      {stage0_5[58]},
      {stage1_5[29]}
   );
   gpc1_1 gpc194 (
      {stage0_5[59]},
      {stage1_5[30]}
   );
   gpc1_1 gpc195 (
      {stage0_5[60]},
      {stage1_5[31]}
   );
   gpc1_1 gpc196 (
      {stage0_5[61]},
      {stage1_5[32]}
   );
   gpc1_1 gpc197 (
      {stage0_5[62]},
      {stage1_5[33]}
   );
   gpc1_1 gpc198 (
      {stage0_5[63]},
      {stage1_5[34]}
   );
   gpc1_1 gpc199 (
      {stage0_6[58]},
      {stage1_6[22]}
   );
   gpc1_1 gpc200 (
      {stage0_6[59]},
      {stage1_6[23]}
   );
   gpc1_1 gpc201 (
      {stage0_6[60]},
      {stage1_6[24]}
   );
   gpc1_1 gpc202 (
      {stage0_6[61]},
      {stage1_6[25]}
   );
   gpc1_1 gpc203 (
      {stage0_6[62]},
      {stage1_6[26]}
   );
   gpc1_1 gpc204 (
      {stage0_6[63]},
      {stage1_6[27]}
   );
   gpc1_1 gpc205 (
      {stage0_8[54]},
      {stage1_8[25]}
   );
   gpc1_1 gpc206 (
      {stage0_8[55]},
      {stage1_8[26]}
   );
   gpc1_1 gpc207 (
      {stage0_8[56]},
      {stage1_8[27]}
   );
   gpc1_1 gpc208 (
      {stage0_8[57]},
      {stage1_8[28]}
   );
   gpc1_1 gpc209 (
      {stage0_8[58]},
      {stage1_8[29]}
   );
   gpc1_1 gpc210 (
      {stage0_8[59]},
      {stage1_8[30]}
   );
   gpc1_1 gpc211 (
      {stage0_8[60]},
      {stage1_8[31]}
   );
   gpc1_1 gpc212 (
      {stage0_8[61]},
      {stage1_8[32]}
   );
   gpc1_1 gpc213 (
      {stage0_8[62]},
      {stage1_8[33]}
   );
   gpc1_1 gpc214 (
      {stage0_8[63]},
      {stage1_8[34]}
   );
   gpc1_1 gpc215 (
      {stage0_9[60]},
      {stage1_9[24]}
   );
   gpc1_1 gpc216 (
      {stage0_9[61]},
      {stage1_9[25]}
   );
   gpc1_1 gpc217 (
      {stage0_9[62]},
      {stage1_9[26]}
   );
   gpc1_1 gpc218 (
      {stage0_9[63]},
      {stage1_9[27]}
   );
   gpc1_1 gpc219 (
      {stage0_10[60]},
      {stage1_10[25]}
   );
   gpc1_1 gpc220 (
      {stage0_10[61]},
      {stage1_10[26]}
   );
   gpc1_1 gpc221 (
      {stage0_10[62]},
      {stage1_10[27]}
   );
   gpc1_1 gpc222 (
      {stage0_10[63]},
      {stage1_10[28]}
   );
   gpc1_1 gpc223 (
      {stage0_11[61]},
      {stage1_11[26]}
   );
   gpc1_1 gpc224 (
      {stage0_11[62]},
      {stage1_11[27]}
   );
   gpc1_1 gpc225 (
      {stage0_11[63]},
      {stage1_11[28]}
   );
   gpc1_1 gpc226 (
      {stage0_12[41]},
      {stage1_12[21]}
   );
   gpc1_1 gpc227 (
      {stage0_12[42]},
      {stage1_12[22]}
   );
   gpc1_1 gpc228 (
      {stage0_12[43]},
      {stage1_12[23]}
   );
   gpc1_1 gpc229 (
      {stage0_12[44]},
      {stage1_12[24]}
   );
   gpc1_1 gpc230 (
      {stage0_12[45]},
      {stage1_12[25]}
   );
   gpc1_1 gpc231 (
      {stage0_12[46]},
      {stage1_12[26]}
   );
   gpc1_1 gpc232 (
      {stage0_12[47]},
      {stage1_12[27]}
   );
   gpc1_1 gpc233 (
      {stage0_12[48]},
      {stage1_12[28]}
   );
   gpc1_1 gpc234 (
      {stage0_12[49]},
      {stage1_12[29]}
   );
   gpc1_1 gpc235 (
      {stage0_12[50]},
      {stage1_12[30]}
   );
   gpc1_1 gpc236 (
      {stage0_12[51]},
      {stage1_12[31]}
   );
   gpc1_1 gpc237 (
      {stage0_12[52]},
      {stage1_12[32]}
   );
   gpc1_1 gpc238 (
      {stage0_12[53]},
      {stage1_12[33]}
   );
   gpc1_1 gpc239 (
      {stage0_12[54]},
      {stage1_12[34]}
   );
   gpc1_1 gpc240 (
      {stage0_12[55]},
      {stage1_12[35]}
   );
   gpc1_1 gpc241 (
      {stage0_12[56]},
      {stage1_12[36]}
   );
   gpc1_1 gpc242 (
      {stage0_12[57]},
      {stage1_12[37]}
   );
   gpc1_1 gpc243 (
      {stage0_12[58]},
      {stage1_12[38]}
   );
   gpc1_1 gpc244 (
      {stage0_12[59]},
      {stage1_12[39]}
   );
   gpc1_1 gpc245 (
      {stage0_12[60]},
      {stage1_12[40]}
   );
   gpc1_1 gpc246 (
      {stage0_12[61]},
      {stage1_12[41]}
   );
   gpc1_1 gpc247 (
      {stage0_12[62]},
      {stage1_12[42]}
   );
   gpc1_1 gpc248 (
      {stage0_12[63]},
      {stage1_12[43]}
   );
   gpc1_1 gpc249 (
      {stage0_14[43]},
      {stage1_14[24]}
   );
   gpc1_1 gpc250 (
      {stage0_14[44]},
      {stage1_14[25]}
   );
   gpc1_1 gpc251 (
      {stage0_14[45]},
      {stage1_14[26]}
   );
   gpc1_1 gpc252 (
      {stage0_14[46]},
      {stage1_14[27]}
   );
   gpc1_1 gpc253 (
      {stage0_14[47]},
      {stage1_14[28]}
   );
   gpc1_1 gpc254 (
      {stage0_14[48]},
      {stage1_14[29]}
   );
   gpc1_1 gpc255 (
      {stage0_14[49]},
      {stage1_14[30]}
   );
   gpc1_1 gpc256 (
      {stage0_14[50]},
      {stage1_14[31]}
   );
   gpc1_1 gpc257 (
      {stage0_14[51]},
      {stage1_14[32]}
   );
   gpc1_1 gpc258 (
      {stage0_14[52]},
      {stage1_14[33]}
   );
   gpc1_1 gpc259 (
      {stage0_14[53]},
      {stage1_14[34]}
   );
   gpc1_1 gpc260 (
      {stage0_14[54]},
      {stage1_14[35]}
   );
   gpc1_1 gpc261 (
      {stage0_14[55]},
      {stage1_14[36]}
   );
   gpc1_1 gpc262 (
      {stage0_14[56]},
      {stage1_14[37]}
   );
   gpc1_1 gpc263 (
      {stage0_14[57]},
      {stage1_14[38]}
   );
   gpc1_1 gpc264 (
      {stage0_14[58]},
      {stage1_14[39]}
   );
   gpc1_1 gpc265 (
      {stage0_14[59]},
      {stage1_14[40]}
   );
   gpc1_1 gpc266 (
      {stage0_14[60]},
      {stage1_14[41]}
   );
   gpc1_1 gpc267 (
      {stage0_14[61]},
      {stage1_14[42]}
   );
   gpc1_1 gpc268 (
      {stage0_14[62]},
      {stage1_14[43]}
   );
   gpc1_1 gpc269 (
      {stage0_14[63]},
      {stage1_14[44]}
   );
   gpc1_1 gpc270 (
      {stage0_15[52]},
      {stage1_15[20]}
   );
   gpc1_1 gpc271 (
      {stage0_15[53]},
      {stage1_15[21]}
   );
   gpc1_1 gpc272 (
      {stage0_15[54]},
      {stage1_15[22]}
   );
   gpc1_1 gpc273 (
      {stage0_15[55]},
      {stage1_15[23]}
   );
   gpc1_1 gpc274 (
      {stage0_15[56]},
      {stage1_15[24]}
   );
   gpc1_1 gpc275 (
      {stage0_15[57]},
      {stage1_15[25]}
   );
   gpc1_1 gpc276 (
      {stage0_15[58]},
      {stage1_15[26]}
   );
   gpc1_1 gpc277 (
      {stage0_15[59]},
      {stage1_15[27]}
   );
   gpc1_1 gpc278 (
      {stage0_15[60]},
      {stage1_15[28]}
   );
   gpc1_1 gpc279 (
      {stage0_15[61]},
      {stage1_15[29]}
   );
   gpc1_1 gpc280 (
      {stage0_15[62]},
      {stage1_15[30]}
   );
   gpc1_1 gpc281 (
      {stage0_15[63]},
      {stage1_15[31]}
   );
   gpc1_1 gpc282 (
      {stage0_16[62]},
      {stage1_16[19]}
   );
   gpc1_1 gpc283 (
      {stage0_16[63]},
      {stage1_16[20]}
   );
   gpc1_1 gpc284 (
      {stage0_17[57]},
      {stage1_17[28]}
   );
   gpc1_1 gpc285 (
      {stage0_17[58]},
      {stage1_17[29]}
   );
   gpc1_1 gpc286 (
      {stage0_17[59]},
      {stage1_17[30]}
   );
   gpc1_1 gpc287 (
      {stage0_17[60]},
      {stage1_17[31]}
   );
   gpc1_1 gpc288 (
      {stage0_17[61]},
      {stage1_17[32]}
   );
   gpc1_1 gpc289 (
      {stage0_17[62]},
      {stage1_17[33]}
   );
   gpc1_1 gpc290 (
      {stage0_17[63]},
      {stage1_17[34]}
   );
   gpc1_1 gpc291 (
      {stage0_18[42]},
      {stage1_18[21]}
   );
   gpc1_1 gpc292 (
      {stage0_18[43]},
      {stage1_18[22]}
   );
   gpc1_1 gpc293 (
      {stage0_18[44]},
      {stage1_18[23]}
   );
   gpc1_1 gpc294 (
      {stage0_18[45]},
      {stage1_18[24]}
   );
   gpc1_1 gpc295 (
      {stage0_18[46]},
      {stage1_18[25]}
   );
   gpc1_1 gpc296 (
      {stage0_18[47]},
      {stage1_18[26]}
   );
   gpc1_1 gpc297 (
      {stage0_18[48]},
      {stage1_18[27]}
   );
   gpc1_1 gpc298 (
      {stage0_18[49]},
      {stage1_18[28]}
   );
   gpc1_1 gpc299 (
      {stage0_18[50]},
      {stage1_18[29]}
   );
   gpc1_1 gpc300 (
      {stage0_18[51]},
      {stage1_18[30]}
   );
   gpc1_1 gpc301 (
      {stage0_18[52]},
      {stage1_18[31]}
   );
   gpc1_1 gpc302 (
      {stage0_18[53]},
      {stage1_18[32]}
   );
   gpc1_1 gpc303 (
      {stage0_18[54]},
      {stage1_18[33]}
   );
   gpc1_1 gpc304 (
      {stage0_18[55]},
      {stage1_18[34]}
   );
   gpc1_1 gpc305 (
      {stage0_18[56]},
      {stage1_18[35]}
   );
   gpc1_1 gpc306 (
      {stage0_18[57]},
      {stage1_18[36]}
   );
   gpc1_1 gpc307 (
      {stage0_18[58]},
      {stage1_18[37]}
   );
   gpc1_1 gpc308 (
      {stage0_18[59]},
      {stage1_18[38]}
   );
   gpc1_1 gpc309 (
      {stage0_18[60]},
      {stage1_18[39]}
   );
   gpc1_1 gpc310 (
      {stage0_18[61]},
      {stage1_18[40]}
   );
   gpc1_1 gpc311 (
      {stage0_18[62]},
      {stage1_18[41]}
   );
   gpc1_1 gpc312 (
      {stage0_18[63]},
      {stage1_18[42]}
   );
   gpc1_1 gpc313 (
      {stage0_20[53]},
      {stage1_20[27]}
   );
   gpc1_1 gpc314 (
      {stage0_20[54]},
      {stage1_20[28]}
   );
   gpc1_1 gpc315 (
      {stage0_20[55]},
      {stage1_20[29]}
   );
   gpc1_1 gpc316 (
      {stage0_20[56]},
      {stage1_20[30]}
   );
   gpc1_1 gpc317 (
      {stage0_20[57]},
      {stage1_20[31]}
   );
   gpc1_1 gpc318 (
      {stage0_20[58]},
      {stage1_20[32]}
   );
   gpc1_1 gpc319 (
      {stage0_20[59]},
      {stage1_20[33]}
   );
   gpc1_1 gpc320 (
      {stage0_20[60]},
      {stage1_20[34]}
   );
   gpc1_1 gpc321 (
      {stage0_20[61]},
      {stage1_20[35]}
   );
   gpc1_1 gpc322 (
      {stage0_20[62]},
      {stage1_20[36]}
   );
   gpc1_1 gpc323 (
      {stage0_20[63]},
      {stage1_20[37]}
   );
   gpc1_1 gpc324 (
      {stage0_23[37]},
      {stage1_23[21]}
   );
   gpc1_1 gpc325 (
      {stage0_23[38]},
      {stage1_23[22]}
   );
   gpc1_1 gpc326 (
      {stage0_23[39]},
      {stage1_23[23]}
   );
   gpc1_1 gpc327 (
      {stage0_23[40]},
      {stage1_23[24]}
   );
   gpc1_1 gpc328 (
      {stage0_23[41]},
      {stage1_23[25]}
   );
   gpc1_1 gpc329 (
      {stage0_23[42]},
      {stage1_23[26]}
   );
   gpc1_1 gpc330 (
      {stage0_23[43]},
      {stage1_23[27]}
   );
   gpc1_1 gpc331 (
      {stage0_23[44]},
      {stage1_23[28]}
   );
   gpc1_1 gpc332 (
      {stage0_23[45]},
      {stage1_23[29]}
   );
   gpc1_1 gpc333 (
      {stage0_23[46]},
      {stage1_23[30]}
   );
   gpc1_1 gpc334 (
      {stage0_23[47]},
      {stage1_23[31]}
   );
   gpc1_1 gpc335 (
      {stage0_23[48]},
      {stage1_23[32]}
   );
   gpc1_1 gpc336 (
      {stage0_23[49]},
      {stage1_23[33]}
   );
   gpc1_1 gpc337 (
      {stage0_23[50]},
      {stage1_23[34]}
   );
   gpc1_1 gpc338 (
      {stage0_23[51]},
      {stage1_23[35]}
   );
   gpc1_1 gpc339 (
      {stage0_23[52]},
      {stage1_23[36]}
   );
   gpc1_1 gpc340 (
      {stage0_23[53]},
      {stage1_23[37]}
   );
   gpc1_1 gpc341 (
      {stage0_23[54]},
      {stage1_23[38]}
   );
   gpc1_1 gpc342 (
      {stage0_23[55]},
      {stage1_23[39]}
   );
   gpc1_1 gpc343 (
      {stage0_23[56]},
      {stage1_23[40]}
   );
   gpc1_1 gpc344 (
      {stage0_23[57]},
      {stage1_23[41]}
   );
   gpc1_1 gpc345 (
      {stage0_23[58]},
      {stage1_23[42]}
   );
   gpc1_1 gpc346 (
      {stage0_23[59]},
      {stage1_23[43]}
   );
   gpc1_1 gpc347 (
      {stage0_23[60]},
      {stage1_23[44]}
   );
   gpc1_1 gpc348 (
      {stage0_23[61]},
      {stage1_23[45]}
   );
   gpc1_1 gpc349 (
      {stage0_23[62]},
      {stage1_23[46]}
   );
   gpc1_1 gpc350 (
      {stage0_23[63]},
      {stage1_23[47]}
   );
   gpc1_1 gpc351 (
      {stage0_24[43]},
      {stage1_24[23]}
   );
   gpc1_1 gpc352 (
      {stage0_24[44]},
      {stage1_24[24]}
   );
   gpc1_1 gpc353 (
      {stage0_24[45]},
      {stage1_24[25]}
   );
   gpc1_1 gpc354 (
      {stage0_24[46]},
      {stage1_24[26]}
   );
   gpc1_1 gpc355 (
      {stage0_24[47]},
      {stage1_24[27]}
   );
   gpc1_1 gpc356 (
      {stage0_24[48]},
      {stage1_24[28]}
   );
   gpc1_1 gpc357 (
      {stage0_24[49]},
      {stage1_24[29]}
   );
   gpc1_1 gpc358 (
      {stage0_24[50]},
      {stage1_24[30]}
   );
   gpc1_1 gpc359 (
      {stage0_24[51]},
      {stage1_24[31]}
   );
   gpc1_1 gpc360 (
      {stage0_24[52]},
      {stage1_24[32]}
   );
   gpc1_1 gpc361 (
      {stage0_24[53]},
      {stage1_24[33]}
   );
   gpc1_1 gpc362 (
      {stage0_24[54]},
      {stage1_24[34]}
   );
   gpc1_1 gpc363 (
      {stage0_24[55]},
      {stage1_24[35]}
   );
   gpc1_1 gpc364 (
      {stage0_24[56]},
      {stage1_24[36]}
   );
   gpc1_1 gpc365 (
      {stage0_24[57]},
      {stage1_24[37]}
   );
   gpc1_1 gpc366 (
      {stage0_24[58]},
      {stage1_24[38]}
   );
   gpc1_1 gpc367 (
      {stage0_24[59]},
      {stage1_24[39]}
   );
   gpc1_1 gpc368 (
      {stage0_24[60]},
      {stage1_24[40]}
   );
   gpc1_1 gpc369 (
      {stage0_24[61]},
      {stage1_24[41]}
   );
   gpc1_1 gpc370 (
      {stage0_24[62]},
      {stage1_24[42]}
   );
   gpc1_1 gpc371 (
      {stage0_24[63]},
      {stage1_24[43]}
   );
   gpc1_1 gpc372 (
      {stage0_26[57]},
      {stage1_26[21]}
   );
   gpc1_1 gpc373 (
      {stage0_26[58]},
      {stage1_26[22]}
   );
   gpc1_1 gpc374 (
      {stage0_26[59]},
      {stage1_26[23]}
   );
   gpc1_1 gpc375 (
      {stage0_26[60]},
      {stage1_26[24]}
   );
   gpc1_1 gpc376 (
      {stage0_26[61]},
      {stage1_26[25]}
   );
   gpc1_1 gpc377 (
      {stage0_26[62]},
      {stage1_26[26]}
   );
   gpc1_1 gpc378 (
      {stage0_26[63]},
      {stage1_26[27]}
   );
   gpc1_1 gpc379 (
      {stage0_27[62]},
      {stage1_27[20]}
   );
   gpc1_1 gpc380 (
      {stage0_27[63]},
      {stage1_27[21]}
   );
   gpc1_1 gpc381 (
      {stage0_29[56]},
      {stage1_29[30]}
   );
   gpc1_1 gpc382 (
      {stage0_29[57]},
      {stage1_29[31]}
   );
   gpc1_1 gpc383 (
      {stage0_29[58]},
      {stage1_29[32]}
   );
   gpc1_1 gpc384 (
      {stage0_29[59]},
      {stage1_29[33]}
   );
   gpc1_1 gpc385 (
      {stage0_29[60]},
      {stage1_29[34]}
   );
   gpc1_1 gpc386 (
      {stage0_29[61]},
      {stage1_29[35]}
   );
   gpc1_1 gpc387 (
      {stage0_29[62]},
      {stage1_29[36]}
   );
   gpc1_1 gpc388 (
      {stage0_29[63]},
      {stage1_29[37]}
   );
   gpc1_1 gpc389 (
      {stage0_30[54]},
      {stage1_30[20]}
   );
   gpc1_1 gpc390 (
      {stage0_30[55]},
      {stage1_30[21]}
   );
   gpc1_1 gpc391 (
      {stage0_30[56]},
      {stage1_30[22]}
   );
   gpc1_1 gpc392 (
      {stage0_30[57]},
      {stage1_30[23]}
   );
   gpc1_1 gpc393 (
      {stage0_30[58]},
      {stage1_30[24]}
   );
   gpc1_1 gpc394 (
      {stage0_30[59]},
      {stage1_30[25]}
   );
   gpc1_1 gpc395 (
      {stage0_30[60]},
      {stage1_30[26]}
   );
   gpc1_1 gpc396 (
      {stage0_30[61]},
      {stage1_30[27]}
   );
   gpc1_1 gpc397 (
      {stage0_30[62]},
      {stage1_30[28]}
   );
   gpc1_1 gpc398 (
      {stage0_30[63]},
      {stage1_30[29]}
   );
   gpc1_1 gpc399 (
      {stage0_31[54]},
      {stage1_31[18]}
   );
   gpc1_1 gpc400 (
      {stage0_31[55]},
      {stage1_31[19]}
   );
   gpc1_1 gpc401 (
      {stage0_31[56]},
      {stage1_31[20]}
   );
   gpc1_1 gpc402 (
      {stage0_31[57]},
      {stage1_31[21]}
   );
   gpc1_1 gpc403 (
      {stage0_31[58]},
      {stage1_31[22]}
   );
   gpc1_1 gpc404 (
      {stage0_31[59]},
      {stage1_31[23]}
   );
   gpc1_1 gpc405 (
      {stage0_31[60]},
      {stage1_31[24]}
   );
   gpc1_1 gpc406 (
      {stage0_31[61]},
      {stage1_31[25]}
   );
   gpc1_1 gpc407 (
      {stage0_31[62]},
      {stage1_31[26]}
   );
   gpc1_1 gpc408 (
      {stage0_31[63]},
      {stage1_31[27]}
   );
   gpc606_5 gpc409 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc410 (
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage2_5[0],stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1]}
   );
   gpc606_5 gpc411 (
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage2_5[1],stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2]}
   );
   gpc606_5 gpc412 (
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage2_5[2],stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3]}
   );
   gpc606_5 gpc413 (
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[0],stage2_6[0],stage2_5[3],stage2_4[4]}
   );
   gpc606_5 gpc414 (
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[1],stage2_6[1],stage2_5[4],stage2_4[5]}
   );
   gpc606_5 gpc415 (
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[2],stage2_6[2],stage2_5[5],stage2_4[6]}
   );
   gpc606_5 gpc416 (
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[3],stage2_6[3],stage2_5[6],stage2_4[7]}
   );
   gpc606_5 gpc417 (
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[4],stage2_7[4],stage2_6[4],stage2_5[7]}
   );
   gpc606_5 gpc418 (
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[5],stage2_7[5],stage2_6[5],stage2_5[8]}
   );
   gpc606_5 gpc419 (
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[6],stage2_7[6],stage2_6[6],stage2_5[9]}
   );
   gpc615_5 gpc420 (
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22]},
      {stage1_8[0]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[0],stage2_9[3],stage2_8[7],stage2_7[7]}
   );
   gpc606_5 gpc421 (
      {stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5], stage1_8[6]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[1],stage2_10[1],stage2_9[4],stage2_8[8]}
   );
   gpc606_5 gpc422 (
      {stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11], stage1_8[12]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[2],stage2_10[2],stage2_9[5],stage2_8[9]}
   );
   gpc606_5 gpc423 (
      {stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17], stage1_8[18]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[3],stage2_10[3],stage2_9[6],stage2_8[10]}
   );
   gpc606_5 gpc424 (
      {stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23], stage1_8[24]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[4],stage2_10[4],stage2_9[7],stage2_8[11]}
   );
   gpc606_5 gpc425 (
      {stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29], stage1_8[30]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], 1'b0},
      {stage2_12[4],stage2_11[5],stage2_10[5],stage2_9[8],stage2_8[12]}
   );
   gpc606_5 gpc426 (
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[5],stage2_11[6],stage2_10[6],stage2_9[9]}
   );
   gpc606_5 gpc427 (
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[6],stage2_11[7],stage2_10[7],stage2_9[10]}
   );
   gpc606_5 gpc428 (
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[7],stage2_11[8],stage2_10[8],stage2_9[11]}
   );
   gpc615_5 gpc429 (
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22]},
      {stage1_12[0]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[0],stage2_13[3],stage2_12[8],stage2_11[9]}
   );
   gpc615_5 gpc430 (
      {stage1_11[23], stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27]},
      {stage1_12[1]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[1],stage2_13[4],stage2_12[9],stage2_11[10]}
   );
   gpc606_5 gpc431 (
      {stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5], stage1_12[6], stage1_12[7]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[2],stage2_14[2],stage2_13[5],stage2_12[10]}
   );
   gpc606_5 gpc432 (
      {stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11], stage1_12[12], stage1_12[13]},
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage2_16[1],stage2_15[3],stage2_14[3],stage2_13[6],stage2_12[11]}
   );
   gpc606_5 gpc433 (
      {stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17], stage1_12[18], stage1_12[19]},
      {stage1_14[12], stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17]},
      {stage2_16[2],stage2_15[4],stage2_14[4],stage2_13[7],stage2_12[12]}
   );
   gpc606_5 gpc434 (
      {stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23], stage1_12[24], stage1_12[25]},
      {stage1_14[18], stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23]},
      {stage2_16[3],stage2_15[5],stage2_14[5],stage2_13[8],stage2_12[13]}
   );
   gpc606_5 gpc435 (
      {stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29], stage1_12[30], stage1_12[31]},
      {stage1_14[24], stage1_14[25], stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29]},
      {stage2_16[4],stage2_15[6],stage2_14[6],stage2_13[9],stage2_12[14]}
   );
   gpc606_5 gpc436 (
      {stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35], stage1_12[36], stage1_12[37]},
      {stage1_14[30], stage1_14[31], stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35]},
      {stage2_16[5],stage2_15[7],stage2_14[7],stage2_13[10],stage2_12[15]}
   );
   gpc606_5 gpc437 (
      {stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41], stage1_12[42], stage1_12[43]},
      {stage1_14[36], stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41]},
      {stage2_16[6],stage2_15[8],stage2_14[8],stage2_13[11],stage2_12[16]}
   );
   gpc606_5 gpc438 (
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[7],stage2_15[9],stage2_14[9],stage2_13[12]}
   );
   gpc615_5 gpc439 (
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10]},
      {stage1_16[0]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[0],stage2_17[1],stage2_16[8],stage2_15[10]}
   );
   gpc615_5 gpc440 (
      {stage1_15[11], stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15]},
      {stage1_16[1]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[1],stage2_17[2],stage2_16[9],stage2_15[11]}
   );
   gpc615_5 gpc441 (
      {stage1_15[16], stage1_15[17], stage1_15[18], stage1_15[19], stage1_15[20]},
      {stage1_16[2]},
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage2_19[2],stage2_18[2],stage2_17[3],stage2_16[10],stage2_15[12]}
   );
   gpc606_5 gpc442 (
      {stage1_16[3], stage1_16[4], stage1_16[5], stage1_16[6], stage1_16[7], stage1_16[8]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[3],stage2_18[3],stage2_17[4],stage2_16[11]}
   );
   gpc606_5 gpc443 (
      {stage1_16[9], stage1_16[10], stage1_16[11], stage1_16[12], stage1_16[13], stage1_16[14]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[4],stage2_18[4],stage2_17[5],stage2_16[12]}
   );
   gpc606_5 gpc444 (
      {stage1_16[15], stage1_16[16], stage1_16[17], stage1_16[18], stage1_16[19], stage1_16[20]},
      {stage1_18[12], stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17]},
      {stage2_20[2],stage2_19[5],stage2_18[5],stage2_17[6],stage2_16[13]}
   );
   gpc606_5 gpc445 (
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[3],stage2_19[6],stage2_18[6],stage2_17[7]}
   );
   gpc606_5 gpc446 (
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[4],stage2_19[7],stage2_18[7],stage2_17[8]}
   );
   gpc615_5 gpc447 (
      {stage1_18[18], stage1_18[19], stage1_18[20], stage1_18[21], stage1_18[22]},
      {stage1_19[12]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[2],stage2_20[5],stage2_19[8],stage2_18[8]}
   );
   gpc615_5 gpc448 (
      {stage1_18[23], stage1_18[24], stage1_18[25], stage1_18[26], stage1_18[27]},
      {stage1_19[13]},
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage2_22[1],stage2_21[3],stage2_20[6],stage2_19[9],stage2_18[9]}
   );
   gpc615_5 gpc449 (
      {stage1_18[28], stage1_18[29], stage1_18[30], stage1_18[31], stage1_18[32]},
      {stage1_19[14]},
      {stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15], stage1_20[16], stage1_20[17]},
      {stage2_22[2],stage2_21[4],stage2_20[7],stage2_19[10],stage2_18[10]}
   );
   gpc615_5 gpc450 (
      {stage1_20[18], stage1_20[19], stage1_20[20], stage1_20[21], stage1_20[22]},
      {stage1_21[0]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[0],stage2_22[3],stage2_21[5],stage2_20[8]}
   );
   gpc606_5 gpc451 (
      {stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5], stage1_21[6]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[1],stage2_23[1],stage2_22[4],stage2_21[6]}
   );
   gpc606_5 gpc452 (
      {stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11], stage1_21[12]},
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage2_25[1],stage2_24[2],stage2_23[2],stage2_22[5],stage2_21[7]}
   );
   gpc606_5 gpc453 (
      {stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17], stage1_21[18]},
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage2_25[2],stage2_24[3],stage2_23[3],stage2_22[6],stage2_21[8]}
   );
   gpc606_5 gpc454 (
      {stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23], stage1_21[24]},
      {stage1_23[18], stage1_23[19], stage1_23[20], stage1_23[21], stage1_23[22], stage1_23[23]},
      {stage2_25[3],stage2_24[4],stage2_23[4],stage2_22[7],stage2_21[9]}
   );
   gpc615_5 gpc455 (
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10]},
      {stage1_23[24]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5]},
      {stage2_26[0],stage2_25[4],stage2_24[5],stage2_23[5],stage2_22[8]}
   );
   gpc615_5 gpc456 (
      {stage1_23[25], stage1_23[26], stage1_23[27], stage1_23[28], stage1_23[29]},
      {stage1_24[6]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[1],stage2_25[5],stage2_24[6],stage2_23[6]}
   );
   gpc615_5 gpc457 (
      {stage1_23[30], stage1_23[31], stage1_23[32], stage1_23[33], stage1_23[34]},
      {stage1_24[7]},
      {stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11]},
      {stage2_27[1],stage2_26[2],stage2_25[6],stage2_24[7],stage2_23[7]}
   );
   gpc615_5 gpc458 (
      {stage1_23[35], stage1_23[36], stage1_23[37], stage1_23[38], stage1_23[39]},
      {stage1_24[8]},
      {stage1_25[12], stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {stage2_27[2],stage2_26[3],stage2_25[7],stage2_24[8],stage2_23[8]}
   );
   gpc606_5 gpc459 (
      {stage1_24[9], stage1_24[10], stage1_24[11], stage1_24[12], stage1_24[13], stage1_24[14]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[3],stage2_26[4],stage2_25[8],stage2_24[9]}
   );
   gpc606_5 gpc460 (
      {stage1_24[15], stage1_24[16], stage1_24[17], stage1_24[18], stage1_24[19], stage1_24[20]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[4],stage2_26[5],stage2_25[9],stage2_24[10]}
   );
   gpc606_5 gpc461 (
      {stage1_24[21], stage1_24[22], stage1_24[23], stage1_24[24], stage1_24[25], stage1_24[26]},
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17]},
      {stage2_28[2],stage2_27[5],stage2_26[6],stage2_25[10],stage2_24[11]}
   );
   gpc606_5 gpc462 (
      {stage1_24[27], stage1_24[28], stage1_24[29], stage1_24[30], stage1_24[31], stage1_24[32]},
      {stage1_26[18], stage1_26[19], stage1_26[20], stage1_26[21], stage1_26[22], stage1_26[23]},
      {stage2_28[3],stage2_27[6],stage2_26[7],stage2_25[11],stage2_24[12]}
   );
   gpc615_5 gpc463 (
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4]},
      {stage1_28[0]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[0],stage2_29[0],stage2_28[4],stage2_27[7]}
   );
   gpc615_5 gpc464 (
      {stage1_27[5], stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9]},
      {stage1_28[1]},
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage2_31[1],stage2_30[1],stage2_29[1],stage2_28[5],stage2_27[8]}
   );
   gpc615_5 gpc465 (
      {stage1_27[10], stage1_27[11], stage1_27[12], stage1_27[13], stage1_27[14]},
      {stage1_28[2]},
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17]},
      {stage2_31[2],stage2_30[2],stage2_29[2],stage2_28[6],stage2_27[9]}
   );
   gpc2135_5 gpc466 (
      {stage1_28[3], stage1_28[4], stage1_28[5], stage1_28[6], stage1_28[7]},
      {stage1_29[18], stage1_29[19], stage1_29[20]},
      {stage1_30[0]},
      {stage1_31[0], stage1_31[1]},
      {stage2_32[0],stage2_31[3],stage2_30[3],stage2_29[3],stage2_28[7]}
   );
   gpc606_5 gpc467 (
      {stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11], stage1_28[12], stage1_28[13]},
      {stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5], stage1_30[6]},
      {stage2_32[1],stage2_31[4],stage2_30[4],stage2_29[4],stage2_28[8]}
   );
   gpc606_5 gpc468 (
      {stage1_28[14], stage1_28[15], stage1_28[16], stage1_28[17], stage1_28[18], stage1_28[19]},
      {stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11], stage1_30[12]},
      {stage2_32[2],stage2_31[5],stage2_30[5],stage2_29[5],stage2_28[9]}
   );
   gpc606_5 gpc469 (
      {stage1_29[21], stage1_29[22], stage1_29[23], stage1_29[24], stage1_29[25], stage1_29[26]},
      {stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5], stage1_31[6], stage1_31[7]},
      {stage2_33[0],stage2_32[3],stage2_31[6],stage2_30[6],stage2_29[6]}
   );
   gpc615_5 gpc470 (
      {stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage1_31[8]},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[1],stage2_32[4],stage2_31[7],stage2_30[7]}
   );
   gpc615_5 gpc471 (
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22]},
      {stage1_31[9]},
      {stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11]},
      {stage2_34[1],stage2_33[2],stage2_32[5],stage2_31[8],stage2_30[8]}
   );
   gpc615_5 gpc472 (
      {stage1_30[23], stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27]},
      {stage1_31[10]},
      {stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16], stage1_32[17]},
      {stage2_34[2],stage2_33[3],stage2_32[6],stage2_31[9],stage2_30[9]}
   );
   gpc606_5 gpc473 (
      {stage1_31[11], stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15], stage1_31[16]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5]},
      {stage2_35[0],stage2_34[3],stage2_33[4],stage2_32[7],stage2_31[10]}
   );
   gpc1_1 gpc474 (
      {stage1_0[6]},
      {stage2_0[1]}
   );
   gpc1_1 gpc475 (
      {stage1_0[7]},
      {stage2_0[2]}
   );
   gpc1_1 gpc476 (
      {stage1_0[8]},
      {stage2_0[3]}
   );
   gpc1_1 gpc477 (
      {stage1_0[9]},
      {stage2_0[4]}
   );
   gpc1_1 gpc478 (
      {stage1_0[10]},
      {stage2_0[5]}
   );
   gpc1_1 gpc479 (
      {stage1_0[11]},
      {stage2_0[6]}
   );
   gpc1_1 gpc480 (
      {stage1_0[12]},
      {stage2_0[7]}
   );
   gpc1_1 gpc481 (
      {stage1_0[13]},
      {stage2_0[8]}
   );
   gpc1_1 gpc482 (
      {stage1_0[14]},
      {stage2_0[9]}
   );
   gpc1_1 gpc483 (
      {stage1_0[15]},
      {stage2_0[10]}
   );
   gpc1_1 gpc484 (
      {stage1_0[16]},
      {stage2_0[11]}
   );
   gpc1_1 gpc485 (
      {stage1_0[17]},
      {stage2_0[12]}
   );
   gpc1_1 gpc486 (
      {stage1_0[18]},
      {stage2_0[13]}
   );
   gpc1_1 gpc487 (
      {stage1_0[19]},
      {stage2_0[14]}
   );
   gpc1_1 gpc488 (
      {stage1_0[20]},
      {stage2_0[15]}
   );
   gpc1_1 gpc489 (
      {stage1_0[21]},
      {stage2_0[16]}
   );
   gpc1_1 gpc490 (
      {stage1_0[22]},
      {stage2_0[17]}
   );
   gpc1_1 gpc491 (
      {stage1_0[23]},
      {stage2_0[18]}
   );
   gpc1_1 gpc492 (
      {stage1_1[18]},
      {stage2_1[4]}
   );
   gpc1_1 gpc493 (
      {stage1_1[19]},
      {stage2_1[5]}
   );
   gpc1_1 gpc494 (
      {stage1_2[6]},
      {stage2_2[4]}
   );
   gpc1_1 gpc495 (
      {stage1_2[7]},
      {stage2_2[5]}
   );
   gpc1_1 gpc496 (
      {stage1_2[8]},
      {stage2_2[6]}
   );
   gpc1_1 gpc497 (
      {stage1_2[9]},
      {stage2_2[7]}
   );
   gpc1_1 gpc498 (
      {stage1_2[10]},
      {stage2_2[8]}
   );
   gpc1_1 gpc499 (
      {stage1_2[11]},
      {stage2_2[9]}
   );
   gpc1_1 gpc500 (
      {stage1_2[12]},
      {stage2_2[10]}
   );
   gpc1_1 gpc501 (
      {stage1_2[13]},
      {stage2_2[11]}
   );
   gpc1_1 gpc502 (
      {stage1_2[14]},
      {stage2_2[12]}
   );
   gpc1_1 gpc503 (
      {stage1_2[15]},
      {stage2_2[13]}
   );
   gpc1_1 gpc504 (
      {stage1_2[16]},
      {stage2_2[14]}
   );
   gpc1_1 gpc505 (
      {stage1_2[17]},
      {stage2_2[15]}
   );
   gpc1_1 gpc506 (
      {stage1_2[18]},
      {stage2_2[16]}
   );
   gpc1_1 gpc507 (
      {stage1_2[19]},
      {stage2_2[17]}
   );
   gpc1_1 gpc508 (
      {stage1_2[20]},
      {stage2_2[18]}
   );
   gpc1_1 gpc509 (
      {stage1_2[21]},
      {stage2_2[19]}
   );
   gpc1_1 gpc510 (
      {stage1_2[22]},
      {stage2_2[20]}
   );
   gpc1_1 gpc511 (
      {stage1_2[23]},
      {stage2_2[21]}
   );
   gpc1_1 gpc512 (
      {stage1_3[18]},
      {stage2_3[4]}
   );
   gpc1_1 gpc513 (
      {stage1_3[19]},
      {stage2_3[5]}
   );
   gpc1_1 gpc514 (
      {stage1_3[20]},
      {stage2_3[6]}
   );
   gpc1_1 gpc515 (
      {stage1_3[21]},
      {stage2_3[7]}
   );
   gpc1_1 gpc516 (
      {stage1_3[22]},
      {stage2_3[8]}
   );
   gpc1_1 gpc517 (
      {stage1_3[23]},
      {stage2_3[9]}
   );
   gpc1_1 gpc518 (
      {stage1_3[24]},
      {stage2_3[10]}
   );
   gpc1_1 gpc519 (
      {stage1_3[25]},
      {stage2_3[11]}
   );
   gpc1_1 gpc520 (
      {stage1_3[26]},
      {stage2_3[12]}
   );
   gpc1_1 gpc521 (
      {stage1_3[27]},
      {stage2_3[13]}
   );
   gpc1_1 gpc522 (
      {stage1_3[28]},
      {stage2_3[14]}
   );
   gpc1_1 gpc523 (
      {stage1_3[29]},
      {stage2_3[15]}
   );
   gpc1_1 gpc524 (
      {stage1_3[30]},
      {stage2_3[16]}
   );
   gpc1_1 gpc525 (
      {stage1_3[31]},
      {stage2_3[17]}
   );
   gpc1_1 gpc526 (
      {stage1_4[24]},
      {stage2_4[8]}
   );
   gpc1_1 gpc527 (
      {stage1_4[25]},
      {stage2_4[9]}
   );
   gpc1_1 gpc528 (
      {stage1_4[26]},
      {stage2_4[10]}
   );
   gpc1_1 gpc529 (
      {stage1_4[27]},
      {stage2_4[11]}
   );
   gpc1_1 gpc530 (
      {stage1_4[28]},
      {stage2_4[12]}
   );
   gpc1_1 gpc531 (
      {stage1_4[29]},
      {stage2_4[13]}
   );
   gpc1_1 gpc532 (
      {stage1_4[30]},
      {stage2_4[14]}
   );
   gpc1_1 gpc533 (
      {stage1_4[31]},
      {stage2_4[15]}
   );
   gpc1_1 gpc534 (
      {stage1_4[32]},
      {stage2_4[16]}
   );
   gpc1_1 gpc535 (
      {stage1_4[33]},
      {stage2_4[17]}
   );
   gpc1_1 gpc536 (
      {stage1_4[34]},
      {stage2_4[18]}
   );
   gpc1_1 gpc537 (
      {stage1_5[18]},
      {stage2_5[10]}
   );
   gpc1_1 gpc538 (
      {stage1_5[19]},
      {stage2_5[11]}
   );
   gpc1_1 gpc539 (
      {stage1_5[20]},
      {stage2_5[12]}
   );
   gpc1_1 gpc540 (
      {stage1_5[21]},
      {stage2_5[13]}
   );
   gpc1_1 gpc541 (
      {stage1_5[22]},
      {stage2_5[14]}
   );
   gpc1_1 gpc542 (
      {stage1_5[23]},
      {stage2_5[15]}
   );
   gpc1_1 gpc543 (
      {stage1_5[24]},
      {stage2_5[16]}
   );
   gpc1_1 gpc544 (
      {stage1_5[25]},
      {stage2_5[17]}
   );
   gpc1_1 gpc545 (
      {stage1_5[26]},
      {stage2_5[18]}
   );
   gpc1_1 gpc546 (
      {stage1_5[27]},
      {stage2_5[19]}
   );
   gpc1_1 gpc547 (
      {stage1_5[28]},
      {stage2_5[20]}
   );
   gpc1_1 gpc548 (
      {stage1_5[29]},
      {stage2_5[21]}
   );
   gpc1_1 gpc549 (
      {stage1_5[30]},
      {stage2_5[22]}
   );
   gpc1_1 gpc550 (
      {stage1_5[31]},
      {stage2_5[23]}
   );
   gpc1_1 gpc551 (
      {stage1_5[32]},
      {stage2_5[24]}
   );
   gpc1_1 gpc552 (
      {stage1_5[33]},
      {stage2_5[25]}
   );
   gpc1_1 gpc553 (
      {stage1_5[34]},
      {stage2_5[26]}
   );
   gpc1_1 gpc554 (
      {stage1_6[24]},
      {stage2_6[7]}
   );
   gpc1_1 gpc555 (
      {stage1_6[25]},
      {stage2_6[8]}
   );
   gpc1_1 gpc556 (
      {stage1_6[26]},
      {stage2_6[9]}
   );
   gpc1_1 gpc557 (
      {stage1_6[27]},
      {stage2_6[10]}
   );
   gpc1_1 gpc558 (
      {stage1_7[23]},
      {stage2_7[8]}
   );
   gpc1_1 gpc559 (
      {stage1_8[31]},
      {stage2_8[13]}
   );
   gpc1_1 gpc560 (
      {stage1_8[32]},
      {stage2_8[14]}
   );
   gpc1_1 gpc561 (
      {stage1_8[33]},
      {stage2_8[15]}
   );
   gpc1_1 gpc562 (
      {stage1_8[34]},
      {stage2_8[16]}
   );
   gpc1_1 gpc563 (
      {stage1_9[24]},
      {stage2_9[12]}
   );
   gpc1_1 gpc564 (
      {stage1_9[25]},
      {stage2_9[13]}
   );
   gpc1_1 gpc565 (
      {stage1_9[26]},
      {stage2_9[14]}
   );
   gpc1_1 gpc566 (
      {stage1_9[27]},
      {stage2_9[15]}
   );
   gpc1_1 gpc567 (
      {stage1_11[28]},
      {stage2_11[11]}
   );
   gpc1_1 gpc568 (
      {stage1_13[18]},
      {stage2_13[13]}
   );
   gpc1_1 gpc569 (
      {stage1_13[19]},
      {stage2_13[14]}
   );
   gpc1_1 gpc570 (
      {stage1_13[20]},
      {stage2_13[15]}
   );
   gpc1_1 gpc571 (
      {stage1_13[21]},
      {stage2_13[16]}
   );
   gpc1_1 gpc572 (
      {stage1_13[22]},
      {stage2_13[17]}
   );
   gpc1_1 gpc573 (
      {stage1_14[42]},
      {stage2_14[10]}
   );
   gpc1_1 gpc574 (
      {stage1_14[43]},
      {stage2_14[11]}
   );
   gpc1_1 gpc575 (
      {stage1_14[44]},
      {stage2_14[12]}
   );
   gpc1_1 gpc576 (
      {stage1_15[21]},
      {stage2_15[13]}
   );
   gpc1_1 gpc577 (
      {stage1_15[22]},
      {stage2_15[14]}
   );
   gpc1_1 gpc578 (
      {stage1_15[23]},
      {stage2_15[15]}
   );
   gpc1_1 gpc579 (
      {stage1_15[24]},
      {stage2_15[16]}
   );
   gpc1_1 gpc580 (
      {stage1_15[25]},
      {stage2_15[17]}
   );
   gpc1_1 gpc581 (
      {stage1_15[26]},
      {stage2_15[18]}
   );
   gpc1_1 gpc582 (
      {stage1_15[27]},
      {stage2_15[19]}
   );
   gpc1_1 gpc583 (
      {stage1_15[28]},
      {stage2_15[20]}
   );
   gpc1_1 gpc584 (
      {stage1_15[29]},
      {stage2_15[21]}
   );
   gpc1_1 gpc585 (
      {stage1_15[30]},
      {stage2_15[22]}
   );
   gpc1_1 gpc586 (
      {stage1_15[31]},
      {stage2_15[23]}
   );
   gpc1_1 gpc587 (
      {stage1_17[30]},
      {stage2_17[9]}
   );
   gpc1_1 gpc588 (
      {stage1_17[31]},
      {stage2_17[10]}
   );
   gpc1_1 gpc589 (
      {stage1_17[32]},
      {stage2_17[11]}
   );
   gpc1_1 gpc590 (
      {stage1_17[33]},
      {stage2_17[12]}
   );
   gpc1_1 gpc591 (
      {stage1_17[34]},
      {stage2_17[13]}
   );
   gpc1_1 gpc592 (
      {stage1_18[33]},
      {stage2_18[11]}
   );
   gpc1_1 gpc593 (
      {stage1_18[34]},
      {stage2_18[12]}
   );
   gpc1_1 gpc594 (
      {stage1_18[35]},
      {stage2_18[13]}
   );
   gpc1_1 gpc595 (
      {stage1_18[36]},
      {stage2_18[14]}
   );
   gpc1_1 gpc596 (
      {stage1_18[37]},
      {stage2_18[15]}
   );
   gpc1_1 gpc597 (
      {stage1_18[38]},
      {stage2_18[16]}
   );
   gpc1_1 gpc598 (
      {stage1_18[39]},
      {stage2_18[17]}
   );
   gpc1_1 gpc599 (
      {stage1_18[40]},
      {stage2_18[18]}
   );
   gpc1_1 gpc600 (
      {stage1_18[41]},
      {stage2_18[19]}
   );
   gpc1_1 gpc601 (
      {stage1_18[42]},
      {stage2_18[20]}
   );
   gpc1_1 gpc602 (
      {stage1_19[15]},
      {stage2_19[11]}
   );
   gpc1_1 gpc603 (
      {stage1_19[16]},
      {stage2_19[12]}
   );
   gpc1_1 gpc604 (
      {stage1_19[17]},
      {stage2_19[13]}
   );
   gpc1_1 gpc605 (
      {stage1_19[18]},
      {stage2_19[14]}
   );
   gpc1_1 gpc606 (
      {stage1_19[19]},
      {stage2_19[15]}
   );
   gpc1_1 gpc607 (
      {stage1_20[23]},
      {stage2_20[9]}
   );
   gpc1_1 gpc608 (
      {stage1_20[24]},
      {stage2_20[10]}
   );
   gpc1_1 gpc609 (
      {stage1_20[25]},
      {stage2_20[11]}
   );
   gpc1_1 gpc610 (
      {stage1_20[26]},
      {stage2_20[12]}
   );
   gpc1_1 gpc611 (
      {stage1_20[27]},
      {stage2_20[13]}
   );
   gpc1_1 gpc612 (
      {stage1_20[28]},
      {stage2_20[14]}
   );
   gpc1_1 gpc613 (
      {stage1_20[29]},
      {stage2_20[15]}
   );
   gpc1_1 gpc614 (
      {stage1_20[30]},
      {stage2_20[16]}
   );
   gpc1_1 gpc615 (
      {stage1_20[31]},
      {stage2_20[17]}
   );
   gpc1_1 gpc616 (
      {stage1_20[32]},
      {stage2_20[18]}
   );
   gpc1_1 gpc617 (
      {stage1_20[33]},
      {stage2_20[19]}
   );
   gpc1_1 gpc618 (
      {stage1_20[34]},
      {stage2_20[20]}
   );
   gpc1_1 gpc619 (
      {stage1_20[35]},
      {stage2_20[21]}
   );
   gpc1_1 gpc620 (
      {stage1_20[36]},
      {stage2_20[22]}
   );
   gpc1_1 gpc621 (
      {stage1_20[37]},
      {stage2_20[23]}
   );
   gpc1_1 gpc622 (
      {stage1_21[25]},
      {stage2_21[10]}
   );
   gpc1_1 gpc623 (
      {stage1_21[26]},
      {stage2_21[11]}
   );
   gpc1_1 gpc624 (
      {stage1_21[27]},
      {stage2_21[12]}
   );
   gpc1_1 gpc625 (
      {stage1_22[11]},
      {stage2_22[9]}
   );
   gpc1_1 gpc626 (
      {stage1_22[12]},
      {stage2_22[10]}
   );
   gpc1_1 gpc627 (
      {stage1_22[13]},
      {stage2_22[11]}
   );
   gpc1_1 gpc628 (
      {stage1_22[14]},
      {stage2_22[12]}
   );
   gpc1_1 gpc629 (
      {stage1_22[15]},
      {stage2_22[13]}
   );
   gpc1_1 gpc630 (
      {stage1_22[16]},
      {stage2_22[14]}
   );
   gpc1_1 gpc631 (
      {stage1_22[17]},
      {stage2_22[15]}
   );
   gpc1_1 gpc632 (
      {stage1_22[18]},
      {stage2_22[16]}
   );
   gpc1_1 gpc633 (
      {stage1_22[19]},
      {stage2_22[17]}
   );
   gpc1_1 gpc634 (
      {stage1_23[40]},
      {stage2_23[9]}
   );
   gpc1_1 gpc635 (
      {stage1_23[41]},
      {stage2_23[10]}
   );
   gpc1_1 gpc636 (
      {stage1_23[42]},
      {stage2_23[11]}
   );
   gpc1_1 gpc637 (
      {stage1_23[43]},
      {stage2_23[12]}
   );
   gpc1_1 gpc638 (
      {stage1_23[44]},
      {stage2_23[13]}
   );
   gpc1_1 gpc639 (
      {stage1_23[45]},
      {stage2_23[14]}
   );
   gpc1_1 gpc640 (
      {stage1_23[46]},
      {stage2_23[15]}
   );
   gpc1_1 gpc641 (
      {stage1_23[47]},
      {stage2_23[16]}
   );
   gpc1_1 gpc642 (
      {stage1_24[33]},
      {stage2_24[13]}
   );
   gpc1_1 gpc643 (
      {stage1_24[34]},
      {stage2_24[14]}
   );
   gpc1_1 gpc644 (
      {stage1_24[35]},
      {stage2_24[15]}
   );
   gpc1_1 gpc645 (
      {stage1_24[36]},
      {stage2_24[16]}
   );
   gpc1_1 gpc646 (
      {stage1_24[37]},
      {stage2_24[17]}
   );
   gpc1_1 gpc647 (
      {stage1_24[38]},
      {stage2_24[18]}
   );
   gpc1_1 gpc648 (
      {stage1_24[39]},
      {stage2_24[19]}
   );
   gpc1_1 gpc649 (
      {stage1_24[40]},
      {stage2_24[20]}
   );
   gpc1_1 gpc650 (
      {stage1_24[41]},
      {stage2_24[21]}
   );
   gpc1_1 gpc651 (
      {stage1_24[42]},
      {stage2_24[22]}
   );
   gpc1_1 gpc652 (
      {stage1_24[43]},
      {stage2_24[23]}
   );
   gpc1_1 gpc653 (
      {stage1_25[18]},
      {stage2_25[12]}
   );
   gpc1_1 gpc654 (
      {stage1_25[19]},
      {stage2_25[13]}
   );
   gpc1_1 gpc655 (
      {stage1_25[20]},
      {stage2_25[14]}
   );
   gpc1_1 gpc656 (
      {stage1_25[21]},
      {stage2_25[15]}
   );
   gpc1_1 gpc657 (
      {stage1_25[22]},
      {stage2_25[16]}
   );
   gpc1_1 gpc658 (
      {stage1_25[23]},
      {stage2_25[17]}
   );
   gpc1_1 gpc659 (
      {stage1_26[24]},
      {stage2_26[8]}
   );
   gpc1_1 gpc660 (
      {stage1_26[25]},
      {stage2_26[9]}
   );
   gpc1_1 gpc661 (
      {stage1_26[26]},
      {stage2_26[10]}
   );
   gpc1_1 gpc662 (
      {stage1_26[27]},
      {stage2_26[11]}
   );
   gpc1_1 gpc663 (
      {stage1_27[15]},
      {stage2_27[10]}
   );
   gpc1_1 gpc664 (
      {stage1_27[16]},
      {stage2_27[11]}
   );
   gpc1_1 gpc665 (
      {stage1_27[17]},
      {stage2_27[12]}
   );
   gpc1_1 gpc666 (
      {stage1_27[18]},
      {stage2_27[13]}
   );
   gpc1_1 gpc667 (
      {stage1_27[19]},
      {stage2_27[14]}
   );
   gpc1_1 gpc668 (
      {stage1_27[20]},
      {stage2_27[15]}
   );
   gpc1_1 gpc669 (
      {stage1_27[21]},
      {stage2_27[16]}
   );
   gpc1_1 gpc670 (
      {stage1_28[20]},
      {stage2_28[10]}
   );
   gpc1_1 gpc671 (
      {stage1_28[21]},
      {stage2_28[11]}
   );
   gpc1_1 gpc672 (
      {stage1_28[22]},
      {stage2_28[12]}
   );
   gpc1_1 gpc673 (
      {stage1_28[23]},
      {stage2_28[13]}
   );
   gpc1_1 gpc674 (
      {stage1_28[24]},
      {stage2_28[14]}
   );
   gpc1_1 gpc675 (
      {stage1_28[25]},
      {stage2_28[15]}
   );
   gpc1_1 gpc676 (
      {stage1_28[26]},
      {stage2_28[16]}
   );
   gpc1_1 gpc677 (
      {stage1_28[27]},
      {stage2_28[17]}
   );
   gpc1_1 gpc678 (
      {stage1_29[27]},
      {stage2_29[7]}
   );
   gpc1_1 gpc679 (
      {stage1_29[28]},
      {stage2_29[8]}
   );
   gpc1_1 gpc680 (
      {stage1_29[29]},
      {stage2_29[9]}
   );
   gpc1_1 gpc681 (
      {stage1_29[30]},
      {stage2_29[10]}
   );
   gpc1_1 gpc682 (
      {stage1_29[31]},
      {stage2_29[11]}
   );
   gpc1_1 gpc683 (
      {stage1_29[32]},
      {stage2_29[12]}
   );
   gpc1_1 gpc684 (
      {stage1_29[33]},
      {stage2_29[13]}
   );
   gpc1_1 gpc685 (
      {stage1_29[34]},
      {stage2_29[14]}
   );
   gpc1_1 gpc686 (
      {stage1_29[35]},
      {stage2_29[15]}
   );
   gpc1_1 gpc687 (
      {stage1_29[36]},
      {stage2_29[16]}
   );
   gpc1_1 gpc688 (
      {stage1_29[37]},
      {stage2_29[17]}
   );
   gpc1_1 gpc689 (
      {stage1_30[28]},
      {stage2_30[10]}
   );
   gpc1_1 gpc690 (
      {stage1_30[29]},
      {stage2_30[11]}
   );
   gpc1_1 gpc691 (
      {stage1_31[17]},
      {stage2_31[11]}
   );
   gpc1_1 gpc692 (
      {stage1_31[18]},
      {stage2_31[12]}
   );
   gpc1_1 gpc693 (
      {stage1_31[19]},
      {stage2_31[13]}
   );
   gpc1_1 gpc694 (
      {stage1_31[20]},
      {stage2_31[14]}
   );
   gpc1_1 gpc695 (
      {stage1_31[21]},
      {stage2_31[15]}
   );
   gpc1_1 gpc696 (
      {stage1_31[22]},
      {stage2_31[16]}
   );
   gpc1_1 gpc697 (
      {stage1_31[23]},
      {stage2_31[17]}
   );
   gpc1_1 gpc698 (
      {stage1_31[24]},
      {stage2_31[18]}
   );
   gpc1_1 gpc699 (
      {stage1_31[25]},
      {stage2_31[19]}
   );
   gpc1_1 gpc700 (
      {stage1_31[26]},
      {stage2_31[20]}
   );
   gpc1_1 gpc701 (
      {stage1_31[27]},
      {stage2_31[21]}
   );
   gpc1_1 gpc702 (
      {stage1_33[6]},
      {stage2_33[5]}
   );
   gpc1_1 gpc703 (
      {stage1_33[7]},
      {stage2_33[6]}
   );
   gpc1_1 gpc704 (
      {stage1_33[8]},
      {stage2_33[7]}
   );
   gpc615_5 gpc705 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4]},
      {stage2_1[0]},
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc615_5 gpc706 (
      {stage2_0[5], stage2_0[6], stage2_0[7], stage2_0[8], stage2_0[9]},
      {stage2_1[1]},
      {stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc615_5 gpc707 (
      {stage2_0[10], stage2_0[11], stage2_0[12], stage2_0[13], stage2_0[14]},
      {stage2_1[2]},
      {stage2_2[12], stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc606_5 gpc708 (
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[0],stage3_5[0],stage3_4[3],stage3_3[3]}
   );
   gpc606_5 gpc709 (
      {stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[1],stage3_5[1],stage3_4[4],stage3_3[4]}
   );
   gpc615_5 gpc710 (
      {stage2_3[12], stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16]},
      {stage2_4[0]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[2],stage3_5[2],stage3_4[5],stage3_3[5]}
   );
   gpc135_4 gpc711 (
      {stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage2_5[18], stage2_5[19], stage2_5[20]},
      {stage2_6[0]},
      {stage3_7[3],stage3_6[3],stage3_5[3],stage3_4[6]}
   );
   gpc135_4 gpc712 (
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10]},
      {stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage2_6[1]},
      {stage3_7[4],stage3_6[4],stage3_5[4],stage3_4[7]}
   );
   gpc135_4 gpc713 (
      {stage2_4[11], stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15]},
      {stage2_5[24], stage2_5[25], stage2_5[26]},
      {stage2_6[2]},
      {stage3_7[5],stage3_6[5],stage3_5[5],stage3_4[8]}
   );
   gpc615_5 gpc714 (
      {stage2_6[3], stage2_6[4], stage2_6[5], stage2_6[6], stage2_6[7]},
      {stage2_7[0]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[0],stage3_8[0],stage3_7[6],stage3_6[6]}
   );
   gpc615_5 gpc715 (
      {stage2_6[8], stage2_6[9], stage2_6[10], 1'b0, 1'b0},
      {stage2_7[1]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[1],stage3_8[1],stage3_7[7],stage3_6[7]}
   );
   gpc615_5 gpc716 (
      {stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5], stage2_7[6]},
      {stage2_8[12]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[2],stage3_9[2],stage3_8[2],stage3_7[8]}
   );
   gpc615_5 gpc717 (
      {stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], 1'b0},
      {stage2_9[6]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[1],stage3_10[3],stage3_9[3],stage3_8[3]}
   );
   gpc606_5 gpc718 (
      {stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11], stage2_9[12]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[1],stage3_11[2],stage3_10[4],stage3_9[4]}
   );
   gpc1163_5 gpc719 (
      {stage2_10[6], stage2_10[7], stage2_10[8]},
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage2_12[0]},
      {stage2_13[0]},
      {stage3_14[0],stage3_13[1],stage3_12[2],stage3_11[3],stage3_10[5]}
   );
   gpc207_4 gpc720 (
      {stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5], stage2_12[6], stage2_12[7]},
      {stage2_14[0], stage2_14[1]},
      {stage3_15[0],stage3_14[1],stage3_13[2],stage3_12[3]}
   );
   gpc207_4 gpc721 (
      {stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11], stage2_12[12], stage2_12[13], stage2_12[14]},
      {stage2_14[2], stage2_14[3]},
      {stage3_15[1],stage3_14[2],stage3_13[3],stage3_12[4]}
   );
   gpc615_5 gpc722 (
      {stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage2_14[4]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[0],stage3_15[2],stage3_14[3],stage3_13[4]}
   );
   gpc615_5 gpc723 (
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10]},
      {stage2_14[5]},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage3_17[1],stage3_16[1],stage3_15[3],stage3_14[4],stage3_13[5]}
   );
   gpc615_5 gpc724 (
      {stage2_13[11], stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15]},
      {stage2_14[6]},
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17]},
      {stage3_17[2],stage3_16[2],stage3_15[4],stage3_14[5],stage3_13[6]}
   );
   gpc615_5 gpc725 (
      {stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage2_15[18]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[3],stage3_16[3],stage3_15[5],stage3_14[6]}
   );
   gpc615_5 gpc726 (
      {stage2_15[19], stage2_15[20], stage2_15[21], stage2_15[22], stage2_15[23]},
      {stage2_16[6]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[1],stage3_17[4],stage3_16[4],stage3_15[6]}
   );
   gpc117_4 gpc727 (
      {stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11], stage2_16[12], stage2_16[13]},
      {stage2_17[6]},
      {stage2_18[0]},
      {stage3_19[1],stage3_18[2],stage3_17[5],stage3_16[5]}
   );
   gpc606_5 gpc728 (
      {stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11], stage2_17[12]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[0],stage3_19[2],stage3_18[3],stage3_17[6]}
   );
   gpc615_5 gpc729 (
      {stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage2_19[6]},
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage3_22[0],stage3_21[1],stage3_20[1],stage3_19[3],stage3_18[4]}
   );
   gpc615_5 gpc730 (
      {stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10]},
      {stage2_19[7]},
      {stage2_20[6], stage2_20[7], stage2_20[8], stage2_20[9], stage2_20[10], stage2_20[11]},
      {stage3_22[1],stage3_21[2],stage3_20[2],stage3_19[4],stage3_18[5]}
   );
   gpc615_5 gpc731 (
      {stage2_18[11], stage2_18[12], stage2_18[13], stage2_18[14], stage2_18[15]},
      {stage2_19[8]},
      {stage2_20[12], stage2_20[13], stage2_20[14], stage2_20[15], stage2_20[16], stage2_20[17]},
      {stage3_22[2],stage3_21[3],stage3_20[3],stage3_19[5],stage3_18[6]}
   );
   gpc615_5 gpc732 (
      {stage2_18[16], stage2_18[17], stage2_18[18], stage2_18[19], stage2_18[20]},
      {stage2_19[9]},
      {stage2_20[18], stage2_20[19], stage2_20[20], stage2_20[21], stage2_20[22], stage2_20[23]},
      {stage3_22[3],stage3_21[4],stage3_20[4],stage3_19[6],stage3_18[7]}
   );
   gpc606_5 gpc733 (
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3], stage2_21[4], stage2_21[5]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[0],stage3_23[0],stage3_22[4],stage3_21[5]}
   );
   gpc615_5 gpc734 (
      {stage2_21[6], stage2_21[7], stage2_21[8], stage2_21[9], stage2_21[10]},
      {stage2_22[0]},
      {stage2_23[6], stage2_23[7], stage2_23[8], stage2_23[9], stage2_23[10], stage2_23[11]},
      {stage3_25[1],stage3_24[1],stage3_23[1],stage3_22[5],stage3_21[6]}
   );
   gpc615_5 gpc735 (
      {stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage2_23[12]},
      {stage2_24[0], stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5]},
      {stage3_26[0],stage3_25[2],stage3_24[2],stage3_23[2],stage3_22[6]}
   );
   gpc615_5 gpc736 (
      {stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10]},
      {stage2_23[13]},
      {stage2_24[6], stage2_24[7], stage2_24[8], stage2_24[9], stage2_24[10], stage2_24[11]},
      {stage3_26[1],stage3_25[3],stage3_24[3],stage3_23[3],stage3_22[7]}
   );
   gpc615_5 gpc737 (
      {stage2_22[11], stage2_22[12], stage2_22[13], stage2_22[14], stage2_22[15]},
      {stage2_23[14]},
      {stage2_24[12], stage2_24[13], stage2_24[14], stage2_24[15], stage2_24[16], stage2_24[17]},
      {stage3_26[2],stage3_25[4],stage3_24[4],stage3_23[4],stage3_22[8]}
   );
   gpc615_5 gpc738 (
      {stage2_24[18], stage2_24[19], stage2_24[20], stage2_24[21], stage2_24[22]},
      {stage2_25[0]},
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage3_28[0],stage3_27[0],stage3_26[3],stage3_25[5],stage3_24[5]}
   );
   gpc606_5 gpc739 (
      {stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5], stage2_25[6]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage3_29[0],stage3_28[1],stage3_27[1],stage3_26[4],stage3_25[6]}
   );
   gpc606_5 gpc740 (
      {stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11], stage2_25[12]},
      {stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11]},
      {stage3_29[1],stage3_28[2],stage3_27[2],stage3_26[5],stage3_25[7]}
   );
   gpc606_5 gpc741 (
      {stage2_25[13], stage2_25[14], stage2_25[15], stage2_25[16], stage2_25[17], 1'b0},
      {stage2_27[12], stage2_27[13], stage2_27[14], stage2_27[15], stage2_27[16], 1'b0},
      {stage3_29[2],stage3_28[3],stage3_27[3],stage3_26[6],stage3_25[8]}
   );
   gpc606_5 gpc742 (
      {stage2_26[6], stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11]},
      {stage2_28[0], stage2_28[1], stage2_28[2], stage2_28[3], stage2_28[4], stage2_28[5]},
      {stage3_30[0],stage3_29[3],stage3_28[4],stage3_27[4],stage3_26[7]}
   );
   gpc606_5 gpc743 (
      {stage2_28[6], stage2_28[7], stage2_28[8], stage2_28[9], stage2_28[10], stage2_28[11]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[0],stage3_30[1],stage3_29[4],stage3_28[5]}
   );
   gpc606_5 gpc744 (
      {stage2_28[12], stage2_28[13], stage2_28[14], stage2_28[15], stage2_28[16], stage2_28[17]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage3_32[1],stage3_31[1],stage3_30[2],stage3_29[5],stage3_28[6]}
   );
   gpc606_5 gpc745 (
      {stage2_29[0], stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5]},
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage3_33[0],stage3_32[2],stage3_31[2],stage3_30[3],stage3_29[6]}
   );
   gpc606_5 gpc746 (
      {stage2_29[6], stage2_29[7], stage2_29[8], stage2_29[9], stage2_29[10], stage2_29[11]},
      {stage2_31[6], stage2_31[7], stage2_31[8], stage2_31[9], stage2_31[10], stage2_31[11]},
      {stage3_33[1],stage3_32[3],stage3_31[3],stage3_30[4],stage3_29[7]}
   );
   gpc606_5 gpc747 (
      {stage2_29[12], stage2_29[13], stage2_29[14], stage2_29[15], stage2_29[16], stage2_29[17]},
      {stage2_31[12], stage2_31[13], stage2_31[14], stage2_31[15], stage2_31[16], stage2_31[17]},
      {stage3_33[2],stage3_32[4],stage3_31[4],stage3_30[5],stage3_29[8]}
   );
   gpc2135_5 gpc748 (
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4]},
      {stage2_34[0], stage2_34[1], stage2_34[2]},
      {stage2_35[0]},
      {1'b0, 1'b0},
      {stage3_37[0],stage3_36[0],stage3_35[0],stage3_34[0],stage3_33[3]}
   );
   gpc1_1 gpc749 (
      {stage2_0[15]},
      {stage3_0[3]}
   );
   gpc1_1 gpc750 (
      {stage2_0[16]},
      {stage3_0[4]}
   );
   gpc1_1 gpc751 (
      {stage2_0[17]},
      {stage3_0[5]}
   );
   gpc1_1 gpc752 (
      {stage2_0[18]},
      {stage3_0[6]}
   );
   gpc1_1 gpc753 (
      {stage2_1[3]},
      {stage3_1[3]}
   );
   gpc1_1 gpc754 (
      {stage2_1[4]},
      {stage3_1[4]}
   );
   gpc1_1 gpc755 (
      {stage2_1[5]},
      {stage3_1[5]}
   );
   gpc1_1 gpc756 (
      {stage2_2[18]},
      {stage3_2[3]}
   );
   gpc1_1 gpc757 (
      {stage2_2[19]},
      {stage3_2[4]}
   );
   gpc1_1 gpc758 (
      {stage2_2[20]},
      {stage3_2[5]}
   );
   gpc1_1 gpc759 (
      {stage2_2[21]},
      {stage3_2[6]}
   );
   gpc1_1 gpc760 (
      {stage2_3[17]},
      {stage3_3[6]}
   );
   gpc1_1 gpc761 (
      {stage2_4[16]},
      {stage3_4[9]}
   );
   gpc1_1 gpc762 (
      {stage2_4[17]},
      {stage3_4[10]}
   );
   gpc1_1 gpc763 (
      {stage2_4[18]},
      {stage3_4[11]}
   );
   gpc1_1 gpc764 (
      {stage2_7[7]},
      {stage3_7[9]}
   );
   gpc1_1 gpc765 (
      {stage2_7[8]},
      {stage3_7[10]}
   );
   gpc1_1 gpc766 (
      {stage2_9[13]},
      {stage3_9[5]}
   );
   gpc1_1 gpc767 (
      {stage2_9[14]},
      {stage3_9[6]}
   );
   gpc1_1 gpc768 (
      {stage2_9[15]},
      {stage3_9[7]}
   );
   gpc1_1 gpc769 (
      {stage2_12[15]},
      {stage3_12[5]}
   );
   gpc1_1 gpc770 (
      {stage2_12[16]},
      {stage3_12[6]}
   );
   gpc1_1 gpc771 (
      {stage2_13[16]},
      {stage3_13[7]}
   );
   gpc1_1 gpc772 (
      {stage2_13[17]},
      {stage3_13[8]}
   );
   gpc1_1 gpc773 (
      {stage2_14[12]},
      {stage3_14[7]}
   );
   gpc1_1 gpc774 (
      {stage2_17[13]},
      {stage3_17[7]}
   );
   gpc1_1 gpc775 (
      {stage2_19[10]},
      {stage3_19[7]}
   );
   gpc1_1 gpc776 (
      {stage2_19[11]},
      {stage3_19[8]}
   );
   gpc1_1 gpc777 (
      {stage2_19[12]},
      {stage3_19[9]}
   );
   gpc1_1 gpc778 (
      {stage2_19[13]},
      {stage3_19[10]}
   );
   gpc1_1 gpc779 (
      {stage2_19[14]},
      {stage3_19[11]}
   );
   gpc1_1 gpc780 (
      {stage2_19[15]},
      {stage3_19[12]}
   );
   gpc1_1 gpc781 (
      {stage2_21[11]},
      {stage3_21[7]}
   );
   gpc1_1 gpc782 (
      {stage2_21[12]},
      {stage3_21[8]}
   );
   gpc1_1 gpc783 (
      {stage2_22[16]},
      {stage3_22[9]}
   );
   gpc1_1 gpc784 (
      {stage2_22[17]},
      {stage3_22[10]}
   );
   gpc1_1 gpc785 (
      {stage2_23[15]},
      {stage3_23[5]}
   );
   gpc1_1 gpc786 (
      {stage2_23[16]},
      {stage3_23[6]}
   );
   gpc1_1 gpc787 (
      {stage2_24[23]},
      {stage3_24[6]}
   );
   gpc1_1 gpc788 (
      {stage2_31[18]},
      {stage3_31[5]}
   );
   gpc1_1 gpc789 (
      {stage2_31[19]},
      {stage3_31[6]}
   );
   gpc1_1 gpc790 (
      {stage2_31[20]},
      {stage3_31[7]}
   );
   gpc1_1 gpc791 (
      {stage2_31[21]},
      {stage3_31[8]}
   );
   gpc1_1 gpc792 (
      {stage2_32[0]},
      {stage3_32[5]}
   );
   gpc1_1 gpc793 (
      {stage2_32[1]},
      {stage3_32[6]}
   );
   gpc1_1 gpc794 (
      {stage2_32[2]},
      {stage3_32[7]}
   );
   gpc1_1 gpc795 (
      {stage2_32[3]},
      {stage3_32[8]}
   );
   gpc1_1 gpc796 (
      {stage2_32[4]},
      {stage3_32[9]}
   );
   gpc1_1 gpc797 (
      {stage2_32[5]},
      {stage3_32[10]}
   );
   gpc1_1 gpc798 (
      {stage2_32[6]},
      {stage3_32[11]}
   );
   gpc1_1 gpc799 (
      {stage2_32[7]},
      {stage3_32[12]}
   );
   gpc1_1 gpc800 (
      {stage2_33[5]},
      {stage3_33[4]}
   );
   gpc1_1 gpc801 (
      {stage2_33[6]},
      {stage3_33[5]}
   );
   gpc1_1 gpc802 (
      {stage2_33[7]},
      {stage3_33[6]}
   );
   gpc1_1 gpc803 (
      {stage2_34[3]},
      {stage3_34[1]}
   );
   gpc606_5 gpc804 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc606_5 gpc805 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc2135_5 gpc806 (
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4]},
      {stage3_5[0], stage3_5[1], stage3_5[2]},
      {stage3_6[0]},
      {stage3_7[0], stage3_7[1]},
      {stage4_8[0],stage4_7[0],stage4_6[0],stage4_5[1],stage4_4[2]}
   );
   gpc606_5 gpc807 (
      {stage3_4[5], stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10]},
      {stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5], stage3_6[6]},
      {stage4_8[1],stage4_7[1],stage4_6[1],stage4_5[2],stage4_4[3]}
   );
   gpc2223_5 gpc808 (
      {stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage3_6[7], 1'b0},
      {stage3_7[2], stage3_7[3]},
      {stage3_8[0], stage3_8[1]},
      {stage4_9[0],stage4_8[2],stage4_7[2],stage4_6[2],stage4_5[3]}
   );
   gpc615_5 gpc809 (
      {stage3_7[4], stage3_7[5], stage3_7[6], stage3_7[7], stage3_7[8]},
      {stage3_8[2]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[0],stage4_9[1],stage4_8[3],stage4_7[3]}
   );
   gpc1163_5 gpc810 (
      {stage3_9[6], stage3_9[7], 1'b0},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage3_11[0]},
      {stage3_12[0]},
      {stage4_13[0],stage4_12[0],stage4_11[1],stage4_10[1],stage4_9[2]}
   );
   gpc1163_5 gpc811 (
      {stage3_11[1], stage3_11[2], stage3_11[3]},
      {stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5], stage3_12[6]},
      {stage3_13[0]},
      {stage3_14[0]},
      {stage4_15[0],stage4_14[0],stage4_13[1],stage4_12[1],stage4_11[2]}
   );
   gpc615_5 gpc812 (
      {stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage3_14[1]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[0],stage4_15[1],stage4_14[1],stage4_13[2]}
   );
   gpc615_5 gpc813 (
      {stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5], stage3_14[6]},
      {stage3_15[6]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[1],stage4_16[1],stage4_15[2],stage4_14[2]}
   );
   gpc606_5 gpc814 (
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[0],stage4_19[0],stage4_18[1],stage4_17[2]}
   );
   gpc135_4 gpc815 (
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4]},
      {stage3_19[6], stage3_19[7], stage3_19[8]},
      {stage3_20[0]},
      {stage4_21[1],stage4_20[1],stage4_19[1],stage4_18[2]}
   );
   gpc615_5 gpc816 (
      {stage3_19[9], stage3_19[10], stage3_19[11], stage3_19[12], 1'b0},
      {stage3_20[1]},
      {stage3_21[0], stage3_21[1], stage3_21[2], stage3_21[3], stage3_21[4], stage3_21[5]},
      {stage4_23[0],stage4_22[0],stage4_21[2],stage4_20[2],stage4_19[2]}
   );
   gpc623_5 gpc817 (
      {stage3_20[2], stage3_20[3], stage3_20[4]},
      {stage3_21[6], stage3_21[7]},
      {stage3_22[0], stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5]},
      {stage4_24[0],stage4_23[1],stage4_22[1],stage4_21[3],stage4_20[3]}
   );
   gpc1325_5 gpc818 (
      {stage3_22[6], stage3_22[7], stage3_22[8], stage3_22[9], stage3_22[10]},
      {stage3_23[0], stage3_23[1]},
      {stage3_24[0], stage3_24[1], stage3_24[2]},
      {stage3_25[0]},
      {stage4_26[0],stage4_25[0],stage4_24[1],stage4_23[2],stage4_22[2]}
   );
   gpc615_5 gpc819 (
      {stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5], stage3_23[6]},
      {stage3_24[3]},
      {stage3_25[1], stage3_25[2], stage3_25[3], stage3_25[4], stage3_25[5], stage3_25[6]},
      {stage4_27[0],stage4_26[1],stage4_25[1],stage4_24[2],stage4_23[3]}
   );
   gpc606_5 gpc820 (
      {stage3_26[0], stage3_26[1], stage3_26[2], stage3_26[3], stage3_26[4], stage3_26[5]},
      {stage3_28[0], stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4], stage3_28[5]},
      {stage4_30[0],stage4_29[0],stage4_28[0],stage4_27[1],stage4_26[2]}
   );
   gpc615_5 gpc821 (
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4]},
      {stage3_28[6]},
      {stage3_29[0], stage3_29[1], stage3_29[2], stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage4_31[0],stage4_30[1],stage4_29[1],stage4_28[1],stage4_27[2]}
   );
   gpc623_5 gpc822 (
      {stage3_30[0], stage3_30[1], stage3_30[2]},
      {stage3_31[0], stage3_31[1]},
      {stage3_32[0], stage3_32[1], stage3_32[2], stage3_32[3], stage3_32[4], stage3_32[5]},
      {stage4_34[0],stage4_33[0],stage4_32[0],stage4_31[1],stage4_30[2]}
   );
   gpc623_5 gpc823 (
      {stage3_30[3], stage3_30[4], stage3_30[5]},
      {stage3_31[2], stage3_31[3]},
      {stage3_32[6], stage3_32[7], stage3_32[8], stage3_32[9], stage3_32[10], stage3_32[11]},
      {stage4_34[1],stage4_33[1],stage4_32[1],stage4_31[2],stage4_30[3]}
   );
   gpc606_5 gpc824 (
      {stage3_31[4], stage3_31[5], stage3_31[6], stage3_31[7], stage3_31[8], 1'b0},
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4], stage3_33[5]},
      {stage4_35[0],stage4_34[2],stage4_33[2],stage4_32[2],stage4_31[3]}
   );
   gpc1_1 gpc825 (
      {stage3_0[6]},
      {stage4_0[1]}
   );
   gpc1_1 gpc826 (
      {stage3_2[6]},
      {stage4_2[2]}
   );
   gpc1_1 gpc827 (
      {stage3_3[6]},
      {stage4_3[2]}
   );
   gpc1_1 gpc828 (
      {stage3_4[11]},
      {stage4_4[4]}
   );
   gpc1_1 gpc829 (
      {stage3_7[9]},
      {stage4_7[4]}
   );
   gpc1_1 gpc830 (
      {stage3_7[10]},
      {stage4_7[5]}
   );
   gpc1_1 gpc831 (
      {stage3_8[3]},
      {stage4_8[4]}
   );
   gpc1_1 gpc832 (
      {stage3_13[6]},
      {stage4_13[3]}
   );
   gpc1_1 gpc833 (
      {stage3_13[7]},
      {stage4_13[4]}
   );
   gpc1_1 gpc834 (
      {stage3_13[8]},
      {stage4_13[5]}
   );
   gpc1_1 gpc835 (
      {stage3_14[7]},
      {stage4_14[3]}
   );
   gpc1_1 gpc836 (
      {stage3_17[6]},
      {stage4_17[3]}
   );
   gpc1_1 gpc837 (
      {stage3_17[7]},
      {stage4_17[4]}
   );
   gpc1_1 gpc838 (
      {stage3_18[5]},
      {stage4_18[3]}
   );
   gpc1_1 gpc839 (
      {stage3_18[6]},
      {stage4_18[4]}
   );
   gpc1_1 gpc840 (
      {stage3_18[7]},
      {stage4_18[5]}
   );
   gpc1_1 gpc841 (
      {stage3_21[8]},
      {stage4_21[4]}
   );
   gpc1_1 gpc842 (
      {stage3_24[4]},
      {stage4_24[3]}
   );
   gpc1_1 gpc843 (
      {stage3_24[5]},
      {stage4_24[4]}
   );
   gpc1_1 gpc844 (
      {stage3_24[6]},
      {stage4_24[5]}
   );
   gpc1_1 gpc845 (
      {stage3_25[7]},
      {stage4_25[2]}
   );
   gpc1_1 gpc846 (
      {stage3_25[8]},
      {stage4_25[3]}
   );
   gpc1_1 gpc847 (
      {stage3_26[6]},
      {stage4_26[3]}
   );
   gpc1_1 gpc848 (
      {stage3_26[7]},
      {stage4_26[4]}
   );
   gpc1_1 gpc849 (
      {stage3_29[6]},
      {stage4_29[2]}
   );
   gpc1_1 gpc850 (
      {stage3_29[7]},
      {stage4_29[3]}
   );
   gpc1_1 gpc851 (
      {stage3_29[8]},
      {stage4_29[4]}
   );
   gpc1_1 gpc852 (
      {stage3_32[12]},
      {stage4_32[3]}
   );
   gpc1_1 gpc853 (
      {stage3_33[6]},
      {stage4_33[3]}
   );
   gpc1_1 gpc854 (
      {stage3_34[0]},
      {stage4_34[3]}
   );
   gpc1_1 gpc855 (
      {stage3_34[1]},
      {stage4_34[4]}
   );
   gpc1_1 gpc856 (
      {stage3_35[0]},
      {stage4_35[1]}
   );
   gpc1_1 gpc857 (
      {stage3_36[0]},
      {stage4_36[0]}
   );
   gpc1_1 gpc858 (
      {stage3_37[0]},
      {stage4_37[0]}
   );
   gpc1423_5 gpc859 (
      {stage4_2[0], stage4_2[1], stage4_2[2]},
      {stage4_3[0], stage4_3[1]},
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3]},
      {stage4_5[0]},
      {stage5_6[0],stage5_5[0],stage5_4[0],stage5_3[0],stage5_2[0]}
   );
   gpc1343_5 gpc860 (
      {stage4_5[1], stage4_5[2], stage4_5[3]},
      {stage4_6[0], stage4_6[1], stage4_6[2], 1'b0},
      {stage4_7[0], stage4_7[1], stage4_7[2]},
      {stage4_8[0]},
      {stage5_9[0],stage5_8[0],stage5_7[0],stage5_6[1],stage5_5[1]}
   );
   gpc1343_5 gpc861 (
      {stage4_7[3], stage4_7[4], stage4_7[5]},
      {stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4]},
      {stage4_9[0], stage4_9[1], stage4_9[2]},
      {stage4_10[0]},
      {stage5_11[0],stage5_10[0],stage5_9[1],stage5_8[1],stage5_7[1]}
   );
   gpc623_5 gpc862 (
      {stage4_11[0], stage4_11[1], stage4_11[2]},
      {stage4_12[0], stage4_12[1]},
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5]},
      {stage5_15[0],stage5_14[0],stage5_13[0],stage5_12[0],stage5_11[1]}
   );
   gpc135_4 gpc863 (
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], 1'b0},
      {stage4_15[0], stage4_15[1], stage4_15[2]},
      {stage4_16[0]},
      {stage5_17[0],stage5_16[0],stage5_15[1],stage5_14[1]}
   );
   gpc215_4 gpc864 (
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4]},
      {stage4_18[0]},
      {stage4_19[0], stage4_19[1]},
      {stage5_20[0],stage5_19[0],stage5_18[0],stage5_17[1]}
   );
   gpc615_5 gpc865 (
      {stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5]},
      {stage4_19[2]},
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], 1'b0, 1'b0},
      {stage5_22[0],stage5_21[0],stage5_20[1],stage5_19[1],stage5_18[1]}
   );
   gpc135_4 gpc866 (
      {stage4_21[0], stage4_21[1], stage4_21[2], stage4_21[3], stage4_21[4]},
      {stage4_22[0], stage4_22[1], stage4_22[2]},
      {stage4_23[0]},
      {stage5_24[0],stage5_23[0],stage5_22[1],stage5_21[1]}
   );
   gpc1163_5 gpc867 (
      {stage4_23[1], stage4_23[2], stage4_23[3]},
      {stage4_24[0], stage4_24[1], stage4_24[2], stage4_24[3], stage4_24[4], stage4_24[5]},
      {stage4_25[0]},
      {stage4_26[0]},
      {stage5_27[0],stage5_26[0],stage5_25[0],stage5_24[1],stage5_23[1]}
   );
   gpc1343_5 gpc868 (
      {stage4_25[1], stage4_25[2], stage4_25[3]},
      {stage4_26[1], stage4_26[2], stage4_26[3], stage4_26[4]},
      {stage4_27[0], stage4_27[1], stage4_27[2]},
      {stage4_28[0]},
      {stage5_29[0],stage5_28[0],stage5_27[1],stage5_26[1],stage5_25[1]}
   );
   gpc2135_5 gpc869 (
      {stage4_29[0], stage4_29[1], stage4_29[2], stage4_29[3], stage4_29[4]},
      {stage4_30[0], stage4_30[1], stage4_30[2]},
      {stage4_31[0]},
      {stage4_32[0], stage4_32[1]},
      {stage5_33[0],stage5_32[0],stage5_31[0],stage5_30[0],stage5_29[1]}
   );
   gpc623_5 gpc870 (
      {stage4_31[1], stage4_31[2], stage4_31[3]},
      {stage4_32[2], stage4_32[3]},
      {stage4_33[0], stage4_33[1], stage4_33[2], stage4_33[3], 1'b0, 1'b0},
      {stage5_35[0],stage5_34[0],stage5_33[1],stage5_32[1],stage5_31[1]}
   );
   gpc2135_5 gpc871 (
      {stage4_34[0], stage4_34[1], stage4_34[2], stage4_34[3], stage4_34[4]},
      {stage4_35[0], stage4_35[1], 1'b0},
      {stage4_36[0]},
      {stage4_37[0], 1'b0},
      {stage5_37[0],stage5_36[0],stage5_35[1],stage5_34[1]}
   );
   gpc1_1 gpc872 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc873 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc874 (
      {stage4_1[0]},
      {stage5_1[0]}
   );
   gpc1_1 gpc875 (
      {stage4_1[1]},
      {stage5_1[1]}
   );
   gpc1_1 gpc876 (
      {stage4_3[2]},
      {stage5_3[1]}
   );
   gpc1_1 gpc877 (
      {stage4_4[4]},
      {stage5_4[1]}
   );
   gpc1_1 gpc878 (
      {stage4_10[1]},
      {stage5_10[1]}
   );
   gpc1_1 gpc879 (
      {stage4_16[1]},
      {stage5_16[1]}
   );
   gpc1_1 gpc880 (
      {stage4_28[1]},
      {stage5_28[1]}
   );
   gpc1_1 gpc881 (
      {stage4_30[3]},
      {stage5_30[1]}
   );
endmodule

module testbench();
    reg [63:0] src0;
    reg [63:0] src1;
    reg [63:0] src2;
    reg [63:0] src3;
    reg [63:0] src4;
    reg [63:0] src5;
    reg [63:0] src6;
    reg [63:0] src7;
    reg [63:0] src8;
    reg [63:0] src9;
    reg [63:0] src10;
    reg [63:0] src11;
    reg [63:0] src12;
    reg [63:0] src13;
    reg [63:0] src14;
    reg [63:0] src15;
    reg [63:0] src16;
    reg [63:0] src17;
    reg [63:0] src18;
    reg [63:0] src19;
    reg [63:0] src20;
    reg [63:0] src21;
    reg [63:0] src22;
    reg [63:0] src23;
    reg [63:0] src24;
    reg [63:0] src25;
    reg [63:0] src26;
    reg [63:0] src27;
    reg [63:0] src28;
    reg [63:0] src29;
    reg [63:0] src30;
    reg [63:0] src31;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [37:0] srcsum;
    wire [37:0] dstsum;
    wire test;
    compressor_CLA64_32 compressor_CLA64_32(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63])<<31);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he1ea970fe3716f84bdb433950a49d463d66b9f3d69f848cbdfdcbc30ff1cdb29a05b696d308f7b2bf0a61817eaba7aafb4569dad1cc8ad998a527bf520c7ae56dbc606d57ff452180cf7565799007b48bc8bb07b878c5126c5fa51c99db64732228b6ae22c4ed26ad94514fc9f303ee2efa6c922384c0409c1260804589a388215ab9a57de6a1dff78abfb9f4cf10124d0ef5d387544625dcdcea12bec392ae2b9dd8a294564cbb857c16729f2ab0dbb34c2e3cf39d7bd5006df1a75f276835b23d57d14fbc13bf98e4c17d640252d83c392189c3612c5759ef157ca5e09ae021d48e0c15a9112109510d24eaf80bd10acd60f58dcb685286d1bdc83cc8aa645;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h4997ce01d279abf281f28dd8e1871831deea3cd88aa0b77c734dee0324272e2a22a5114a678106ba0bb922f97b593a1c1da7952be503c76fabc021e435a24be3395b1ebc70e36ee65908a3a5000b2fb8cd05ee9766df0bfe308fe988a3da2bece73267015a05ced5eaf0dab4c240de4a027708f95a4fd0a2d901e45dfdd83af4e31a843dac5671248fbc635340a12cbba325caf1c418bc7583603f621962e01a14b082bb669f49132982cb437c079f0db76f68b3ce2db968d0fd34398ef32154acde02c076765f98fa65dd65ab277dd34a9a74e7dd677605de04fa358c888eea9bf420238d6a77c8af3185b59014f3c9713aef31c6d96d6955a905c426019c17;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h6bd04bd155ddb6b8c4986493a0fc3d419f0a4bc873f335a5a8d9d7b7823eaa2b5df54e03678699a482b82d59f62a120377eb866074908c26bb10cd976597b4d22bf92ec8fc02648fad8aaab103c8ba9bcee216788a57c9bd993850d8ee56e8bd88bbd4e2671bd368326a17142f0cb4fe665f49b758c545f19b8af267c5334584efe43e086bce3db66c72bcb0f07909c169ff232af44d741a0c6874ec0985636d77f043a8a436f52cb06ba07496063bf0fdcbc22e0e16cb78dac4cc80101a6ab08d130ea5cf6a7e37511d1c280520183b96892eacc6a379ed4bc949a564dc36101008464be1a943899e65b0acf231acd0b5987f66f0a564cf9e49a41539d30658;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'ha60ad78634509f362e7853c6cc4f280bd556882105fda7d2991c57199202b3d1ab070f059e03597b1e41a063034627d843cbf2bbb73db2c62a5d37eb5b9cb2dc5a1a0cb858f45461741cc5005a1d0f76958d9e4e3a72919bb23ba0d7dc44509e8deea51d86c37ed734f470f9c2490714432371660cda27c7a43c53315f09918ad21aa37fdb23d09d88c17439d141fda4fec87657ce25183a0c40fd0cc9b716a480683526215570fc0de64c26cdfe17ef592e916cfc80b844351f95e95b4e73a039831a4af2425f199ffce9889fc12c3cfe4784e315225b1531c416c45af55126e245aa39e6f56cfe64c9dec0591dfb45977eaf18388f086c111295bda7239e32;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h36b6467f4d716011b07092bf7aedb03694a38995d267ebf839f5f8964140aca1dd5020a607d17ce899e10b1ca5c83daac9d1aee798aaa8b8b091af6005eef86a2385c7f0958910a04dd3fa3f3c838120193f0aab5e24a9885b7caf487b19f6b6db1aee4838f37a117bf0e2368c6e258b5a9000265ce718ca101a05f23ca0dae98ae721dd4a259d526f1aab26d42a54c58d34dd1a9ff0dad57a0b2c0cc71666d3f969d2f07fc317e025d1a99b926ca471e527264c0119544421cf6bc62dd503b8dba69f73eb1bc685156a336b8784b2a80eda930ed000b63c5a178c2e4c1e1dcacadf19a3463c3322fa61a34ec291572ca57d831acf9871afd3e3882d180c9beb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hf7249486b28d539711cb5dca47f5e97fc8a58ecc1d4b0f6f3ddf90ced814585641817ff4239a48bac5d2be3baa346dadc22e1d4c6c5f207cd207fa0adf6600172cb71da7b368d28454bd0eaa3bda846853bc802aa6282ee09320be43770c01fc27e98eb8a1cfec11c696c8d7175993c45aff2ecd01aa1e9067d9efe76942befd63ab2b043bf9d8ad4e28df576bc1a5480972c4a5e9beb0b2fbe18889ce5f75ee32281fcc9e392a2a69ffe4d9698e0d06530301b7921eabdb53b178cc3b2f7b3817e25df5d2d8173419b08c687fbd8e9fe3911a4d0893763cd49581bdc8c59760c21361c86e4f6649d197b9e052e15d122a2f5d95c5a657ee7d559542cd6f549b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h32d0ceade77215c9a60671d9e032b91976f1b9dc58fead5a966ac8a96b09da2d2a5485048d7ebd4192f15c37a1bb133e4af558b300901a8a87d808f52867f97ba445a78e71a3d061f58b08d63bf514e7fbbaaefdffee19147804e4d03559390c46332fd027f1d9692823557a9f2d2401d9629cae68282e897bf3581a7e19f9fdf56e51a7f3ca25bb83ace267c56e2af28b3ffbab09d44bd442ddad6f255578e2f85af0687a3e469087b79496987f789bc3ea29b4ed19d3bb0880320962f33c4625e41e274ea911e8850326c5185763c7407de8abc77de8620608873e20240053992e31bf1ef328e6225a74dc68b06b0b9959a4fd4e5ce413c630defda275bc9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he7a7be5fa93206768717a989d21002d31a183f0dfd2a082f9c82a0c1ee3b2913a29bdfc1971df046ffc0371d7756e400b60ac5c77734fe1a8c0471714228b7800afbb7fd2d7c36aedcbdaab6b34fdb588f0bd966bf4d7ee60bf9dc1edf3b6fbfab8b2d4bfaf8e8ea0eedcc80ae1e2b4db6e41d2f9dfa7e057525dd80d9e4c8eb2100d2edaf5e574ef53da6b5e91c0f5dba84be421f8a47697d2c9780acc4fb2e8afa53cddfa95a1dd96d2a78460de55d5365fcc21d7e24feec69f7261f3bd9864e5e354265c86a87716846263ca83fd2c48627ad6dabcd0fa9ce9b8cafa1c95198046274455403ac8fc9eaff18dfab14c00eda116a980def96aee939f70ae478;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h4607755a89ea2906c42fd7287023b1a1300d248dca379b110995e645b7964e062e25fba48b625e2d78fb2c52d735d867b1092d28af9e4a65bdd2d65f28963c8dad5379fbc4bc9bef4bd7346241dc7ce363a9301d64e3270c978f74be5b19d5ec3ea8964b56a29456f8a233c9bb5ee6761fae99245509dc46dfcc17757cd9aee5dc74c2e2cf89855c40762f15c45ce302234204617c6396488116b5d6da7c86fcacc657e041e5526988385bfdb7882f5d06f654415d70f1a54d08a02ba4e0a81297633d9706ecc1c3575f3496e06765f3af1c5c8068d02a6c7e02469de8844f4b2319515fa5a78e3ee876cf65943c1e0d22069a4e510dd59698b30604cc6aa4a1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h50069436402c4e3e68767ae773e8b3d56bb91b0145b0e81302985bc7b26ab40fb48728a10821d842601b1a6d0966d06564e3ab296890e10fa41a46e5ff65b02e31b0f53b19856e75a73444efa2bb6bbecaca05bb1ce90e6a75c5b3b4771aeddaff94567a924efd91ca32572ab8ebf9504279f4557380bdc91756275b3650eeb11595cbc230325e2b6e4452d504f390669fdc71d04bf6f5c117ef920bac3b05a7ae1d2badde4c571c99a4971d5b1fa763931ef645c99d62210ae2717329f64c2409b64b85aaa2610cd099a397a29143f4d02ccbc9f28c8ff8236011a41620aa5d1d841f72f6870cf3a6ea92e4f8cf3e291b9d882284240aff58edbe18c9395823;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h73c5343a35e8f03509c250bf244df19e83a8b19aa40928c8109b9c708fd3e149ab4f28659c45097038ae5c038c4d163a2645d20c0bf62f56a272f4c213123ff4e27add18032c9679ea3d1c19bf91d32b920dc4fb38f81d058433ffdce8b4e416862fd751c7c44357a19f9d74cbf3261d7d0c84a8b18c8f6216f8ae8b31d6a9145e15c092f42a65301544b8a6d7efbbfb8783730123bca06bade774b1edc62f7d7701361e05b28fed822cf0c5a84ec5008b389c39f8036da2a4cd27313a496f1293c9dedff4a25d579cdef130fa09923f3287845f32f71c83417708f12c8a2648299d451ffa9ecd034d7c135b188fa653238c8562b198ddd6bb99804c85b878ee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8e9654197587f3fc7293118cfaf322db38155384d8a2db27ae914ccf1dec87799d061850bfeb748d6907e0e7474b83fb8a15fb421c37f3ac825867b535818282993d02ba9f7d88bb299e9ba74b649a80a47b734dd0448b17e6b2404f365a7ed48926e8bbf943efc6746be675c177bcd4ca64c962fdcbceddb4be7b74a1d69ae08045d61e6b93759800c36a667af86b4ee1fdb0f1ca9cff104e0a34af67f59ae72a186d79dc500f53038e97d2d434c2270ba6a68099740f113f7cbd61291ecd4848f31732f92c526ad476dda6e5b76b1da0b73ae8608d7d71b07c51c81488bbd0d79460cd0bf2c0e5ac829aac2c33c000ebc2064a7c6545b07a6be373d4caa2a1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h815e76ac622d0d7e34f5f4b3a5db990487f800873c60bd3af5a46725f046a4c4030ac0026802beec1a3905a390007ae03b93802d0dfca1e8aea0daa528a26c935d743d062e6e96f8734e00e7281066cca9d7f204f8fd45194719adaaca49b155e6043430e1d5cb8c95a390e80f9def4a78247f7580c1a61aa6a63e4f92e5c7485bd499fca27ee434dd980d84474b7ff68511f57ef1407cee598bc32be5bb2b610a3a7e4619f6329d24bdde6d9ea2b6a84f536e8b57ebecad4339b336cc4676b54a4ec67a58623cf50a3913a6b1acdf64bcacc0e73b0b0c79a3f97a435bdfee93e1cfd58bdfe9d7f99ddbf73bb0ab876bf93fffa0e0a65792c24b11fd2610c444;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hf10ac444d5dd3afa421650fba7892c533a00337ec63df0a773d46c2622c631de913bb70c47d7f4ee2873f583e3e966a51391406d2e3a21fe672c345ff2ed22d1837d6c1f7d3e115bd95be328ea0e1bd14ca7f219f846d30b7bbe3b9f951b2e1e5445d82df29c2cea1a35f883d0aa84344d02e02e08da58f029a10c23db33281344cf7fc5030433ba91505515d0f131c90ed351b9f26bb0dc6f3d33afd835eb39931cc251f6510a1a923119e88923da013ad5792441829438101647e26a7c12932db9f584421bf739353f0b854a58ff94f2476b3d0c8abd4ecb90c473d234d796b010770bb0a52ad7cdefcf5d8b9b26aa43ea3e173ac424276b46e7dd92f2df38;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h6768f6efbb8bc74a4ea060ff7d88ab33bd82adffda4436ad2a1771de8b20b4c06de95c3f79882b5c1d7c55dbaec59a45d11da13b466eff48a81a0ea31e27735a0d242c2f8510fe8750bf71dd28f196b41c8596f42713265ba5098496a356dc618625472e0c947f511e0f6215020080b49fe6d4c49214541ecb5947e6886434789bc293f2556498f549b495c1c73f38f8e8fd0562e97e32a1dc7244469b55998b9f5c22ddd59acb6b498faf09d4c8ba4a3307fb881e8c9da69e6915381e7c1c4e9c773ae5d6e819e843891693775f4dee237768b21d17d6efdd71e44a4a39e083517a17d7edb9c05f5ffc9f09d6933cbdc1719f4395dd810858c8abd720b9546d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he0f3fcdad1457061baa5f504460c1a5a90c06c7713470aca08100abd1bd7688243a00cedbee4c2e4f919ad2223cabaec14d5e77288d342d407a8e15c88dfbbfccd4910ca4bce74fa8c36710e451330b918f2da6157e7c6160466263adaacfcd902c5215ae371c91688bbc2a081dcfcaa1df40ec7c512f604db61cad37dc43e574f64e8d5299f667d45ff3dd5fc20709dc2cff0861d0e91a84e36f82f44b265bdb596b53725d38e765fe95885e591b8ee5c8770108318bb9b4bbc143d68e327c6157b5033be9c225275547234c9f6966da16665b7fae316d2066fc5cce336535612d2fe936faa08299c73d45e8136a692da393cf767876380f7bc8c490797559a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h7da11d92e144ffa09afa298748ffffc6470a2b25c5ff5d1a2aaae57866ca1f4f134abdb4cfedda9ae2f6d9232232cb26af4f5b020645af751635384e7bd1fd01b3c060b6d468ceab0d1d2dff29d89666c6e559f90b2b82a4b023fc75bc54b5639fe10de91926710e9b638689d92ecf2ad90d78467ff8d18281c7c4939ada4312b5debed8290fbbad2dfb31024c43b96f7dea3cd05471e1bd86391309421af807b75451d934ee18a3030a4e43ea1490dad2d78ea13612e128dcb342a2455e9c78ec53ab54e4b5993fb9a8891d45bfd4c1959784261151dd1f58e7d60ec68bb219ea01442d1d47d7bf8b1b58cb547e03b5c70ef0d1555e81b46f5fd2ebb5f2d6ef;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hfb6f6a48129e38f9f78e7f76fbcc89cc9c2315ac8b6c872577c2496fb9031f77a27dc41239225e4470ce4502450d8e99af6a34762e5725f040468ee1adf1f0ab7b32208a258e676f2e8606548fabc2b67621bce926d6501047ef32388836ec829d757bced99cffe47ce524d479be1c151e31d7db8600b60f3c814380aa676a5e66f0ebe08576c4590fb350c7bd7cf9f1184b29882423e1d307fee32d45d8cda0040a736b063517e9fbdb36d78f825123982c46f84f09cd52f40a86e3b4da498af4f1aa8540403d295e0b36adce7d8096f34734215d4f7995862ac8429161e485450373e7f3ea35c6845ef4e952ce5f35ec0a348db6aa60b8bd95993b63b1bfdd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'heae07f6b4520e3afbd6a65b04422667ed75698c6b7c7496aadb2503c13cfb2375956ca6dd78d39801d19e594e17357ced7281f249e759844b17b17ab429938aed8c8d4f3f65d376719b6744ee11ebe16b9ed60c769186aa88fc224039e847491680fd3bfe0d82772501402bc707a4fccccdd5667402923eb56a86dcf55dfd0de31709293e64d543364cdc6b9cb8874b0ea10d43ec80a7b4235ae7999dd647a658548a7222c45fe55f7e45f3e6a225f6dc570bb903150f2bccc8f6f764ccb5259e9ea06f257d9bbf8eacf9ca406b1be00d7fafe9babba3cd36de185cd202329e2507a76dbcc9c47d008878ab86f81bf73a15edaf5e4abe83cc42b2a8d65bf913;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h5c84f61650b5d366e08696e7d68f530d725b3b0a9731c36fdb2c9986f25fe6a6ab15d12d350bbbadab5522ad9a59714f64930c07186af5305afa1b037a8ecc5fd30be1eed8913a5298d6db4d1b0917b706686875520daeacfe47cf458ec817de1bcdf6ad7b755e5d6e526985859cc12e921444d98c2647c76dc0db33ffb6bd0d2733bbfbce97a2a416982331364b81c50be65f34f73c6732bb71e4db63e4631d16f99c3ff0162beae6f56a84657a088d5fdcef7fd1c2c819259b1d3d13291bacf73d2d73988d840e9cb45932487585163de49fc1c681b3b4076446128d75ef3fdd368fe5b79def4ac44585b14d173a17a8735a75a7f0f3047d257dccf8a47d94;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hd265bd11c6a9615fb13d6afb6edee594b713705378c2991836e6bc5bd6ab393bd9181bf0c7dc3f0b806455809c9839d10d1055d9783695bf5fb25bde3010f50eeec4c53be7dfa618ff2e71670b9998c496492596b36441769686574cca99db476e68b20435d778dbcbb9f6391d1995c577d03858a79cbd49e9a27548792cb1b1d7644239a966872a0cb98f4e57f3ce4836c32cc234cd85988a40c8c83f3af9555707f8876ddc84301f16c07cd1cd2e6b418a58fb94ad58f13a9c64eb9ba90482ba2cc751a56959a43d1a65af6193be0f046b0c691ed78d1a01660473109f07d32b2f0deeba6a14a5527592f876fa79e120f7ba737099849138c2934cf869fafc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hc819dd653d660363dc0884642f30beb40a63d1a342b8f8ea7f8c2db12ab8a3632828e9424417745c0900c890a8fbe4af85b492c6ac2408cd2f3814aa43fc7bbbd7b211edf1e8c1993ab6071b33f17b60d96da76e7610b4fe171d25e4cb67b6d5fb3790765d45146711c31980dc4a88be37dec4e8b247c5f9587d0f8687dd25bbec53daf4854a5722967fe9fad324cb222fe7f1b7d8629bcbc28f9dda163c0d7ffc7c3d95d4f6b7f589adad2c24d5332d2e3dd4174990c8b3527331b3c7c9c6e2e316aa78648f8b40601659c8a9d55a61f63d6d55ae40d07d4cf295f27267467362d20e4bc256663884bb6dc318b354a64384de57f1ab8fc34eb4a17227c96306;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h1f3ee527af2b4458249a91fed40e2c2045d12f47270b2383d9563cdf4d6b32c2ad4531d55577d3df3459843a6468964fecbb305dc86ce2c1f8c2f17624678a3473981706e4c4f49f6c152910c4ca4dbe9ef52f72163adde997a331d51971302fc61ded08f3b4efcb2b23173b5a4c3fe4318959521e5af26e6a3f571026d454068616ccf22f6825c44fe8abd4f73505b1395a37f38ad46f3b08c7717c862fa9bad051ceb5af7206334b67a2214df470dcfba1c8194a0c8e9fbf4ff47bcdac724f8641ea413effa46639ad7b2d5571ff84a54179d8d4cc73f69597309a803deaf7f5a8c097d4b7c3d44133f780d0812cbc5d8d7cb31aaa9f86fddb2ef3aaf38de;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hdb80987334c119c0b4be602eb792f73544cb21b488fd7cc22b07112a2b3ef4c3f2aec26d44a44496ee011fc80fbf6b6ae7fa1a898799c5de19c369f3dea59add9fedaafbbf84d2ba9bae0dd083eaef8bd38559a57742193e4f22a60dbe6132118dc561d43ccabebd87545e3da0165602991acda1960e8c28a6fc341579842b31e3ba0c477f459a9f97b36fa8a78a0cf5165204eac61f09059e72bcba2cdf21d84175595209736fab9c747850af64306671c6c855d3d04646aa29a5a7e3f0a30b9466d0639c975b7434addec7e277b96159b3424e7848ba3edcf098a8762ccfed34b15a70025a5d7867a05a1e7c588380cf944c4f0f67c2fcb9f97a4b34f71787;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h471a15ceaec25d8ef6c3cb7d62cca3d89d87135048e3ce38f7d1f7448de831fbe9b6e9ee899d495f689aea7e003a117693ba9e52ec7523b5ae405a667b36ff44fbdb1ca6fa24f8e95e7d33ecfd3159af1156a94f9af920065a137792e5cf9e7e2fa39291fee6cc7062bc9ba586d19362d9c0ea974e1f089d1984c2ed7cc0079d582265195f69cc58c43788f79aebae353f2c2d7e06a2dc88e78b4a3bc0bcd6d10c86c64b3b581f6fab3202da08aa0a881dbb1aec7a48b044850dc4d99ccab70e9e7a055424857af6ef102211775d6d7555ec01d216fb1cad9189f57fe36a69b9a810d9a5cca5c7bd24120b71a93b10e70983a42aa0aead2d94c7cefac0dc090c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h563189214bc47195308de1a0da0c212efe92f45d8815d78f83ded364c1e6c3bea7a2a2bdc88e889f38c1eaeab215d558ee325ffeba374ee2499b51066614aa50ae2a68bf3c023fb31ddab2c73f8414dbb78bc9eb288ca31eaad1222d514e73010c99fba7dd489334711bbd793098cb21fa72bf1e3412ffe4e2a22c2e56fe9a05c7a862da275eadc4457568b580ff73cecb748774cffc1740cc9660b8f5714677a2111e9ab81546816fcc57164984f241a155e3cabd482c6609d12ea0af647ed1695f27f3243fce08e50088bfc0cd89692606d76b3954cc2b1d4b11f0e6fe36d2b4739e4fd76114797e4e312cf2c006af2acda0ffdf50cb37eb2b5b099fc2c4dc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he29d7d7d7d7813f95f36744a45c9d65236aa85c439b7d7a8e96d67e0f196a8912e87e262b365162682d2eaea038072b220bfd07adce2130f29dfe6d5fad1c1a29758185bb8966a64bc1e4742edd7ab9b27c0aef3d4fff51b0a61e3872bcab502d0d7ea7ec67da2c66740df1b22ddf17d902e8ac4c0daa5c98cb11e67ace54b78ca61b5e677c9d8c61c8b6ef5e1eb19b4577b5a197afe944565249373c35d1292bd1092694db753fa87e116aa065cbd94b48a4c0a5292973486f813d5f42cbf99e4a5ca0705c89a2c17facfd3dc1e64f81cb513756b21277f9d3ae1f411d5e9bc1c168ba99efe399aab5972f390df95cc9e441fefcdf64aa7b02d80cc88f8a8d8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8d1c85ebf9941a7e73bc1fb36c3f7b940ba384b0cfa6d2d4355cba4f5b0706d02d8fd955263867680bfecc944dc8d495a609e68f6161676ffd3089edc62ccf97d9e8460be1427017077fb766c97f77e80c5e0bdf24e633714a8d3b306aa5df80cf146d7d94e05d7e141219168bff26acc9bec95caec87eeac928cb6571e3470dadba6e84456e8f21f82ba1f28c36f787ecd2c6a3133b68cd3a8ea02a0df1bbf8a1a1e63e9a30e347574f4a85ab68e0efdf5e71779d56b4b5e590d2c76581b105b3eb0d61ff8e6c4fde8dec8687f2b935c208cf152d585467e35d1b1f47fe6e8e75f0321887cae3f9afb7b7d90a193f41cfd0e613b39fff86ec1149cfb0256523;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h6f42ecf68934f31a137dd806ff9f5fa2ebb06a2a74ce14fa141d3c5b502cc5de8f3093892ef4dab9c4b349b83943aa8a55a09a6d84f91b9fb3159698d07bfa53b0412f468ef62120168fdc8b9951072761922c901b19e73c3e5a04d7e739c5a66adb31a367262a67e568bdda797536d4b2bbc28fdd0f4fd49da1d14457a1edc0f734ccf628f7efb2282c9aad98be4ab6c1adf8e1c237a8d51f1be5fa12a46af0812d7cc9348589686cc369778e84471d25fec180c1eda12097dc77e4f07c1838c6cd1c360bff533b8e61a158ffd7341a1651ef65eb23095e0f113b7af7c021dd2a8e21f9a80bfdf6b6d713656488741c0d23b25fefba97a4387546d2d58b8ba1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'ha10f0d8451c30b29c436f50755cb9312ce77ca8943820348f538867a24919a6b6a8670ec8f9acba25af6c36f4ca407b1723ecb2cd00199c8e86dd670d8900a9fe3fe4bb94ec8417390d38ca7825a6ff95ec4006d100e99934a217da46de4a8722489a289e872eb338c47665c73b21d0017f947e287860ef9be2ede1de8fdea76df70c106aa8a3f99d0fd475bde7b9a2fa54ac9a8602e3862a15a0c361ee5e78fa280c6ae3d8ab4bfbeeb44b5633c3fdd8617427619248c2efacbf5e4988daf3f4122e25e9a14b09cc412c528cf99e06244538d8bf1fdae6701a2b8be1f199f69900e1a1d8ed9e6c6305cbfd987a2ee1e1a3354d66396c2a6ce03aa70c9e73276;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h9ed9eb90dea538690fe9da2aed9f39c3353c0101ebc77a4784d28c2c2ca679494152d819e48721229bfff555c535539c3cb1c3154b86789a0e545e02e78837346828efbba26cdcd4cb5e2f6899d895994c2e203ad98693dc6d3356b2c081d61fc137ef26b2df5866a99fe12c2bc0c4efc768390885757f264581f45d518d30aed34b9b9b5e0521da46ddc7695f84b28cd7e8a488fe71ebed424a561f40de79f333d8ebce012cc227a10627c1588749e54e3ee34b9b5147aa44cc70e03837c4478bb2c6ec204c8d04cd67d695c51fdd1c81a1bc0dc089b829d86698d80e756106a4891274ff5691503117c1b8535e10ad0516605ad54b2bd16e8a489c712fbc37;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h67bebf89629bee55ad1a383db020cee96f697c1dc958bdfc5f3d7f5a93be5ea6dc4276e21de918cb600010efc57d67400046e8fba25a48db1777460d0fae7e5fdfb93e9e29e71d085a2352fd32ac3ef8e1976fd2cea9df8c911138cb7152e0cbe65761ed6fc794effe721139f299df864276b9a0c3ebd4553c5b0803f00150d64aad832581152352b189db56a2c1f64df47c0b4c91a91ad896f5d370b010d4861940076112d0ad2fb6f8f646106b8a56373decf604528f4cdca4c5beecd7fe5a6a584cf0b242bdf3a828d16658dfcc9681ae4cab8d90a8804d3bbe373cb93237ce62272398fa4c1bb21cebc8f1c5f4309fe41caf017a4b8f85d3afa832ce2a03;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h7f530f130c49a855e16c7351f8b875f2a3a62f08102374fc369f6380ed1a5cfe68a90b98996511cd082569e9abd606d5fbbdeccbc786b930a8d761c9f9c1f189eb3b38338b6ff87e933a55f78ef0d35ae7a7c4de464a9081353b395e73d74110633c1e406afd915488e5687b238811ad0c8d77326e35ba8c25bfb6cbe6664d72819a1b77bf5f97187e509a7002a35de9232c8f78b278fb022bfec634afa9a3c7df7ec390b488eaa128e4aaa918e2885df4058ab609679f077532659d699f9f6985ecbb7b359b7a6e0408fae1adfbce3d4bcf52e4b81d44c20182f6b01d5d22fb7df510a666782a73d200e5a6fef6d55daf9d37dbb7079ad5f0468c9c7477922b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hd5be570165da46df788bc1953a9c51ad428ab956be5042a55d7e5530a72ea23454d213e7e9d913daf481f0aff9b7962f28e0fdd8184949b4a92b8b60769d02a477835f47910256c1080c382ac106b4c05aae56aa8f5a3d45cb0c552d1e10abffceb6ed355824c4c89c53c8cd7a4125eca35174533bf298d45e9f84e1c6654dc2d335b85e135b4196fe56305ea035104cac9b22f14d55442f894f87afd4b5dc54cf24861b76da843f577974e880f97ba085683eff295c03b9da28bf916e5d4c0e3d89b8fc96e6ad0056109c4f44f31e7a3be114ad3966417c0f9daed917aa7311682392a768b4f0abdacc1b0cb7c739238199031c5e562818b670dd21586d6b63;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hd9e00bd1cfff82aa021ef6cdbfb96d505916e1414eaa1826f349a293d74f5b4e9e1c2df4522976c57d850385a8062f46ee2e9e657728d50d8049fc1bfc807f594ebb566a239e52d94a8a51463b42591b7ca377616d3cca72e80d8974f2eb812ae1a59b5b9f684d38aa834d08c133757301d6dd2367417f8e687aa2d674745fb5548bfa1cc918dda1f96d220523f46b04f4938f537f1e43781ec3a7b2000f85ef6dd69f7312ba5bb2f0330df8b9e42dfc6378f4b68f8d139f7bffd2085c4e413dc10b1e4535b04ef5d02f6ed2f141adb027abdbccaceea7e684bc4ab07f8824977d2067686d3c51baf3885afc102b25f6a8249e2dd8c9b53a44e7f03398241e5b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hc434ed5a58c73c72ddfceb65aa302af9dd15b1edcfc4d0a39d65e6dc1ebcf456c084c5fdec5ad37968d7fda51ac0e4d1496f94fd13781a8762ef522e6a7f15f4ec933b1d4c4cfb61aa9bbaedde270aef21f8b6f6405384b27a8f29eca0f81d3b3b3d79bffacc5aa4416fdef4e919d7feff79c2935ebdc1ddeb1348052709d9a1e171bb58cd07f4fbe46256454b0c1f984858efa846a9712acd5e7a63e74de3502fc8d333e87d5b0af9de450169c944c3695720bc8c5e301a83a2ca34f5e8a5eacdce983e128dcb8d6a0bf83c80e91dcbb54e4e4d2fce57d8e9e25be0da3f61c20f32e70378fe33796376d496261f77d2cd056e66e4150d698f91ce81ffdbd13;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h87edc67225d5643ba45d81b013985a8df958a99973b1bd67216a17721a60ad6c19a5fe438ade7bf82e63947a9b79a68a91e1319b2fe7f3b6ece978ee59eb7c69dddaf0d49a8f87e4e61b3aa1eb4d9e8b1d0d8ad7247e2279414dacc5e566953eba8f0d7d0e4a184de392b435105fa141dd498d392b8fe19186f1725a60af95ad6da7950144de48ddd7aa89dbd4d39f07146b843c49e22d826e519ed7da37317041e37f83aa0bf51939513fc147c000e58769d365212de79617bd3588137f3ecdfc3055afaecf34b9c3e8114b7637ee557b4ecb1708397455ac4043bdce166c6574588e584b15573de00fd10a451b0ae09c7b532361277385a836be6dc118a767;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hd92809eb766cefb91280ba7ada1ade2dced5d484551eb86f8087b408bfff8ccae72cb05376cccc2224a647cf71a9386e49fe3fc256df36a29319fc17a7eccda70d49d0fb3180e920b5071d4717399039afbf6a2d3591a7cfbdf715063b072a0bd720257655ea76e17df1509513f20c8f30e38e71a109568b112ca445243f42082fb9adaa599f8820c1ca0c320e67757c88cef36a9cd24ae18f59c9bed8d9f4dc6b4c53dbd258a4b6050f16ce7b9641006ef600ca986c270241d02d4d2d35a3512ae6591c41abcd14e3a236253312ff830fffe3cbcc33604b24058d1345f279e669bade712d6716053a113423dfe8c6d3b9aee3f6bd2db371ad2863c404cde587;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h6602247faf1be3a7cdf43d137fdfdc2a6d731a4194b38154f27e2c2ed40643448c9cc5a516cf5c7efb53f9ff24bf80adcbd05a51e4eef8b2c7958c49814239634f34882b354d01f49ce1fa6da9d28d112bda280f98e630c6a392e5538d02034322245c55d92e2e47664b60ae69786e0aae054e57b6ca05cad078e5730aa37b675b9d1f8b54cdb598bf16629bc44388d2cb65bfca35d781872bfdaa025d4ecb5a0858e9ffab7e8ade1a1431b2c7d1b97ce13906241983a922f6dce473ef8c8fae64937ef7a466908891814400f46f56f79f91b727258982ce3e744c52edafcf0215f6409d748ccfa3a9bcda8dc7dacc55fb21627a4b7f0de0ccc42d44dfcf400f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hc98b3bd806eb17016d9bdc0655886f0337b0f4e7905e54c4aace8649db9b5c32e22651cc69d5b0909e015b0b75630aa1032bdad143d6c7cffba06ef22d9a38e17cd002c78f82d9237bef08e88f0384448df698561e24ea27078d48cc457a2742d7005188a44fd6f364cff90412f901a0534a42819f1b7c3928a816917d757a4093285d0bdf62ba20ac19e19b1e1dd5d98d6a8e46b8d68250976fe680f9de2612eda2148d2332587f271225808b738af1c94933c50b9e78c4b8b741a0d5f2014fa1af03b5c928a1bb77c3e1f69400223a7cb6a2820261c0f482a7f83a12cd1cb874f08d03c293f8ddcf1be157155ac7d59da3fea4c843c59cdaffb3035cfdcd1c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he0908ab758444964912a489c686003881028c9d89d61c96e4839b966f8c88688530dae3e6b85277b8ab9c694ca51b71bce85718943d351377ca05e909a665148239c57a8a5e7e63b5243db743a55bef084047c366b9f4598e1e7793016fead901d28165065de2b5e8e0ab16a03d7913480af7b336832a590c5234513a7527969a0c24ea5bf5e088120a3377ccc9a4f1cb852ee206e598ee913b0b82c60ff8fe63c27b7261e51161969d824a6dd9ed112b79830e202e2185127dc68e25751180c23a7e73c7231501b7efe900253da6fbc3433e1db9700c7ae7ab674b83b249b3149c1a0e7118e8cfe8d091f7db8ba76074e583c0ca222fde4f309ee6bc419956a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h5d17b6540e66c3a5bd63c3f97a85c03478a6cb465b3160200a74ab2de489f9b4de76273c35647ab11a71ee1c920f2665fe777216f6c3c7976eff8553ad71a2a64fff527e760d961b9cd0dc43b5193ebcedaca3a6c6579ce89ecb5a6d4032b326de8b53011e50032d73025c4aeec00e914d4ececd1bab968f0be8f9ccd64f490546d2d93f04eac5809d96a8123e628a51a871d04bfb33aead84b1548e5358b79b4914e7b2408e5ffcad53ab62466f6671908ed1229530072274f28adeb29de7b69308fdd493404ac573e69df636df5099462efb8e0a136e881b7f16c4f7f456a0f9168f352e7597d7c57d2c5015592b3b1bc9b5127989638ed48762739fe3a0f1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hc14c15ec35c6103e4b22f93b3ff91f6e5e5f274650d427afb38afc722f7acc5f6975483f23ac4373f70e082e20d219a8436326b6c0c7cf75062fbe3a50d2d20f46660e0691c88fe32c4118999de3a1f8fcd294eb8acf5e6b1ca0e1f49293582d69e9aecd37164ed585c5b829d6287d2a28785ed9a3e48886c3097065749955416f397c49bd9e83166d47469d48db8c3bd99dcec3c01fa07e2bd79651c7db4024ca0087f647b524f8f2f7d4b8855a516adbbf51fd255067f1925c9c9fef56ddca5946f64e89b199384addb626b9c3285946ede0120cf981fee4f74e41adacd7382a7a76a41f73efed407a54e2bcb727c12012220f8908a142d3886ce8aea13011;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h862f0f2257d451516a2c39f1bbebc7b7508378de1828006558999849cde43348177b6e477981e2ad7d73d9f99c243f4aba5b2788a14033def5b41801bc8cc92a654f44aef12f91ca7d0e8ba842cff5e63f4045c2a133c8cc0a5dab3760c7b166190cb8089f8dad77e5239a447ce8f696a3decf4f4b9a099ee6d0276af85d596fb900b92f1cfeba73dbf09464a8ee1ea78d7c2ded3619831b9bd1fc52d12f817303f75bb0ca5014176c188aff3fe9aecac9393a0130bba240c7e209a1b930a7786f7b75ab27298a378dcaa69cd1c9d0fd7edb63031142af052d1701de3ae56998d89869518fdac177ae8d2d9b4c78a5c99bf62a812a4e0a8aca8eacfaaf5844b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'haf3f19a1ef52cce67a603f8a7da94b45840ce53a02b66f3176c5e392a0c3d3d4629e5262a5cdaad3b6ad44f6cbce53e3659180a72fb7521cf5c24ab7f89650f9dd940d4f1018259ea3fb9818854c51be7a97a760d53c68c5f92dfb12bd4986d69a167c5be2b431419fefa590629bc63012bdad97615cf7fe790c122a0c64648fcdc8684598b03f990cffb9463e990b385d7821cce0e01cb98b04a44cf16c553d2d06c0f5e5e58d743405364e0fefe64de70bbc1836f2a6e71e5899cd3b9eb8e1d45990ba27549f277b6fbad6422aecfee89b9b97499241274b5d9fe6d96b9412fd303186bc6033a491997096625627712e032cc80d25212546fa7ccf18230cce;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h4c167d8ed74f8c45b431d191fa48b72588e8853a0867e640796a8feaceb92c1e98ad1d2981b39d50ca7621cab4e7efe82e6d9d5096d2dc58bc93d8f02ef75dc7803741b8deddc2ae0d4d343b39624ceb0c8c7d511cb9a454bdde59dfac72b3af787d4435203654e96bfb0f03a85c6b27d2812be241df8fe7f55d5ec4473e84d856f8b0dd1bd9198d2de357b0c2ae23c5f12cc52b1fad2c2d8be3f724db405c3390cb41ab4304a547b3e14200790723e217dac1bef83d73ac57731450ba11dcbdb3cb9825dbce000324ebd2f740656bc670b7192de10af16f616b5c82af5a1f4a0ff741534d13f0bb42afa6800de941cf127fd4d88801ee00b897747fc5ad1524;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h52b9fe231c692024cdcd75b6f2b36fcf0cdf03b2692ca7a373e885b608083ddfa6f30f3655500856f839cb5ba8cba7f32647a424ea4ea27f1bbcdad8b49df2a87d35ab4b36f891cb5003c6df3edec66cdf8695c5ba9a36a6ea40f04a4802abdeac1b8c5f80162ade6161d14d034d03d086488424170adca7739ca905d918027d5217d18a0966a41eda7b4cda726226ab2a1f2958a460845a0df84362a21a6448ecdeb01e56b30d392cc3af4c3b8e13e396d44cfab1cf268b8291f964da0ad276d6117602740befe661873e6b66accc3deca1e2e098f678101ce80708740dd58541b0f68b10c79cbc64775a7e72003ee008813a4022b6270fa9d24a16272481ef;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h622771a5c9b1e7b0cb9a8fa40ec12dad523f2216554fd1851f077645bcff784bfd02a8f098a3c4ea524b7a12548fad7635fe8be43d830f6f39a9f5ec33fa4b98fa20a8d3e7e4e5e2a28cbe33faa2cfcd5703ab0f087aec2b97869d15fbc79d39fe39c888e3813089a8d5d3e0858149cf9e37f98d541eddcb38fd57e19d198617203ebb6cb5509eacc9367e695a15f1cdbd97554ba0b364b10b54de7eda7a2413b0c4770b6d12e25acd931752a7a071b56a2e6816d797edaee5c086e125cec00fdd026e654e2f370920404d3906b6084bfd40b180ba3cd2ec6a997a8e665cd321b300aae1bcd9f7f1151cfb97a8994d481592c5c799e5caadc0dd35edab8a5c91;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h5647bb85c33e5f23fbc0385f8cbe0be8da69ecfd172c802ad9c6b747fceebfdc964ae6ccc527ed6451a5a6cb5c34dd745e1d20d57251d9ce9b7a4644c82a8fcf2596d9ddd8169f21aa056c2fa9c9d7763f22837cd0ed144240c094c0c89c57ad6ed16f15e4d188ef29ffab83bdb5e78e0dd8791f72d12cc4655fef4513b179c2602dbe080ae9a9d5f4e83cc1f9157bafcd5926b58922a5c777621f8abc2a86d7221b5dc0679815f2cc48ff6ff4791e4cee2c4b13aa0eaf8d65dea3c6ad6c5cb3d4c004c96a56b3986d7c518a65d5ab41ed532e314153313d3b0a5f184bf7394ebcceeb48ffe3ccb505bb9571060271e87ee2ab56212aabdd6b15ce63dfc1eecb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'had57ec211a19814e45a78a718b9ec1baf8f966d0a2903c88ace220d00bc1ae3e8afc2a5e7ee420721021a88a3384f6d714f6f04e30dc8de603127c295b4a8e71560c63fce40ad49cd7340e27af37d088ff4d00103912e67c7868ac4316a97ed9492b4c59ae71cc4cddf61a0597fb1463e3063a8ac4010905b85d82fb8db12bb995f5f32411b892b1881ee51a3332a3dbf4a3b69a2616a3a9a50fbe57644475d4ff56c13409703d47187599eff8366ba2d21d0cf7b1f04e8965b243094c71ee8aad7bf73c953462db11d7ee64c4da621de044bd604e39671052d444044c6bb95a0a4bf708ee240939622cd2193758b33846e3e7fd3aefaea6bf663bb81d4ca838;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h830261922b1875c72004fb23874354c796d13c7ae2ed0948e3c4ba31f29991421e4cb41ac8cfdc5cc6410d1afec6fd94fe3d0c91e6117d406bfbfbf11cb85aedd9bf1ea1203b66998f69fa24829c8654685d4006b445d202f730dace951884df33ee47eb0c8ab1e1d063ce8385081b8f02517d96f3b3d9ccefe46e878346415b0c25e20e589eeee1352640618f7aa5734107d9bd3faac0f2a9b50a4ad97f16054558a467c317f6adb203209da0d48b21fb96bfdc4531a165942b934a6f44433b7c60af42089fb1bb8d70b4be0098ee619d1f21cafaa439317eb017ef8e56ae6e98ed7636f007f55e9255f808fa905936836950b5653d44f4da3e75b7809990e5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h31531d140370effd086cb7aecb13e82a7854cd9e7c784bcf390bbe4bf4b17143eb1a1317120058db07fd18e822cfbe9cc79523592fbd61c4c87918ba182b8dff9ac74f3bb4d25b6bebf1c7ad0b78219f00e4dfc505ac0fc3c565686365ffebd5f04391e51b61575d68d33cf76ffe9ea1fc86234ccda54095c05d7a34c052461e5378e752717efff30873660c9f2cb49b9f77825764173d809de01335490b17460ab47edccaaf61e95dd44a4a7d874e7932ce68495acff53d060e78826b9590f8327a1900564b70b975f5b07aac58b569338fe0d41d8a3a56b4bf7cc6c0f5880caa472f63b066524a548408f386fa26b758d6019c55ca5c144b977ad748664f0c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hb265cf659cb86fdf77f7344c03b2b385521ce9d5fa6183af3c4694ce7f2d99bf58e332c13bb32d53fd76fd7e89e6e7902aa60dc3fd4bc8a5abf3845ac9be9ce376a5c4ea4b1d8f15b92693abf0dba0e550761a00843c48e75a8c00fcb52f9562ea8b3c4747b45ecfd25137eab37ef9dc58ea4f6555d483cda5bc91b790ae7884868ad7a40a189363224b3f061b17037be04ebe58c8ffc320abd4dafdd38fcbb3ae741f64250702ab1ac2e355971231c1a8529018d107ef095d6222003267ff26723540b1281e3e71fd9dc0b3110201df6a3dbcffc31e3ed48e7007a92c7b52717235d4f5f28d8f1d7f207988b5a4a81d29964d028aa6bfc86b7134bd1e3f4208;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h808aaee0ac4ed2abd11c986416e37ef6940ef6789993ea76df71d1da4e3a60f610056118e2f85ebeebd0ad88b0e8e77bb0b40b126069d2fc32a5785ace501c61b6b61bd4650772c2d8c7131091ed3c6f25179c6128b372f09ab4cafff586451d20cf0fe4a49a38f50f21a6b1ea4975e983baea3f4cefd6e66c16f707ab267c59fe828c8cc219fe171b1ed93c260ce5ba9b41292363dd446433227cb9415e82ab8d854905321ef0f576cac682078070c0d4fda4d97f63b68b903d9cfe313b93a0ab91bd0c3eb78b65807671bad6f7bac26f0a7c7b603ca66ec402986f6354436c0272075587d1ab230bc934b4a523b84b9cb40229f3352b536f606d55f8669d59;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h92c575b7112d5655f3d7b6684e348a3b5ff0ea88d2121f6bd49215a04c553aa09e7e19547f162a1adaaec38574b4fad318d91bcdd13162e9855b82c7601b17c0d5f4e17a08228593dfd67e697c1a4266252d2f441c07ffe78a20ec4ad0728e375936c2cf7b93e3d747b8fd949d137f6b9939b2fff06e41b79a8bb7098ca1b03ab71d6ee51459a95855603abee0c2f3cde8ff82100d689027a223d9101b7c89af6691324e4d5b21880c8b682debe78119a67928a80d55f0b8ee577fa69a139fb5a0de04375f36cedc757fade72bdd4e97d6e1091b4f5b8170cf07530727b6d7bfcf129db8f894170214bec5a88a07d4c372a61d03e47d662c7af804050138d7ec;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h3edd55d955e06be8cfb9408e7296b086b473febc07bca7e0c0161d025bac7613fce4f5fe20f7ca43e00cac91db12964fac85c0197ef2a4c682f93d7d55e28b896290b90a2bb33b30e981b16ce50cc6f3442e59454082373b8cfec586b1d3f785f198221e2762f6cd6e3ae88a5fb6f44bfa7fff53cb6457b11ec2605b6c51ff7730e9f64170f7c216b8df609e9cc5d056848523d86bbad7d5dc11827239568fe8ec8f3373cb24b51f4072b029ec3a58a163a8bae89d848dc4cb5d92654f80532ddde70425e3ce5263c5aa80f894de4cb16231ae66d79a10dbf8df0e51b32ff8805b811a2f9753788f7352dff63a1d59dfba49df07c36f9738c78bc22fa889a26;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h432c8cb40f643349d2bd9618c7f28612c835cd0c4a7a57f1ff094dfdffd73b18782db1bf036341ef5333980f7f3502f8136c3df7141fcb69cc7a2bcf1e10305452b441b775f9377ce51bebcf7b87d59cff3d79c5f3fb3ead303aebc82b74f16b5213c45f464912141c57b15d4a6a8f56fd23f5625baa98d6c2e5c67c1f6da38942975e5bda1daa49d2e767ad98c56927868b90e339291cdc4ba07d08d093b7bf5ed82eae95dda0e0abbbc24039ca529f5942c385846d4fe22cd60114ff8e607ae8aad3f8e380db73af95dc147ad53c78ff35c15da5a8045f9e9f38aa6ce0c0c2c11febbbd3c3c2eb365a7d8e74f5178de097a5bd809d778e70d28524a64eba32;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h2a4f9aa9a006ebee06a1272575093e1fefb1fe138b3e4b585396679d358c00c96aab4843551735f02a1aeb9e384b543207aec6dc40e0a9d2adbda8b8b68a3a3b1088473b034fe98f38ca7741e0e315bbfcc2c8e172e87a24f87b23e94c25babb2d7a9b9d8441088554dfd29a29e91af20be619d942728a8f8d080bf36200aa63d1c5c45838e5081f335e44991aaf2d086aece2f5a6c813866cc4b71a2006fcf47b2fa817d2b0e9918babc60a644b8cc29d74a9929c3b73a599cd8034d9ed9e9e49b15ac1eb44c7741995aa4b0dd40a83363c06ba1587ab8d35f3bdc762e9d62f72c81dd8b6591f3da3e31a2ba151999cf9088328018800678643ff0e795ce98a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h36864601c895113f287185e5e5f6eea87c97d73c59d50523b4bc473fa7ca1c643267f9313ee5c1a02849b3c51b8e274301e09d9190c8029526874b6b19746b6456b88426f4406730f25208e8c9e4e18375a5c5619ac53b81ed5d97fdc6013ec845a81ef89a1c7fcaf51a957d7c3ea59bae9a4d2ad8c2ae9f21da7b6db6f4490d5bf872a6b0a455dd0c64ac14015e63b593a41e3c9f6dee2b76f68d47d7ef5c036213fd76e3d17c264d0b55887b7206fbf77134e55b3e91c89979982c80550f020ffd0eb634d214b89f1f34d7f370015c96b773fa9cc2549cd8ff49d876262cf8b8dbd156d17979f7153f927c506560fd158679bd5131a04110f87e3360f31e15;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h3aaaa83879d81af12f6943327709813e1cbd7b83974c5d058eeaa30d66ed4ca95ae86dc106d47952151830e01a9f76d6d2c6fe1891ee8665bb856bd6d932d428c6fe2091f2c0a0baf8854a5a73c5c38ecd0b1b4d834c70858b0b33409c1bb8520e98dfff0e48682a53a86b8c2701d046de52cabebaf32a5679139f1fbeadabb4dceeba612e8e031b7213707272c315ab3429ca4ff4bb5c6f61a0560f14ef4efa101ad3b7f07948cc127429b7ce04cb25340d629a517132b996f49dabd3b6824a4f38c6d77b3d3cfd8e3912519ec60b8330881f10b19884341b292753ec5be9fc23dbfa92401acebe191d3e54e27aeda130f3468b258986d6983f1a8b54e54dc5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hd9fa1ba3833c42838d5e612f6006d70cab22c45a7093a56de910b2ec9fc33bf7d0fc5f14856ed55147ee4131204718fe055afc33fd57d72bbb6b06392129c78e57004c230168b73646a69dce6161588b9f39101a0e319b8169cbd8891ec920d305c9ff8fcd3aa8ff51de28bb0541fe0b6ce6412fdea5436895b40a5f543accf822414aea39718d26e3437f75ece04b6f44961f4776cc8afd22c860e08a74633994e60c81063a3c1e79a474075b1de81abae1cbbb9a66528349466ec6b795adb90349c5644445ecda876b6acb9fdf76a01a236a4596155ea22db882ac87c53064b77cc3a3b92f9beb0b533776afa96a8166a830256c71937dad7f4bbbe8880671;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hde4dae4548ddd30328b2f45f233bfa34b395b47b6bb7a46a42509e059b17b36af9b2a738169651439a9a253bfbe8e77720bba8b1ee612be999e933f8db46e83ddfaff888678edf8bd03f8e5f245786991a205eda2d10f0adad1f10ff423063e30d9b9e04931f1c7e717816d9e7ec438036bf446b961a27d9cd4b29bedf918faabf5a898be56638d0a6a819ce8707ecb51f557c2dc73313a3cae32d0dad737539c1a48da94d81c61ca8e8ad4d884d1fe76733b3e9b818ede6da41ca7090c22b6550dd8b4c831a42733addbf7d4ffea6e66e9923a3496915e779edecae28e73aef5ba1f72475fc40ad5c79dbe9929069a8a134b88a6136065b199d198aa52cfe98;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h896147000c60c1e60aa1f94691ab9e0ac3d2401ed2debb2d16e8f7b1686d9323a7d6c58803d0e12bb0ce0887fe13b04d9d70f5934ec4a0e7940b5aeb6cc0a7cc526baa6600f8051ee2119fba0d4a83afa6fdc1eb1ae2e66504c168776d236462816fccb9e0e52b92e35340ba398b6d969dc8e7e569571bc72d4c75b01dc09fe09779207208d47c50619bfac5d176b540801e738a75c1c51cf819ae28faf3552062250a270bd8ae8ff53f7b326d8fe0f35f946de792199c97bfb1400431743c6f454f9f1e6ebcd14094cb6372e8ac81204043f03f9b15a07398e9032bc074b4e3c4678a254023b3908f10fe499a0299a3ba17e88bac5dd10f05de13c2e74ff37b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h7c1d5875256423ffd3fa96f23790dffa338649cca967e661d7fe177cc5b6227cf50d52de403f1ba3608020339a4ee18e18858734a0ef743a58544803b91c70d979685856ec4b394fb31c4685c79b45dfa1ed809d3a43157d8152127fd3bbbdc836c588eeb115771b15be9fbce97bf82774e9fcf459c18894955fc9eec331681daaf29fc26341652c470a354902104baafa57af02379d24d84cdee833b49f4d5fb6dbfbaa9974fc98442ab237ba233886d785cdc09720f8f5ec21f04b025ea87f75ae209ec38fb0f58a8b4ad1d76b2a8e0561c37a87e697b5e58fdbbae6ad165ea4d2ebb761ed3f707b86d8ba999012bb6c2420231c6a93f97781d2539b44d17d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'ha6de58e6aa1a49560ec1ba23bef2384857e400d8633c3039cd289ef10a0a9e14bbf7ffea8f3aa8b577447801efca78ed3797ba6f3a041d1917b021a646b47149dfcb5f8c88ac5975ab14cb35302a5995d1bfa650a2062d4553853a9e594abca3fe8f4d9067ca113e1f11ec312556a7a2c0cdce0a722c749520d02b263dc27ae71b6d9e8c811adc2ca76986bb565f5ad010156be5df249bdbb408369588f577be25a26dfb562918f5fe7724f7594585495ff86fdd27873c4ef7fafb8e6d8bf4017b5fd6f44a7d0ec739ca7043f4dd0a8fc9506c523a49291f3cdc5c9a986658318c68ecf5aeae7b987657649d55b2cfbf12482133e4c3455359301c4bb946591a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hd687cfe9fae47fb9bcfc4180ab3684910d36440cdbc652a779cb25b0759d0e2589255074499ce8cfeb883a4292aad958e11e09301e7a784b3b6f55829485f73dd0af5c040f2d5fb5fe211394027eeec9b1bf19da2340d53114c52ab7bfa4c3c5e15f375b1e21375114122bce0794111262ae7ada05c2748067025cc76a92a4a5f06c0b575b69c743578b0ebef1a52fc3368a0bf34b9f4ef583e340cfa1ada39d2f7725f42e2b86958fb7874d415ec3c85298b930d4303e8507ab235037c467b53ac6a8f170890a2b1652b9471b3d81b7d4fc248528e842a3a6a960da2ba86e605813bdd7a4eaf3ca6b3245f352c864087f603f3185e250fd8187ee58e2e800b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8947189d96d1ed877ca7805dab901c88009082453e7e6d13dd6211b706883950623cd09b39122dd11494c2db2ec96b1bd050460a59fff66ce33a22c55843288ce77e3a991a200447264fca21532ae1b58da1bf60b5f50a06bf364b37a1196928652c3a20e361fb3ed78fb394de8c9a7784b7c56f9fbd5ec163b26009fed161522cea2310c771ea237846de881aa45e073776396ac321d3bfbb9f443e1061017e912593fe8122c290444f1135d9f4fa1c97f15109a2b6db01bb54ebfca38cc43484552ede57c80f2ba25f5ca31d1e002b857e239839c315b8ba7bbd6c7a0975fff6eb6948053fed0e7dbc10056707c1b7bb7a9d674029c5b20fe23bdeeddcbcf0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8b579a2bb3019978ba3b2c7aaefc1e304103865ecf22a0bdc110b992b78593a69df6786543cec8a249968654c83d0f32835c4c7583adc82f40cfa42c5ec22c8052d9e8f4d62d3110a54b3d5d2d4d5b726001b4576e4a31238b74f13e4ffb44ef8f7e654259b46cb7fb0535862eac73f8d252c7ff95ca102cbaabd7d3bc3bcf1372ac685dd7f2a0efd8456be204909e530b61e9c1eafdf8647dded2c1f7e319fe4e1b6eb0c82b773b9b5456a9dfbd5c996efe5f5cca94c1ea800808e68f1e023afdf636bcf4959e827844d14d5d04719b22b075fca10bfbdd4a1a309cda4f212f82245ea1df3aa8a0e064acaa636c41ff3a88180d535c33a3a205df08811f5a76;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hc9c18711aeb3bb3803b12881eddd1b3511eca45536b456be36d928c835d1d13a73e1ae3a714a98b398df75641b27c441d09c16ad93b0eae6afc0dac3ad5e3138099efd6e9cf2fb6465d846b4381e085839bc89f041f0f4b247e0d1658357ce653ff1a087438097932bbaa517dc82022607446fad50eb70b708c3e50d8d8ab09cd8d16044eb69431eeb9371c0974e764453ade43df870f8f3739953ec90fad75eaba4a663ceb811fbb7a58d4387a1796785b63af0c4765f6254d086a889ebd591d04efa720847f08bb4eebacab5ffadb5bd949f4f767e8514bddadcb94ac2a3a8dd56979df3ad7ebf345dd61f999fc67eb6001599d5e2d0085e1e005a61a9743a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hc6c074f74c9fa21eaef009a163cb555ffd1d6ee8362b8ac93681b5f82b0e761d7a24fec1598af2f9804aab78ef033ae3744b010b0e0d115010084aa2bf43af56f5cc55fdb58b721bcffe17997741ed5b001e03ed9bd941495b90cd58df4bb6ded5214bc95727fb7c766fbbee64c9a9d66168a22658515381b5f958f286cfc8ac767c5162494bf369f419002252e8887926d6cc5cd2d19df0f63eec17aa6e0ea35f1d70e24bd67f10892e4c2ddaab95ac82d682511b31f471341a6db5178650d43eb984f94f65ffb162f13e7b4ba91d5dc7c8758fd5733cbcaab519afab5249f59cac94734baa73c6acddecec1588e5f3d05a9f7e2e47016b8fc43361de1da678;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hb86af6504fcc7655177b58f8d11b87f00d7369e0a7db5fc4eee7677ceabef5d856af60299b6fa033e70d64dd27fec3a9dbf46262c1600459042d66176fabf429c0184cf969dc24d2ace081dd5051a0e93b3901dbee99690b8a49a17fed12a19d0e1355ca2e1e99e3e9ac8c6e510dbc1ed1193bc684a71701979e13195cbbdd1cd2d08006f712d2484b865e2fbf761f6dd8ea11222aa6cbf1effc6db328c517ee53bda3278c9c8d28707ea8ea6741e4303f7c39fce06b3275cec958e597c6863892042d246ece54f8bdbaaec4ecaf4deb1dbbbd3531e826a3b8bade8792b63a4d1b695dbbcf0152605cb9f62b2cc4b85a846eff092c1c1baae3364afe3bc11897;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8b2de9f9e2f47e31f3be4142520dbc6b555c30b41a6198b229b084feffd01f83e07a1ee5c99f9f43707fa52db999ecc52a4ad71e162c9c283723b0d78579d17ac28e4b1d49eed7f58a818b6649fb4324a92d66e52fee3f902249748483fec25f7495992ecdc63a400d0b996001df36ce0f93d12d662e099a3cff827e325ec2e70693b83627f4560df41de7bb12552dbdaca0d99f6098f037a71ee0b0fef7658bcf15b973efcb0ca8ccf9bb5d31b4ace89aa6ce04589c2c258c7a47dc873bf097c943b3f5e5cb574e0205409d49035d7e5bc8e0e473faf50f065d2b29c22578165f4543682f31a68c1131d7ed4f1e999f38cd930ea94cd65cb37710880ca5fc2b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h6b24b2bc7f938140468ab7773017d0ee4c7971528ffd0a671e3bc2736d7393382ed017449f4940658874bf00bf0f9e7508daa73d4592e96bd7cc0a442a4917a3e443fbcc260d7786408973b262d8d35fd3e87ff7a89f0682cb18c40aa56ecabf03455a718dbaa6cb600e5d086163b4215b6c2d12c461a3ebfa0058eac4f7c2122d093792af8c51d6fc69c445fba79bcf80be39105962f09ea49c367b6d55502726706d573971be3bebae623131e5f69556b16a429e8ddc982850ab117975def87f73a318a10b7db433d19994bdcc30217bd7f885adbcd103939c8a92143fc3871d890d14ab4205eb5b0b3bf3c2ecb3e0306a8ae09f5d3312ef905c43e6e31175;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h302c6b8bfa5b27ac1058f8f8fe530d2d198004a0878ef480b3060a4e134b83ca5a2ab14e1ae17c5c5ea8cb69f4b705bb8db3f96f0ae5ea1f52abcf89f46b404ca18abc4aa851a2f6a4928b65f6eab1fa1621604e645f9574c8701a35e211ebe8645ff62af73801d6dceb738ff691ced3085482b8872f9a3767be278cbc4a7c29a714c7f0ebad3d5f9dfe6220cccdda56f73fdaf391e385f2d3102fabf10589420ba5195767e041bfc56ed8b495ecfd0f7787c710ff17e603638ffed43a4072c1c50531ffa1f08f378401e69200b116f51ba82a64a19c0cc035c87c35dde256342708b34540eeb60e768acc7c2313a2544ce20b5ac1398e8bcc9600da3d5ffb7b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hdbf6b7470791d409adf3aabe2fbc67416d851b2dba21296a1e1900bec56780465176c34746d72a062b6f695eedbd9096aa367295db495d014dedca205afeb85a9c341e340519b19b99cb14fe9f97e70c42fe331070a6924eb0f16149e4259c15f9b2893e101f5fb8cacab920ad8c2a4739f304fae3a6e7742a6a2375dbb4149b73c184c7de32a91e57ea6d7e12e3412f52a9ce95bdabc1b11daa5e94276f65ecb621f404f6c7c5711e6c6a65da403142d704148fcf5bbfcad3df6a2640cb50d9c2ac3b7942da8920cdca30931b8245ae1224451ba106b682e4bb789928b7a0bca22702d27a9e4a55c2a27d6938a8f3ca8fc135024a6624344fa20d556d28f875;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h521dc8febff7dcb0dd7614c7551b0d00c82af8aa6adfc3f31af38014a86640acc4d00644aa5a04ad5f7c7409090307f9baeb36ba2f3822ed3525bbeb40bd20fb54a6e8f903aa6e646a32bd7a647abbed60b49927cf60167ae6d670be6d3881f336aae9831bbbd7ba8601b5f29e0fd44bcf00838903d4f54ce600b9f7a0c8bd31ea18e72d47a41abba85eface125b78cdc9194caeb6bcb4adfbe73065d7d80ec81a486062da740f74146f2676940120cde2d31e28ae3deb72c15560e34eaac9e06ef2259ba417c4b10efe06dc4e791b42764fc9ce78edb51fb794c2f93bd1db3d8ea9fefdbd8c2b8d4ecd7d1e9ed7bc4c7815ad6484415e17d8c6727ae78abb83;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hc2561c9d25de387b575db2238f835a73a900f4730f080533d19a31e0cc6e820f2cf4d2b19c396ca9ef5b770138e1b79f8d6d309f851a485fef633d553bc879bf03e030c5bbdae8e0a0ed2fd1bf580cc170ea26e9ba2ce24e32793da88aca33654297442b4e25824146c57ad2db77dcbde3891811da04bb079020538a43f655e7cef7946066926452eac0dc2deff82ef134e1b0f8fe2be023340acc6c3bafcce8f07e09cba7ae9a76ad0ab01867c5daf6f2787e24bca27f0320a8032a7a38c3a2c5da0fc72bf02e93cbe3b40b358bd11741c176000be5b9caa0d7ff550ecd01a4eb428ff3c99b438572bfc181c40817c64c99f8fa7091a55281ea22c4b3b20a2d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h6da10c724131cd6875d77c8d22e25154c603fd7765ce4eae180e21c79905d28c0715563eec77dd76dbbc3bb0bad24a0f83368bd1cb8a5180588dd38eeed5265f1d1bd74b29b0a13fca215d81c5c6a5323f7884b277e4b6d629204e4129e8b1b797c8e3825fa1a1c5d97eeb4b0e3332ed89394d0afeae567b9000aba6b072853c296aa58eb8c6799d296453d844c8279c1c5f9b6fce556d3d92927f66ca2f16cedad6600c9823a7c67d3ab4d7e523ae0ef71ca79947205166540a7a115caf97cbbe2612452af8d8c6ab476b8fc1bb2dc042be380dc20bbb6cbb692232a46f0af1ae98f1e8197a30938c72347801b2615b9f3fe17e5b8cc7c7a693915d2324f1ee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h3c6126fc770fd012ac52c8b83b8c02b952850f78f20937c9e71524c67868ea7a214ce16435b9e67ba9bb2c22492c4293afa58fb54e5c81c24dffbb3dd13ffb7b93a42d3cd20925972697e7d28a1f81d1cd37f5300efbf08bb06bc36d3b750b2dcbfba9f48422b25e0227b834d5d08ef48af1114cbe97a59f5feda1c4e048542a2c1872e7ea5b0e5906578b46818a7ae10b6d41a9556412c6c2e300f3ba9cc18c0575d62c3da7e1778048568c9d01e0dc4af27fa731d4cfe3660d1e567cbb0d2b42fec39c3a8ef53a65df092dc18dced571e0ecdf6c0ef4f51d90de4071965a88dbabacdda845ba75e65da13dbfae09cad6c7603113d5011cb52abe961021c47c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h53177389e2908f145ed4f840f9059108c4bc8270dfc6535eef150dbb4be1aa0f253cdea5c9b285fab27014f2653c0079be0cf0c4f5ab1229bed1f4cc8ee75eee75ff199881a603ea76bbc3b99cb097a1932fcb52e58c0db923b077f0987a434a1df7eca17d3247749584022691e6edf487e59be7f48746d571d617487d633f43dee4a15e70dfc2b36d1284e4b7da83d97fe4f943834ffff6f02e54a97d24976dd626d0574e5987ba280e1d4bdcf02349a298a2eeccd098cd2b300e4c5276b7fc7304337055e1ddea38246410e288b20ed962a41257c428788ff58a1a5f2844f95005367d7ad2c8910d59e9261209eb40340feeb3f7ed9bf68f416717b38f8070;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h5ced8dc99c8363252d9933134c5fc5f073bda92bfa754cd6ad57c14f6e8137a00a8efac5edcf29959af6543265d0b53cd6a27b16695bda32b9c2bffe4f9061ebaeae1fc33d35fd4f6255c47c2bd3135b339cde4357dfa16ede2f5036205186037a50e400382ec2b117208a1eb40db3919aaefac61c8dfd17b9ab0a5a3dbb9c34308557224df57938456358f2088fa28e8ee3d38dc515ad8ee5fab91cf8af0661a344eba44cd25ab961953689c49d52f32f34cb2cdc18f088d7e6323fe8baac830e17fe18414b15822387c7971cb3e5e19e651a1c4e819677b8cefba8604f5ab4f75a24650f74ab7244c7ed15f316eda617758511ada29ad32633a11a6de7c762;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hfaa0d9e01aad090044f001ea82ae73385e7d2307f1721331280424f5ca2b085e7c9edd26720dc8fc041365c5b0feee7f17d7f0333a6d7b96c8dce70b6dc589146bafdc74ddd3441b63cb6fdc0eac3a39564402b30da97504338cf4a7fca945f4cc28e8cb91ff9c1c9581e5f5e85589f7ffa9f7ddd21a0661174d30e1beefd24b947a1e8f39694398966bdc4edce1a87e4b78b018ff6cb5efe90bf6bb588f05a3d41ac652d2bf6e33435eb87ee215c57db64c0fe7be07681c6b602447e3f7a0ed4cb2797257d037ede3238f646e76ba37d41cd964b98afa197310aa5ed02f8a030240dda67d86a9d1bffd8f0cb76f3c740dad500324db38d766c0574cd1fecdaf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h7ba73612f2e043528becee5e8d2683438fd00275fa5d2665b043059ea62dae2b671e64588b5400b1b4c686e8044593bedadad47d6c5c305276d044d49e7afb0e752b2d96db83e4612d6f07ec56c17ad21d5c6757e9f3efbcf2ba7600f5e927710e9902e1b5dc79ee82238f3c135703950c7deccbf59a48ce9e3a19d382d81b71015f5be0630a50bc85c824f24aa1659abd4348781dd603878e75f547bb51a244f42d2e574132cdc42ec442f7083b915cbae8df2e042c70466ec503d8c924a1f24967595224034d8bfa1d2227c2106c60ef8b3c515515bddff19e71275bd1f2fb8faa81a0063593a5e02538d8a6e64edf137211ec01c934d0df4c373a56b6eb1f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he2dbabc25d4545c63bf560d1a75a91561031b8052c7ed2acd82b7df7b3203b031a31237252e4332e45c1b8886e530aa9e0f053acd686a0e77556871077378fa609de98f2e1aa20454f0944b55deab2abdef7ea42915a1e34afdb57ac0d7ab2abd9df02e6a9a361e215ba17db20fbd69ce6911817ee94c6b83585c32241bfc74da36cd1d15bf2db9ed6350663cb2ae761533a1b8aec844f32bd6563b08bfc8d291b2d74b843ca9f7c88f8e3d139f31ddb905a10d6b49e9ab98da14798c58bdcfe71d28b7944f9c0ba321eb65a5459033532741c6c8a71fb3c26557228f71e56524930b77150600f55df695165cf756fad1e25f603e97c39f8875c249209d34b91;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h848d2da80fe45dfaf0b834040980353b70d9836b141daaa560f5165ea5ffc39f3e31a969d97ed7e4e06996401252b7fb1d2ea2fbf95ffe2e2939e0f53b00ca1bd9b92bb075efb64687cd30905f800c0dd5222445a8c6ddef7bd32259e0ab7ff435444725c6903ea42e93eb30801a0bc2e5f658e21185977932480c2812ea5fb8a29d9e55cb863a4c4960a29ab6146942b502e1421651ed642bb18b55f79184fe6e71c3a275688a1e56c7ea34ac94ffbc1e4ca6e2798073e9bab5e032fc269460aa987a17a6eb2dd0ebcb099b4cfb0aaed494cb31e72fb4f2e9a4cb80772360e9c4edb87a7f4f4fdcbbbea1a11ae41985b7595c1fa2e265b048cca3f9dc111891;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h36499f7b24887c0992d276cb84019d5a3afa4e1ffdd5e3249f78913bac68992c5a1639f5857d3c2c15badee6dee883f883e0a333416ce28bc0355ca14b3933807d13eb4c41ecee0e749d1c369234773365ca67dc14ac4a867bcbece9f01372ba712544bfd2b39ad59851985f20091ad76cb116deb553b18a753ebc0038cfd9791b02d65679f564234d68fc1cd819c29fe22e07706c3f45cb561a2bc7f8545508328938a2c97fd4aae5e17e493e7c0a93093ea4de16a29be097b7b6404fa98dab2ff8ac18629c4e30b8cb8f457817e3290ccf8f8d16b3a8dde1e4446783066ee1a02baecb143a9313d71f63c8853a9ab63be0758dd9cca3b205ef5c08e0ebd200;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hc86a163a12a00f587be72c22ba242d68c4c720de40a8d72596d1153c31346e7868c1b11a7376719284c6432c963314149c7318e2bdc49a464105521516a09afb2f87575b143810cbbefb57426ac23a7043d20b4fdaff1f4f7bfb4452a4b85fbd23d22854393ed73a8a0d3b196c082f19f187ca848e1a58becc6a08743e9d247adf8465adb1c15055deb38df775cd1b1c37b61c803cfabd75340a60bd6f906dcecf27e837d21cf32f293cebd0e14c8f9d8c5858c0055aaaa02c941c5a821c77f89eff6a49be35e9efc87beb982bf23f90e4a499f5b4c32d08c0cba376b50d6ba144da00c19863d1a61a26892359c39c0e7bba6e3f684f62f812470c835b3a6557;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h99a243285ce0f57c0c5b805199aac323f8bac2389000f126560bb4a85218a52fd3b1ef6de5cdbe8aea2e5949a7119830d2001f87c90c6a7597b24866bd31f7def616b495e214b64590a4d19259f54e39c7d990987c0d8ebe55f0b105d2a3c5029e96c3277472fadddc76de94479baa6b2a05a9662036b23adc6c88d77ead0f8ff4621a0f5558d4d7d0494cb000b58183dc01851f4203774697ce678e79cccca6b6816e8a183a9fe7635edf20da0c5dad9e0ca1c806eea9e7d6b0ca1556f08fdffbdfe0b42ed14eeb296ced9cba17f52234abba7c233d2ccf93a00c9a453ef709cd00a5b75697a61586143b6905760ecf7d9c3c2cd397ff3fde4b79c4bf8fd09a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'haf6453e31632802cc507213b906fca318acaa1b6ba9e48879133bf3686800f15d110628b20aac64c91fd22ddfb33ec1b7f6b5f217d931c067d47ab2a44d6ae5dbe02f6cb4ba7acadf33eeb9479d92cd72e88389d9f20b36d9c3fdbfa8fe753b4ee20c17c5225d54abd7504e40d253a51d06e15dfeab7b30730fa28e7de8f281ad5403c37e3ddb018b01f37136c44e0c654e9d9c41a6ec8ca35c8329e84eea8095df9ac82c67e4c2e0811087d81396ff93963897507ef02a80120565efae83835135bcf8b810960224b525e6ebdef9a3406e33b8464f188447045e29ab80b960241aaad43cd3cc9c5ea86eb516f54930246c6ee8761010d70fa506df6a89f6529;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h54789d1146b9da5a21ffa489c5d5f11082d0019e0d59db1fa80759c325634766078b938153f8cb6f42a4ef45c8b8306dede5764cdd5bac54cdb131bc2ea51204e292173cb7e0717cebba06fc0435f60de18550d9f42bbc1575020b276b44f0fd4f717028990417591f75126b2119480e0107a8e2b5c5a4561d71a35a2c681d9710f26226420cd09adab012517b1a03db5242f579bcf79b6cc77a574f3069b7162d905aba86caed34c5ddc954367de7fdb25122345ef0ee68d3a6ec0e417efc19192a94cadebd229f8495e93ecc0a1122f54472ce82f8c49fb04f99ae1c54d4c98279453f9f8487242712b738adb75bd5934359e03a4c364ba571bc37c7faad2d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h31f37e37e40773b8752ea324c9be921015829c36613821eb2b3d24df80730229ec41bfbf5a17c3185c3f0d73c20055760f8a3fa5a8f29e2bcdfabed68d631619a50c3be3907af6750f268366cdedb85f52bf6b59f3b98a299b2db11d327e06b84c6510738fedca1af14b07aa298fb4314e58794ca84af732211c15cc121f29416db342249ea5979a03e28ded8b0f5d74efef1308021b690f9d99ffead8841462233f672cb24c5b0554fa48de44d67e6c5e020987c1d14f730c10e9e7aa90aa9609490f78d7bb813ddf77b7527ca8139ded104a1e4702115592f9cac6ea926557bb4ba3a80d58d6a678ea41f01242828d4c3bc87a1625074f120a3d2e560b3649;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h73fef105976068afd2fb3b03a2831e1a3c2af86d4125090beb0c9dba8a4bd3e46554444ecf18162c11f68f20ddf344fa9817bc86e6191b114111c5fa33fbddae07b3c8fa5afa20ccca03d66fa1a730d0ae0c10d63897bd761611780d9862fd7dea5e578a8ae9a7b3b5910bf3a61f3bfe8f3c0b0e7699a209d5c3efbc1ed937ec51b7b6d1c29950b12a1a80dd644b656b381ba5edd586263069be712646235f1ade6b52ce98f790da49bde763d0b2995de3584bfc51ce6fe22c40ed0b9c817a1de97d704fb0a46567b609abc13bc70395d7a348e35512f455eb8b9ccc510cc2999da71c5ecc6a49aa5373861d125eb4b705adfdb9811fe44e357b7d8e21121f9a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'habf3c00b2a34b2a73796f547148e080ce3f9a971db67600272916efee6afee8173fa5d96b2ce8ceb0b671a9e1c4ad07b55d2d4e72bd7de9595e65f841d53c693ae39d921f88b83b89510931f577444af0940b2bb3ee75e879b6dfab83c16966e90ac0d29105be2a84256e2e02a03ee3d1ce569262ef1b91993e0caf90b368fc4b2c2a405df11c6b00013b3f3b2704b927eec04164b6c71ed7cfe02ad521815b1d50751a6871e5344a6a67b433f55c6a56515a97f8c51e8c50bdcb262fae985dc843fac2a9da2c9f13601914a6bb13fc82e4b9e04b17d50b84ee122bb20253848fc735cd5314ce5c9f69dc254f7b8c8817cd8bd59c7905fab2d08a81c7ee16258;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h502954f7268ef5322f2809b7ca7adc6dae0081f34ecaed528933331ca2cbba83c1f4f5d37ab3cfe82f2742cc9ae84d53f67c8e78ff4b5d53619d9c7395dd221ae3403017068b54027192b5fe21044407d2b52bd873f2bcf80db457db758b369d326f85d96059380f1c816065cebab31342bb13e56d584be270b693682c49c9079d4928a1691b2c7980f7a5d712df807fbe872424d80c0484d07cf111b1e36b9c1472fe18801642574dd6c15c3dd4096c5fe76964366efbf820a9f8644d7c3fe112fa72edd513119715005e4d7f39df1b09a7396c212bae2026bab2acd0a3c21c30f7aa4faf2bfbc5ef93c4d09e27b44b112a67afce4f448a2e37fe86abb839d3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hce763659d158affa43caf79fad6862e2c4c4f277d975add5aa6795c9f448f3ae0795d98553d85975a373aa21e0bd3bb65ed9cb3ba01ac8c23fd97ff233685c37ee17d78d1d98f9df48146d026f8fbc22de2b29883eafa4752e7d5341e68040c68bf19bebf7ae256dfdee756a97c04d0474e4bd463611e1b7477e8397e760b5d8f1da095e3e8afe70450ef6ab61593353b8693328b873df8d91bed9850366b933510c6834e72f04f117f630c8da01ce11ebb79360dc9b62655b338fdb38f543df968c84f50b7c2c73646b537e99960e70c121747d42cbccbc37030eb732c778e0ce6c90e446107a53636b429c48a3d67be9aab91673413b2f2983de0175ed3a4a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h6198dc8b447892bc3a55f0b23a10e982fba6d187bc21c7e6f6cad46a1de8b64d0aba30f3a956f5f1143ad9d4132a0dd07e42c5fce4a935d64554e4da97596056d2aa578ac85e95af7b03fd5d1c98a23f518ae85360184cf13be0d3faa4728cc7b1366696e0baeef79a60c1965a8e0b2b6a30e64d77aa598d678594783ea2c26186c620d6538c19daf89f421a56572698947a1e7eb1fffe34ade5570fb8227ef857ce4ea0f28cf4c5c6087db9527913adc8f2653c16ee1c84fe8644424f40ab9527e57b3d1911c43ecc8f05103a0c4216635d4d7fe821de9aa6f63ed43dc2d0ef4fd2231572567006a947c0ce1c5897ee833ded99046efa13be15b13789946539;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h3631b1c1d1ef404def660415d4a33039540b4f57e978501e615503c310d8e4596d6f93ec9c6ca95626dde010522b0cc625a29d3496932391cd3cab1a4fa5d8aaaf1fc463f4f4f0c32c1cc619a931f5ee58ab783e2ab5eaf9956ae4d2a73e70e3570793f72640f80cbf1286db0b15357b9c5a5f7484d19b2faaaac6aac52d8cc1ba26a95b5b5521e2aacd5445983ab7c93835f72da85d6b49630b3467145ce0e80c2ed3e53dcbb5d73d339f1be35636538c79b9ecf785cc73eb6916617e66a62560d345bfffc693406d1728f53bf655a0bf50af254c33d0d507336841ec3ea1fab0efbfb4e6a5330d51b32575cf8388fc8cdcc80f46977f9b587045483726f00f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'ha405efd68c8963f6f2c5235dad659ffe656c232a792339e21099a0b850b891538e0976ef74d72b194b03ade0cdc2cb0a2643aeab5d5973c31b17a4c241e7082680c5b70d12857c160605733c7681b7ef01053e5ff32eb40661c1b83b36297271fdb0fb48037c053833eb041e6cf7f78b11961c1922e08152b40411006e9fe4b88620a03353e34eebf4f61330223d1ecfcfd3ccdfe195a519ebc27e971d3962d53b9e099107b3b206a292b7844a6f748e12362326cee7eddb972f15e1d7c55283fca8738efd854f244124284aaf7295ecc0df18f5f17590e80ec26cbb59e7b2cf2aca2f818ec400a025037f6577b5c81920b7b060f6329faaa52e6cce3001ba80;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h18383edcea9bb58343bfc5aad6459dd7dd190ada5bc1ef165be5eec16d6a4f0dfc5a67bb77d42363db9f09625d86bfa28d2b475d6c5431159a91a55474ab0325fdfb9ab45653c40c1809015fa489b77b5ed7e1343a191b61ac262a731bb59aff4706866112681d87c44a3fc8059058ca579784299dcb96c7ff04ee4c7972252d20ee8514073bceb0a82867863468d991859c2377ad1a1b20629fae0884ed2aad9886a6afe92229ea8dcc574947fcb632a3dd3cbebb3af59789189644f46a23b631a3cfc34ea961ea9adc6ca4844defab87bbb505c585d29a96a00e626820d9f85864aba1ed45c3acf61bd9221fd2e4a05475f722af2464e638f0c6e20db560b3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'ha599c06d484ae0c8fed241c75b0b57c3043fc7265cc50cc4ba65532473904261fddf0389e059dcb9988d2211d594719ce17eb7e462c341ae78f1c8cb4b677cbaffcd8c7e7a7f7b787b5d873374c1430f9d37c313020a6c855eecc7ecd829a2ca46c9825eead38f3c37ed8213a3c0d25c3a74e0726613915b26ab60a41858e24546665f2b96aa710de73652bf0f4e9a24832397270f80a3334c7e911fab3a444cbd9adc24a95cc03ea4a42035c6bb2f118ea6faafab4d86e2d929c2f3224b47624f7eb8ac2d3a920da10ee5831369eae9aa8cf89048deebb31402dc005b7561fcaa37c77daf9c8f1bd741a02550fd42a087741dbcca7319c36ce9d3a2e6bda89d;
        #1
        $finish();
    end
endmodule
