module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19);
    reg [255:0] src0;
    reg [255:0] src1;
    reg [255:0] src2;
    reg [255:0] src3;
    reg [255:0] src4;
    reg [255:0] src5;
    reg [255:0] src6;
    reg [255:0] src7;
    reg [255:0] src8;
    reg [255:0] src9;
    reg [255:0] src10;
    reg [255:0] src11;
    compressor2_1_256_12 compressor2_1_256_12(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19));
    initial begin
        src0 <= 256'h0;
        src1 <= 256'h0;
        src2 <= 256'h0;
        src3 <= 256'h0;
        src4 <= 256'h0;
        src5 <= 256'h0;
        src6 <= 256'h0;
        src7 <= 256'h0;
        src8 <= 256'h0;
        src9 <= 256'h0;
        src10 <= 256'h0;
        src11 <= 256'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
    end
endmodule
module compressor2_1_256_12(
    input [255:0]src0,
    input [255:0]src1,
    input [255:0]src2,
    input [255:0]src3,
    input [255:0]src4,
    input [255:0]src5,
    input [255:0]src6,
    input [255:0]src7,
    input [255:0]src8,
    input [255:0]src9,
    input [255:0]src10,
    input [255:0]src11,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19);

    wire [1:0] comp_out0;
    wire [0:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [0:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [0:0] comp_out19;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19)
    );
    rowadder2_1_20 rowadder2_1inst(
        .src0({comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], 1'h0, comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], 1'h0, comp_out0[1]}),
        .dst0({dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [255:0] src0,
      input wire [255:0] src1,
      input wire [255:0] src2,
      input wire [255:0] src3,
      input wire [255:0] src4,
      input wire [255:0] src5,
      input wire [255:0] src6,
      input wire [255:0] src7,
      input wire [255:0] src8,
      input wire [255:0] src9,
      input wire [255:0] src10,
      input wire [255:0] src11,
      output wire [1:0] dst0,
      output wire [0:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [0:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [0:0] dst19);

   wire [255:0] stage0_0;
   wire [255:0] stage0_1;
   wire [255:0] stage0_2;
   wire [255:0] stage0_3;
   wire [255:0] stage0_4;
   wire [255:0] stage0_5;
   wire [255:0] stage0_6;
   wire [255:0] stage0_7;
   wire [255:0] stage0_8;
   wire [255:0] stage0_9;
   wire [255:0] stage0_10;
   wire [255:0] stage0_11;
   wire [47:0] stage1_0;
   wire [89:0] stage1_1;
   wire [84:0] stage1_2;
   wire [96:0] stage1_3;
   wire [126:0] stage1_4;
   wire [128:0] stage1_5;
   wire [88:0] stage1_6;
   wire [90:0] stage1_7;
   wire [154:0] stage1_8;
   wire [119:0] stage1_9;
   wire [121:0] stage1_10;
   wire [82:0] stage1_11;
   wire [71:0] stage1_12;
   wire [41:0] stage1_13;
   wire [18:0] stage2_0;
   wire [24:0] stage2_1;
   wire [25:0] stage2_2;
   wire [41:0] stage2_3;
   wire [49:0] stage2_4;
   wire [41:0] stage2_5;
   wire [53:0] stage2_6;
   wire [47:0] stage2_7;
   wire [70:0] stage2_8;
   wire [42:0] stage2_9;
   wire [49:0] stage2_10;
   wire [46:0] stage2_11;
   wire [35:0] stage2_12;
   wire [35:0] stage2_13;
   wire [15:0] stage2_14;
   wire [4:0] stage2_15;
   wire [18:0] stage3_0;
   wire [4:0] stage3_1;
   wire [12:0] stage3_2;
   wire [10:0] stage3_3;
   wire [18:0] stage3_4;
   wire [17:0] stage3_5;
   wire [22:0] stage3_6;
   wire [20:0] stage3_7;
   wire [23:0] stage3_8;
   wire [27:0] stage3_9;
   wire [19:0] stage3_10;
   wire [21:0] stage3_11;
   wire [18:0] stage3_12;
   wire [12:0] stage3_13;
   wire [11:0] stage3_14;
   wire [12:0] stage3_15;
   wire [2:0] stage3_16;
   wire [13:0] stage4_0;
   wire [5:0] stage4_1;
   wire [3:0] stage4_2;
   wire [3:0] stage4_3;
   wire [6:0] stage4_4;
   wire [6:0] stage4_5;
   wire [12:0] stage4_6;
   wire [6:0] stage4_7;
   wire [11:0] stage4_8;
   wire [10:0] stage4_9;
   wire [8:0] stage4_10;
   wire [11:0] stage4_11;
   wire [8:0] stage4_12;
   wire [8:0] stage4_13;
   wire [4:0] stage4_14;
   wire [11:0] stage4_15;
   wire [3:0] stage4_16;
   wire [1:0] stage4_17;
   wire [5:0] stage5_0;
   wire [1:0] stage5_1;
   wire [3:0] stage5_2;
   wire [1:0] stage5_3;
   wire [4:0] stage5_4;
   wire [1:0] stage5_5;
   wire [4:0] stage5_6;
   wire [2:0] stage5_7;
   wire [3:0] stage5_8;
   wire [5:0] stage5_9;
   wire [4:0] stage5_10;
   wire [2:0] stage5_11;
   wire [3:0] stage5_12;
   wire [5:0] stage5_13;
   wire [5:0] stage5_14;
   wire [1:0] stage5_15;
   wire [5:0] stage5_16;
   wire [3:0] stage5_17;
   wire [1:0] stage6_0;
   wire [0:0] stage6_1;
   wire [1:0] stage6_2;
   wire [1:0] stage6_3;
   wire [1:0] stage6_4;
   wire [1:0] stage6_5;
   wire [0:0] stage6_6;
   wire [1:0] stage6_7;
   wire [1:0] stage6_8;
   wire [1:0] stage6_9;
   wire [1:0] stage6_10;
   wire [1:0] stage6_11;
   wire [1:0] stage6_12;
   wire [1:0] stage6_13;
   wire [1:0] stage6_14;
   wire [1:0] stage6_15;
   wire [1:0] stage6_16;
   wire [1:0] stage6_17;
   wire [1:0] stage6_18;
   wire [0:0] stage6_19;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage6_0;
   assign dst1 = stage6_1;
   assign dst2 = stage6_2;
   assign dst3 = stage6_3;
   assign dst4 = stage6_4;
   assign dst5 = stage6_5;
   assign dst6 = stage6_6;
   assign dst7 = stage6_7;
   assign dst8 = stage6_8;
   assign dst9 = stage6_9;
   assign dst10 = stage6_10;
   assign dst11 = stage6_11;
   assign dst12 = stage6_12;
   assign dst13 = stage6_13;
   assign dst14 = stage6_14;
   assign dst15 = stage6_15;
   assign dst16 = stage6_16;
   assign dst17 = stage6_17;
   assign dst18 = stage6_18;
   assign dst19 = stage6_19;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc1163_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12]},
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[2]},
      {stage0_3[4]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc1163_5 gpc3 (
      {stage0_0[13], stage0_0[14], stage0_0[15]},
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[3]},
      {stage0_3[5]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc1163_5 gpc4 (
      {stage0_0[16], stage0_0[17], stage0_0[18]},
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[4]},
      {stage0_3[6]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc1163_5 gpc5 (
      {stage0_0[19], stage0_0[20], stage0_0[21]},
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_2[5]},
      {stage0_3[7]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc1163_5 gpc6 (
      {stage0_0[22], stage0_0[23], stage0_0[24]},
      {stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_2[6]},
      {stage0_3[8]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30]},
      {stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34], stage0_0[35], stage0_0[36]},
      {stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_0[37], stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42]},
      {stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc606_5 gpc10 (
      {stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48]},
      {stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc606_5 gpc11 (
      {stage0_0[49], stage0_0[50], stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54]},
      {stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc606_5 gpc12 (
      {stage0_0[55], stage0_0[56], stage0_0[57], stage0_0[58], stage0_0[59], stage0_0[60]},
      {stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc606_5 gpc13 (
      {stage0_0[61], stage0_0[62], stage0_0[63], stage0_0[64], stage0_0[65], stage0_0[66]},
      {stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc606_5 gpc14 (
      {stage0_0[67], stage0_0[68], stage0_0[69], stage0_0[70], stage0_0[71], stage0_0[72]},
      {stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc606_5 gpc15 (
      {stage0_0[73], stage0_0[74], stage0_0[75], stage0_0[76], stage0_0[77], stage0_0[78]},
      {stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc606_5 gpc16 (
      {stage0_0[79], stage0_0[80], stage0_0[81], stage0_0[82], stage0_0[83], stage0_0[84]},
      {stage0_2[61], stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc606_5 gpc17 (
      {stage0_0[85], stage0_0[86], stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90]},
      {stage0_2[67], stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc606_5 gpc18 (
      {stage0_0[91], stage0_0[92], stage0_0[93], stage0_0[94], stage0_0[95], stage0_0[96]},
      {stage0_2[73], stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc606_5 gpc19 (
      {stage0_0[97], stage0_0[98], stage0_0[99], stage0_0[100], stage0_0[101], stage0_0[102]},
      {stage0_2[79], stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc606_5 gpc20 (
      {stage0_0[103], stage0_0[104], stage0_0[105], stage0_0[106], stage0_0[107], stage0_0[108]},
      {stage0_2[85], stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc606_5 gpc21 (
      {stage0_0[109], stage0_0[110], stage0_0[111], stage0_0[112], stage0_0[113], stage0_0[114]},
      {stage0_2[91], stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc606_5 gpc22 (
      {stage0_0[115], stage0_0[116], stage0_0[117], stage0_0[118], stage0_0[119], stage0_0[120]},
      {stage0_2[97], stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc606_5 gpc23 (
      {stage0_0[121], stage0_0[122], stage0_0[123], stage0_0[124], stage0_0[125], stage0_0[126]},
      {stage0_2[103], stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108]},
      {stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc606_5 gpc24 (
      {stage0_0[127], stage0_0[128], stage0_0[129], stage0_0[130], stage0_0[131], stage0_0[132]},
      {stage0_2[109], stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114]},
      {stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc606_5 gpc25 (
      {stage0_0[133], stage0_0[134], stage0_0[135], stage0_0[136], stage0_0[137], stage0_0[138]},
      {stage0_2[115], stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120]},
      {stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc606_5 gpc26 (
      {stage0_0[139], stage0_0[140], stage0_0[141], stage0_0[142], stage0_0[143], stage0_0[144]},
      {stage0_2[121], stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126]},
      {stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc606_5 gpc27 (
      {stage0_0[145], stage0_0[146], stage0_0[147], stage0_0[148], stage0_0[149], stage0_0[150]},
      {stage0_2[127], stage0_2[128], stage0_2[129], stage0_2[130], stage0_2[131], stage0_2[132]},
      {stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc606_5 gpc28 (
      {stage0_0[151], stage0_0[152], stage0_0[153], stage0_0[154], stage0_0[155], stage0_0[156]},
      {stage0_2[133], stage0_2[134], stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138]},
      {stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc606_5 gpc29 (
      {stage0_0[157], stage0_0[158], stage0_0[159], stage0_0[160], stage0_0[161], stage0_0[162]},
      {stage0_2[139], stage0_2[140], stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144]},
      {stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc606_5 gpc30 (
      {stage0_0[163], stage0_0[164], stage0_0[165], stage0_0[166], stage0_0[167], stage0_0[168]},
      {stage0_2[145], stage0_2[146], stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150]},
      {stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc606_5 gpc31 (
      {stage0_0[169], stage0_0[170], stage0_0[171], stage0_0[172], stage0_0[173], stage0_0[174]},
      {stage0_2[151], stage0_2[152], stage0_2[153], stage0_2[154], stage0_2[155], stage0_2[156]},
      {stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc606_5 gpc32 (
      {stage0_0[175], stage0_0[176], stage0_0[177], stage0_0[178], stage0_0[179], stage0_0[180]},
      {stage0_2[157], stage0_2[158], stage0_2[159], stage0_2[160], stage0_2[161], stage0_2[162]},
      {stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc606_5 gpc33 (
      {stage0_0[181], stage0_0[182], stage0_0[183], stage0_0[184], stage0_0[185], stage0_0[186]},
      {stage0_2[163], stage0_2[164], stage0_2[165], stage0_2[166], stage0_2[167], stage0_2[168]},
      {stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc606_5 gpc34 (
      {stage0_0[187], stage0_0[188], stage0_0[189], stage0_0[190], stage0_0[191], stage0_0[192]},
      {stage0_2[169], stage0_2[170], stage0_2[171], stage0_2[172], stage0_2[173], stage0_2[174]},
      {stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc606_5 gpc35 (
      {stage0_0[193], stage0_0[194], stage0_0[195], stage0_0[196], stage0_0[197], stage0_0[198]},
      {stage0_2[175], stage0_2[176], stage0_2[177], stage0_2[178], stage0_2[179], stage0_2[180]},
      {stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc606_5 gpc36 (
      {stage0_0[199], stage0_0[200], stage0_0[201], stage0_0[202], stage0_0[203], stage0_0[204]},
      {stage0_2[181], stage0_2[182], stage0_2[183], stage0_2[184], stage0_2[185], stage0_2[186]},
      {stage1_4[36],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc606_5 gpc37 (
      {stage0_0[205], stage0_0[206], stage0_0[207], stage0_0[208], stage0_0[209], stage0_0[210]},
      {stage0_2[187], stage0_2[188], stage0_2[189], stage0_2[190], stage0_2[191], stage0_2[192]},
      {stage1_4[37],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc606_5 gpc38 (
      {stage0_0[211], stage0_0[212], stage0_0[213], stage0_0[214], stage0_0[215], stage0_0[216]},
      {stage0_2[193], stage0_2[194], stage0_2[195], stage0_2[196], stage0_2[197], stage0_2[198]},
      {stage1_4[38],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc606_5 gpc39 (
      {stage0_0[217], stage0_0[218], stage0_0[219], stage0_0[220], stage0_0[221], stage0_0[222]},
      {stage0_2[199], stage0_2[200], stage0_2[201], stage0_2[202], stage0_2[203], stage0_2[204]},
      {stage1_4[39],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc606_5 gpc40 (
      {stage0_0[223], stage0_0[224], stage0_0[225], stage0_0[226], stage0_0[227], stage0_0[228]},
      {stage0_2[205], stage0_2[206], stage0_2[207], stage0_2[208], stage0_2[209], stage0_2[210]},
      {stage1_4[40],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc606_5 gpc41 (
      {stage0_0[229], stage0_0[230], stage0_0[231], stage0_0[232], stage0_0[233], stage0_0[234]},
      {stage0_2[211], stage0_2[212], stage0_2[213], stage0_2[214], stage0_2[215], stage0_2[216]},
      {stage1_4[41],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc606_5 gpc42 (
      {stage0_0[235], stage0_0[236], stage0_0[237], stage0_0[238], stage0_0[239], stage0_0[240]},
      {stage0_2[217], stage0_2[218], stage0_2[219], stage0_2[220], stage0_2[221], stage0_2[222]},
      {stage1_4[42],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc606_5 gpc43 (
      {stage0_0[241], stage0_0[242], stage0_0[243], stage0_0[244], stage0_0[245], stage0_0[246]},
      {stage0_2[223], stage0_2[224], stage0_2[225], stage0_2[226], stage0_2[227], stage0_2[228]},
      {stage1_4[43],stage1_3[43],stage1_2[43],stage1_1[43],stage1_0[43]}
   );
   gpc606_5 gpc44 (
      {stage0_0[247], stage0_0[248], stage0_0[249], stage0_0[250], stage0_0[251], stage0_0[252]},
      {stage0_2[229], stage0_2[230], stage0_2[231], stage0_2[232], stage0_2[233], stage0_2[234]},
      {stage1_4[44],stage1_3[44],stage1_2[44],stage1_1[44],stage1_0[44]}
   );
   gpc606_5 gpc45 (
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12], stage0_3[13], stage0_3[14]},
      {stage1_5[0],stage1_4[45],stage1_3[45],stage1_2[45],stage1_1[45]}
   );
   gpc606_5 gpc46 (
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19], stage0_3[20]},
      {stage1_5[1],stage1_4[46],stage1_3[46],stage1_2[46],stage1_1[46]}
   );
   gpc606_5 gpc47 (
      {stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26]},
      {stage1_5[2],stage1_4[47],stage1_3[47],stage1_2[47],stage1_1[47]}
   );
   gpc606_5 gpc48 (
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59]},
      {stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32]},
      {stage1_5[3],stage1_4[48],stage1_3[48],stage1_2[48],stage1_1[48]}
   );
   gpc606_5 gpc49 (
      {stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65]},
      {stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38]},
      {stage1_5[4],stage1_4[49],stage1_3[49],stage1_2[49],stage1_1[49]}
   );
   gpc606_5 gpc50 (
      {stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71]},
      {stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44]},
      {stage1_5[5],stage1_4[50],stage1_3[50],stage1_2[50],stage1_1[50]}
   );
   gpc606_5 gpc51 (
      {stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77]},
      {stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50]},
      {stage1_5[6],stage1_4[51],stage1_3[51],stage1_2[51],stage1_1[51]}
   );
   gpc606_5 gpc52 (
      {stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83]},
      {stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56]},
      {stage1_5[7],stage1_4[52],stage1_3[52],stage1_2[52],stage1_1[52]}
   );
   gpc606_5 gpc53 (
      {stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89]},
      {stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62]},
      {stage1_5[8],stage1_4[53],stage1_3[53],stage1_2[53],stage1_1[53]}
   );
   gpc606_5 gpc54 (
      {stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95]},
      {stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68]},
      {stage1_5[9],stage1_4[54],stage1_3[54],stage1_2[54],stage1_1[54]}
   );
   gpc606_5 gpc55 (
      {stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101]},
      {stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74]},
      {stage1_5[10],stage1_4[55],stage1_3[55],stage1_2[55],stage1_1[55]}
   );
   gpc606_5 gpc56 (
      {stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107]},
      {stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80]},
      {stage1_5[11],stage1_4[56],stage1_3[56],stage1_2[56],stage1_1[56]}
   );
   gpc606_5 gpc57 (
      {stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113]},
      {stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86]},
      {stage1_5[12],stage1_4[57],stage1_3[57],stage1_2[57],stage1_1[57]}
   );
   gpc606_5 gpc58 (
      {stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119]},
      {stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92]},
      {stage1_5[13],stage1_4[58],stage1_3[58],stage1_2[58],stage1_1[58]}
   );
   gpc606_5 gpc59 (
      {stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125]},
      {stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98]},
      {stage1_5[14],stage1_4[59],stage1_3[59],stage1_2[59],stage1_1[59]}
   );
   gpc606_5 gpc60 (
      {stage0_1[126], stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131]},
      {stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104]},
      {stage1_5[15],stage1_4[60],stage1_3[60],stage1_2[60],stage1_1[60]}
   );
   gpc606_5 gpc61 (
      {stage0_1[132], stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137]},
      {stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110]},
      {stage1_5[16],stage1_4[61],stage1_3[61],stage1_2[61],stage1_1[61]}
   );
   gpc606_5 gpc62 (
      {stage0_1[138], stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143]},
      {stage0_3[111], stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116]},
      {stage1_5[17],stage1_4[62],stage1_3[62],stage1_2[62],stage1_1[62]}
   );
   gpc606_5 gpc63 (
      {stage0_1[144], stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149]},
      {stage0_3[117], stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121], stage0_3[122]},
      {stage1_5[18],stage1_4[63],stage1_3[63],stage1_2[63],stage1_1[63]}
   );
   gpc606_5 gpc64 (
      {stage0_1[150], stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155]},
      {stage0_3[123], stage0_3[124], stage0_3[125], stage0_3[126], stage0_3[127], stage0_3[128]},
      {stage1_5[19],stage1_4[64],stage1_3[64],stage1_2[64],stage1_1[64]}
   );
   gpc606_5 gpc65 (
      {stage0_1[156], stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161]},
      {stage0_3[129], stage0_3[130], stage0_3[131], stage0_3[132], stage0_3[133], stage0_3[134]},
      {stage1_5[20],stage1_4[65],stage1_3[65],stage1_2[65],stage1_1[65]}
   );
   gpc606_5 gpc66 (
      {stage0_1[162], stage0_1[163], stage0_1[164], stage0_1[165], stage0_1[166], stage0_1[167]},
      {stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138], stage0_3[139], stage0_3[140]},
      {stage1_5[21],stage1_4[66],stage1_3[66],stage1_2[66],stage1_1[66]}
   );
   gpc606_5 gpc67 (
      {stage0_1[168], stage0_1[169], stage0_1[170], stage0_1[171], stage0_1[172], stage0_1[173]},
      {stage0_3[141], stage0_3[142], stage0_3[143], stage0_3[144], stage0_3[145], stage0_3[146]},
      {stage1_5[22],stage1_4[67],stage1_3[67],stage1_2[67],stage1_1[67]}
   );
   gpc606_5 gpc68 (
      {stage0_1[174], stage0_1[175], stage0_1[176], stage0_1[177], stage0_1[178], stage0_1[179]},
      {stage0_3[147], stage0_3[148], stage0_3[149], stage0_3[150], stage0_3[151], stage0_3[152]},
      {stage1_5[23],stage1_4[68],stage1_3[68],stage1_2[68],stage1_1[68]}
   );
   gpc606_5 gpc69 (
      {stage0_1[180], stage0_1[181], stage0_1[182], stage0_1[183], stage0_1[184], stage0_1[185]},
      {stage0_3[153], stage0_3[154], stage0_3[155], stage0_3[156], stage0_3[157], stage0_3[158]},
      {stage1_5[24],stage1_4[69],stage1_3[69],stage1_2[69],stage1_1[69]}
   );
   gpc606_5 gpc70 (
      {stage0_1[186], stage0_1[187], stage0_1[188], stage0_1[189], stage0_1[190], stage0_1[191]},
      {stage0_3[159], stage0_3[160], stage0_3[161], stage0_3[162], stage0_3[163], stage0_3[164]},
      {stage1_5[25],stage1_4[70],stage1_3[70],stage1_2[70],stage1_1[70]}
   );
   gpc606_5 gpc71 (
      {stage0_1[192], stage0_1[193], stage0_1[194], stage0_1[195], stage0_1[196], stage0_1[197]},
      {stage0_3[165], stage0_3[166], stage0_3[167], stage0_3[168], stage0_3[169], stage0_3[170]},
      {stage1_5[26],stage1_4[71],stage1_3[71],stage1_2[71],stage1_1[71]}
   );
   gpc606_5 gpc72 (
      {stage0_1[198], stage0_1[199], stage0_1[200], stage0_1[201], stage0_1[202], stage0_1[203]},
      {stage0_3[171], stage0_3[172], stage0_3[173], stage0_3[174], stage0_3[175], stage0_3[176]},
      {stage1_5[27],stage1_4[72],stage1_3[72],stage1_2[72],stage1_1[72]}
   );
   gpc606_5 gpc73 (
      {stage0_1[204], stage0_1[205], stage0_1[206], stage0_1[207], stage0_1[208], stage0_1[209]},
      {stage0_3[177], stage0_3[178], stage0_3[179], stage0_3[180], stage0_3[181], stage0_3[182]},
      {stage1_5[28],stage1_4[73],stage1_3[73],stage1_2[73],stage1_1[73]}
   );
   gpc606_5 gpc74 (
      {stage0_1[210], stage0_1[211], stage0_1[212], stage0_1[213], stage0_1[214], stage0_1[215]},
      {stage0_3[183], stage0_3[184], stage0_3[185], stage0_3[186], stage0_3[187], stage0_3[188]},
      {stage1_5[29],stage1_4[74],stage1_3[74],stage1_2[74],stage1_1[74]}
   );
   gpc606_5 gpc75 (
      {stage0_1[216], stage0_1[217], stage0_1[218], stage0_1[219], stage0_1[220], stage0_1[221]},
      {stage0_3[189], stage0_3[190], stage0_3[191], stage0_3[192], stage0_3[193], stage0_3[194]},
      {stage1_5[30],stage1_4[75],stage1_3[75],stage1_2[75],stage1_1[75]}
   );
   gpc606_5 gpc76 (
      {stage0_1[222], stage0_1[223], stage0_1[224], stage0_1[225], stage0_1[226], stage0_1[227]},
      {stage0_3[195], stage0_3[196], stage0_3[197], stage0_3[198], stage0_3[199], stage0_3[200]},
      {stage1_5[31],stage1_4[76],stage1_3[76],stage1_2[76],stage1_1[76]}
   );
   gpc606_5 gpc77 (
      {stage0_1[228], stage0_1[229], stage0_1[230], stage0_1[231], stage0_1[232], stage0_1[233]},
      {stage0_3[201], stage0_3[202], stage0_3[203], stage0_3[204], stage0_3[205], stage0_3[206]},
      {stage1_5[32],stage1_4[77],stage1_3[77],stage1_2[77],stage1_1[77]}
   );
   gpc606_5 gpc78 (
      {stage0_1[234], stage0_1[235], stage0_1[236], stage0_1[237], stage0_1[238], stage0_1[239]},
      {stage0_3[207], stage0_3[208], stage0_3[209], stage0_3[210], stage0_3[211], stage0_3[212]},
      {stage1_5[33],stage1_4[78],stage1_3[78],stage1_2[78],stage1_1[78]}
   );
   gpc606_5 gpc79 (
      {stage0_1[240], stage0_1[241], stage0_1[242], stage0_1[243], stage0_1[244], stage0_1[245]},
      {stage0_3[213], stage0_3[214], stage0_3[215], stage0_3[216], stage0_3[217], stage0_3[218]},
      {stage1_5[34],stage1_4[79],stage1_3[79],stage1_2[79],stage1_1[79]}
   );
   gpc615_5 gpc80 (
      {stage0_2[235], stage0_2[236], stage0_2[237], stage0_2[238], stage0_2[239]},
      {stage0_3[219]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[35],stage1_4[80],stage1_3[80],stage1_2[80]}
   );
   gpc615_5 gpc81 (
      {stage0_2[240], stage0_2[241], stage0_2[242], stage0_2[243], stage0_2[244]},
      {stage0_3[220]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[36],stage1_4[81],stage1_3[81],stage1_2[81]}
   );
   gpc615_5 gpc82 (
      {stage0_2[245], stage0_2[246], stage0_2[247], stage0_2[248], stage0_2[249]},
      {stage0_3[221]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[37],stage1_4[82],stage1_3[82],stage1_2[82]}
   );
   gpc615_5 gpc83 (
      {stage0_2[250], stage0_2[251], stage0_2[252], stage0_2[253], stage0_2[254]},
      {stage0_3[222]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[38],stage1_4[83],stage1_3[83],stage1_2[83]}
   );
   gpc615_5 gpc84 (
      {stage0_3[223], stage0_3[224], stage0_3[225], stage0_3[226], stage0_3[227]},
      {stage0_4[24]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[4],stage1_5[39],stage1_4[84],stage1_3[84]}
   );
   gpc615_5 gpc85 (
      {stage0_3[228], stage0_3[229], stage0_3[230], stage0_3[231], stage0_3[232]},
      {stage0_4[25]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[5],stage1_5[40],stage1_4[85],stage1_3[85]}
   );
   gpc615_5 gpc86 (
      {stage0_3[233], stage0_3[234], stage0_3[235], stage0_3[236], stage0_3[237]},
      {stage0_4[26]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[6],stage1_5[41],stage1_4[86],stage1_3[86]}
   );
   gpc615_5 gpc87 (
      {stage0_3[238], stage0_3[239], stage0_3[240], stage0_3[241], stage0_3[242]},
      {stage0_4[27]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[7],stage1_5[42],stage1_4[87],stage1_3[87]}
   );
   gpc615_5 gpc88 (
      {stage0_3[243], stage0_3[244], stage0_3[245], stage0_3[246], stage0_3[247]},
      {stage0_4[28]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[8],stage1_5[43],stage1_4[88],stage1_3[88]}
   );
   gpc606_5 gpc89 (
      {stage0_4[29], stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[5],stage1_6[9],stage1_5[44],stage1_4[89]}
   );
   gpc606_5 gpc90 (
      {stage0_4[35], stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[6],stage1_6[10],stage1_5[45],stage1_4[90]}
   );
   gpc606_5 gpc91 (
      {stage0_4[41], stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[7],stage1_6[11],stage1_5[46],stage1_4[91]}
   );
   gpc606_5 gpc92 (
      {stage0_4[47], stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[8],stage1_6[12],stage1_5[47],stage1_4[92]}
   );
   gpc606_5 gpc93 (
      {stage0_4[53], stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[9],stage1_6[13],stage1_5[48],stage1_4[93]}
   );
   gpc606_5 gpc94 (
      {stage0_4[59], stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[10],stage1_6[14],stage1_5[49],stage1_4[94]}
   );
   gpc606_5 gpc95 (
      {stage0_4[65], stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[11],stage1_6[15],stage1_5[50],stage1_4[95]}
   );
   gpc606_5 gpc96 (
      {stage0_4[71], stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[12],stage1_6[16],stage1_5[51],stage1_4[96]}
   );
   gpc606_5 gpc97 (
      {stage0_4[77], stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[13],stage1_6[17],stage1_5[52],stage1_4[97]}
   );
   gpc606_5 gpc98 (
      {stage0_4[83], stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[14],stage1_6[18],stage1_5[53],stage1_4[98]}
   );
   gpc606_5 gpc99 (
      {stage0_4[89], stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[15],stage1_6[19],stage1_5[54],stage1_4[99]}
   );
   gpc606_5 gpc100 (
      {stage0_4[95], stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[16],stage1_6[20],stage1_5[55],stage1_4[100]}
   );
   gpc606_5 gpc101 (
      {stage0_4[101], stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[17],stage1_6[21],stage1_5[56],stage1_4[101]}
   );
   gpc606_5 gpc102 (
      {stage0_4[107], stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[18],stage1_6[22],stage1_5[57],stage1_4[102]}
   );
   gpc606_5 gpc103 (
      {stage0_4[113], stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[19],stage1_6[23],stage1_5[58],stage1_4[103]}
   );
   gpc606_5 gpc104 (
      {stage0_4[119], stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[20],stage1_6[24],stage1_5[59],stage1_4[104]}
   );
   gpc606_5 gpc105 (
      {stage0_4[125], stage0_4[126], stage0_4[127], stage0_4[128], stage0_4[129], stage0_4[130]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[21],stage1_6[25],stage1_5[60],stage1_4[105]}
   );
   gpc606_5 gpc106 (
      {stage0_4[131], stage0_4[132], stage0_4[133], stage0_4[134], stage0_4[135], stage0_4[136]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[22],stage1_6[26],stage1_5[61],stage1_4[106]}
   );
   gpc606_5 gpc107 (
      {stage0_4[137], stage0_4[138], stage0_4[139], stage0_4[140], stage0_4[141], stage0_4[142]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[23],stage1_6[27],stage1_5[62],stage1_4[107]}
   );
   gpc606_5 gpc108 (
      {stage0_4[143], stage0_4[144], stage0_4[145], stage0_4[146], stage0_4[147], stage0_4[148]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[24],stage1_6[28],stage1_5[63],stage1_4[108]}
   );
   gpc606_5 gpc109 (
      {stage0_4[149], stage0_4[150], stage0_4[151], stage0_4[152], stage0_4[153], stage0_4[154]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[25],stage1_6[29],stage1_5[64],stage1_4[109]}
   );
   gpc606_5 gpc110 (
      {stage0_4[155], stage0_4[156], stage0_4[157], stage0_4[158], stage0_4[159], stage0_4[160]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[21],stage1_7[26],stage1_6[30],stage1_5[65],stage1_4[110]}
   );
   gpc606_5 gpc111 (
      {stage0_4[161], stage0_4[162], stage0_4[163], stage0_4[164], stage0_4[165], stage0_4[166]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[22],stage1_7[27],stage1_6[31],stage1_5[66],stage1_4[111]}
   );
   gpc606_5 gpc112 (
      {stage0_4[167], stage0_4[168], stage0_4[169], stage0_4[170], stage0_4[171], stage0_4[172]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[23],stage1_7[28],stage1_6[32],stage1_5[67],stage1_4[112]}
   );
   gpc606_5 gpc113 (
      {stage0_4[173], stage0_4[174], stage0_4[175], stage0_4[176], stage0_4[177], stage0_4[178]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[24],stage1_7[29],stage1_6[33],stage1_5[68],stage1_4[113]}
   );
   gpc606_5 gpc114 (
      {stage0_4[179], stage0_4[180], stage0_4[181], stage0_4[182], stage0_4[183], stage0_4[184]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[25],stage1_7[30],stage1_6[34],stage1_5[69],stage1_4[114]}
   );
   gpc606_5 gpc115 (
      {stage0_4[185], stage0_4[186], stage0_4[187], stage0_4[188], stage0_4[189], stage0_4[190]},
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage1_8[26],stage1_7[31],stage1_6[35],stage1_5[70],stage1_4[115]}
   );
   gpc606_5 gpc116 (
      {stage0_4[191], stage0_4[192], stage0_4[193], stage0_4[194], stage0_4[195], stage0_4[196]},
      {stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167]},
      {stage1_8[27],stage1_7[32],stage1_6[36],stage1_5[71],stage1_4[116]}
   );
   gpc606_5 gpc117 (
      {stage0_4[197], stage0_4[198], stage0_4[199], stage0_4[200], stage0_4[201], stage0_4[202]},
      {stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173]},
      {stage1_8[28],stage1_7[33],stage1_6[37],stage1_5[72],stage1_4[117]}
   );
   gpc606_5 gpc118 (
      {stage0_4[203], stage0_4[204], stage0_4[205], stage0_4[206], stage0_4[207], stage0_4[208]},
      {stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179]},
      {stage1_8[29],stage1_7[34],stage1_6[38],stage1_5[73],stage1_4[118]}
   );
   gpc606_5 gpc119 (
      {stage0_4[209], stage0_4[210], stage0_4[211], stage0_4[212], stage0_4[213], stage0_4[214]},
      {stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184], stage0_6[185]},
      {stage1_8[30],stage1_7[35],stage1_6[39],stage1_5[74],stage1_4[119]}
   );
   gpc606_5 gpc120 (
      {stage0_4[215], stage0_4[216], stage0_4[217], stage0_4[218], stage0_4[219], stage0_4[220]},
      {stage0_6[186], stage0_6[187], stage0_6[188], stage0_6[189], stage0_6[190], stage0_6[191]},
      {stage1_8[31],stage1_7[36],stage1_6[40],stage1_5[75],stage1_4[120]}
   );
   gpc606_5 gpc121 (
      {stage0_4[221], stage0_4[222], stage0_4[223], stage0_4[224], stage0_4[225], stage0_4[226]},
      {stage0_6[192], stage0_6[193], stage0_6[194], stage0_6[195], stage0_6[196], stage0_6[197]},
      {stage1_8[32],stage1_7[37],stage1_6[41],stage1_5[76],stage1_4[121]}
   );
   gpc606_5 gpc122 (
      {stage0_4[227], stage0_4[228], stage0_4[229], stage0_4[230], stage0_4[231], stage0_4[232]},
      {stage0_6[198], stage0_6[199], stage0_6[200], stage0_6[201], stage0_6[202], stage0_6[203]},
      {stage1_8[33],stage1_7[38],stage1_6[42],stage1_5[77],stage1_4[122]}
   );
   gpc606_5 gpc123 (
      {stage0_4[233], stage0_4[234], stage0_4[235], stage0_4[236], stage0_4[237], stage0_4[238]},
      {stage0_6[204], stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208], stage0_6[209]},
      {stage1_8[34],stage1_7[39],stage1_6[43],stage1_5[78],stage1_4[123]}
   );
   gpc606_5 gpc124 (
      {stage0_4[239], stage0_4[240], stage0_4[241], stage0_4[242], stage0_4[243], stage0_4[244]},
      {stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214], stage0_6[215]},
      {stage1_8[35],stage1_7[40],stage1_6[44],stage1_5[79],stage1_4[124]}
   );
   gpc606_5 gpc125 (
      {stage0_4[245], stage0_4[246], stage0_4[247], stage0_4[248], stage0_4[249], stage0_4[250]},
      {stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219], stage0_6[220], stage0_6[221]},
      {stage1_8[36],stage1_7[41],stage1_6[45],stage1_5[80],stage1_4[125]}
   );
   gpc615_5 gpc126 (
      {stage0_4[251], stage0_4[252], stage0_4[253], stage0_4[254], stage0_4[255]},
      {stage0_5[30]},
      {stage0_6[222], stage0_6[223], stage0_6[224], stage0_6[225], stage0_6[226], stage0_6[227]},
      {stage1_8[37],stage1_7[42],stage1_6[46],stage1_5[81],stage1_4[126]}
   );
   gpc606_5 gpc127 (
      {stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35], stage0_5[36]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[38],stage1_7[43],stage1_6[47],stage1_5[82]}
   );
   gpc606_5 gpc128 (
      {stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41], stage0_5[42]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[39],stage1_7[44],stage1_6[48],stage1_5[83]}
   );
   gpc606_5 gpc129 (
      {stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47], stage0_5[48]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[40],stage1_7[45],stage1_6[49],stage1_5[84]}
   );
   gpc606_5 gpc130 (
      {stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53], stage0_5[54]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[41],stage1_7[46],stage1_6[50],stage1_5[85]}
   );
   gpc606_5 gpc131 (
      {stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59], stage0_5[60]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[42],stage1_7[47],stage1_6[51],stage1_5[86]}
   );
   gpc606_5 gpc132 (
      {stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65], stage0_5[66]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[43],stage1_7[48],stage1_6[52],stage1_5[87]}
   );
   gpc606_5 gpc133 (
      {stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71], stage0_5[72]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[44],stage1_7[49],stage1_6[53],stage1_5[88]}
   );
   gpc606_5 gpc134 (
      {stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77], stage0_5[78]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[45],stage1_7[50],stage1_6[54],stage1_5[89]}
   );
   gpc606_5 gpc135 (
      {stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83], stage0_5[84]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[46],stage1_7[51],stage1_6[55],stage1_5[90]}
   );
   gpc606_5 gpc136 (
      {stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89], stage0_5[90]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[47],stage1_7[52],stage1_6[56],stage1_5[91]}
   );
   gpc606_5 gpc137 (
      {stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95], stage0_5[96]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[48],stage1_7[53],stage1_6[57],stage1_5[92]}
   );
   gpc606_5 gpc138 (
      {stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101], stage0_5[102]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[49],stage1_7[54],stage1_6[58],stage1_5[93]}
   );
   gpc606_5 gpc139 (
      {stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107], stage0_5[108]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[50],stage1_7[55],stage1_6[59],stage1_5[94]}
   );
   gpc606_5 gpc140 (
      {stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113], stage0_5[114]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[51],stage1_7[56],stage1_6[60],stage1_5[95]}
   );
   gpc606_5 gpc141 (
      {stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119], stage0_5[120]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[52],stage1_7[57],stage1_6[61],stage1_5[96]}
   );
   gpc606_5 gpc142 (
      {stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125], stage0_5[126]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[53],stage1_7[58],stage1_6[62],stage1_5[97]}
   );
   gpc606_5 gpc143 (
      {stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131], stage0_5[132]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[54],stage1_7[59],stage1_6[63],stage1_5[98]}
   );
   gpc606_5 gpc144 (
      {stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137], stage0_5[138]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[55],stage1_7[60],stage1_6[64],stage1_5[99]}
   );
   gpc606_5 gpc145 (
      {stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143], stage0_5[144]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[56],stage1_7[61],stage1_6[65],stage1_5[100]}
   );
   gpc606_5 gpc146 (
      {stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149], stage0_5[150]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[57],stage1_7[62],stage1_6[66],stage1_5[101]}
   );
   gpc606_5 gpc147 (
      {stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155], stage0_5[156]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[58],stage1_7[63],stage1_6[67],stage1_5[102]}
   );
   gpc606_5 gpc148 (
      {stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161], stage0_5[162]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[59],stage1_7[64],stage1_6[68],stage1_5[103]}
   );
   gpc606_5 gpc149 (
      {stage0_5[163], stage0_5[164], stage0_5[165], stage0_5[166], stage0_5[167], stage0_5[168]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[60],stage1_7[65],stage1_6[69],stage1_5[104]}
   );
   gpc606_5 gpc150 (
      {stage0_5[169], stage0_5[170], stage0_5[171], stage0_5[172], stage0_5[173], stage0_5[174]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[61],stage1_7[66],stage1_6[70],stage1_5[105]}
   );
   gpc606_5 gpc151 (
      {stage0_5[175], stage0_5[176], stage0_5[177], stage0_5[178], stage0_5[179], stage0_5[180]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[62],stage1_7[67],stage1_6[71],stage1_5[106]}
   );
   gpc606_5 gpc152 (
      {stage0_5[181], stage0_5[182], stage0_5[183], stage0_5[184], stage0_5[185], stage0_5[186]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[63],stage1_7[68],stage1_6[72],stage1_5[107]}
   );
   gpc606_5 gpc153 (
      {stage0_5[187], stage0_5[188], stage0_5[189], stage0_5[190], stage0_5[191], stage0_5[192]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[64],stage1_7[69],stage1_6[73],stage1_5[108]}
   );
   gpc606_5 gpc154 (
      {stage0_5[193], stage0_5[194], stage0_5[195], stage0_5[196], stage0_5[197], stage0_5[198]},
      {stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167]},
      {stage1_9[27],stage1_8[65],stage1_7[70],stage1_6[74],stage1_5[109]}
   );
   gpc606_5 gpc155 (
      {stage0_5[199], stage0_5[200], stage0_5[201], stage0_5[202], stage0_5[203], stage0_5[204]},
      {stage0_7[168], stage0_7[169], stage0_7[170], stage0_7[171], stage0_7[172], stage0_7[173]},
      {stage1_9[28],stage1_8[66],stage1_7[71],stage1_6[75],stage1_5[110]}
   );
   gpc606_5 gpc156 (
      {stage0_5[205], stage0_5[206], stage0_5[207], stage0_5[208], stage0_5[209], stage0_5[210]},
      {stage0_7[174], stage0_7[175], stage0_7[176], stage0_7[177], stage0_7[178], stage0_7[179]},
      {stage1_9[29],stage1_8[67],stage1_7[72],stage1_6[76],stage1_5[111]}
   );
   gpc606_5 gpc157 (
      {stage0_5[211], stage0_5[212], stage0_5[213], stage0_5[214], stage0_5[215], stage0_5[216]},
      {stage0_7[180], stage0_7[181], stage0_7[182], stage0_7[183], stage0_7[184], stage0_7[185]},
      {stage1_9[30],stage1_8[68],stage1_7[73],stage1_6[77],stage1_5[112]}
   );
   gpc606_5 gpc158 (
      {stage0_5[217], stage0_5[218], stage0_5[219], stage0_5[220], stage0_5[221], stage0_5[222]},
      {stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189], stage0_7[190], stage0_7[191]},
      {stage1_9[31],stage1_8[69],stage1_7[74],stage1_6[78],stage1_5[113]}
   );
   gpc606_5 gpc159 (
      {stage0_5[223], stage0_5[224], stage0_5[225], stage0_5[226], stage0_5[227], stage0_5[228]},
      {stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195], stage0_7[196], stage0_7[197]},
      {stage1_9[32],stage1_8[70],stage1_7[75],stage1_6[79],stage1_5[114]}
   );
   gpc606_5 gpc160 (
      {stage0_5[229], stage0_5[230], stage0_5[231], stage0_5[232], stage0_5[233], stage0_5[234]},
      {stage0_7[198], stage0_7[199], stage0_7[200], stage0_7[201], stage0_7[202], stage0_7[203]},
      {stage1_9[33],stage1_8[71],stage1_7[76],stage1_6[80],stage1_5[115]}
   );
   gpc615_5 gpc161 (
      {stage0_5[235], stage0_5[236], stage0_5[237], stage0_5[238], stage0_5[239]},
      {stage0_6[228]},
      {stage0_7[204], stage0_7[205], stage0_7[206], stage0_7[207], stage0_7[208], stage0_7[209]},
      {stage1_9[34],stage1_8[72],stage1_7[77],stage1_6[81],stage1_5[116]}
   );
   gpc615_5 gpc162 (
      {stage0_5[240], stage0_5[241], stage0_5[242], stage0_5[243], stage0_5[244]},
      {stage0_6[229]},
      {stage0_7[210], stage0_7[211], stage0_7[212], stage0_7[213], stage0_7[214], stage0_7[215]},
      {stage1_9[35],stage1_8[73],stage1_7[78],stage1_6[82],stage1_5[117]}
   );
   gpc615_5 gpc163 (
      {stage0_6[230], stage0_6[231], stage0_6[232], stage0_6[233], stage0_6[234]},
      {stage0_7[216]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[36],stage1_8[74],stage1_7[79],stage1_6[83]}
   );
   gpc615_5 gpc164 (
      {stage0_6[235], stage0_6[236], stage0_6[237], stage0_6[238], stage0_6[239]},
      {stage0_7[217]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[37],stage1_8[75],stage1_7[80],stage1_6[84]}
   );
   gpc615_5 gpc165 (
      {stage0_6[240], stage0_6[241], stage0_6[242], stage0_6[243], stage0_6[244]},
      {stage0_7[218]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[38],stage1_8[76],stage1_7[81],stage1_6[85]}
   );
   gpc615_5 gpc166 (
      {stage0_6[245], stage0_6[246], stage0_6[247], stage0_6[248], stage0_6[249]},
      {stage0_7[219]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[39],stage1_8[77],stage1_7[82],stage1_6[86]}
   );
   gpc615_5 gpc167 (
      {stage0_6[250], stage0_6[251], stage0_6[252], stage0_6[253], stage0_6[254]},
      {stage0_7[220]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[40],stage1_8[78],stage1_7[83],stage1_6[87]}
   );
   gpc615_5 gpc168 (
      {stage0_7[221], stage0_7[222], stage0_7[223], stage0_7[224], stage0_7[225]},
      {stage0_8[30]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[5],stage1_9[41],stage1_8[79],stage1_7[84]}
   );
   gpc615_5 gpc169 (
      {stage0_7[226], stage0_7[227], stage0_7[228], stage0_7[229], stage0_7[230]},
      {stage0_8[31]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[6],stage1_9[42],stage1_8[80],stage1_7[85]}
   );
   gpc615_5 gpc170 (
      {stage0_7[231], stage0_7[232], stage0_7[233], stage0_7[234], stage0_7[235]},
      {stage0_8[32]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[7],stage1_9[43],stage1_8[81],stage1_7[86]}
   );
   gpc615_5 gpc171 (
      {stage0_7[236], stage0_7[237], stage0_7[238], stage0_7[239], stage0_7[240]},
      {stage0_8[33]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[8],stage1_9[44],stage1_8[82],stage1_7[87]}
   );
   gpc615_5 gpc172 (
      {stage0_7[241], stage0_7[242], stage0_7[243], stage0_7[244], stage0_7[245]},
      {stage0_8[34]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[9],stage1_9[45],stage1_8[83],stage1_7[88]}
   );
   gpc615_5 gpc173 (
      {stage0_7[246], stage0_7[247], stage0_7[248], stage0_7[249], stage0_7[250]},
      {stage0_8[35]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[10],stage1_9[46],stage1_8[84],stage1_7[89]}
   );
   gpc615_5 gpc174 (
      {stage0_7[251], stage0_7[252], stage0_7[253], stage0_7[254], stage0_7[255]},
      {stage0_8[36]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[11],stage1_9[47],stage1_8[85],stage1_7[90]}
   );
   gpc606_5 gpc175 (
      {stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41], stage0_8[42]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[7],stage1_10[12],stage1_9[48],stage1_8[86]}
   );
   gpc606_5 gpc176 (
      {stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47], stage0_8[48]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[8],stage1_10[13],stage1_9[49],stage1_8[87]}
   );
   gpc606_5 gpc177 (
      {stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53], stage0_8[54]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[9],stage1_10[14],stage1_9[50],stage1_8[88]}
   );
   gpc606_5 gpc178 (
      {stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59], stage0_8[60]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[10],stage1_10[15],stage1_9[51],stage1_8[89]}
   );
   gpc606_5 gpc179 (
      {stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65], stage0_8[66]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[11],stage1_10[16],stage1_9[52],stage1_8[90]}
   );
   gpc606_5 gpc180 (
      {stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71], stage0_8[72]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[12],stage1_10[17],stage1_9[53],stage1_8[91]}
   );
   gpc606_5 gpc181 (
      {stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77], stage0_8[78]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[13],stage1_10[18],stage1_9[54],stage1_8[92]}
   );
   gpc606_5 gpc182 (
      {stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83], stage0_8[84]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[14],stage1_10[19],stage1_9[55],stage1_8[93]}
   );
   gpc606_5 gpc183 (
      {stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89], stage0_8[90]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[15],stage1_10[20],stage1_9[56],stage1_8[94]}
   );
   gpc606_5 gpc184 (
      {stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95], stage0_8[96]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[16],stage1_10[21],stage1_9[57],stage1_8[95]}
   );
   gpc606_5 gpc185 (
      {stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101], stage0_8[102]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[17],stage1_10[22],stage1_9[58],stage1_8[96]}
   );
   gpc606_5 gpc186 (
      {stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107], stage0_8[108]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[18],stage1_10[23],stage1_9[59],stage1_8[97]}
   );
   gpc606_5 gpc187 (
      {stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113], stage0_8[114]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[19],stage1_10[24],stage1_9[60],stage1_8[98]}
   );
   gpc606_5 gpc188 (
      {stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119], stage0_8[120]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[20],stage1_10[25],stage1_9[61],stage1_8[99]}
   );
   gpc606_5 gpc189 (
      {stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125], stage0_8[126]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[21],stage1_10[26],stage1_9[62],stage1_8[100]}
   );
   gpc606_5 gpc190 (
      {stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131], stage0_8[132]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[22],stage1_10[27],stage1_9[63],stage1_8[101]}
   );
   gpc606_5 gpc191 (
      {stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137], stage0_8[138]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[23],stage1_10[28],stage1_9[64],stage1_8[102]}
   );
   gpc606_5 gpc192 (
      {stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143], stage0_8[144]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[24],stage1_10[29],stage1_9[65],stage1_8[103]}
   );
   gpc606_5 gpc193 (
      {stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149], stage0_8[150]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[25],stage1_10[30],stage1_9[66],stage1_8[104]}
   );
   gpc606_5 gpc194 (
      {stage0_8[151], stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155], stage0_8[156]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[26],stage1_10[31],stage1_9[67],stage1_8[105]}
   );
   gpc606_5 gpc195 (
      {stage0_8[157], stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161], stage0_8[162]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[27],stage1_10[32],stage1_9[68],stage1_8[106]}
   );
   gpc606_5 gpc196 (
      {stage0_8[163], stage0_8[164], stage0_8[165], stage0_8[166], stage0_8[167], stage0_8[168]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[28],stage1_10[33],stage1_9[69],stage1_8[107]}
   );
   gpc606_5 gpc197 (
      {stage0_8[169], stage0_8[170], stage0_8[171], stage0_8[172], stage0_8[173], stage0_8[174]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[29],stage1_10[34],stage1_9[70],stage1_8[108]}
   );
   gpc606_5 gpc198 (
      {stage0_8[175], stage0_8[176], stage0_8[177], stage0_8[178], stage0_8[179], stage0_8[180]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[30],stage1_10[35],stage1_9[71],stage1_8[109]}
   );
   gpc606_5 gpc199 (
      {stage0_8[181], stage0_8[182], stage0_8[183], stage0_8[184], stage0_8[185], stage0_8[186]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[31],stage1_10[36],stage1_9[72],stage1_8[110]}
   );
   gpc606_5 gpc200 (
      {stage0_8[187], stage0_8[188], stage0_8[189], stage0_8[190], stage0_8[191], stage0_8[192]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[32],stage1_10[37],stage1_9[73],stage1_8[111]}
   );
   gpc606_5 gpc201 (
      {stage0_8[193], stage0_8[194], stage0_8[195], stage0_8[196], stage0_8[197], stage0_8[198]},
      {stage0_10[156], stage0_10[157], stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161]},
      {stage1_12[26],stage1_11[33],stage1_10[38],stage1_9[74],stage1_8[112]}
   );
   gpc606_5 gpc202 (
      {stage0_8[199], stage0_8[200], stage0_8[201], stage0_8[202], stage0_8[203], stage0_8[204]},
      {stage0_10[162], stage0_10[163], stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167]},
      {stage1_12[27],stage1_11[34],stage1_10[39],stage1_9[75],stage1_8[113]}
   );
   gpc606_5 gpc203 (
      {stage0_8[205], stage0_8[206], stage0_8[207], stage0_8[208], stage0_8[209], stage0_8[210]},
      {stage0_10[168], stage0_10[169], stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173]},
      {stage1_12[28],stage1_11[35],stage1_10[40],stage1_9[76],stage1_8[114]}
   );
   gpc606_5 gpc204 (
      {stage0_8[211], stage0_8[212], stage0_8[213], stage0_8[214], stage0_8[215], stage0_8[216]},
      {stage0_10[174], stage0_10[175], stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179]},
      {stage1_12[29],stage1_11[36],stage1_10[41],stage1_9[77],stage1_8[115]}
   );
   gpc606_5 gpc205 (
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[30],stage1_11[37],stage1_10[42],stage1_9[78]}
   );
   gpc606_5 gpc206 (
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[31],stage1_11[38],stage1_10[43],stage1_9[79]}
   );
   gpc606_5 gpc207 (
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[32],stage1_11[39],stage1_10[44],stage1_9[80]}
   );
   gpc606_5 gpc208 (
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[33],stage1_11[40],stage1_10[45],stage1_9[81]}
   );
   gpc615_5 gpc209 (
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70]},
      {stage0_10[180]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[34],stage1_11[41],stage1_10[46],stage1_9[82]}
   );
   gpc615_5 gpc210 (
      {stage0_9[71], stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75]},
      {stage0_10[181]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[35],stage1_11[42],stage1_10[47],stage1_9[83]}
   );
   gpc615_5 gpc211 (
      {stage0_9[76], stage0_9[77], stage0_9[78], stage0_9[79], stage0_9[80]},
      {stage0_10[182]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[36],stage1_11[43],stage1_10[48],stage1_9[84]}
   );
   gpc615_5 gpc212 (
      {stage0_9[81], stage0_9[82], stage0_9[83], stage0_9[84], stage0_9[85]},
      {stage0_10[183]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[37],stage1_11[44],stage1_10[49],stage1_9[85]}
   );
   gpc615_5 gpc213 (
      {stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89], stage0_9[90]},
      {stage0_10[184]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[38],stage1_11[45],stage1_10[50],stage1_9[86]}
   );
   gpc615_5 gpc214 (
      {stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage0_10[185]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[39],stage1_11[46],stage1_10[51],stage1_9[87]}
   );
   gpc615_5 gpc215 (
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100]},
      {stage0_10[186]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[40],stage1_11[47],stage1_10[52],stage1_9[88]}
   );
   gpc615_5 gpc216 (
      {stage0_9[101], stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105]},
      {stage0_10[187]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[41],stage1_11[48],stage1_10[53],stage1_9[89]}
   );
   gpc615_5 gpc217 (
      {stage0_9[106], stage0_9[107], stage0_9[108], stage0_9[109], stage0_9[110]},
      {stage0_10[188]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[42],stage1_11[49],stage1_10[54],stage1_9[90]}
   );
   gpc615_5 gpc218 (
      {stage0_9[111], stage0_9[112], stage0_9[113], stage0_9[114], stage0_9[115]},
      {stage0_10[189]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[43],stage1_11[50],stage1_10[55],stage1_9[91]}
   );
   gpc615_5 gpc219 (
      {stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119], stage0_9[120]},
      {stage0_10[190]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[44],stage1_11[51],stage1_10[56],stage1_9[92]}
   );
   gpc615_5 gpc220 (
      {stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage0_10[191]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[45],stage1_11[52],stage1_10[57],stage1_9[93]}
   );
   gpc615_5 gpc221 (
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130]},
      {stage0_10[192]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[46],stage1_11[53],stage1_10[58],stage1_9[94]}
   );
   gpc615_5 gpc222 (
      {stage0_9[131], stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135]},
      {stage0_10[193]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[47],stage1_11[54],stage1_10[59],stage1_9[95]}
   );
   gpc615_5 gpc223 (
      {stage0_9[136], stage0_9[137], stage0_9[138], stage0_9[139], stage0_9[140]},
      {stage0_10[194]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[48],stage1_11[55],stage1_10[60],stage1_9[96]}
   );
   gpc615_5 gpc224 (
      {stage0_9[141], stage0_9[142], stage0_9[143], stage0_9[144], stage0_9[145]},
      {stage0_10[195]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[49],stage1_11[56],stage1_10[61],stage1_9[97]}
   );
   gpc615_5 gpc225 (
      {stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149], stage0_9[150]},
      {stage0_10[196]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[50],stage1_11[57],stage1_10[62],stage1_9[98]}
   );
   gpc615_5 gpc226 (
      {stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage0_10[197]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[51],stage1_11[58],stage1_10[63],stage1_9[99]}
   );
   gpc615_5 gpc227 (
      {stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160]},
      {stage0_10[198]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[52],stage1_11[59],stage1_10[64],stage1_9[100]}
   );
   gpc615_5 gpc228 (
      {stage0_9[161], stage0_9[162], stage0_9[163], stage0_9[164], stage0_9[165]},
      {stage0_10[199]},
      {stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage1_13[23],stage1_12[53],stage1_11[60],stage1_10[65],stage1_9[101]}
   );
   gpc615_5 gpc229 (
      {stage0_9[166], stage0_9[167], stage0_9[168], stage0_9[169], stage0_9[170]},
      {stage0_10[200]},
      {stage0_11[144], stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage1_13[24],stage1_12[54],stage1_11[61],stage1_10[66],stage1_9[102]}
   );
   gpc615_5 gpc230 (
      {stage0_9[171], stage0_9[172], stage0_9[173], stage0_9[174], stage0_9[175]},
      {stage0_10[201]},
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154], stage0_11[155]},
      {stage1_13[25],stage1_12[55],stage1_11[62],stage1_10[67],stage1_9[103]}
   );
   gpc615_5 gpc231 (
      {stage0_9[176], stage0_9[177], stage0_9[178], stage0_9[179], stage0_9[180]},
      {stage0_10[202]},
      {stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159], stage0_11[160], stage0_11[161]},
      {stage1_13[26],stage1_12[56],stage1_11[63],stage1_10[68],stage1_9[104]}
   );
   gpc615_5 gpc232 (
      {stage0_9[181], stage0_9[182], stage0_9[183], stage0_9[184], stage0_9[185]},
      {stage0_10[203]},
      {stage0_11[162], stage0_11[163], stage0_11[164], stage0_11[165], stage0_11[166], stage0_11[167]},
      {stage1_13[27],stage1_12[57],stage1_11[64],stage1_10[69],stage1_9[105]}
   );
   gpc615_5 gpc233 (
      {stage0_9[186], stage0_9[187], stage0_9[188], stage0_9[189], stage0_9[190]},
      {stage0_10[204]},
      {stage0_11[168], stage0_11[169], stage0_11[170], stage0_11[171], stage0_11[172], stage0_11[173]},
      {stage1_13[28],stage1_12[58],stage1_11[65],stage1_10[70],stage1_9[106]}
   );
   gpc615_5 gpc234 (
      {stage0_9[191], stage0_9[192], stage0_9[193], stage0_9[194], stage0_9[195]},
      {stage0_10[205]},
      {stage0_11[174], stage0_11[175], stage0_11[176], stage0_11[177], stage0_11[178], stage0_11[179]},
      {stage1_13[29],stage1_12[59],stage1_11[66],stage1_10[71],stage1_9[107]}
   );
   gpc615_5 gpc235 (
      {stage0_9[196], stage0_9[197], stage0_9[198], stage0_9[199], stage0_9[200]},
      {stage0_10[206]},
      {stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183], stage0_11[184], stage0_11[185]},
      {stage1_13[30],stage1_12[60],stage1_11[67],stage1_10[72],stage1_9[108]}
   );
   gpc615_5 gpc236 (
      {stage0_9[201], stage0_9[202], stage0_9[203], stage0_9[204], stage0_9[205]},
      {stage0_10[207]},
      {stage0_11[186], stage0_11[187], stage0_11[188], stage0_11[189], stage0_11[190], stage0_11[191]},
      {stage1_13[31],stage1_12[61],stage1_11[68],stage1_10[73],stage1_9[109]}
   );
   gpc615_5 gpc237 (
      {stage0_9[206], stage0_9[207], stage0_9[208], stage0_9[209], stage0_9[210]},
      {stage0_10[208]},
      {stage0_11[192], stage0_11[193], stage0_11[194], stage0_11[195], stage0_11[196], stage0_11[197]},
      {stage1_13[32],stage1_12[62],stage1_11[69],stage1_10[74],stage1_9[110]}
   );
   gpc615_5 gpc238 (
      {stage0_9[211], stage0_9[212], stage0_9[213], stage0_9[214], stage0_9[215]},
      {stage0_10[209]},
      {stage0_11[198], stage0_11[199], stage0_11[200], stage0_11[201], stage0_11[202], stage0_11[203]},
      {stage1_13[33],stage1_12[63],stage1_11[70],stage1_10[75],stage1_9[111]}
   );
   gpc615_5 gpc239 (
      {stage0_9[216], stage0_9[217], stage0_9[218], stage0_9[219], stage0_9[220]},
      {stage0_10[210]},
      {stage0_11[204], stage0_11[205], stage0_11[206], stage0_11[207], stage0_11[208], stage0_11[209]},
      {stage1_13[34],stage1_12[64],stage1_11[71],stage1_10[76],stage1_9[112]}
   );
   gpc615_5 gpc240 (
      {stage0_9[221], stage0_9[222], stage0_9[223], stage0_9[224], stage0_9[225]},
      {stage0_10[211]},
      {stage0_11[210], stage0_11[211], stage0_11[212], stage0_11[213], stage0_11[214], stage0_11[215]},
      {stage1_13[35],stage1_12[65],stage1_11[72],stage1_10[77],stage1_9[113]}
   );
   gpc615_5 gpc241 (
      {stage0_9[226], stage0_9[227], stage0_9[228], stage0_9[229], stage0_9[230]},
      {stage0_10[212]},
      {stage0_11[216], stage0_11[217], stage0_11[218], stage0_11[219], stage0_11[220], stage0_11[221]},
      {stage1_13[36],stage1_12[66],stage1_11[73],stage1_10[78],stage1_9[114]}
   );
   gpc615_5 gpc242 (
      {stage0_9[231], stage0_9[232], stage0_9[233], stage0_9[234], stage0_9[235]},
      {stage0_10[213]},
      {stage0_11[222], stage0_11[223], stage0_11[224], stage0_11[225], stage0_11[226], stage0_11[227]},
      {stage1_13[37],stage1_12[67],stage1_11[74],stage1_10[79],stage1_9[115]}
   );
   gpc615_5 gpc243 (
      {stage0_9[236], stage0_9[237], stage0_9[238], stage0_9[239], stage0_9[240]},
      {stage0_10[214]},
      {stage0_11[228], stage0_11[229], stage0_11[230], stage0_11[231], stage0_11[232], stage0_11[233]},
      {stage1_13[38],stage1_12[68],stage1_11[75],stage1_10[80],stage1_9[116]}
   );
   gpc615_5 gpc244 (
      {stage0_9[241], stage0_9[242], stage0_9[243], stage0_9[244], stage0_9[245]},
      {stage0_10[215]},
      {stage0_11[234], stage0_11[235], stage0_11[236], stage0_11[237], stage0_11[238], stage0_11[239]},
      {stage1_13[39],stage1_12[69],stage1_11[76],stage1_10[81],stage1_9[117]}
   );
   gpc615_5 gpc245 (
      {stage0_9[246], stage0_9[247], stage0_9[248], stage0_9[249], stage0_9[250]},
      {stage0_10[216]},
      {stage0_11[240], stage0_11[241], stage0_11[242], stage0_11[243], stage0_11[244], stage0_11[245]},
      {stage1_13[40],stage1_12[70],stage1_11[77],stage1_10[82],stage1_9[118]}
   );
   gpc615_5 gpc246 (
      {stage0_9[251], stage0_9[252], stage0_9[253], stage0_9[254], stage0_9[255]},
      {stage0_10[217]},
      {stage0_11[246], stage0_11[247], stage0_11[248], stage0_11[249], stage0_11[250], stage0_11[251]},
      {stage1_13[41],stage1_12[71],stage1_11[78],stage1_10[83],stage1_9[119]}
   );
   gpc1_1 gpc247 (
      {stage0_0[253]},
      {stage1_0[45]}
   );
   gpc1_1 gpc248 (
      {stage0_0[254]},
      {stage1_0[46]}
   );
   gpc1_1 gpc249 (
      {stage0_0[255]},
      {stage1_0[47]}
   );
   gpc1_1 gpc250 (
      {stage0_1[246]},
      {stage1_1[80]}
   );
   gpc1_1 gpc251 (
      {stage0_1[247]},
      {stage1_1[81]}
   );
   gpc1_1 gpc252 (
      {stage0_1[248]},
      {stage1_1[82]}
   );
   gpc1_1 gpc253 (
      {stage0_1[249]},
      {stage1_1[83]}
   );
   gpc1_1 gpc254 (
      {stage0_1[250]},
      {stage1_1[84]}
   );
   gpc1_1 gpc255 (
      {stage0_1[251]},
      {stage1_1[85]}
   );
   gpc1_1 gpc256 (
      {stage0_1[252]},
      {stage1_1[86]}
   );
   gpc1_1 gpc257 (
      {stage0_1[253]},
      {stage1_1[87]}
   );
   gpc1_1 gpc258 (
      {stage0_1[254]},
      {stage1_1[88]}
   );
   gpc1_1 gpc259 (
      {stage0_1[255]},
      {stage1_1[89]}
   );
   gpc1_1 gpc260 (
      {stage0_2[255]},
      {stage1_2[84]}
   );
   gpc1_1 gpc261 (
      {stage0_3[248]},
      {stage1_3[89]}
   );
   gpc1_1 gpc262 (
      {stage0_3[249]},
      {stage1_3[90]}
   );
   gpc1_1 gpc263 (
      {stage0_3[250]},
      {stage1_3[91]}
   );
   gpc1_1 gpc264 (
      {stage0_3[251]},
      {stage1_3[92]}
   );
   gpc1_1 gpc265 (
      {stage0_3[252]},
      {stage1_3[93]}
   );
   gpc1_1 gpc266 (
      {stage0_3[253]},
      {stage1_3[94]}
   );
   gpc1_1 gpc267 (
      {stage0_3[254]},
      {stage1_3[95]}
   );
   gpc1_1 gpc268 (
      {stage0_3[255]},
      {stage1_3[96]}
   );
   gpc1_1 gpc269 (
      {stage0_5[245]},
      {stage1_5[118]}
   );
   gpc1_1 gpc270 (
      {stage0_5[246]},
      {stage1_5[119]}
   );
   gpc1_1 gpc271 (
      {stage0_5[247]},
      {stage1_5[120]}
   );
   gpc1_1 gpc272 (
      {stage0_5[248]},
      {stage1_5[121]}
   );
   gpc1_1 gpc273 (
      {stage0_5[249]},
      {stage1_5[122]}
   );
   gpc1_1 gpc274 (
      {stage0_5[250]},
      {stage1_5[123]}
   );
   gpc1_1 gpc275 (
      {stage0_5[251]},
      {stage1_5[124]}
   );
   gpc1_1 gpc276 (
      {stage0_5[252]},
      {stage1_5[125]}
   );
   gpc1_1 gpc277 (
      {stage0_5[253]},
      {stage1_5[126]}
   );
   gpc1_1 gpc278 (
      {stage0_5[254]},
      {stage1_5[127]}
   );
   gpc1_1 gpc279 (
      {stage0_5[255]},
      {stage1_5[128]}
   );
   gpc1_1 gpc280 (
      {stage0_6[255]},
      {stage1_6[88]}
   );
   gpc1_1 gpc281 (
      {stage0_8[217]},
      {stage1_8[116]}
   );
   gpc1_1 gpc282 (
      {stage0_8[218]},
      {stage1_8[117]}
   );
   gpc1_1 gpc283 (
      {stage0_8[219]},
      {stage1_8[118]}
   );
   gpc1_1 gpc284 (
      {stage0_8[220]},
      {stage1_8[119]}
   );
   gpc1_1 gpc285 (
      {stage0_8[221]},
      {stage1_8[120]}
   );
   gpc1_1 gpc286 (
      {stage0_8[222]},
      {stage1_8[121]}
   );
   gpc1_1 gpc287 (
      {stage0_8[223]},
      {stage1_8[122]}
   );
   gpc1_1 gpc288 (
      {stage0_8[224]},
      {stage1_8[123]}
   );
   gpc1_1 gpc289 (
      {stage0_8[225]},
      {stage1_8[124]}
   );
   gpc1_1 gpc290 (
      {stage0_8[226]},
      {stage1_8[125]}
   );
   gpc1_1 gpc291 (
      {stage0_8[227]},
      {stage1_8[126]}
   );
   gpc1_1 gpc292 (
      {stage0_8[228]},
      {stage1_8[127]}
   );
   gpc1_1 gpc293 (
      {stage0_8[229]},
      {stage1_8[128]}
   );
   gpc1_1 gpc294 (
      {stage0_8[230]},
      {stage1_8[129]}
   );
   gpc1_1 gpc295 (
      {stage0_8[231]},
      {stage1_8[130]}
   );
   gpc1_1 gpc296 (
      {stage0_8[232]},
      {stage1_8[131]}
   );
   gpc1_1 gpc297 (
      {stage0_8[233]},
      {stage1_8[132]}
   );
   gpc1_1 gpc298 (
      {stage0_8[234]},
      {stage1_8[133]}
   );
   gpc1_1 gpc299 (
      {stage0_8[235]},
      {stage1_8[134]}
   );
   gpc1_1 gpc300 (
      {stage0_8[236]},
      {stage1_8[135]}
   );
   gpc1_1 gpc301 (
      {stage0_8[237]},
      {stage1_8[136]}
   );
   gpc1_1 gpc302 (
      {stage0_8[238]},
      {stage1_8[137]}
   );
   gpc1_1 gpc303 (
      {stage0_8[239]},
      {stage1_8[138]}
   );
   gpc1_1 gpc304 (
      {stage0_8[240]},
      {stage1_8[139]}
   );
   gpc1_1 gpc305 (
      {stage0_8[241]},
      {stage1_8[140]}
   );
   gpc1_1 gpc306 (
      {stage0_8[242]},
      {stage1_8[141]}
   );
   gpc1_1 gpc307 (
      {stage0_8[243]},
      {stage1_8[142]}
   );
   gpc1_1 gpc308 (
      {stage0_8[244]},
      {stage1_8[143]}
   );
   gpc1_1 gpc309 (
      {stage0_8[245]},
      {stage1_8[144]}
   );
   gpc1_1 gpc310 (
      {stage0_8[246]},
      {stage1_8[145]}
   );
   gpc1_1 gpc311 (
      {stage0_8[247]},
      {stage1_8[146]}
   );
   gpc1_1 gpc312 (
      {stage0_8[248]},
      {stage1_8[147]}
   );
   gpc1_1 gpc313 (
      {stage0_8[249]},
      {stage1_8[148]}
   );
   gpc1_1 gpc314 (
      {stage0_8[250]},
      {stage1_8[149]}
   );
   gpc1_1 gpc315 (
      {stage0_8[251]},
      {stage1_8[150]}
   );
   gpc1_1 gpc316 (
      {stage0_8[252]},
      {stage1_8[151]}
   );
   gpc1_1 gpc317 (
      {stage0_8[253]},
      {stage1_8[152]}
   );
   gpc1_1 gpc318 (
      {stage0_8[254]},
      {stage1_8[153]}
   );
   gpc1_1 gpc319 (
      {stage0_8[255]},
      {stage1_8[154]}
   );
   gpc1_1 gpc320 (
      {stage0_10[218]},
      {stage1_10[84]}
   );
   gpc1_1 gpc321 (
      {stage0_10[219]},
      {stage1_10[85]}
   );
   gpc1_1 gpc322 (
      {stage0_10[220]},
      {stage1_10[86]}
   );
   gpc1_1 gpc323 (
      {stage0_10[221]},
      {stage1_10[87]}
   );
   gpc1_1 gpc324 (
      {stage0_10[222]},
      {stage1_10[88]}
   );
   gpc1_1 gpc325 (
      {stage0_10[223]},
      {stage1_10[89]}
   );
   gpc1_1 gpc326 (
      {stage0_10[224]},
      {stage1_10[90]}
   );
   gpc1_1 gpc327 (
      {stage0_10[225]},
      {stage1_10[91]}
   );
   gpc1_1 gpc328 (
      {stage0_10[226]},
      {stage1_10[92]}
   );
   gpc1_1 gpc329 (
      {stage0_10[227]},
      {stage1_10[93]}
   );
   gpc1_1 gpc330 (
      {stage0_10[228]},
      {stage1_10[94]}
   );
   gpc1_1 gpc331 (
      {stage0_10[229]},
      {stage1_10[95]}
   );
   gpc1_1 gpc332 (
      {stage0_10[230]},
      {stage1_10[96]}
   );
   gpc1_1 gpc333 (
      {stage0_10[231]},
      {stage1_10[97]}
   );
   gpc1_1 gpc334 (
      {stage0_10[232]},
      {stage1_10[98]}
   );
   gpc1_1 gpc335 (
      {stage0_10[233]},
      {stage1_10[99]}
   );
   gpc1_1 gpc336 (
      {stage0_10[234]},
      {stage1_10[100]}
   );
   gpc1_1 gpc337 (
      {stage0_10[235]},
      {stage1_10[101]}
   );
   gpc1_1 gpc338 (
      {stage0_10[236]},
      {stage1_10[102]}
   );
   gpc1_1 gpc339 (
      {stage0_10[237]},
      {stage1_10[103]}
   );
   gpc1_1 gpc340 (
      {stage0_10[238]},
      {stage1_10[104]}
   );
   gpc1_1 gpc341 (
      {stage0_10[239]},
      {stage1_10[105]}
   );
   gpc1_1 gpc342 (
      {stage0_10[240]},
      {stage1_10[106]}
   );
   gpc1_1 gpc343 (
      {stage0_10[241]},
      {stage1_10[107]}
   );
   gpc1_1 gpc344 (
      {stage0_10[242]},
      {stage1_10[108]}
   );
   gpc1_1 gpc345 (
      {stage0_10[243]},
      {stage1_10[109]}
   );
   gpc1_1 gpc346 (
      {stage0_10[244]},
      {stage1_10[110]}
   );
   gpc1_1 gpc347 (
      {stage0_10[245]},
      {stage1_10[111]}
   );
   gpc1_1 gpc348 (
      {stage0_10[246]},
      {stage1_10[112]}
   );
   gpc1_1 gpc349 (
      {stage0_10[247]},
      {stage1_10[113]}
   );
   gpc1_1 gpc350 (
      {stage0_10[248]},
      {stage1_10[114]}
   );
   gpc1_1 gpc351 (
      {stage0_10[249]},
      {stage1_10[115]}
   );
   gpc1_1 gpc352 (
      {stage0_10[250]},
      {stage1_10[116]}
   );
   gpc1_1 gpc353 (
      {stage0_10[251]},
      {stage1_10[117]}
   );
   gpc1_1 gpc354 (
      {stage0_10[252]},
      {stage1_10[118]}
   );
   gpc1_1 gpc355 (
      {stage0_10[253]},
      {stage1_10[119]}
   );
   gpc1_1 gpc356 (
      {stage0_10[254]},
      {stage1_10[120]}
   );
   gpc1_1 gpc357 (
      {stage0_10[255]},
      {stage1_10[121]}
   );
   gpc1_1 gpc358 (
      {stage0_11[252]},
      {stage1_11[79]}
   );
   gpc1_1 gpc359 (
      {stage0_11[253]},
      {stage1_11[80]}
   );
   gpc1_1 gpc360 (
      {stage0_11[254]},
      {stage1_11[81]}
   );
   gpc1_1 gpc361 (
      {stage0_11[255]},
      {stage1_11[82]}
   );
   gpc1163_5 gpc362 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc363 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc364 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc365 (
      {stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[3]},
      {stage1_3[3]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc366 (
      {stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[4]},
      {stage1_3[4]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc1163_5 gpc367 (
      {stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_2[5]},
      {stage1_3[5]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc1163_5 gpc368 (
      {stage1_0[18], stage1_0[19], stage1_0[20]},
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_2[6]},
      {stage1_3[6]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc1163_5 gpc369 (
      {stage1_0[21], stage1_0[22], stage1_0[23]},
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_2[7]},
      {stage1_3[7]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc1163_5 gpc370 (
      {stage1_0[24], stage1_0[25], stage1_0[26]},
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_2[8]},
      {stage1_3[8]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc1163_5 gpc371 (
      {stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59]},
      {stage1_2[9]},
      {stage1_3[9]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc1163_5 gpc372 (
      {stage1_0[30], stage1_0[31], stage1_0[32]},
      {stage1_1[60], stage1_1[61], stage1_1[62], stage1_1[63], stage1_1[64], stage1_1[65]},
      {stage1_2[10]},
      {stage1_3[10]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc1163_5 gpc373 (
      {stage1_0[33], stage1_0[34], stage1_0[35]},
      {stage1_1[66], stage1_1[67], stage1_1[68], stage1_1[69], stage1_1[70], stage1_1[71]},
      {stage1_2[11]},
      {stage1_3[11]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc606_5 gpc374 (
      {stage1_0[36], stage1_0[37], stage1_0[38], stage1_0[39], stage1_0[40], stage1_0[41]},
      {stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17]},
      {stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12],stage2_0[12]}
   );
   gpc7_3 gpc375 (
      {stage1_1[72], stage1_1[73], stage1_1[74], stage1_1[75], stage1_1[76], stage1_1[77], stage1_1[78]},
      {stage2_3[13],stage2_2[13],stage2_1[13]}
   );
   gpc606_5 gpc376 (
      {stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[0],stage2_4[13],stage2_3[14],stage2_2[14]}
   );
   gpc606_5 gpc377 (
      {stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27], stage1_2[28], stage1_2[29]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[1],stage2_4[14],stage2_3[15],stage2_2[15]}
   );
   gpc606_5 gpc378 (
      {stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33], stage1_2[34], stage1_2[35]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[2],stage2_4[15],stage2_3[16],stage2_2[16]}
   );
   gpc606_5 gpc379 (
      {stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39], stage1_2[40], stage1_2[41]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[3],stage2_4[16],stage2_3[17],stage2_2[17]}
   );
   gpc606_5 gpc380 (
      {stage1_2[42], stage1_2[43], stage1_2[44], stage1_2[45], stage1_2[46], stage1_2[47]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[4],stage2_4[17],stage2_3[18],stage2_2[18]}
   );
   gpc606_5 gpc381 (
      {stage1_2[48], stage1_2[49], stage1_2[50], stage1_2[51], stage1_2[52], stage1_2[53]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[5],stage2_4[18],stage2_3[19],stage2_2[19]}
   );
   gpc606_5 gpc382 (
      {stage1_2[54], stage1_2[55], stage1_2[56], stage1_2[57], stage1_2[58], stage1_2[59]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[6],stage2_4[19],stage2_3[20],stage2_2[20]}
   );
   gpc606_5 gpc383 (
      {stage1_2[60], stage1_2[61], stage1_2[62], stage1_2[63], stage1_2[64], stage1_2[65]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[7],stage2_4[20],stage2_3[21],stage2_2[21]}
   );
   gpc606_5 gpc384 (
      {stage1_2[66], stage1_2[67], stage1_2[68], stage1_2[69], stage1_2[70], stage1_2[71]},
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage2_6[8],stage2_5[8],stage2_4[21],stage2_3[22],stage2_2[22]}
   );
   gpc606_5 gpc385 (
      {stage1_2[72], stage1_2[73], stage1_2[74], stage1_2[75], stage1_2[76], stage1_2[77]},
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage2_6[9],stage2_5[9],stage2_4[22],stage2_3[23],stage2_2[23]}
   );
   gpc606_5 gpc386 (
      {stage1_2[78], stage1_2[79], stage1_2[80], stage1_2[81], stage1_2[82], stage1_2[83]},
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage2_6[10],stage2_5[10],stage2_4[23],stage2_3[24],stage2_2[24]}
   );
   gpc615_5 gpc387 (
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16]},
      {stage1_4[66]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[11],stage2_5[11],stage2_4[24],stage2_3[25]}
   );
   gpc615_5 gpc388 (
      {stage1_3[17], stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21]},
      {stage1_4[67]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[12],stage2_5[12],stage2_4[25],stage2_3[26]}
   );
   gpc615_5 gpc389 (
      {stage1_3[22], stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26]},
      {stage1_4[68]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[13],stage2_5[13],stage2_4[26],stage2_3[27]}
   );
   gpc615_5 gpc390 (
      {stage1_3[27], stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31]},
      {stage1_4[69]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[14],stage2_5[14],stage2_4[27],stage2_3[28]}
   );
   gpc615_5 gpc391 (
      {stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35], stage1_3[36]},
      {stage1_4[70]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[15],stage2_5[15],stage2_4[28],stage2_3[29]}
   );
   gpc615_5 gpc392 (
      {stage1_3[37], stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41]},
      {stage1_4[71]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[16],stage2_5[16],stage2_4[29],stage2_3[30]}
   );
   gpc615_5 gpc393 (
      {stage1_3[42], stage1_3[43], stage1_3[44], stage1_3[45], stage1_3[46]},
      {stage1_4[72]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[17],stage2_5[17],stage2_4[30],stage2_3[31]}
   );
   gpc615_5 gpc394 (
      {stage1_3[47], stage1_3[48], stage1_3[49], stage1_3[50], stage1_3[51]},
      {stage1_4[73]},
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage2_7[7],stage2_6[18],stage2_5[18],stage2_4[31],stage2_3[32]}
   );
   gpc615_5 gpc395 (
      {stage1_3[52], stage1_3[53], stage1_3[54], stage1_3[55], stage1_3[56]},
      {stage1_4[74]},
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage2_7[8],stage2_6[19],stage2_5[19],stage2_4[32],stage2_3[33]}
   );
   gpc615_5 gpc396 (
      {stage1_3[57], stage1_3[58], stage1_3[59], stage1_3[60], stage1_3[61]},
      {stage1_4[75]},
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage2_7[9],stage2_6[20],stage2_5[20],stage2_4[33],stage2_3[34]}
   );
   gpc615_5 gpc397 (
      {stage1_3[62], stage1_3[63], stage1_3[64], stage1_3[65], stage1_3[66]},
      {stage1_4[76]},
      {stage1_5[60], stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65]},
      {stage2_7[10],stage2_6[21],stage2_5[21],stage2_4[34],stage2_3[35]}
   );
   gpc615_5 gpc398 (
      {stage1_3[67], stage1_3[68], stage1_3[69], stage1_3[70], stage1_3[71]},
      {stage1_4[77]},
      {stage1_5[66], stage1_5[67], stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71]},
      {stage2_7[11],stage2_6[22],stage2_5[22],stage2_4[35],stage2_3[36]}
   );
   gpc615_5 gpc399 (
      {stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75], stage1_3[76]},
      {stage1_4[78]},
      {stage1_5[72], stage1_5[73], stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77]},
      {stage2_7[12],stage2_6[23],stage2_5[23],stage2_4[36],stage2_3[37]}
   );
   gpc615_5 gpc400 (
      {stage1_3[77], stage1_3[78], stage1_3[79], stage1_3[80], stage1_3[81]},
      {stage1_4[79]},
      {stage1_5[78], stage1_5[79], stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83]},
      {stage2_7[13],stage2_6[24],stage2_5[24],stage2_4[37],stage2_3[38]}
   );
   gpc615_5 gpc401 (
      {stage1_3[82], stage1_3[83], stage1_3[84], stage1_3[85], stage1_3[86]},
      {stage1_4[80]},
      {stage1_5[84], stage1_5[85], stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89]},
      {stage2_7[14],stage2_6[25],stage2_5[25],stage2_4[38],stage2_3[39]}
   );
   gpc615_5 gpc402 (
      {stage1_3[87], stage1_3[88], stage1_3[89], stage1_3[90], stage1_3[91]},
      {stage1_4[81]},
      {stage1_5[90], stage1_5[91], stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95]},
      {stage2_7[15],stage2_6[26],stage2_5[26],stage2_4[39],stage2_3[40]}
   );
   gpc615_5 gpc403 (
      {stage1_3[92], stage1_3[93], stage1_3[94], stage1_3[95], stage1_3[96]},
      {stage1_4[82]},
      {stage1_5[96], stage1_5[97], stage1_5[98], stage1_5[99], stage1_5[100], stage1_5[101]},
      {stage2_7[16],stage2_6[27],stage2_5[27],stage2_4[40],stage2_3[41]}
   );
   gpc606_5 gpc404 (
      {stage1_4[83], stage1_4[84], stage1_4[85], stage1_4[86], stage1_4[87], stage1_4[88]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[17],stage2_6[28],stage2_5[28],stage2_4[41]}
   );
   gpc606_5 gpc405 (
      {stage1_4[89], stage1_4[90], stage1_4[91], stage1_4[92], stage1_4[93], stage1_4[94]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[18],stage2_6[29],stage2_5[29],stage2_4[42]}
   );
   gpc606_5 gpc406 (
      {stage1_4[95], stage1_4[96], stage1_4[97], stage1_4[98], stage1_4[99], stage1_4[100]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[19],stage2_6[30],stage2_5[30],stage2_4[43]}
   );
   gpc606_5 gpc407 (
      {stage1_4[101], stage1_4[102], stage1_4[103], stage1_4[104], stage1_4[105], stage1_4[106]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[20],stage2_6[31],stage2_5[31],stage2_4[44]}
   );
   gpc606_5 gpc408 (
      {stage1_4[107], stage1_4[108], stage1_4[109], stage1_4[110], stage1_4[111], stage1_4[112]},
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage2_8[4],stage2_7[21],stage2_6[32],stage2_5[32],stage2_4[45]}
   );
   gpc606_5 gpc409 (
      {stage1_4[113], stage1_4[114], stage1_4[115], stage1_4[116], stage1_4[117], stage1_4[118]},
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage2_8[5],stage2_7[22],stage2_6[33],stage2_5[33],stage2_4[46]}
   );
   gpc606_5 gpc410 (
      {stage1_4[119], stage1_4[120], stage1_4[121], stage1_4[122], stage1_4[123], stage1_4[124]},
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage2_8[6],stage2_7[23],stage2_6[34],stage2_5[34],stage2_4[47]}
   );
   gpc606_5 gpc411 (
      {stage1_5[102], stage1_5[103], stage1_5[104], stage1_5[105], stage1_5[106], stage1_5[107]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[7],stage2_7[24],stage2_6[35],stage2_5[35]}
   );
   gpc606_5 gpc412 (
      {stage1_5[108], stage1_5[109], stage1_5[110], stage1_5[111], stage1_5[112], stage1_5[113]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[8],stage2_7[25],stage2_6[36],stage2_5[36]}
   );
   gpc606_5 gpc413 (
      {stage1_5[114], stage1_5[115], stage1_5[116], stage1_5[117], stage1_5[118], stage1_5[119]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[9],stage2_7[26],stage2_6[37],stage2_5[37]}
   );
   gpc606_5 gpc414 (
      {stage1_5[120], stage1_5[121], stage1_5[122], stage1_5[123], stage1_5[124], stage1_5[125]},
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage2_9[3],stage2_8[10],stage2_7[27],stage2_6[38],stage2_5[38]}
   );
   gpc615_5 gpc415 (
      {stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46]},
      {stage1_7[24]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[4],stage2_8[11],stage2_7[28],stage2_6[39]}
   );
   gpc615_5 gpc416 (
      {stage1_6[47], stage1_6[48], stage1_6[49], stage1_6[50], stage1_6[51]},
      {stage1_7[25]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[5],stage2_8[12],stage2_7[29],stage2_6[40]}
   );
   gpc615_5 gpc417 (
      {stage1_6[52], stage1_6[53], stage1_6[54], stage1_6[55], stage1_6[56]},
      {stage1_7[26]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[6],stage2_8[13],stage2_7[30],stage2_6[41]}
   );
   gpc615_5 gpc418 (
      {stage1_6[57], stage1_6[58], stage1_6[59], stage1_6[60], stage1_6[61]},
      {stage1_7[27]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[7],stage2_8[14],stage2_7[31],stage2_6[42]}
   );
   gpc615_5 gpc419 (
      {stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65], stage1_6[66]},
      {stage1_7[28]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[8],stage2_8[15],stage2_7[32],stage2_6[43]}
   );
   gpc615_5 gpc420 (
      {stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71]},
      {stage1_7[29]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[9],stage2_8[16],stage2_7[33],stage2_6[44]}
   );
   gpc615_5 gpc421 (
      {stage1_6[72], stage1_6[73], stage1_6[74], stage1_6[75], stage1_6[76]},
      {stage1_7[30]},
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage2_10[6],stage2_9[10],stage2_8[17],stage2_7[34],stage2_6[45]}
   );
   gpc615_5 gpc422 (
      {stage1_6[77], stage1_6[78], stage1_6[79], stage1_6[80], stage1_6[81]},
      {stage1_7[31]},
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage2_10[7],stage2_9[11],stage2_8[18],stage2_7[35],stage2_6[46]}
   );
   gpc615_5 gpc423 (
      {stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35], stage1_7[36]},
      {stage1_8[48]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[8],stage2_9[12],stage2_8[19],stage2_7[36]}
   );
   gpc615_5 gpc424 (
      {stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage1_8[49]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[9],stage2_9[13],stage2_8[20],stage2_7[37]}
   );
   gpc615_5 gpc425 (
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46]},
      {stage1_8[50]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[10],stage2_9[14],stage2_8[21],stage2_7[38]}
   );
   gpc615_5 gpc426 (
      {stage1_7[47], stage1_7[48], stage1_7[49], stage1_7[50], stage1_7[51]},
      {stage1_8[51]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[11],stage2_9[15],stage2_8[22],stage2_7[39]}
   );
   gpc615_5 gpc427 (
      {stage1_7[52], stage1_7[53], stage1_7[54], stage1_7[55], stage1_7[56]},
      {stage1_8[52]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[12],stage2_9[16],stage2_8[23],stage2_7[40]}
   );
   gpc615_5 gpc428 (
      {stage1_7[57], stage1_7[58], stage1_7[59], stage1_7[60], stage1_7[61]},
      {stage1_8[53]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[13],stage2_9[17],stage2_8[24],stage2_7[41]}
   );
   gpc615_5 gpc429 (
      {stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65], stage1_7[66]},
      {stage1_8[54]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[14],stage2_9[18],stage2_8[25],stage2_7[42]}
   );
   gpc615_5 gpc430 (
      {stage1_7[67], stage1_7[68], stage1_7[69], stage1_7[70], stage1_7[71]},
      {stage1_8[55]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[15],stage2_9[19],stage2_8[26],stage2_7[43]}
   );
   gpc615_5 gpc431 (
      {stage1_7[72], stage1_7[73], stage1_7[74], stage1_7[75], stage1_7[76]},
      {stage1_8[56]},
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage2_11[8],stage2_10[16],stage2_9[20],stage2_8[27],stage2_7[44]}
   );
   gpc615_5 gpc432 (
      {stage1_7[77], stage1_7[78], stage1_7[79], stage1_7[80], stage1_7[81]},
      {stage1_8[57]},
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage2_11[9],stage2_10[17],stage2_9[21],stage2_8[28],stage2_7[45]}
   );
   gpc615_5 gpc433 (
      {stage1_7[82], stage1_7[83], stage1_7[84], stage1_7[85], stage1_7[86]},
      {stage1_8[58]},
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage2_11[10],stage2_10[18],stage2_9[22],stage2_8[29],stage2_7[46]}
   );
   gpc615_5 gpc434 (
      {stage1_7[87], stage1_7[88], stage1_7[89], stage1_7[90], 1'b0},
      {stage1_8[59]},
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage2_11[11],stage2_10[19],stage2_9[23],stage2_8[30],stage2_7[47]}
   );
   gpc606_5 gpc435 (
      {stage1_8[60], stage1_8[61], stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[12],stage2_10[20],stage2_9[24],stage2_8[31]}
   );
   gpc606_5 gpc436 (
      {stage1_8[66], stage1_8[67], stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[13],stage2_10[21],stage2_9[25],stage2_8[32]}
   );
   gpc606_5 gpc437 (
      {stage1_8[72], stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[14],stage2_10[22],stage2_9[26],stage2_8[33]}
   );
   gpc606_5 gpc438 (
      {stage1_8[78], stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[15],stage2_10[23],stage2_9[27],stage2_8[34]}
   );
   gpc606_5 gpc439 (
      {stage1_8[84], stage1_8[85], stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[16],stage2_10[24],stage2_9[28],stage2_8[35]}
   );
   gpc606_5 gpc440 (
      {stage1_8[90], stage1_8[91], stage1_8[92], stage1_8[93], stage1_8[94], stage1_8[95]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[17],stage2_10[25],stage2_9[29],stage2_8[36]}
   );
   gpc606_5 gpc441 (
      {stage1_8[96], stage1_8[97], stage1_8[98], stage1_8[99], stage1_8[100], stage1_8[101]},
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage2_12[6],stage2_11[18],stage2_10[26],stage2_9[30],stage2_8[37]}
   );
   gpc606_5 gpc442 (
      {stage1_8[102], stage1_8[103], stage1_8[104], stage1_8[105], stage1_8[106], stage1_8[107]},
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage2_12[7],stage2_11[19],stage2_10[27],stage2_9[31],stage2_8[38]}
   );
   gpc606_5 gpc443 (
      {stage1_8[108], stage1_8[109], stage1_8[110], stage1_8[111], stage1_8[112], stage1_8[113]},
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage2_12[8],stage2_11[20],stage2_10[28],stage2_9[32],stage2_8[39]}
   );
   gpc606_5 gpc444 (
      {stage1_8[114], stage1_8[115], stage1_8[116], stage1_8[117], stage1_8[118], stage1_8[119]},
      {stage1_10[54], stage1_10[55], stage1_10[56], stage1_10[57], stage1_10[58], stage1_10[59]},
      {stage2_12[9],stage2_11[21],stage2_10[29],stage2_9[33],stage2_8[40]}
   );
   gpc606_5 gpc445 (
      {stage1_8[120], stage1_8[121], stage1_8[122], stage1_8[123], stage1_8[124], stage1_8[125]},
      {stage1_10[60], stage1_10[61], stage1_10[62], stage1_10[63], stage1_10[64], stage1_10[65]},
      {stage2_12[10],stage2_11[22],stage2_10[30],stage2_9[34],stage2_8[41]}
   );
   gpc606_5 gpc446 (
      {stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[11],stage2_11[23],stage2_10[31],stage2_9[35]}
   );
   gpc606_5 gpc447 (
      {stage1_9[78], stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[12],stage2_11[24],stage2_10[32],stage2_9[36]}
   );
   gpc606_5 gpc448 (
      {stage1_9[84], stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[13],stage2_11[25],stage2_10[33],stage2_9[37]}
   );
   gpc606_5 gpc449 (
      {stage1_9[90], stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[14],stage2_11[26],stage2_10[34],stage2_9[38]}
   );
   gpc606_5 gpc450 (
      {stage1_9[96], stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100], stage1_9[101]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[15],stage2_11[27],stage2_10[35],stage2_9[39]}
   );
   gpc606_5 gpc451 (
      {stage1_9[102], stage1_9[103], stage1_9[104], stage1_9[105], stage1_9[106], stage1_9[107]},
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage2_13[5],stage2_12[16],stage2_11[28],stage2_10[36],stage2_9[40]}
   );
   gpc606_5 gpc452 (
      {stage1_9[108], stage1_9[109], stage1_9[110], stage1_9[111], stage1_9[112], stage1_9[113]},
      {stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41]},
      {stage2_13[6],stage2_12[17],stage2_11[29],stage2_10[37],stage2_9[41]}
   );
   gpc606_5 gpc453 (
      {stage1_9[114], stage1_9[115], stage1_9[116], stage1_9[117], stage1_9[118], stage1_9[119]},
      {stage1_11[42], stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage2_13[7],stage2_12[18],stage2_11[30],stage2_10[38],stage2_9[42]}
   );
   gpc606_5 gpc454 (
      {stage1_10[66], stage1_10[67], stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[8],stage2_12[19],stage2_11[31],stage2_10[39]}
   );
   gpc615_5 gpc455 (
      {stage1_10[72], stage1_10[73], stage1_10[74], stage1_10[75], stage1_10[76]},
      {stage1_11[48]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[9],stage2_12[20],stage2_11[32],stage2_10[40]}
   );
   gpc615_5 gpc456 (
      {stage1_10[77], stage1_10[78], stage1_10[79], stage1_10[80], stage1_10[81]},
      {stage1_11[49]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[10],stage2_12[21],stage2_11[33],stage2_10[41]}
   );
   gpc615_5 gpc457 (
      {stage1_10[82], stage1_10[83], stage1_10[84], stage1_10[85], stage1_10[86]},
      {stage1_11[50]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[11],stage2_12[22],stage2_11[34],stage2_10[42]}
   );
   gpc615_5 gpc458 (
      {stage1_10[87], stage1_10[88], stage1_10[89], stage1_10[90], stage1_10[91]},
      {stage1_11[51]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[12],stage2_12[23],stage2_11[35],stage2_10[43]}
   );
   gpc615_5 gpc459 (
      {stage1_10[92], stage1_10[93], stage1_10[94], stage1_10[95], stage1_10[96]},
      {stage1_11[52]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[13],stage2_12[24],stage2_11[36],stage2_10[44]}
   );
   gpc615_5 gpc460 (
      {stage1_10[97], stage1_10[98], stage1_10[99], stage1_10[100], stage1_10[101]},
      {stage1_11[53]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[14],stage2_12[25],stage2_11[37],stage2_10[45]}
   );
   gpc615_5 gpc461 (
      {stage1_10[102], stage1_10[103], stage1_10[104], stage1_10[105], stage1_10[106]},
      {stage1_11[54]},
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage2_14[7],stage2_13[15],stage2_12[26],stage2_11[38],stage2_10[46]}
   );
   gpc615_5 gpc462 (
      {stage1_10[107], stage1_10[108], stage1_10[109], stage1_10[110], stage1_10[111]},
      {stage1_11[55]},
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage2_14[8],stage2_13[16],stage2_12[27],stage2_11[39],stage2_10[47]}
   );
   gpc615_5 gpc463 (
      {stage1_10[112], stage1_10[113], stage1_10[114], stage1_10[115], stage1_10[116]},
      {stage1_11[56]},
      {stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage2_14[9],stage2_13[17],stage2_12[28],stage2_11[40],stage2_10[48]}
   );
   gpc615_5 gpc464 (
      {stage1_10[117], stage1_10[118], stage1_10[119], stage1_10[120], stage1_10[121]},
      {stage1_11[57]},
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64], stage1_12[65]},
      {stage2_14[10],stage2_13[18],stage2_12[29],stage2_11[41],stage2_10[49]}
   );
   gpc615_5 gpc465 (
      {stage1_11[58], stage1_11[59], stage1_11[60], stage1_11[61], stage1_11[62]},
      {stage1_12[66]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[11],stage2_13[19],stage2_12[30],stage2_11[42]}
   );
   gpc615_5 gpc466 (
      {stage1_11[63], stage1_11[64], stage1_11[65], stage1_11[66], stage1_11[67]},
      {stage1_12[67]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[12],stage2_13[20],stage2_12[31],stage2_11[43]}
   );
   gpc615_5 gpc467 (
      {stage1_11[68], stage1_11[69], stage1_11[70], stage1_11[71], stage1_11[72]},
      {stage1_12[68]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[13],stage2_13[21],stage2_12[32],stage2_11[44]}
   );
   gpc615_5 gpc468 (
      {stage1_11[73], stage1_11[74], stage1_11[75], stage1_11[76], stage1_11[77]},
      {stage1_12[69]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[14],stage2_13[22],stage2_12[33],stage2_11[45]}
   );
   gpc615_5 gpc469 (
      {stage1_11[78], stage1_11[79], stage1_11[80], stage1_11[81], stage1_11[82]},
      {stage1_12[70]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[15],stage2_13[23],stage2_12[34],stage2_11[46]}
   );
   gpc1_1 gpc470 (
      {stage1_0[42]},
      {stage2_0[13]}
   );
   gpc1_1 gpc471 (
      {stage1_0[43]},
      {stage2_0[14]}
   );
   gpc1_1 gpc472 (
      {stage1_0[44]},
      {stage2_0[15]}
   );
   gpc1_1 gpc473 (
      {stage1_0[45]},
      {stage2_0[16]}
   );
   gpc1_1 gpc474 (
      {stage1_0[46]},
      {stage2_0[17]}
   );
   gpc1_1 gpc475 (
      {stage1_0[47]},
      {stage2_0[18]}
   );
   gpc1_1 gpc476 (
      {stage1_1[79]},
      {stage2_1[14]}
   );
   gpc1_1 gpc477 (
      {stage1_1[80]},
      {stage2_1[15]}
   );
   gpc1_1 gpc478 (
      {stage1_1[81]},
      {stage2_1[16]}
   );
   gpc1_1 gpc479 (
      {stage1_1[82]},
      {stage2_1[17]}
   );
   gpc1_1 gpc480 (
      {stage1_1[83]},
      {stage2_1[18]}
   );
   gpc1_1 gpc481 (
      {stage1_1[84]},
      {stage2_1[19]}
   );
   gpc1_1 gpc482 (
      {stage1_1[85]},
      {stage2_1[20]}
   );
   gpc1_1 gpc483 (
      {stage1_1[86]},
      {stage2_1[21]}
   );
   gpc1_1 gpc484 (
      {stage1_1[87]},
      {stage2_1[22]}
   );
   gpc1_1 gpc485 (
      {stage1_1[88]},
      {stage2_1[23]}
   );
   gpc1_1 gpc486 (
      {stage1_1[89]},
      {stage2_1[24]}
   );
   gpc1_1 gpc487 (
      {stage1_2[84]},
      {stage2_2[25]}
   );
   gpc1_1 gpc488 (
      {stage1_4[125]},
      {stage2_4[48]}
   );
   gpc1_1 gpc489 (
      {stage1_4[126]},
      {stage2_4[49]}
   );
   gpc1_1 gpc490 (
      {stage1_5[126]},
      {stage2_5[39]}
   );
   gpc1_1 gpc491 (
      {stage1_5[127]},
      {stage2_5[40]}
   );
   gpc1_1 gpc492 (
      {stage1_5[128]},
      {stage2_5[41]}
   );
   gpc1_1 gpc493 (
      {stage1_6[82]},
      {stage2_6[47]}
   );
   gpc1_1 gpc494 (
      {stage1_6[83]},
      {stage2_6[48]}
   );
   gpc1_1 gpc495 (
      {stage1_6[84]},
      {stage2_6[49]}
   );
   gpc1_1 gpc496 (
      {stage1_6[85]},
      {stage2_6[50]}
   );
   gpc1_1 gpc497 (
      {stage1_6[86]},
      {stage2_6[51]}
   );
   gpc1_1 gpc498 (
      {stage1_6[87]},
      {stage2_6[52]}
   );
   gpc1_1 gpc499 (
      {stage1_6[88]},
      {stage2_6[53]}
   );
   gpc1_1 gpc500 (
      {stage1_8[126]},
      {stage2_8[42]}
   );
   gpc1_1 gpc501 (
      {stage1_8[127]},
      {stage2_8[43]}
   );
   gpc1_1 gpc502 (
      {stage1_8[128]},
      {stage2_8[44]}
   );
   gpc1_1 gpc503 (
      {stage1_8[129]},
      {stage2_8[45]}
   );
   gpc1_1 gpc504 (
      {stage1_8[130]},
      {stage2_8[46]}
   );
   gpc1_1 gpc505 (
      {stage1_8[131]},
      {stage2_8[47]}
   );
   gpc1_1 gpc506 (
      {stage1_8[132]},
      {stage2_8[48]}
   );
   gpc1_1 gpc507 (
      {stage1_8[133]},
      {stage2_8[49]}
   );
   gpc1_1 gpc508 (
      {stage1_8[134]},
      {stage2_8[50]}
   );
   gpc1_1 gpc509 (
      {stage1_8[135]},
      {stage2_8[51]}
   );
   gpc1_1 gpc510 (
      {stage1_8[136]},
      {stage2_8[52]}
   );
   gpc1_1 gpc511 (
      {stage1_8[137]},
      {stage2_8[53]}
   );
   gpc1_1 gpc512 (
      {stage1_8[138]},
      {stage2_8[54]}
   );
   gpc1_1 gpc513 (
      {stage1_8[139]},
      {stage2_8[55]}
   );
   gpc1_1 gpc514 (
      {stage1_8[140]},
      {stage2_8[56]}
   );
   gpc1_1 gpc515 (
      {stage1_8[141]},
      {stage2_8[57]}
   );
   gpc1_1 gpc516 (
      {stage1_8[142]},
      {stage2_8[58]}
   );
   gpc1_1 gpc517 (
      {stage1_8[143]},
      {stage2_8[59]}
   );
   gpc1_1 gpc518 (
      {stage1_8[144]},
      {stage2_8[60]}
   );
   gpc1_1 gpc519 (
      {stage1_8[145]},
      {stage2_8[61]}
   );
   gpc1_1 gpc520 (
      {stage1_8[146]},
      {stage2_8[62]}
   );
   gpc1_1 gpc521 (
      {stage1_8[147]},
      {stage2_8[63]}
   );
   gpc1_1 gpc522 (
      {stage1_8[148]},
      {stage2_8[64]}
   );
   gpc1_1 gpc523 (
      {stage1_8[149]},
      {stage2_8[65]}
   );
   gpc1_1 gpc524 (
      {stage1_8[150]},
      {stage2_8[66]}
   );
   gpc1_1 gpc525 (
      {stage1_8[151]},
      {stage2_8[67]}
   );
   gpc1_1 gpc526 (
      {stage1_8[152]},
      {stage2_8[68]}
   );
   gpc1_1 gpc527 (
      {stage1_8[153]},
      {stage2_8[69]}
   );
   gpc1_1 gpc528 (
      {stage1_8[154]},
      {stage2_8[70]}
   );
   gpc1_1 gpc529 (
      {stage1_12[71]},
      {stage2_12[35]}
   );
   gpc1_1 gpc530 (
      {stage1_13[30]},
      {stage2_13[24]}
   );
   gpc1_1 gpc531 (
      {stage1_13[31]},
      {stage2_13[25]}
   );
   gpc1_1 gpc532 (
      {stage1_13[32]},
      {stage2_13[26]}
   );
   gpc1_1 gpc533 (
      {stage1_13[33]},
      {stage2_13[27]}
   );
   gpc1_1 gpc534 (
      {stage1_13[34]},
      {stage2_13[28]}
   );
   gpc1_1 gpc535 (
      {stage1_13[35]},
      {stage2_13[29]}
   );
   gpc1_1 gpc536 (
      {stage1_13[36]},
      {stage2_13[30]}
   );
   gpc1_1 gpc537 (
      {stage1_13[37]},
      {stage2_13[31]}
   );
   gpc1_1 gpc538 (
      {stage1_13[38]},
      {stage2_13[32]}
   );
   gpc1_1 gpc539 (
      {stage1_13[39]},
      {stage2_13[33]}
   );
   gpc1_1 gpc540 (
      {stage1_13[40]},
      {stage2_13[34]}
   );
   gpc1_1 gpc541 (
      {stage1_13[41]},
      {stage2_13[35]}
   );
   gpc606_5 gpc542 (
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0]}
   );
   gpc606_5 gpc543 (
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11]},
      {stage3_5[1],stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1]}
   );
   gpc606_5 gpc544 (
      {stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15], stage2_1[16], stage2_1[17]},
      {stage2_3[12], stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17]},
      {stage3_5[2],stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2]}
   );
   gpc606_5 gpc545 (
      {stage2_1[18], stage2_1[19], stage2_1[20], stage2_1[21], stage2_1[22], stage2_1[23]},
      {stage2_3[18], stage2_3[19], stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23]},
      {stage3_5[3],stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3]}
   );
   gpc606_5 gpc546 (
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[4],stage3_4[4],stage3_3[4],stage3_2[4]}
   );
   gpc615_5 gpc547 (
      {stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10]},
      {stage2_3[24]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[5],stage3_4[5],stage3_3[5],stage3_2[5]}
   );
   gpc615_5 gpc548 (
      {stage2_2[11], stage2_2[12], stage2_2[13], stage2_2[14], stage2_2[15]},
      {stage2_3[25]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage3_6[2],stage3_5[6],stage3_4[6],stage3_3[6],stage3_2[6]}
   );
   gpc615_5 gpc549 (
      {stage2_2[16], stage2_2[17], stage2_2[18], stage2_2[19], stage2_2[20]},
      {stage2_3[26]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage3_6[3],stage3_5[7],stage3_4[7],stage3_3[7],stage3_2[7]}
   );
   gpc615_5 gpc550 (
      {stage2_3[27], stage2_3[28], stage2_3[29], stage2_3[30], stage2_3[31]},
      {stage2_4[24]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[4],stage3_5[8],stage3_4[8],stage3_3[8]}
   );
   gpc615_5 gpc551 (
      {stage2_3[32], stage2_3[33], stage2_3[34], stage2_3[35], stage2_3[36]},
      {stage2_4[25]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[5],stage3_5[9],stage3_4[9],stage3_3[9]}
   );
   gpc615_5 gpc552 (
      {stage2_3[37], stage2_3[38], stage2_3[39], stage2_3[40], stage2_3[41]},
      {stage2_4[26]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[6],stage3_5[10],stage3_4[10],stage3_3[10]}
   );
   gpc606_5 gpc553 (
      {stage2_4[27], stage2_4[28], stage2_4[29], stage2_4[30], stage2_4[31], stage2_4[32]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[3],stage3_6[7],stage3_5[11],stage3_4[11]}
   );
   gpc606_5 gpc554 (
      {stage2_4[33], stage2_4[34], stage2_4[35], stage2_4[36], stage2_4[37], stage2_4[38]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[4],stage3_6[8],stage3_5[12],stage3_4[12]}
   );
   gpc606_5 gpc555 (
      {stage2_4[39], stage2_4[40], stage2_4[41], stage2_4[42], stage2_4[43], stage2_4[44]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[5],stage3_6[9],stage3_5[13],stage3_4[13]}
   );
   gpc606_5 gpc556 (
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[3],stage3_7[6],stage3_6[10],stage3_5[14]}
   );
   gpc606_5 gpc557 (
      {stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[4],stage3_7[7],stage3_6[11],stage3_5[15]}
   );
   gpc606_5 gpc558 (
      {stage2_5[30], stage2_5[31], stage2_5[32], stage2_5[33], stage2_5[34], stage2_5[35]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[5],stage3_7[8],stage3_6[12],stage3_5[16]}
   );
   gpc606_5 gpc559 (
      {stage2_5[36], stage2_5[37], stage2_5[38], stage2_5[39], stage2_5[40], stage2_5[41]},
      {stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage3_9[3],stage3_8[6],stage3_7[9],stage3_6[13],stage3_5[17]}
   );
   gpc606_5 gpc560 (
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[4],stage3_8[7],stage3_7[10],stage3_6[14]}
   );
   gpc606_5 gpc561 (
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[5],stage3_8[8],stage3_7[11],stage3_6[15]}
   );
   gpc606_5 gpc562 (
      {stage2_6[30], stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[6],stage3_8[9],stage3_7[12],stage3_6[16]}
   );
   gpc615_5 gpc563 (
      {stage2_6[36], stage2_6[37], stage2_6[38], stage2_6[39], stage2_6[40]},
      {stage2_7[24]},
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23]},
      {stage3_10[3],stage3_9[7],stage3_8[10],stage3_7[13],stage3_6[17]}
   );
   gpc615_5 gpc564 (
      {stage2_6[41], stage2_6[42], stage2_6[43], stage2_6[44], stage2_6[45]},
      {stage2_7[25]},
      {stage2_8[24], stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29]},
      {stage3_10[4],stage3_9[8],stage3_8[11],stage3_7[14],stage3_6[18]}
   );
   gpc615_5 gpc565 (
      {stage2_6[46], stage2_6[47], stage2_6[48], stage2_6[49], stage2_6[50]},
      {stage2_7[26]},
      {stage2_8[30], stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35]},
      {stage3_10[5],stage3_9[9],stage3_8[12],stage3_7[15],stage3_6[19]}
   );
   gpc615_5 gpc566 (
      {stage2_7[27], stage2_7[28], stage2_7[29], stage2_7[30], stage2_7[31]},
      {stage2_8[36]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[6],stage3_9[10],stage3_8[13],stage3_7[16]}
   );
   gpc615_5 gpc567 (
      {stage2_7[32], stage2_7[33], stage2_7[34], stage2_7[35], stage2_7[36]},
      {stage2_8[37]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[7],stage3_9[11],stage3_8[14],stage3_7[17]}
   );
   gpc615_5 gpc568 (
      {stage2_7[37], stage2_7[38], stage2_7[39], stage2_7[40], stage2_7[41]},
      {stage2_8[38]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[8],stage3_9[12],stage3_8[15],stage3_7[18]}
   );
   gpc615_5 gpc569 (
      {stage2_7[42], stage2_7[43], stage2_7[44], stage2_7[45], stage2_7[46]},
      {stage2_8[39]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[9],stage3_9[13],stage3_8[16],stage3_7[19]}
   );
   gpc615_5 gpc570 (
      {stage2_8[40], stage2_8[41], stage2_8[42], stage2_8[43], stage2_8[44]},
      {stage2_9[24]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[4],stage3_10[10],stage3_9[14],stage3_8[17]}
   );
   gpc615_5 gpc571 (
      {stage2_8[45], stage2_8[46], stage2_8[47], stage2_8[48], stage2_8[49]},
      {stage2_9[25]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[5],stage3_10[11],stage3_9[15],stage3_8[18]}
   );
   gpc615_5 gpc572 (
      {stage2_8[50], stage2_8[51], stage2_8[52], stage2_8[53], stage2_8[54]},
      {stage2_9[26]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[6],stage3_10[12],stage3_9[16],stage3_8[19]}
   );
   gpc615_5 gpc573 (
      {stage2_8[55], stage2_8[56], stage2_8[57], stage2_8[58], stage2_8[59]},
      {stage2_9[27]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage3_12[3],stage3_11[7],stage3_10[13],stage3_9[17],stage3_8[20]}
   );
   gpc615_5 gpc574 (
      {stage2_8[60], stage2_8[61], stage2_8[62], stage2_8[63], stage2_8[64]},
      {stage2_9[28]},
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage3_12[4],stage3_11[8],stage3_10[14],stage3_9[18],stage3_8[21]}
   );
   gpc615_5 gpc575 (
      {stage2_8[65], stage2_8[66], stage2_8[67], stage2_8[68], stage2_8[69]},
      {stage2_9[29]},
      {stage2_10[30], stage2_10[31], stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35]},
      {stage3_12[5],stage3_11[9],stage3_10[15],stage3_9[19],stage3_8[22]}
   );
   gpc606_5 gpc576 (
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[6],stage3_11[10],stage3_10[16],stage3_9[20]}
   );
   gpc615_5 gpc577 (
      {stage2_10[36], stage2_10[37], stage2_10[38], stage2_10[39], stage2_10[40]},
      {stage2_11[6]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[1],stage3_12[7],stage3_11[11],stage3_10[17]}
   );
   gpc615_5 gpc578 (
      {stage2_10[41], stage2_10[42], stage2_10[43], stage2_10[44], stage2_10[45]},
      {stage2_11[7]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[2],stage3_12[8],stage3_11[12],stage3_10[18]}
   );
   gpc615_5 gpc579 (
      {stage2_10[46], stage2_10[47], stage2_10[48], stage2_10[49], 1'b0},
      {stage2_11[8]},
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage3_14[2],stage3_13[3],stage3_12[9],stage3_11[13],stage3_10[19]}
   );
   gpc606_5 gpc580 (
      {stage2_11[9], stage2_11[10], stage2_11[11], stage2_11[12], stage2_11[13], stage2_11[14]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[3],stage3_13[4],stage3_12[10],stage3_11[14]}
   );
   gpc606_5 gpc581 (
      {stage2_11[15], stage2_11[16], stage2_11[17], stage2_11[18], stage2_11[19], stage2_11[20]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[4],stage3_13[5],stage3_12[11],stage3_11[15]}
   );
   gpc606_5 gpc582 (
      {stage2_11[21], stage2_11[22], stage2_11[23], stage2_11[24], stage2_11[25], stage2_11[26]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[5],stage3_13[6],stage3_12[12],stage3_11[16]}
   );
   gpc606_5 gpc583 (
      {stage2_11[27], stage2_11[28], stage2_11[29], stage2_11[30], stage2_11[31], stage2_11[32]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[6],stage3_13[7],stage3_12[13],stage3_11[17]}
   );
   gpc606_5 gpc584 (
      {stage2_11[33], stage2_11[34], stage2_11[35], stage2_11[36], stage2_11[37], stage2_11[38]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[7],stage3_13[8],stage3_12[14],stage3_11[18]}
   );
   gpc606_5 gpc585 (
      {stage2_11[39], stage2_11[40], stage2_11[41], stage2_11[42], stage2_11[43], stage2_11[44]},
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage3_15[5],stage3_14[8],stage3_13[9],stage3_12[15],stage3_11[19]}
   );
   gpc1406_5 gpc586 (
      {stage2_12[18], stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3]},
      {stage2_15[0]},
      {stage3_16[0],stage3_15[6],stage3_14[9],stage3_13[10],stage3_12[16]}
   );
   gpc606_5 gpc587 (
      {stage2_12[24], stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29]},
      {stage2_14[4], stage2_14[5], stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9]},
      {stage3_16[1],stage3_15[7],stage3_14[10],stage3_13[11],stage3_12[17]}
   );
   gpc606_5 gpc588 (
      {stage2_12[30], stage2_12[31], stage2_12[32], stage2_12[33], stage2_12[34], stage2_12[35]},
      {stage2_14[10], stage2_14[11], stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15]},
      {stage3_16[2],stage3_15[8],stage3_14[11],stage3_13[12],stage3_12[18]}
   );
   gpc1_1 gpc589 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc590 (
      {stage2_0[1]},
      {stage3_0[1]}
   );
   gpc1_1 gpc591 (
      {stage2_0[2]},
      {stage3_0[2]}
   );
   gpc1_1 gpc592 (
      {stage2_0[3]},
      {stage3_0[3]}
   );
   gpc1_1 gpc593 (
      {stage2_0[4]},
      {stage3_0[4]}
   );
   gpc1_1 gpc594 (
      {stage2_0[5]},
      {stage3_0[5]}
   );
   gpc1_1 gpc595 (
      {stage2_0[6]},
      {stage3_0[6]}
   );
   gpc1_1 gpc596 (
      {stage2_0[7]},
      {stage3_0[7]}
   );
   gpc1_1 gpc597 (
      {stage2_0[8]},
      {stage3_0[8]}
   );
   gpc1_1 gpc598 (
      {stage2_0[9]},
      {stage3_0[9]}
   );
   gpc1_1 gpc599 (
      {stage2_0[10]},
      {stage3_0[10]}
   );
   gpc1_1 gpc600 (
      {stage2_0[11]},
      {stage3_0[11]}
   );
   gpc1_1 gpc601 (
      {stage2_0[12]},
      {stage3_0[12]}
   );
   gpc1_1 gpc602 (
      {stage2_0[13]},
      {stage3_0[13]}
   );
   gpc1_1 gpc603 (
      {stage2_0[14]},
      {stage3_0[14]}
   );
   gpc1_1 gpc604 (
      {stage2_0[15]},
      {stage3_0[15]}
   );
   gpc1_1 gpc605 (
      {stage2_0[16]},
      {stage3_0[16]}
   );
   gpc1_1 gpc606 (
      {stage2_0[17]},
      {stage3_0[17]}
   );
   gpc1_1 gpc607 (
      {stage2_0[18]},
      {stage3_0[18]}
   );
   gpc1_1 gpc608 (
      {stage2_1[24]},
      {stage3_1[4]}
   );
   gpc1_1 gpc609 (
      {stage2_2[21]},
      {stage3_2[8]}
   );
   gpc1_1 gpc610 (
      {stage2_2[22]},
      {stage3_2[9]}
   );
   gpc1_1 gpc611 (
      {stage2_2[23]},
      {stage3_2[10]}
   );
   gpc1_1 gpc612 (
      {stage2_2[24]},
      {stage3_2[11]}
   );
   gpc1_1 gpc613 (
      {stage2_2[25]},
      {stage3_2[12]}
   );
   gpc1_1 gpc614 (
      {stage2_4[45]},
      {stage3_4[14]}
   );
   gpc1_1 gpc615 (
      {stage2_4[46]},
      {stage3_4[15]}
   );
   gpc1_1 gpc616 (
      {stage2_4[47]},
      {stage3_4[16]}
   );
   gpc1_1 gpc617 (
      {stage2_4[48]},
      {stage3_4[17]}
   );
   gpc1_1 gpc618 (
      {stage2_4[49]},
      {stage3_4[18]}
   );
   gpc1_1 gpc619 (
      {stage2_6[51]},
      {stage3_6[20]}
   );
   gpc1_1 gpc620 (
      {stage2_6[52]},
      {stage3_6[21]}
   );
   gpc1_1 gpc621 (
      {stage2_6[53]},
      {stage3_6[22]}
   );
   gpc1_1 gpc622 (
      {stage2_7[47]},
      {stage3_7[20]}
   );
   gpc1_1 gpc623 (
      {stage2_8[70]},
      {stage3_8[23]}
   );
   gpc1_1 gpc624 (
      {stage2_9[36]},
      {stage3_9[21]}
   );
   gpc1_1 gpc625 (
      {stage2_9[37]},
      {stage3_9[22]}
   );
   gpc1_1 gpc626 (
      {stage2_9[38]},
      {stage3_9[23]}
   );
   gpc1_1 gpc627 (
      {stage2_9[39]},
      {stage3_9[24]}
   );
   gpc1_1 gpc628 (
      {stage2_9[40]},
      {stage3_9[25]}
   );
   gpc1_1 gpc629 (
      {stage2_9[41]},
      {stage3_9[26]}
   );
   gpc1_1 gpc630 (
      {stage2_9[42]},
      {stage3_9[27]}
   );
   gpc1_1 gpc631 (
      {stage2_11[45]},
      {stage3_11[20]}
   );
   gpc1_1 gpc632 (
      {stage2_11[46]},
      {stage3_11[21]}
   );
   gpc1_1 gpc633 (
      {stage2_15[1]},
      {stage3_15[9]}
   );
   gpc1_1 gpc634 (
      {stage2_15[2]},
      {stage3_15[10]}
   );
   gpc1_1 gpc635 (
      {stage2_15[3]},
      {stage3_15[11]}
   );
   gpc1_1 gpc636 (
      {stage2_15[4]},
      {stage3_15[12]}
   );
   gpc606_5 gpc637 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc615_5 gpc638 (
      {stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9], stage3_2[10]},
      {stage3_3[0]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1]}
   );
   gpc2135_5 gpc639 (
      {stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage3_4[6], stage3_4[7], stage3_4[8]},
      {stage3_5[0]},
      {stage3_6[0], stage3_6[1]},
      {stage4_7[0],stage4_6[1],stage4_5[1],stage4_4[2],stage4_3[2]}
   );
   gpc2135_5 gpc640 (
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10]},
      {stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage3_5[1]},
      {stage3_6[2], stage3_6[3]},
      {stage4_7[1],stage4_6[2],stage4_5[2],stage4_4[3],stage4_3[3]}
   );
   gpc615_5 gpc641 (
      {stage3_4[12], stage3_4[13], stage3_4[14], stage3_4[15], stage3_4[16]},
      {stage3_5[2]},
      {stage3_6[4], stage3_6[5], stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9]},
      {stage4_8[0],stage4_7[2],stage4_6[3],stage4_5[3],stage4_4[4]}
   );
   gpc615_5 gpc642 (
      {stage3_5[3], stage3_5[4], stage3_5[5], stage3_5[6], stage3_5[7]},
      {stage3_6[10]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[1],stage4_7[3],stage4_6[4],stage4_5[4]}
   );
   gpc615_5 gpc643 (
      {stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11], stage3_5[12]},
      {stage3_6[11]},
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage4_9[1],stage4_8[2],stage4_7[4],stage4_6[5],stage4_5[5]}
   );
   gpc615_5 gpc644 (
      {stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17]},
      {stage3_6[12]},
      {stage3_7[12], stage3_7[13], stage3_7[14], stage3_7[15], stage3_7[16], stage3_7[17]},
      {stage4_9[2],stage4_8[3],stage4_7[5],stage4_6[6],stage4_5[6]}
   );
   gpc2135_5 gpc645 (
      {stage3_6[13], stage3_6[14], stage3_6[15], stage3_6[16], stage3_6[17]},
      {stage3_7[18], stage3_7[19], stage3_7[20]},
      {stage3_8[0]},
      {stage3_9[0], stage3_9[1]},
      {stage4_10[0],stage4_9[3],stage4_8[4],stage4_7[6],stage4_6[7]}
   );
   gpc135_4 gpc646 (
      {stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage3_9[2], stage3_9[3], stage3_9[4]},
      {stage3_10[0]},
      {stage4_11[0],stage4_10[1],stage4_9[4],stage4_8[5]}
   );
   gpc135_4 gpc647 (
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10]},
      {stage3_9[5], stage3_9[6], stage3_9[7]},
      {stage3_10[1]},
      {stage4_11[1],stage4_10[2],stage4_9[5],stage4_8[6]}
   );
   gpc615_5 gpc648 (
      {stage3_8[11], stage3_8[12], stage3_8[13], stage3_8[14], stage3_8[15]},
      {stage3_9[8]},
      {stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5], stage3_10[6], stage3_10[7]},
      {stage4_12[0],stage4_11[2],stage4_10[3],stage4_9[6],stage4_8[7]}
   );
   gpc615_5 gpc649 (
      {stage3_8[16], stage3_8[17], stage3_8[18], stage3_8[19], stage3_8[20]},
      {stage3_9[9]},
      {stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11], stage3_10[12], stage3_10[13]},
      {stage4_12[1],stage4_11[3],stage4_10[4],stage4_9[7],stage4_8[8]}
   );
   gpc606_5 gpc650 (
      {stage3_9[10], stage3_9[11], stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[2],stage4_11[4],stage4_10[5],stage4_9[8]}
   );
   gpc606_5 gpc651 (
      {stage3_9[16], stage3_9[17], stage3_9[18], stage3_9[19], stage3_9[20], stage3_9[21]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[3],stage4_11[5],stage4_10[6],stage4_9[9]}
   );
   gpc606_5 gpc652 (
      {stage3_9[22], stage3_9[23], stage3_9[24], stage3_9[25], stage3_9[26], stage3_9[27]},
      {stage3_11[12], stage3_11[13], stage3_11[14], stage3_11[15], stage3_11[16], stage3_11[17]},
      {stage4_13[2],stage4_12[4],stage4_11[6],stage4_10[7],stage4_9[10]}
   );
   gpc606_5 gpc653 (
      {stage3_10[14], stage3_10[15], stage3_10[16], stage3_10[17], stage3_10[18], stage3_10[19]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[3],stage4_12[5],stage4_11[7],stage4_10[8]}
   );
   gpc606_5 gpc654 (
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[0],stage4_14[1],stage4_13[4],stage4_12[6]}
   );
   gpc606_5 gpc655 (
      {stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15], stage3_12[16], stage3_12[17]},
      {stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10], stage3_14[11]},
      {stage4_16[1],stage4_15[1],stage4_14[2],stage4_13[5],stage4_12[7]}
   );
   gpc1406_5 gpc656 (
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3]},
      {stage3_16[0]},
      {stage4_17[0],stage4_16[2],stage4_15[2],stage4_14[3],stage4_13[6]}
   );
   gpc2116_5 gpc657 (
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11]},
      {1'b0},
      {stage3_15[4]},
      {stage3_16[1], stage3_16[2]},
      {stage4_17[1],stage4_16[3],stage4_15[3],stage4_14[4],stage4_13[7]}
   );
   gpc1_1 gpc658 (
      {stage3_0[6]},
      {stage4_0[1]}
   );
   gpc1_1 gpc659 (
      {stage3_0[7]},
      {stage4_0[2]}
   );
   gpc1_1 gpc660 (
      {stage3_0[8]},
      {stage4_0[3]}
   );
   gpc1_1 gpc661 (
      {stage3_0[9]},
      {stage4_0[4]}
   );
   gpc1_1 gpc662 (
      {stage3_0[10]},
      {stage4_0[5]}
   );
   gpc1_1 gpc663 (
      {stage3_0[11]},
      {stage4_0[6]}
   );
   gpc1_1 gpc664 (
      {stage3_0[12]},
      {stage4_0[7]}
   );
   gpc1_1 gpc665 (
      {stage3_0[13]},
      {stage4_0[8]}
   );
   gpc1_1 gpc666 (
      {stage3_0[14]},
      {stage4_0[9]}
   );
   gpc1_1 gpc667 (
      {stage3_0[15]},
      {stage4_0[10]}
   );
   gpc1_1 gpc668 (
      {stage3_0[16]},
      {stage4_0[11]}
   );
   gpc1_1 gpc669 (
      {stage3_0[17]},
      {stage4_0[12]}
   );
   gpc1_1 gpc670 (
      {stage3_0[18]},
      {stage4_0[13]}
   );
   gpc1_1 gpc671 (
      {stage3_1[0]},
      {stage4_1[1]}
   );
   gpc1_1 gpc672 (
      {stage3_1[1]},
      {stage4_1[2]}
   );
   gpc1_1 gpc673 (
      {stage3_1[2]},
      {stage4_1[3]}
   );
   gpc1_1 gpc674 (
      {stage3_1[3]},
      {stage4_1[4]}
   );
   gpc1_1 gpc675 (
      {stage3_1[4]},
      {stage4_1[5]}
   );
   gpc1_1 gpc676 (
      {stage3_2[11]},
      {stage4_2[2]}
   );
   gpc1_1 gpc677 (
      {stage3_2[12]},
      {stage4_2[3]}
   );
   gpc1_1 gpc678 (
      {stage3_4[17]},
      {stage4_4[5]}
   );
   gpc1_1 gpc679 (
      {stage3_4[18]},
      {stage4_4[6]}
   );
   gpc1_1 gpc680 (
      {stage3_6[18]},
      {stage4_6[8]}
   );
   gpc1_1 gpc681 (
      {stage3_6[19]},
      {stage4_6[9]}
   );
   gpc1_1 gpc682 (
      {stage3_6[20]},
      {stage4_6[10]}
   );
   gpc1_1 gpc683 (
      {stage3_6[21]},
      {stage4_6[11]}
   );
   gpc1_1 gpc684 (
      {stage3_6[22]},
      {stage4_6[12]}
   );
   gpc1_1 gpc685 (
      {stage3_8[21]},
      {stage4_8[9]}
   );
   gpc1_1 gpc686 (
      {stage3_8[22]},
      {stage4_8[10]}
   );
   gpc1_1 gpc687 (
      {stage3_8[23]},
      {stage4_8[11]}
   );
   gpc1_1 gpc688 (
      {stage3_11[18]},
      {stage4_11[8]}
   );
   gpc1_1 gpc689 (
      {stage3_11[19]},
      {stage4_11[9]}
   );
   gpc1_1 gpc690 (
      {stage3_11[20]},
      {stage4_11[10]}
   );
   gpc1_1 gpc691 (
      {stage3_11[21]},
      {stage4_11[11]}
   );
   gpc1_1 gpc692 (
      {stage3_12[18]},
      {stage4_12[8]}
   );
   gpc1_1 gpc693 (
      {stage3_13[12]},
      {stage4_13[8]}
   );
   gpc1_1 gpc694 (
      {stage3_15[5]},
      {stage4_15[4]}
   );
   gpc1_1 gpc695 (
      {stage3_15[6]},
      {stage4_15[5]}
   );
   gpc1_1 gpc696 (
      {stage3_15[7]},
      {stage4_15[6]}
   );
   gpc1_1 gpc697 (
      {stage3_15[8]},
      {stage4_15[7]}
   );
   gpc1_1 gpc698 (
      {stage3_15[9]},
      {stage4_15[8]}
   );
   gpc1_1 gpc699 (
      {stage3_15[10]},
      {stage4_15[9]}
   );
   gpc1_1 gpc700 (
      {stage3_15[11]},
      {stage4_15[10]}
   );
   gpc1_1 gpc701 (
      {stage3_15[12]},
      {stage4_15[11]}
   );
   gpc2135_5 gpc702 (
      {stage4_0[0], stage4_0[1], stage4_0[2], stage4_0[3], stage4_0[4]},
      {stage4_1[0], stage4_1[1], stage4_1[2]},
      {stage4_2[0]},
      {stage4_3[0], stage4_3[1]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc2135_5 gpc703 (
      {stage4_0[5], stage4_0[6], stage4_0[7], stage4_0[8], stage4_0[9]},
      {stage4_1[3], stage4_1[4], stage4_1[5]},
      {stage4_2[1]},
      {stage4_3[2], stage4_3[3]},
      {stage5_4[1],stage5_3[1],stage5_2[1],stage5_1[1],stage5_0[1]}
   );
   gpc615_5 gpc704 (
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4]},
      {stage4_5[0]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage5_8[0],stage5_7[0],stage5_6[0],stage5_5[0],stage5_4[2]}
   );
   gpc606_5 gpc705 (
      {stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5], stage4_5[6]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5]},
      {stage5_9[0],stage5_8[1],stage5_7[1],stage5_6[1],stage5_5[1]}
   );
   gpc615_5 gpc706 (
      {stage4_6[6], stage4_6[7], stage4_6[8], stage4_6[9], stage4_6[10]},
      {stage4_7[6]},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage5_10[0],stage5_9[1],stage5_8[2],stage5_7[2],stage5_6[2]}
   );
   gpc7_3 gpc707 (
      {stage4_8[6], stage4_8[7], stage4_8[8], stage4_8[9], stage4_8[10], stage4_8[11], 1'b0},
      {stage5_10[1],stage5_9[2],stage5_8[3]}
   );
   gpc1343_5 gpc708 (
      {stage4_9[0], stage4_9[1], stage4_9[2]},
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3]},
      {stage4_11[0], stage4_11[1], stage4_11[2]},
      {stage4_12[0]},
      {stage5_13[0],stage5_12[0],stage5_11[0],stage5_10[2],stage5_9[3]}
   );
   gpc1343_5 gpc709 (
      {stage4_9[3], stage4_9[4], stage4_9[5]},
      {stage4_10[4], stage4_10[5], stage4_10[6], stage4_10[7]},
      {stage4_11[3], stage4_11[4], stage4_11[5]},
      {stage4_12[1]},
      {stage5_13[1],stage5_12[1],stage5_11[1],stage5_10[3],stage5_9[4]}
   );
   gpc615_5 gpc710 (
      {stage4_9[6], stage4_9[7], stage4_9[8], stage4_9[9], stage4_9[10]},
      {stage4_10[8]},
      {stage4_11[6], stage4_11[7], stage4_11[8], stage4_11[9], stage4_11[10], stage4_11[11]},
      {stage5_13[2],stage5_12[2],stage5_11[2],stage5_10[4],stage5_9[5]}
   );
   gpc7_3 gpc711 (
      {stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5], stage4_12[6], stage4_12[7], stage4_12[8]},
      {stage5_14[0],stage5_13[3],stage5_12[3]}
   );
   gpc615_5 gpc712 (
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3], stage4_13[4]},
      {stage4_14[0]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5]},
      {stage5_17[0],stage5_16[0],stage5_15[0],stage5_14[1],stage5_13[4]}
   );
   gpc615_5 gpc713 (
      {stage4_13[5], stage4_13[6], stage4_13[7], stage4_13[8], 1'b0},
      {stage4_14[1]},
      {stage4_15[6], stage4_15[7], stage4_15[8], stage4_15[9], stage4_15[10], stage4_15[11]},
      {stage5_17[1],stage5_16[1],stage5_15[1],stage5_14[2],stage5_13[5]}
   );
   gpc1_1 gpc714 (
      {stage4_0[10]},
      {stage5_0[2]}
   );
   gpc1_1 gpc715 (
      {stage4_0[11]},
      {stage5_0[3]}
   );
   gpc1_1 gpc716 (
      {stage4_0[12]},
      {stage5_0[4]}
   );
   gpc1_1 gpc717 (
      {stage4_0[13]},
      {stage5_0[5]}
   );
   gpc1_1 gpc718 (
      {stage4_2[2]},
      {stage5_2[2]}
   );
   gpc1_1 gpc719 (
      {stage4_2[3]},
      {stage5_2[3]}
   );
   gpc1_1 gpc720 (
      {stage4_4[5]},
      {stage5_4[3]}
   );
   gpc1_1 gpc721 (
      {stage4_4[6]},
      {stage5_4[4]}
   );
   gpc1_1 gpc722 (
      {stage4_6[11]},
      {stage5_6[3]}
   );
   gpc1_1 gpc723 (
      {stage4_6[12]},
      {stage5_6[4]}
   );
   gpc1_1 gpc724 (
      {stage4_14[2]},
      {stage5_14[3]}
   );
   gpc1_1 gpc725 (
      {stage4_14[3]},
      {stage5_14[4]}
   );
   gpc1_1 gpc726 (
      {stage4_14[4]},
      {stage5_14[5]}
   );
   gpc1_1 gpc727 (
      {stage4_16[0]},
      {stage5_16[2]}
   );
   gpc1_1 gpc728 (
      {stage4_16[1]},
      {stage5_16[3]}
   );
   gpc1_1 gpc729 (
      {stage4_16[2]},
      {stage5_16[4]}
   );
   gpc1_1 gpc730 (
      {stage4_16[3]},
      {stage5_16[5]}
   );
   gpc1_1 gpc731 (
      {stage4_17[0]},
      {stage5_17[2]}
   );
   gpc1_1 gpc732 (
      {stage4_17[1]},
      {stage5_17[3]}
   );
   gpc1325_5 gpc733 (
      {stage5_0[0], stage5_0[1], stage5_0[2], stage5_0[3], stage5_0[4]},
      {stage5_1[0], stage5_1[1]},
      {stage5_2[0], stage5_2[1], stage5_2[2]},
      {stage5_3[0]},
      {stage6_4[0],stage6_3[0],stage6_2[0],stage6_1[0],stage6_0[0]}
   );
   gpc615_5 gpc734 (
      {stage5_4[0], stage5_4[1], stage5_4[2], stage5_4[3], stage5_4[4]},
      {stage5_5[0]},
      {stage5_6[0], stage5_6[1], stage5_6[2], stage5_6[3], stage5_6[4], 1'b0},
      {stage6_8[0],stage6_7[0],stage6_6[0],stage6_5[0],stage6_4[1]}
   );
   gpc1343_5 gpc735 (
      {stage5_7[0], stage5_7[1], stage5_7[2]},
      {stage5_8[0], stage5_8[1], stage5_8[2], stage5_8[3]},
      {stage5_9[0], stage5_9[1], stage5_9[2]},
      {stage5_10[0]},
      {stage6_11[0],stage6_10[0],stage6_9[0],stage6_8[1],stage6_7[1]}
   );
   gpc1343_5 gpc736 (
      {stage5_9[3], stage5_9[4], stage5_9[5]},
      {stage5_10[1], stage5_10[2], stage5_10[3], stage5_10[4]},
      {stage5_11[0], stage5_11[1], stage5_11[2]},
      {stage5_12[0]},
      {stage6_13[0],stage6_12[0],stage6_11[1],stage6_10[1],stage6_9[1]}
   );
   gpc1163_5 gpc737 (
      {stage5_12[1], stage5_12[2], stage5_12[3]},
      {stage5_13[0], stage5_13[1], stage5_13[2], stage5_13[3], stage5_13[4], stage5_13[5]},
      {stage5_14[0]},
      {stage5_15[0]},
      {stage6_16[0],stage6_15[0],stage6_14[0],stage6_13[1],stage6_12[1]}
   );
   gpc615_5 gpc738 (
      {stage5_14[1], stage5_14[2], stage5_14[3], stage5_14[4], stage5_14[5]},
      {stage5_15[1]},
      {stage5_16[0], stage5_16[1], stage5_16[2], stage5_16[3], stage5_16[4], stage5_16[5]},
      {stage6_18[0],stage6_17[0],stage6_16[1],stage6_15[1],stage6_14[1]}
   );
   gpc117_4 gpc739 (
      {stage5_17[0], stage5_17[1], stage5_17[2], stage5_17[3], 1'b0, 1'b0, 1'b0},
      {1'b0},
      {1'b0},
      {stage6_19[0],stage6_18[1],stage6_17[1]}
   );
   gpc1_1 gpc740 (
      {stage5_0[5]},
      {stage6_0[1]}
   );
   gpc1_1 gpc741 (
      {stage5_2[3]},
      {stage6_2[1]}
   );
   gpc1_1 gpc742 (
      {stage5_3[1]},
      {stage6_3[1]}
   );
   gpc1_1 gpc743 (
      {stage5_5[1]},
      {stage6_5[1]}
   );
endmodule
module rowadder2_1_20(input [19:0] src0, input [19:0] src1, output [20:0] dst0);
    wire [19:0] gene;
    wire [19:0] prop;
    wire [19:0] out;
    wire [19:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_19_gene (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(gene[19])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_19_prop (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(prop[19])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    assign dst0 = {carryout[19], out[19:0]};
endmodule


module testbench();
    reg [255:0] src0;
    reg [255:0] src1;
    reg [255:0] src2;
    reg [255:0] src3;
    reg [255:0] src4;
    reg [255:0] src5;
    reg [255:0] src6;
    reg [255:0] src7;
    reg [255:0] src8;
    reg [255:0] src9;
    reg [255:0] src10;
    reg [255:0] src11;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [19:0] srcsum;
    wire [19:0] dstsum;
    wire test;
    compressor2_1_256_12 compressor2_1_256_12(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255])<<11);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hae86b577a10332b71c4e953bae7e4d2188dbb11ed64d12d075ad124a0b3bf072bf033a233b25b5380fd0f997601e403ca85544f255accaf27a6554395f3b3e86148e011abe5938222362354b3878da2628515ae7b6086be459e47dad925ccd81267daa54a19c3bc1a699f6a51f9afa2fb5ffb66c8b3ae28fced12c4926015cd0b7dec7578b41a01af70f7790f8627fdb88982b6b026c951dc2869ad0367051fca4c5a4f178e5bad0cd4851c5965fc1fa4d0abf55ac08d6cc3143b4afa5b61366daa28904ef4f2080d2483a31095c4ecf65f4d3a4e89420d2f610378bc53b0578694211fd2f3365741c6f4b85844b517dd235958738f4478cfca0cd9cdd6da67907b509231b9eca98f6c6f68d39c16fb0ad1886a48205cb1cb0794109aa902195e172382af41628755360f22adc596aca1c9548bcef868383d0883c57a98abee2bdb3ea419bdba1e927a054e1dc80baf282988e4528c26defbefc1e06e08168e0e3b5d1489032c65a8e12a48304b21f677877f068a86b089c4b014a455834dd0a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h70d16d9cce1305661d807fd71aa4ce64d6baa3aba1767f54b7e82e68b19ceeeac76c7f6de887f4135479f292018fac54afa07d3cadba72afc0087f65de3f83e196ea7f3c48fc40f7c7174519d75eab75366e8f874179aefab98637d8ab7a0d1a97a53804d629d7fad943f621bfd0e168b524484c3a8a22833a63cbe57cf2a82e613725a387674410a73d1bc55f1aacf94413d8298b31aded6902b8652702f2b843bbd5c6e674ebbf52dab54488b40fb2170fdee91b8a8063c357dc1a74ff98b0c4c98eb346b48a45a2c9f0496f06c18ee23a630bf3734bd2d247c7fbe3b448b03f4852a1131614619eadf497792a18ecc1a3ef4c86614e89220dd995b5dfe2c6f134c8dc62a4c578673a860baf4f3d5049f8210c03515d984a0b73ffe45f19b9c7eeefc727809e0532a48c27c0d792fad3edbd2d3f5270937d461b73f93e445631dcb81c1213ecacfb26a3a1f7852044dbd9ff5ff64118884001df5bcf7c932fec960f5ac63a67cb18044765b195acbebcd18932e224ae87ee781b360166417a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'he70709ea0ad811199998d461316fae7aefc44f45a77f0be4380cd60205d013c3d816d875764caefdca5a40f05ce769d613169ea986f8fa978fbbdd066fee67852ec5253473324a58e1485854c56e296d1611d52b1d36797df23a1b66b252a9348ffc203899467f04f3c3e7ba4bf05653ba963d876162e3c90899073dc39dcf5518d263c461bdd698a5b9139ee5bad2fd2f356795bbd5cfe9165eaa5157b1e11e5ba8973fa39fb3746e2525e0e46c5c536094b6ab3ac1fdb884f07989b8ccb0761533ae5bb2dc71f2aecfac60c5254766f3c798063cc8258826cee21d344349e8ba6cb761faa7a00e5e921723b340ff95040ec9c3d3592c18ff8f48c97ae94d6df2cf73bd8cdd3a6ca5fe424e2cf1173cdd476e9c180fa0b93fb76d6c4e22e862602f5c2915045f692ddadafb710d44fb22bb5a84f72f49b0900bb818bb6cd365dac61eddf3dfb7285ed55adf0a7c936894f5afd177449287e11887b29acb3f0ac7a56d8fc49697a6340e38819ede28bde13671a8e7b805e933fcf719efd71aab;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h6fcec99f96c4310fac847d8b226cd44fe3f220d4b0ccc374e75e4bb6a5d467c60bede733e62033a6a70488d60abd41e4e54c167f9ba417d7b7a5f38584d824fa94edcd4ffc1cb5f5185af756c9a7db1a5bf9fa44c6c7a5cb4251968c9ab20fb3eb92ab2a13c5f7801129159e30bd3c6938058d9d9b62094e83bf426691336d16249caa1ee2673a60683b179b49eec0424a3f882c8b79f47b03b07cf14797812c82ae70f8d272395658ecef0bf9e50eb87b47aa2b36751393715122f997ee423f941247cf2791c2a654537e5419aca03d49073d2ed410e0c02bca5dc4cbe15de68d2c9743fe6e8580d457b83e9740d89b8d1cad0c26d17eb2a410c7c218758fed0c0aa90591c7c46633fc9696e9ab23255ea8558f9b85cc5508c39fd8057b26197417a6f4dcf3424f14599bec454b2a19fe5d631e2ce70a3aa00270206c769f52dd4edbb5decace2404e12b20c1fabdca80ca14b957f2696a937392ffc6a328077398256817b1ec1e30869bfdbb489f15b56da40bf56cc024eb5aa9860ca0829a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h97fb0afc4cd1912dcb148f32b91a3e926e80aa4f251cd157e96d37318ef99b3056737944384b556623898824989f05cab6378ab34de08887b50b89b8838df14f2f8cec5cd335e78f01f56e9c633e6f2b666e5cf26d337fbb996bc66a081aea856bc80c40ac0ca4a07b4e8a8ac0b36e38e8e19f7b72c63c1fac3fc41bcb234042f63f29bbb864c4d360459dc192d328f2560363dfffcbe6184287af38035abc8b03836b2aadb8067bf215f03ad3a462f002603dcf0bdb119a541f93ed4bf8acc7dfc36247e925b9e4fde5f549f5adee373b4b4129e802d4d0032e1a07e5066271182595108177f273dd5812ccbcbfb8a0bc3e86adf3244cf892644afbbff430772dd52d927ba70894d84003eaa43933bc06a84262cb5fc92f48a7d505e15a43b4cc1817e77315d0d80ef26272b6405964fa77e17d1a3cddb2a336cbd71ff21600c6ffb2594ba1c5adc6dfd6132b6d8c43c35562bdc3e7daa9eafc38a56409aaea8850f45637218364059f833b6b119ba1cd59c0391a2889ce8cd06a03bf7a05ce;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hb32acd24735e814b432b04fbdf3aacd3eec439f268d1d52148e79666e7a6cad767c834cbfe72bcd6069aa5a0b1903d6b87ff8b6b67dc0bdb857f444f95b7841eddf2a77d251f2fc44242c43c2f5e3c6434606b64919999526366925c5a930616552bf6004e1c32bfe63aad2998e84bde3508eb0b954cb47397a90471354706101cf0c37be0c5f96b61b652c3c3b4870e1bf9061c087d610ef0af288f1989503cf378f5c0562b9d7cf7a02223cf69f406a1afa8c4f50fe29d82f3bc5bdd197645b1a3e8f6b0cd66bd5639ca6c03a958bc0599c3394ade9ec5adc90015d69a331df8831f5d08970f4c899cada577e587b98f5e5196e01394bc296224a8766e858d5592a62910c9a29c7b61dae7f322fe032ba5a977e23ba8e2f6a03ddf0eb0e1d30254892dbb84115c270bb8e1239c795b246d3113d4a3abf932f2ae050f908c70448bc01eda1b576ebc74d4dd03dfd8bc5643dad897b3511d4a1045def91df6e858164e7ac101b89863c638ee52be7d693e8a4c268da10066e50d1873f84b9288;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h7aff74a6d9d19c0285609e6c25e447c870a24a47cfbf180d0aa6699c2cc476a65ae7e92aef176ae3c83a827a58a131491c330847071196ff48460102fa94e065c1e9d452348eb7a2f4b71c92f49c9f513c78f3744cfbf653f5853a4f3b97245e4fff32d06c62de926b89b4854e99fef2bf26f560d29e1843f3c570ba8f37d8d7fe2f8d7a0ebedae9e7d050b010d765a1182ab10eeb351bd4d7e46463d38a7ab322a2800637cfe91abea9baac2cd72bed0490914ad31ec0c10e5d4dd32cc4a14fcf863416ebb77afa50790b9a0f11d6e19ac8d956b1a9dbaff68ff5732c80a7dd89fe8a485f46e54cffd60672801039f6296d5a11a05e62f742970ce15d4250e9aa980cfb1fac4b9d928929f91cd6e2f1192b8a48f924601bcbf654f728127481d918c57338e8dcd6c7d538c11cc5d5c4dd9812c6ef6737408eb452a652b09636f9edb597e06604372e134efbbb6caa2eb16f0923f74773264b3aece5db39206cde3f968f9353a627e3004863c66fca970c87d5d4759b29e5ed78e18c58a5b913;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h4db567de08567c920ac49422db29eee5f9b8c48662857ce55aecedf3c9833d42358cb936cd35722d4246f0140b38dbe320afce0fde9489f8df9b7d61878e81f9a93d8747e291b41e04f77da91bb887ad61dd6fc11d0203f35e200f72d83cce8eb486c5087147bf46571538654bed3780417a0e7ce19db09fc9d081c548afdbd0c5f34dd1bde011c9f9e7ba5af3954b507d1fdaba2b8cb6bfff67b5743df3e4666043f28bd34d0014e67e9fefabe06d308e59c9ae98b26b0175f0e46e396963fcd6158ba2252cdf99e565ee0260b17a5eb571b3804e750c53c42546f763b8b22de8810c5f73bcf6ef2027cf232a8da8fdaf3cc2c1dfdf8b07bca5a54e8f1424cb7dff2243ec6b61d6706287861d0281474754d9a543002b1db9687edbf19c156fe774f85179f5f67a1af219f8f4088dd8878c745cf57505dd30d036768fdc5cfff079ffef685d7ace17ac5a38ffcde2c6f8706017bf69f360a5b24981af714deb3165aa6cdb8563c7b4b735a21e337d7b3b7d8fd029266791959f27e966ba5c93;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hcbb26ded06474da561903870ad92d4e386583f28340ef94587e40a782391338877430360cb09f7bce09200709a51306571d1496227211ae1ebd5fa371ecf66f7760c4fa01a2711dc5af95a315f9f331c99800ca909628357a216ed4fb8a172db59a34da3cb37e46b335a26477c5bf38dcd86e507e653d01e72710f07abcbd2446f424ce9aae821606610cd3337ae17403957da6d652f9633e874db453d994dab3439be41d4bfd610ef789f0d1165fd04fa5be6514f357af05c17ed01099ce226203cfa28a7f78bdb8610661439d6594bf25f9b079609f367fc4229127cabae8d4a9b3ae6ecf4842003075efa09e167bbc233efa086fa04a6b718c3eb3e012a9f9fd18f753becfc61ed533a3589518e05f42b589d0aae2e1610bd8efb47a9b8bb219abf49238af924941ebd00a0cea95ac81c672c24847287556f5e9afa1fbd29004710c0036391252a261210cd85d581731c090240807c0cfda7112586272d0b0ac0122807884b20f275a077a52d278e387e17e75804387ec961c9dd932b9983;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h1461a8d956359b7af12b03ea6dab5a0acafdb44057d10bbba6f8a4ac0827c42d2c4525c8673877737187b4b167845b72024ad493ba82658a2c9e297d07104f07e269eb712c73b4b170392eea55c3ef19efb7a4a74049b291a2dcd414da0b30959f3277b0a49e6c12246ab2c85b5cfff89c0c0e76ac7b679eb17759473a4b55b4ff78945953f4cbd59fb064747b4cc1b3c1dc849aa54176831773f41e48ced6073e06565bd5a237e5e32abbe6ee882c4dd755e2a33351854113b00205a11141e9c38331f3f5a622098100081322f04a57d085fa060baa8775dec339957f8fb5014d8b38cb31c7f0a17995504f807e4145dd9cd244a46314746923fedefbcb8bef1d31791fd1b713e9ae88db7779dc0b90c8bd5ac18f10ee46e95240cdd532c779d7fad67a0d96d22c1431eb9b1212493d746dcd8959b5cf3ad605aa7df7569a85629639eac3ed78d5fff750bb0cb0bc69148c7d1fc00166415334e93d7c22303494ba2257511115c50555224f522f29fa042a09695242cffbfe03c8240dd645cd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hb2c63a372ff660d6d7bfa02751983bef3e4ac52b8d363d96553359f79aef928aed13e44a39cfa31502ac637f76da06fb0411784e4b29e075360219ab62a81baf9c0243ca7fcd55b4119aca71a44f9418a85dd7f08dd9cd5a615cc72a4aea5301386fc353e8cc106f8bbab04618920e4d510a90af0b60ca0da91c28691da4e2a7ce1b9e2b33d237784a8a6a3847209f0c647af64559315d253e25140198af7f3729de36253d1b446d062c0d52a97ac37115988a2de2361b6e7f80acabacad7e05c14dc6501d69fde8050226aa52d92f6543abfc7bca88c14ac6149ba54b0407b1c3362f0eaf57fee6824fd5039590a493955cc6abc6f9cd323358022a1847dc815872fc0dd048d0292597315038c29f9f027c76535ab2250ed05438f0c8cde9372fa407b94f9dbd52a4ddb4a901b8a788e98a02de1081a5bc5fabfee478d4bf6f695a642b25b34082a170ae870038b9c182ebd145e4738a9c8dfc038d0918f657a3d727cfd899e427a52b93b4df18c5f6bd046afff8362be63a4a6cf2f874f665;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hda3eb219e3c04264a1ffcc17b4807f0dd5ba8ac67b4da7290e0b2ad01069acb4125ba3183af9a285e85b729144a15760b9da35e55d43f4c79ffb1aa4a9e2068385329ed0c99f8fb536715b83124308293651393b0fcc61d0c4074c7b69badb04103a314e5069a6a7dab5a964ec0e95163099c20dc7f15213e29b2e48b56fe525d2388ebf909ffe469a7f66d67f7886176fbcaf27342f8ca41878752d1226c9f6867ec0ec92fc0c3a8a79a9aa65794c4865eacb63521eb5ca5ade66b25df6659499e6d9ce0b38c2320bb27c8a80fe8f14a53e18f877002e864503d73b78ef803c0aca9f73e697284121d5ef4fbe81815485f2c301f5bc34ac57a48811b3f5a08d16e1de68c8cc03fb7e7afc5d9030271d2cd7b7881fc62d230a525f675a4ee45c7a9ce4e6fd297a54ca803df7dea7fb87a0372c618bca489f6bc2ff862aa1239bdaddcd30f6b6959a64323ae07738152a1485e8d8f135dfc2c01fd4e0acb629a80b1f1567a303c9d1d137e804e9fe038c3c8c15034bd510805dee9384abbec1ef;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h93625c9603bc6cf18653cc8913f098e337c75c8ba82f4772bcaef1a6e5460529de72104aaf0b19b880e9527c203ac9100532a5a96b8fdad00ae58d2d8d36347ffea7dec0abcaadb10098c40d1d10c32853fb3701b3058b5f21b195244e303c4e1e4530adbe7cf7b55026e8879dd851ab6e032cb65f1f9d4baeb73cf31b3ce5bd180eb71729aa285dc7afe7f670fab52e3e3c1e549040f03ce3d16852db518f08af1ca50b56b47c68213e4f47f2307b4856b60b7d58ad00ba2e2a900ee1b7d4749ce6de58709b8c1dbb20a028a4b8d914d2b3be2b61b61966e2a40727c347d7359af18d6d3c9110d67be643e70599ac696d1393e519daf916aa7533ddd3e1598e1929f4978defb92824796cd636fb8e79259ee1402c426f502b139f7831e8f5c9aba35236d7682a8b243e2bd74f5ef24ca94a1e2d32b4c35bc068c6aedbcbf57481877eb6ad6f96870929aae7d9ad3feefb67a245f19f85db7dd4e94e110e6bd0354bbe41ab057f7c2c25fe521d2f3d740b260a054fd0e0d9094ba68a86b38a78;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h52da3687139bda6db8dfd510447463b4eee76e1ff52976d8db75a7de129ebb6bbe72c4a066e87e5b86a78a916c9fcb242cbd1ab1ac47cb8e8aaa2342fc16ceb98661ae82aa27deb5facc7fedbf826a7f870ce77ea6671495c51f696d412f307313643ca06ebf2b9bac890057882e275d3f10f6e5426a30d65942fa358c55c10a8b1b7538dba974e025d335660cec27d5fcf7c216ff06188347783a8cc4a6fdd9b3cd9e357b1eda3c2e35c4f48084f00976239c578ffcd7b3f7c271a15ed1e3d6b1cf512f8b508a3d502cff7670a8bc474ec36a3090cb95924341701f048bde4a073c91c55b1de682617f3ca26823664a21d23e4244e1fd42d789426a584dc9fc3792a19765f2d6d4cd0fd847aae3f282eb72492bb3451cb04a7d5dff42d1630015b2465561055be3bb0b8a28f8c02344f4e02f1e2bf9b5eeca13f7ef1b96e9b49a607b1056997f628d37541ef47973a794ee3dd09bae00e9d13e1e4fa58f65014af975e9852e7b899f2741644b9f83ad9e4987b3345f80c62128ec04fe7989b9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h29dcf3cd2df8f2af4331b57e604ddc0b9da923823ef626dff532f9e99113215a58f4848d97ff2fa8642dbc0466ea3ee82f68e0a29541c4e86a16314a676115e113ef6a174c4b6dd63b16a175544f6aecf374dd17e831d7d103adfaf44fe2657b58c6567f25594f5c38de1607bfa9140db7b32f7f842019ca81f824a6660c5c42e1dffcf0d089bac9c2718b1f23904ef174f6a905feff3c77e60243f758b066f542de00ad94dcb440e41d2ca076c5ac0e92ebd32f5942ce673b3a948fe6c6a635dc44967475bfc60a70f5dee68fe22648e978f161dd51e4aa68486d8e5533d3209284b92f2a1c08568204a1fef40938d822f9b51154ace793b46d285eac137dd00266fbfb0088836b68061774e74e8045f64226aa7923cb6d2a2dd1ab5523cbd8ea89790811b1a0809453226974eecc182394e66cbb7cea2445d1e8711a79622e2aa3defff49f20f74fe42bf2e34234a2bfea65ff0c05f796af419ddcb4c6e6e00ab22193f6bcc21106456d9aca4473fcb27b8dd7f0c14d95d3ceabcc027159bd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h7afda2b17092a8d0bd87c5b74386ed7b254b33ebd8e87c43bcb793ff9071db0a8d3835df9e9f6fb9a95662ac16c5288d61c9fb2fdbf23ef2ea352ecc509811b66f6f2374f8e1dddbeabe5f441a0d16ee45eefe04bc8b3e8b29445f9ea4912c1c8346fd45a03f4d3ea9bc501dff2b674cd6b9a10ac9fa239be31d1ed74852bd70d630e02e59fcfe4db11af594b2c0e8e819c21bd879d5154e0ab604359bd402762ce15f285bacbe9ffd2c93dcb99edb4ee70594ebf252c344b7b7d15c1dc82e7e7bb5c12bdf155a7e5bcb35a73dad2ff73cf5ea23359e5eb5ecf0210dffbafc23c78c277ba9c0158a45d08495810d2a053e44703c058f5de6d8f8235c886a07ce2b031681c09d4048999d76fb5638c167b52923b37a37e8c7a5782125cfc439091c9c849c5a0d4845deff83c694c0194f46e400ba02834e52e751606cf756b864269bbd5da7afb99bc0029139dcb4df05724670e91d90262ae78298b966b0c1b0eec8833b6241fc915e762674420282acb85c7a554792114325da16f10432099b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'haaeff7f2f07d26de5d709352d4bd4344ec04a4a81a917d5c74b3c224f1f2419e1bd83a70259d85141ed39c45cf4143ec27b76242fcb69d52ece8e80085acd1ea57376d5e882be969004a03aa87ca53fbad53f893cdd7daa6db89be0ca64d1a3a782bc55ddd44d94aa2eacefe37ab335a332806d4c54b54e9a775c74145b0113121cb46222e21a5eacfa7e751536eb86fc3426d6ed22c747bdcd4a395efbfb2f65af4b293dcc06ac578a738ef200dc80b09d4b30c954f73a417a3b1f1308811cf71be9e4070f5fe88939f953958c3daac675e1c424505470e7815d7804184f55d55b0cc352df600588e11f0b27cc1af2f0500c2b43a20d0469af88668be02b8f32ef335297e752a59afc455839f8c3bf52b4844f94971121292b347f971f5cb8d71f5ad0b52f390e439d2d3dd34a9f9466ec2dc993bf43d3401898f92c9020ae31bf062ce430e3da27b6f4796edd1b49f9c0adfda0088a508fa7d16109c726ffca9e0eb5f39d793f3b23cd18031c79e98c1e2aea76849e257fc1bcee7605329fb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'he25f4ec33f7ae17bd024f9b784b76b46cbc2423d74192538084489f2d8b0565bad96ade4b3fd475c6e909d063bee273630c343be679528778edcd34207b137f4c240cf8386853e9bf701580172d35addbe38c9d6e3573ab076ba707047518f9756ec35395fe9349c3fe848c7f6aefcbfbbc29eccae497bd6c94bf1ecf401ade9bda476e95bfe2a8e9c7dcfc2afcd07a57d82d8f8670436e078fc5073bb58b517a40ac13ee48ecdec98c122a975d219ca77a18390d7522a83c4630597cce2673b6030981e26c0bd6963692fe5cfe2bf18e780dc4b907c2f3cff2b9fc4332ebe6a2c427169a46bb3a5dcd66212e20e5b81ba3bccfc2fa071d9481dfa1dffe102de250c88aafe8fb645f36d5dc48fbb700b8ae87019b16fd7d0cc2beaccc4bb17271365e77955a8cc9efb4b22462df49de884eb465e1be8de357e1c57978efb5268730aa942595d827feb64c2452aed16e3584cc2d8d91bb92be2ca89417f2877e2474dbc6eac88ea7f57e1b7512e75a162c08338b3605c398527c76449ebe7d879;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h4ed72f8c5aa8bd8898049a8a1ca7af887f3237582dedd0ce688303f35bd30f835434046167c5645f4cf7ea4e931fecf1ac720f0496ffc72bb4f833742f5879a4f73af329662834e256d993ad055de9c7c1bac09f04bb30e07d7752649979b02dc68696798c78f782ca4bdf0acd887777a277b1b4acc9b495d69d17df0f0db8d9b326a85346c7212c91076c2636d309b1d97bb41735d46138e15e08195426bbc8276a955b0aaf282583dc0e6f50274ee3f4c87fc79f6ab312b8ccefd8cfa70ecd243da70cab0aac7a73872f3e34c20916a46585338962ff4e45cb1e71bcc554731bae2cdaa95dc759958faef1841a360d68f051c9a814d5d3cbfeccf8193c3dc772948babb42abf7d9ca9801ffb22c04c931c7ef5ea32b82473b856e4bc2e23832938eb1bd4366718cf16f5fc5d28844e61c53b5b6e50023063fa6384fcb47781390a6f59a6c0311b760731fbc575dc366c4733aadb53f7b09bcac5e5dcb6ed324e4843f4ae6b26dd7de22ab74c1c7ece61b19ba61f23c9fdb1a70603bebf85d1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hc5fd4e9f8a48d106f2b30ba4806d453ade98d6779cf96e6dc8886635e4d678e0d4e554bbe13c00edf7fa38b274cd1eb0fa5421129020fc5642403488257b3afccdb422ec30dee1e7a280c1c0f9b2be962310336f86e1edd0f08a93d8a3385a769241892108c74f0075bc44cc662241c4e30e2e1594ae83d5f53d2a8e6a6319446df81db20dcb06dd282a595c55291d5a705be1953e70bbc514297c28930bad7e3147e35df7caa1d88d46fb2322ce2b7499b7188137094f85336ef190cb86808ee09c070d69c8917dc97c6fba6ac56d49f0d5e8585766d3b4273eb32d91168d058b6a3c85d5fc6a1216f5ae78b84cf8797a1945f7e3a52a3662bcc55cd2a8f3a034d7db86c218615dfce3120bce85fb57798d1fa9e9dc58748514c8c214156472cdce4fdf9e32c753eb66ae769972f72e3e9d46d542ca520f8167c3e428c97c9df4c06bbc397ba5b2bb821f90873e7a0722f62d8ae37d22454f5d59e9ce2345dc9ff5330d2295c6c19183daed103fee090fae0cd4b46c7b8d79ef5e531d6c1c8d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h4946aac8dc582112b00140540a69d5216a741d1c5b35a5a0f7bf4f680ce8c5bff296006e1483c6d1ac2a94cd0a382d254bfdc25451a8ad103f2a6a837a3cc6bb2a63413274a2fd109143cea687f9a3397605b155bb790e0ccb0499552192579d9d870fe3c3296bd2532282cc489b57962d6ecc7b7c4ebe5ed16ddaf614836195d28613437c8c45c75fab970d21e75f067f600721bbae643e0e9bf588c1e9e5a46d3a4292b1f4d330fe30dc0e9a024125e7ce7f3c23764de1c154b980f4389d38d7f55943ef1f4ecf0b207255dc70b95dfbe0e0fdd25f43bb52c1a779565de778e16936becde273ab9972473d6729ee020af05ed37ccd52a2f8d14541e707b0d87cc1c3c04d79b22503b13c4f83c9437e364dc64ba4db9b0646ea4266eb32d178d76eb3f31833ff290fde8530ea91a023016759fa142c2726176ecea04785b90501990691e414e367d701912e81a1a4578b706794e6fbc0e46709c3d36fd3225c79c3044cf5618c393a413eef094565c9c34f48a83e94783865c58802953acfc5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h20a8b33a7df19c6e2ca009fe277dc41b23adb49b6504121b2957c28050d0a1cdcf69b6e342cd0a826279fa2bb85ea8de6a0ec0862e6d5004b69ca7ba92403b83b05b663882cb81ab62241b32bbe0c51c5c0adaf8f76eb3e2594c4cb66ac39f18d4a11f9fd914aa912d0c386b17dfba6da848baa89038aa7c6a7ff5144e3d919a5569e8856e2d18b25278596e44ba27749671b37c4305dae1dcb64247ab7c568b927f853f2ea5f08dc7c80dd3ee50813ae822a756991db0f7f608883e74921aa40d3337e9bf0e0f85d94d2852a670c0fa7d0a1a83b05357b278bd24564797522928020d0bef2cb110e5a7036e283eb75e2b3251dff0113927678dc0efc2f98f4b97e0381853aab626a76dbda3ff04d98aec408195e41d73551f50d2491bc8569e5475fa070c2a453dafe817914c92136c8cc5a3eaaeb25578f81321e2c4e36ae34dcba9df31bf5a63ee3f25604fb52c63bd2484f2af673e775e1a1b856c2e2c78bce2616dfa7bc3f1e0839b9e62fb867e6108f1800ffa50687870668a56acb46d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hbc33a24376f5b5b4fd942e27377b8391adda0f956e8e614eced23d4ebca44851a5623b79df1d1474c3e364570f11f6c70b6750af8f10a34506b41dfb5c78b662bf42e555891a22e284173f363571dc0237a29341e90067bdae015e922b6fedc31869ba716cbf03d32267dcd75ea9286a4017f9e0f37353e5a58877cfb5e7e9d4ee0468726a1c5475a379c8ec2fd767210ff0f24fac56c6510b0b36b221b091fcfed7df2a7e85c2e4cdf35516e8439735f45cb6edd924589e59907972da9245cc6fd2bb66b525d586cefa65117eb612cbcd23534d86a8888077bae62aba99746d193a16f505a0452e8ef924fdfe7c258fb1d8fc409495b57f3c1b2b57f733e4c76e7c3931aad3e584d532b9de4adb6045aa48c04bb64fc2b962dfd3b99e94b6d555635056b89fb808280033a3e0143b5efc9912a69c4b0b82ccc1dce45dbbdf1376f8d4ef18ad07bfc43055a579cb0e1f37eb019843dbbf10558e65ae89aa4c1fde04fb1318950f0ed409660bc57e2b5774cf0c2f715e6fb5c6f46b8f3814063e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hab6bf24c3bbf8717230a440a01f07172c8bc42d8521370441f0d260c9a7dc9a9e1b239cccb6533f6a7cd3174ec6e3d4e2434b86286ffc8eeb7721fa2ce236c16bd9ceec1337c5a2e4a7ba5554aa6d5d67a0b87ac5d4d389953aaf7ea33fb0cc4beec091d038a793d56fb782937851257844f2461bf5daa355ee7b0969268a72726103e9a55d406e72390f7651c095996d88d916e859638cc6a19a7980adc7316dcc5d1feada629bcf7a007361af2218abf31f93558b1c0822127720f67ad23587b3fe833e04a8302b533c50e27daf7f918106d24138cbc9956f6820225c183aafac514145de8587e5ae687e9ec7ab9b0f900fab0b67e908115b2c2a58576aec6532f415e7b0c1710abbdc73a957bea8ffb89b2a7d9d403607467e5182807c4854a1078cd5b46db83b57c7906bf346043fb3ddc2ea4acee07d393e4134bfec1c5064e18c1a2e6e930e71b0ec004a5f9973f7987a1b47889593b7ab1e67471b89ddd42737943cb0a835eed7687f06a8015f0ad2d4269c48a6071ca48726e9101f1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h119ce4d97cc720281ca61ab1d64afc3793487e23d9b504adb8cdc88aa46d887ed5dc2ed2645ad3c3b4b3123ce3e2d85e20855eeba8241a2b3eeffed56b7b122a307e38efea6a8742b59b3f4f81dfa85920255fac19f356a8b45a2b168403d57d009303436e94fe742d1879b1540da533ba1c276dc12c8da99dd955f59776721daf386623b0f65a4b9d4322428b03429d60ae3ed1b87da93a59be6d2e74aac6a4883aa27aa9d99c25fc26ec177ed88a7d736a003724061fae3c0c2d7c0c37aa104ad92827f0f8bde50758e2c0cf514688d1b8de7d771f3b075d5fea9a6b4ddb22f1b06d4b54b3996e74fe7154be304cc49fdbc2dd71c033fdca328234faa32f9230966cd99f2c196131e1d5c4e4947ebd6a9c930b9321fae63fd5508dc76e3071122d99aee1285e678588de650b7c81fcc71b08a9f7a5c29fed09819556a0ac4e6662e777afdeb62b49145bfc4396e09095921647bff880216ce1bfcbec3f01bdb085b8ae697192fa9a10cc1fa9e9439f59de96f1ffc754e032cb11ae5184091b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hfa596d4d2d558b69f0829d289dc91b60d4a1958db057e46dbcef03e7634658a4223a41695724f0e5901282c3707cef20708a5242bccecd3736bd2b721d630c77ee1814d5c98e00f62cabcec78d5f5cb13d1e6c73dbba915b6c126654bbc34ee76febf11336ea8b00ba4a903c5b84bddc610bfa7d0a83571ab533419f5266607f2a25d4c0507f0f3d882c8acc87d82067ae91554a3c42ea65777fd123d7b5633b00b61cdfb7074e5f145c3fee1c8189f3e7fdb863f4c6ddea55aa20be9f4a955fe8f42511ecf71a0507a80905b8a63094021d237099322778ec2d6f8237e1180db90507bb6e0cddd8cc80d69af68934588f51d0c7fd1cb49817fd0805b0be14b3b4f7176d1b595f709166c7e4992c9871166b7f27ff3810dcfc5a3d0c53f55b57e4cab0bb684800df7c021610482af58390517e64626bc30abcc6989b6b50b659e47dd4c7dbdc2b9819b7a52ab9556fabe2b49ae39746d1933770e974ed7d7a1a10a1d7d8814d89f8f541c1079c1e29b471ec2d27f9e0e24c9fbcb5d20e25de4c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hd8a824956d68718f0c0f54f2d6e88aeb130fd55a7d7adbb2cdf744efa181c646aec7638df71c89025f1f3c2d6899a05a904c1099872cdafda17116554dcfc3ed6a25fb5898ee69cce8a2115bd691311072b140527240b98cc725a9aba72e963a67081696c1a416a41ce4f9a22900c56cebd3e48b1df6bb9d4bb649e730d986666c74affbfbf45df51210b0001be6d2c70e752c5a0a94a7ae0ae9b5d523f4ae38d8b6d54cf76e55656c7c0a25f950a6d9aab1fec7bd235441b26958f34cd3ac0eaa711e3bedc8273a884c6fc294325fed717a00414efa749562107a78e58409b908cfbcb8c8c5bccedc307f364dfd2cc437b57eedce9c7120d585693c55e45cf0d0bbfc89d1adc303e80a5f9ba3b789b0f9d70b1ce1e169d596372cfb6c074efa1492c9b48e81a915c4f02ef648f2406a50bfb36672827ef035b6e70c892d493813ea9f7d590dead1e835da0c763fe33b387def199470814d20610a3f548983267827111ee37940bdcc48153f1524007b6c827daaa6fa269b925d3fd221a21e73;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h96efd17086caa57a2b6bc427d9875fb9bea8c84855bb2024be19c89eaafcaf4518a8a4d0c512eaff60abac1ed247e4c4e266ae6b8a9eb8d5ef67e0a59ef2ac8a35d32fa4c282e3f316a67ab0a41090a68df174ce6c37ee91697ccbb71f7cf6123ee0fe36d8e88717dc78ac61cf0ced069e689f9b2701f786b3f17c355bd28b76c853a4adaac9d74c6dea8c11933dbb058c027b60a70636390dfe69a6c728def4eeafcfc1c329840f04d3768ec8d7cc5d99d0ffcbb4658143c5b92c3aee7e1dc0d2a8115f60761f9e1c92ab688d8ae0ef7cbcefec1c922802d46ef32a28b02784f9a88b439300606b0739191924da942458c3efbfcc82f63477c201126eaf95493c9960cc0f1241b3041a22925c572903d5b0ab7e41e26d53e1b0634bedb28815ca475a7c61b759afcf60bc61581822fa80e5f22db877deddc560300cd23bb651994a69a34d549f5ec80e758af574abf676fd7045b92788a2e3f436a67c1853fed16741c1dc6c876202c5ec4662f2a5b4ce765a0159b629b75059efe406d02c8f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h6516f7928413cf60bab2a6ef7873476368441c25dad99c721a428a10a11c2aeff591e892391e2870f5b472dad25418adefda6e2e5fba941f98e5973dd5b04f47c99fcdce7c7644ae389c4a481104555274631d38a17654b04d90070fa23ffa98aebe5910a8f7f75c2dc4cdd20da1df5a7485e65df22e655e42d51a525e1856b2301d8db417a8c49ced84a42df76289767882a0869bf5c7f67179c75b2779138b649b9d9fda6285f1a5ca70453152cab9af57fed219328287b25651038030a8c3699c19d3d07d41bd6ee904d181115902b34121a0c87ae36f9c2390a5e1cddf4fc534a6e4b4f84669c1afca08559435a97bfbca1f3e2c200af8f93a23e10881adeaacc4fb4d833aa0828edb8dd3dc4f290fe1b7b719ff69e7e3f88065792f726514d096f81fa18d3a143a30f7e987efa7b6ce8d36baaf7765ef36692a54c069425058bb09e34c5cb1de95af12a4a24eff5131f917fd49e4445a5069b3f658bbdb31b3de93543a1ca3b6834640aa43752bfa2161baf19027c0a508f51db9ee5c1e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h2c953c649a26fe67df56374e44c4f5a0445d70327938c1ac5ebd3d53366e094a8c4df062be943083a27f8ebafbe767b39fcf0dca5e99ca0b715d3e31f0500a5a8ca433b9533ebb618bffc5e935b99f5666c98d556e577a38fac4f130b6c79c51eefc49d48c2283b4391af1494d9c207694be241c5ff730ad431e37464d22d5026f7945dbf392a2fcbaf16ad77e7f841377ea660b3a026395c80f97dbc3f166d85f141c08cfe1fc72d3613e34a70ccac5b2fa618f9b3ef1dcac4cdf83376079d4171887295a205c301d3d3d3cf8dccd2d97907e60aedc354336ba0d4e9996a3418d91f0719408bc032263b299a5206a5359f0eb4b0311532cab936abc50f928a3800a2d4297bde9a275cf8e4d40121fe88d7e584014bc844e92db46fe5da1b14512056155f3fe9ffc66d276114190707b287e141a92adbd66efe73f8d0fe4afa76f1478c34812ca25773e0f7343b899bb23544870a8ca4a89783f15fbaf09c10544fa7e936a7443af30089d4b0dfcb190d59f76faaed1810e3e6db0464178006d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h3dbb5a0fea9a65e4d15948a6680fefcd651a19df737d2577091986e2247402d282f4c77b397d4a1f5ea3f532fc0607cd8fb820e31d8ab2ebd253deb9912096d4920b426e26ad2ceeac476cceae209f0b365d79d58ddeac302c823a9202587d2ee21189477c08a2a736ff794d9cdc8d44c6124311581187c410dbbf08cd32194a86003580d36ffa080007edf058f087da4abd20b005866b2ab083c281dd093eaba803ae5d039d9f20cf622ef1a7c69d5d998f8e4c06443c604f63ffbd063b124a3cf0e8f07b352306ff5adac712ba1dc770a58e6ff1504bf9b64bf345815b27cb4b44740ffcf5dc1042d658641af285cd2f527f56357878a66748be6d2431b8ce84817743bad3348442424fc9dcfdb32a96a3546529ef244fc2460caf1b820c5369cc6aedda24d89e036114a3f90e262a5b4e84523fbbc69896538464508892e6e9aedc85ab3340a95048b54b040efb7b18f2af15db1271c375c76477d2931dbb778c7d09f74bb68520c9fde47d6d7c0c11811e651a132cadd19c1fac796cb039;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hdb996bdf8c2699bfa05fd296d03af1be9635fb3955f5885891f530f585a30110873a72de50da69ebbb2120a19703817a880d898918eb52b79e8600a799f9c9af0ee1035cc32732c096c64645b75cdb6a019d143c87c8777d99aea42804c17026e5742e5bedd8e4bd641d8cf2b6fbc7ec884e398eeee43574a7e0262acb363534b99bc89d3c3235d4a755b952e1778e7fd399ae7706dc272067e4a88388fcfd0bdbf544816b115a01993049d9af42c61a552a09f31631ca1371b82bd1308b76e9cba58c3daa299ef818d37d07a77988be1b402fcc2e9a524a67a416099e915b34d101f443c516ebbe697fd48658cfcd2fdae50da36ab57eba25c9cca334fd9829ba207f8b7d7168897347d4cb4d1d5c2c50f1d65c9bb64560c36794e938a59ca024f5e785f2e48456ba568da6852cd1a128b0cde4805fb7870f2a4edba0b1759f44f3d36611bfb1379084ca36e26350f823a0c4269336273199fd1ec744842075a98852eda46dd153aedce715cb1e623e6ac5117d214c67f547a7bc099cbe7027;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h553ecc6c174a0355c75dfd9efe8ffde656abd5058e4d50076a75fcec659967150e0e055b8488a1a5b4cd9296502bef6fcefdcbb3ac50a53bc9701255e1b1fb2a5bd77543bb33c0f8818609ef8a7a70383edd89e42cc200e3696e7fea468808da0d9130534c7eb6869fb0ceb9d97d5d9e5ae4c8f359e544fcbbf417e6bd300ae84a629204b5029a1fdc5f59f38ef215967c971e05d84cea088b09d89c94c2b129500fbe69e987cb82c0672b2e2625e61c2223e4602f10c9621eef53cd95b0c3f371b22aa35746fbadb98e11b79b7ffbe7e46be6bbd5961a0820a3bab5725853998b92817c0fd4c9d8f63b668603a58553fd05a9aa0bdff58a0f24420817d9dc99dd979fc0865a4678bc96a4400385177cf4f60c599f84eb3a6bfba48c9531a35b6842605e31261c03cbcc4f34543082670cc93e6ce57fae385c3d8afc72fa2ad5668e66c1a1509837963370e278335e8262551ff1e52db56351dd56f4f4e210967bfa561df0f2a9b2e9e7539f9d116eb93682e7e34cbcc4dfc732c1b9233af331;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hd11f5c933a49f72ac988b44393f521fd0238fc19eec6d483a2ca19c98d38098582276910d7f8fb9247c7147f39c95e0933ff24538ccaf9b4dfe946a383dfc7a0c11fa8f5eccf68097c322e68a248c79c38ad537a29f9b1b2fcc2d8ae041142ee51e319e599eab9f5867584770d0ab55eb34ca57d91ab95d6ab8390e9ae9868063b7e484b7b9da86f4c079cec6aca23d955743e3f538efaa0e830eb2a6a2684324747ed6eebeb68de8dc7e271d0bc0fbcf5514310098ab7894af97ee7de3d8b4382d3f5f51b2f0571984bdb8c2dd22334f69712cd25c4bb67306c19960a5d254eaea6640381f1d7a59bbd02f7c2a43f53fefc8b4a934fb818ae9acfa71efead9c302bad12eca5eb3f826133ff97089dae70b26619a4dc10fdb0110c803fa0aa81dd668976580b20db707fe2d006bb787810cc5e0a5df17ea177f021086b1a964cc05f9adfb5e52048011c9ff12040e5e48a300ff222cf7888bb38124564c9b74211531d44ca7c803cf898b23eb1b88fda008b7c42a3aabc65964547a3154cf739;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h388ff3c125bb351e31b846531040d2a57682b15b76bdd6b26f1da8d76836e4541f844ea95ac6c179b77362bb026aa67db6843f950e03957285aa8e613114dfeb8f74b8b1a79ee4511c1f12bf3fde3a5eca54c67f1212da5fd48a6fd38a392b9ccb1e4406a885809cb9e7c6c9521c49d41937009cd076c383fc4649e2daa88a7d5fd09529988d83b9641d951fa60acffefe696a22dbacba97b76a2f9897e704689a199c2d6967c07a2b9dc7441c98b482ba26d05e27c8c805ec8446e4856e562f89204a5b63350810ffbb167105eb8046215cc5385a03ba67881dc3c6055f68446df2ecbca39a24b6419eabd7ea0010354810ab91a2810ca849ff52c8af7383d7d8ae40911eb865cc612d4abe056fa1041989d00cc7daea85f6b084102942ae77b103e8c3e6f250bf0fd6217e12231a16e462a6a9cd1de76b84731c337297c68d05cbaaf696d19e705dd68751640293bfb80d2e17e13dd77246c5042dd7c75cbacd3cae0cda3112853d03faa17fd526fb33d6fd43eb8e685a7581f87b4b6ade44;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h8b73c9afb89ad92faf1de1102eb5c5db9108bd74f70262e58914ffcb54525a78d2d8162c73b9e986ff48c8c35df3e9c78f7cd76e4bea942bf87d8c3073d7427671f4f92106826e2cd7004257e311b2a9cc4419156be3537f41877870fe3571e132e9e3a5a125d05719b3ece9da26fb79dbf4ccf39e51aa945c86179057d653e58123a63cc61fd801c7b2ffb6ac49a92514c542f497105ad0088fa21a4f1eb71999f8be482746dc0eb7fe738ba7a27157c762132948c2b6b12e5fc14b225024b6ccf7899b0a26ad2e58e7697099b202d6f4bb29fa87ebc648de0140d67b7a0d4c3141a2aa40bbbaee05967b0a92d61f0c8fbf55eca699cb6dc863d201dd00dfcf0986920bbf697804623aedc77c82e20149de0bc951e6a12b4997f37695d4788412cdf489c15a939309bd01f27b4e1b6382895932620171bcfc1a34a525bef283341009222d28f9d9531496c7655dcd57a9dc9613ec43f3ed1693f975570e436d9407bc7d26228a595393e09ec5d06aff1d6a1dcae0ea0c66c74f9654bae1b0f5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h480108f7a2ea6890f6e1a13bd9daecef37a6f4a8bf16eb97581c1d062340759fd80f7e5768fde697be9ae3d0a0fa4f584e3cc27773501599bc767eb2356c15eeab165b9c4ce33bb746ef4b7d3783fbb413e96133da7ab3586a035c8d99e82feacf38822fb6bdcac1765431646d1e0ac10384d26ff0f6c606f136aa5449191749bf8f258f98d3c959ea17c2d8cebc8af086f36237e113deaa502d57af8176b6b7270eb701d39f71f0bf5a9d624e0a931dd5584f7d3bc2eb103a84f5730c200f14ce195f87e8be1a609750d0835c1ae95f0d1782654cb6d87f08f01ec07526576db351c23d44942347264c26236c91280d8bbd24da9d498bea2b84896a5d6441cf2c1fe2630f7aa68ef1a8ac7992302cdbaaf131d1d425f07c8fe3bf248a358a94452b580eddde4c650bc9693aa028c7a34f71b0ba17e415d66a13e4eeed573a464847e87b8fc20bfe4bea7f330dbd47d436bbd2e54cefa5b9222c8ef2b66bf60787ec3d5e0aa3c186286439c7ebdbc63136d9fdc1f411af55c7302f3dd0171b8e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h8e501af81016c00a83559b2df0548ebaccd66580efc31d60954ade8b90746d3efeaa23b1595166f061b70e92f0cb052afc739f9d6ef6320e48dd823a7b9b18131623106715264f1502d5c00eca2b7c865837167419834dffc35efbf37c099091f454fa23850d1accf0ef0b41a7c15baaf0c95584afece69213f2a3719dc6931a8559e284eda6907524122d76743c5b4044cb8cc9e199f8b611d316555eb6035f25b82f6d850c858eb3c25e178bb3fd1949c840f9358ebee1e806cc74fb22e8e1e7ce5f6e929bb46d9da33a8fb2d90480b32e7e3c8eb509ce454a572d83c44f070e02013b0c2eb2e4dbb3d37edb073b98d43eaf9158da8aa8da50cca420c12b7679063f3c5eea4257b8ecf82c2b651cc9a6a7ba8c5fe2da2f393f9bde0bded45d884ede505a89ef455f0bb82d76d684eb7c7e51f6eb14415f02acfbd898a0578fbea1580f3aacda1f6b5199133848447ec8e1244357a5f75e8da8ed7f75c6eb201f92361de4824c1056dbab896de73fa95b130f7bf45231136148584eb50fc338;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hc4dcfaa55330e37c886488679b3fccfad08e7ac9c2ad96a4f14163cedc2965043bf0aec3db83e1bf1e38309505854af8be41b7e17ed8ddca4a30d31a8f1553638a75e258ef5a3232e59577f1ecc8cc82a550135f9a1a70481a8c6b01686d7961f21957706f1e87e0bc1aa9b9a971d4b1761deb7528a4604753ac39128127ebe1f04c49534bd03b23de1f6a4d5bc7c65a0f1e6c86cfc8cffa3af2b2fe6ed20fdb6d8284f12b3fa20c46cbe162f2bf047982167e78c69383b4041e8e3a276fcc8ed39ecb3c43364ac0218673fa9da4c7b007b46b7c5e7a8ac83cf3d2e5b457d8507a1c61f2b5a39de8c6e353c4c1714ce55279370cffe3674cb91463a862ce2d373262e419aab22629313687a3d10fd9f62c22c4fd92b9afdbaa2378dc33660f6748e13b343ea9ad619a3eab02b56c1ddf850e829534013b9331b729d67a15c81f2a148bf45dc53f9a1ac3fe7e257066a2e07012df074f781d71f42155083fc30e252eab037afd285bae9f9922c005d04ac21ab909ca4a014013ed483535f37402;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hd9fa935a296dd7787d36ba03c033d0a021b7d1ce528a6f81063c2688dc1fb4c809afd8713c4d82e1403857c1468f3713e68674ec3f89e9990111a4d2c41dca2ef8ae503917db6a4c0edc290695397aa0f9d9a0379e6f90b56babee6c45135dae887997529664d5ee55f2781405ca9510c0a1944e06a12b5cdb8752e8276052fcee824dcbd7fe802b46575b556152ba31c0c3380e9be264237c01c1a0a584e3bc819dfef23a10963d5316c5da940166cf9b37cdfb0b0fa4f3eb4689ad157590abe4b03edc143a4a3bb751247204609a1321d7a9c4f5325b1f834c53280e6b85933c44c4ef0d33b5eb5f003de964cfb2298b0fd22311cc9570fb922fffcac94f3d5164d0c2f39d97bba4b09eb30f424ff170ed1b463b159d4a74c383acf3358e577db5affc8815046a154bacabd2158b6afdbdc88c0e75fca8d6d3c024cabb6ad0d7c8e69c9cc22ea07f428ca2c3b2f2968e128da151b06de82b0968450aa8701bd8faf7b189545c10f33209328c84fd7d11df618aa687bf80cfd6f03f123762ab;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hc8bac04b9880ff9930e5bcca6ff0ec00b38026a4b0dc722b3d7eeb4549cbc8dffc60a794b29d846dda8d9f554f272188a00fba28fb25e6db6edb508dfd682b9c2244244c985c69dd4cd438a1cc35c45474e88d2fcb50a81a4cfc329a7b3766e619d17ab9205a45ea52ddd12f530279aabf5bb11f153b557b5bd8c0fa861f9c2321b1ffe80d2e55d543d86b28f8c02cb04c2e5e984f4a977dbc1538d4edabfe2004c4de9b780e06c66093a8c8d7c77a535f204e3e276aa21935bd6164cf0da7185c51e6874a55d65cb1d8aa39b6050643e83f9c91da29805bacb8f3b968b5f00c1553d70337c0af44f8994155bab4e603a9365c6780105b0c6a61722fae71190263a0b378684809708454d0f7ebec10dfde6af8d4a3047fcb7ea0e192e884de60b93a8c3afc9d9a08022aa25e10c475d9b3b9b189e94adfef63ddbbfb8dacac44ddea4285c0c873c636b743d1eaf6d0fbef2a70993c76bb5bac73816578033febd05c6a59126397d4a5677b104b3b3370b2f930daec8330ea4f1d84f5a163121a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'he340203317050f32fb763f1e3d1bb30de879c06e03044def35a232a7105fbd34b02fa6f00681a0322b97b7e43c8f29d3b83247367610fd44de3d0a17625a4f7f6edc832b00ae70187bb4454e56ad0716a9192e9c9415c01d29278f51c50c10beea56eba5a5c81cd76cbf28a63b54356e8c0db95e90ef58fbf62dd3fc06881aeb10b0f89f480b7429f7f7a85def9162f1320fcbfd301c4c97641404c2d8996f0820ef27bf1e27ecc7811bb55ad39883d0765f6de80053bdc0b4ea92526e48d761160bec79962383624c8b09e563d629d8e795583dc9a1c08ec4766394e385bca7991833e0a4da812499fb6edd0c2c30b72cb50d7204305001dc9d7325a1e30618f80e114a4a3c6579e596c031aa11a58d0a6994a24ef7f124327f909da9775a1f6812fe5f0111f6d5b462578928e1d8c535964dbfe8dd0181956e77aba5e2a3578a654924fd0ff81840f4e598bcb4cdead14b55d481cb9631c574ad3ebab4d96da9bd462bbbfd18dc1eb54e73ee046a2e66d3842bb49744b622ddff578200a2d2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h3ebf16ab218bc401a83b41707d2000a39809370badc420ed0c50903a5dd5c6336416b882ea9a4db23a3027245545838d61af00f0cdfefd5e40979d4e1f48fd7186db4f88a02a9af1bb004f91ee33d1e873000da0441184e0f53c2baf8f7911ffac477ae2e1eb2e65c5faf161c5a7638f72023e6c6cad6299253dca3b80eb8145f6debeae7bdd52538961dfda71b09c151c9bb726d8c023fe9176c9fb7a35edbe4437c9d8142b56ff7735be0fc49dabaa293f44aa8c28e0f20fa954f99ee67b5f866028480494a0880b14577c83a68fbfecdc64c9af208eaf729098dfa86399598ffa3b9a366a33c6474dbfc1c7af5aeb0ccc8a8a2ff81fe79215c4a60305f6c9a334ad4228c9dd4fec12c4251b89cd08f0ffa11520dec428df702b516bc807e951a2e18afb4f8e4c0d95559551a0daf97f4a4721a6dde647d4eaf2f934280e28bc457bd2eab551e7a2722ef7070e8b368d6ee1144653852baa455832996c1d38622f8a91a5b7f37b42dadefba855dd266a2a03263089b48c5e06630e2807c61a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h6d810dd873d7c285c0a4b2b057cac7eca5d7e1fcfa4027158483e7e5b1d077ff146a4efd573288b495fa1d70d0086df5732ffa87b2802e1bc9da2bec78b5461dbc21e86d3c4c2c76f3ce8c3980d35493db62f9a09e5477bf7a911ea80c6e08f70c6d6a3a9378c25a08df6da6f1979e782094f07e2457e6d69d9ea6d4e03a5d5311f6a6e372351fc785498c3e48254a22e1ba4db7c986d50bf22f4314263846a41708cea13a1b84ef48f3df6ec4192f9348e4cb1e8eb65ff037ca1cbde3b3b9ac5055492ac74ceec727d5a879610d597270eff9aa5fe3d16263638618bba3cdf38dcbaa389e64dbe5d2137a3597a3d65b4e46bd1388968ed92a8717db78a64dc362a54f67014231e8c71fc5214a74efa25b6cdb91def5516ffeed419fcdb4759e9e3d01bd8af13c1a1e2bade8814164b1f918c3197053b1f3025e3eadc6b4c5696af2c59319d32d1d47a74b7a32b5da5e6b71fafcef90a22ceff254d8c251538aefed68f1581f5bc61e49144a9e41919315e2f0baa4978e4107a512762c2718d1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'haa2ae4105963df74955dc66709d0dba9e85a32c98b3df733fed8f11eaa44e049c0d9ba2c6a0a9f9d34ee001416c8776a5be5d09d6c96637e5a60d44e27cfa7acc58284a1a557ea369fe044a29b3d915b4bbdc0ec87a5af04a2892287e540136a846ab12f1dc5268725091a42715dc998b314e52e520bdac66e0eb2f3cfb2e8b5d0b121507473f403741bdc7be0190e01ecf66d5aa0be4115d8006f8a59b8461785c58ef122709d43483a41a46c9582a701ab5f152719495ff83f5d8644fab0f3d1e7ddec88e22bffa584e0d7d29fdebef891ce34d2bf143cd206d9cda10eca1aaf562bf925a8ebee276fc8b46984cf83eab88d48d80fe414a5fa80af690bede68d2de7cecc3d47cfe6c2188351fa0bda24563b7b31d42d3b9a84ad7dce1679ba08b8d307af8b89ff5f9255086ae3b6634a37869e505b6e78bc4dd21a359a53a08780437e434c1baf57808c479f90c7b031d3430f920f20cc0374381fa6736fbc982f291b735f321bdd04321930e7664323ff9c452094c962df9ba8a756a4472b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h6b97cbef5ece802061f9714b75b1f946c8fc95d924809d7ec59cf6611067e09466bb7ab4d3fe13788db725e790dec56a5386835203761655205a7bd2edd2fb6d316d7311e5369f37548019a57950a27dcba955ac967e07c166a05e93fb576ac5acea297368e0081cce9a05c36793e7ad0a2ae83bf88be86b65cf51037843e3df7f91c32c7c7ef2553ac1fe37cec792fd20d06d5c4ad14cf7a2c8ef14901bd69ad52e75cd343b0d9f4e7d83265aef8dd4915473e509c8626046b67de11379dabca07298c8f918f4f2aa8d4ac21a88a581d29395c870b6fd0a0f2eed9cd7528acc5b79ab13ddbafcb69323691b787b1f40383f78b5efaaa55a1bc1abd4a3be41314439fed5bae2a9c69207de0b18f86c0deadd39fc7e8302a47933ce24e3757f9c63dd03fe9b3609183100e36a5c35a1e91fbb394f362076ba1005ed78faf4c6ca42a56a740a1227e7c2ee1dcba93ae68da705c6de247e1a4c6e0265a141e7c291658fe0c4aee2c04336ae0b84405afde2f53ebf97cd56054ee044bbb6db3b3f7d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hafc301a65209621d24f5fa5f42ec1a2538bfde88c2dc6672a8be69ac4fccd6de8d340721e417841d8e19699565bd97f5022b93f3f95f26955e61d9c954cc458c60a47c8f19c94ab951f6c82d79a89a38b19f906dab4a108bff800552b292e20ead0d9282137f215209730c53d7cc2c67179f82f75af73a32dc952f090de89e237d244cda9e0f3da47887dd63fc205f2d7f2852f1ffbe5b28340a9b9d498d59896f6fa2ee7855ffe21a8974a0fc701b70879b7c0c059b38dc12e69a400384622645c439774360011e14c75ce61842130aa6f150c817ddea8397a36e3592e63c62e80a198a29f302a3edb64e810a0ec8f2eca12738cc57a9c748bbaaf0aeb20403202a3b127debd478796cf0e7c4601373e251871c79102763307babe5c540630c7e02ed0582c47e3db270f00fbef7a496be87192603007c9566b86a0b35930a643ee825570d5921716b865ab2bab1a7358cde2292f19393b9c8389e2c0f14d8db6737ca862164835125f3a2ef5e7d0d53da8cc987afc5acaf47468329bb577714;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h83b684ff4e86585ac70d42dd873e8156a77e0c0fe9b86dfac4e36c83d9109be7ade17a0dc67ee1ffcffb25cfe86ba5ada62d0dc09f4d9712c6cd126db8cad63586359d7b43a39eca8832b493dd12d89a83a68d58ffd952f75051bd01c0de30bca8cc8524580ea473ae18e917dd573007e0e7aad1f1fcd89a3b67404f32c88cfb30a1c213d0aa9513ec5f6a0a90cdc1d0a9899de0eda07b83ecbfeaf4ef256f62feb487b79b20c050fa90d9b84069d9d5305d2305a0860b32d3faf3268bb85a85a828b18cce8a4f43974aba505d093ed158ce2221cf436dd1e60083d0c83ec1238b25b7cabeeb161123e85d124a7dbae4acd1d6dfe1c278378e526ca662aca78b766b8b12756f846cd8c8d20757eeaaa2531b68d56b100a61e9fbc13d192d3f978e6af8a819d33a240711eb25af4c6c75e8e52d97d16ab25156f3a4fcb68126264389a30ef98075b8e1a3e6260b63af86ed743507ca54b041141649a23ce24e66965a3e1e90dc850d73c194a9fa82b4ede18ef5eee8cd453452de451581cd9432;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h9b7cd235db6b6b758fc0c2572146e76ed6772b75775acefd8bd9639036836bc10707e91d47878aa56eb1987d7794da471c3129b2b7581dfaf0cd865493d151c673c9d307e1f0266fd01ba6347320eeafb2633bff2d93a632104868f4a56b97f993af08973cce9bcbae02a28e9a491f9e0e0e9cf5e025b724334063c20338bc7787359d8907b16e774ac5c00dca42a68616422a1c156f078c7eef1494b4bd4fe4b58ede2649afecd2201084bcf9aebbcd7f84c08eb47a38fc7b6539de13c5caefbdf4ceec3d2ef3a266b8e6f1b90c0061e3276cd7beae2ccf8c7dc0d40219647af391ca3ced9f558246ae4be5280054ab061c31d102f903a8b9bd0de65dab8add42297a48ce2eb746b724f5c571978188677125668e6a7c39895b2b805a960eb44bd22dd25f789f83a0a02c431f0e0406ed5693ddaf6f724c95781bae962084fc35c48fd233801fdcd1146b595189cc8fa832239a818af31506512457d2706abc365ae6c440dfa5891b1c5b829466c2b64ff3544f962eb2ba3495b31f3df95e25;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h751e8f569e592aa1de9d577c58ddb5c74dc9f514035159e48ca5ca8c07d75a67ea01310cb1b9eb923187dcc818a610e939820f7c3dc3c634ecd07e58ce698df74283302639943133514eb895e481b0b606df6bd4789361e269f19ef50ed24f2cb23ab9a7df1ab74028896ef607affe26e8e83e0531ad9f61510c8c153bad61b52dbb14048346319f5cc1a1bed3cc63cb687701ad9342b79cd8b69ef666d36f6b2170967a8cdbbc786aff0aa102b47f616c36b6551841d798039c006d3287584ceb3a9d663914a89b956a1b10e2a114f114f0dfb8e254b98d01989c58d79c901f4a1376531d7a1526380baf2a01958659eca2b156409a1d2556e708260f3604c704c859bda1ed719f1cfcbbb276c9cc3358d2fad1cf8cc9118ad3f12ad00b429f8a68de14706b87cb38cefed917772329e0713031a83a18f8c04aa16e6f783054b620bd1b8091e79878830ec16ce888047039e69d3267e80ea1bc11a21fdab1b7f60b7e5e1bb6ae0b39fec4dd1f0a58468b3e426f4e0ba761073dda8d41ce53a7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h8900c9d35360d731a259ddbee9cc5227e348dbc5f6b0c4ecb273b9e6a122b667f2248a6a5ac1c731a20d413db1647a804d5fcaaf6c1d7eebc4cae4a0744b7325bb75c3d83e40d7af42633edc494b04d858e576057abe62f6b2290919cf44b36d339ca974406f979095a5b7528922e37be0ac21f65c9cc49a41195e113c425d5f0b8511cfab411880f00b96d40d997d8594b3dedff07fbd35db1cba649528670b063636e873515207bed68f9801b33aab0684255f3ff3265c6a536a94d347d628502f2e0a340dad8138bc0871f4ae9498fbf5d2476bade27232944fd5e311e548fdfd66417ef88bf656fa6a4ac8e0349ef88241a9a6d07d13b51396e3dc4a5cc46291959b8897110ad1f638b7e62c0ab4f06f92d881c05658cf75cc2cebd2582efc8cfc91014e9663dbcebd03e6ae535cbdcc2fc128e73c94743198c6daf7afbabfbaf9fc041fd2bcd5716802a48ac72994aa99e9c8f4d817c6ef38cf83fd79b0025df90b5fb13c16b1480e35b23898174c7e031fd45abc078358cd81636dffc9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hb4a6441589dd2d78046a885dc150fd916979794f1a4bfd7562604ee49bd9ad53c312d6e9586bff2f81c6c4f91c594bf4f59046561c6d2276761a51c69e1824a3670a2eb3f98f9696f9004b611d318289b63680357312691500b92e88f18a053984759664e12d167470f5b3f44d0ff3b095415d00d38973091e1ce9eaf1501cd98d3ba1a5109ad222a4df80aa1870707a5f03e65897b686e1aa429f8d9137d4f5aa9e09a5e85e0b5d42b6639c39209abed8e35329d7ab2f4ea31afe0a01ccdccca101ea78c5bcb087b472d70d5dd30e3c6177bfac88836e9178c354d1db92f3e7588516c20fc213123a665d8e2a9690900f2c9d5b181082e9147964c91982b64f91fd259867eac31f677c8ef44984f8b008701bedb451d57beb5d3353c3ce12defae3394135f8d987eb456b4b69917edbcfb4ff709635c4470c462362d5713b2ffa24c018bf16e48d0f5866df92431993467faaa9f2e99fc1ac39ffd06f990a62a26dda832503bb9d17aca02fb314412647e931713490c8a1d66550d8ba279b37;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h134ab487727680c5d7fefe3b30db24ccb17f0d754b65899642b65619a77932f82d39b6e4ea3660a8ecc604b68fb8ccd0214f7bfa26eae5db8de9f115885a671f059275f356684130fc71ab1b19c74cfe1785ec9bd06b1c7342fa0feb0350b2aece2fd3d130bb2c80ee3ec38c0ec9e6f2c3716569de93d42b63e39ac00052ac3295f09c7beffb0f4d44eb6856a06c648fba853b4c6833b81481e1a6e110ceb23e13a0c334cf7b93c0d5f8dca65030071302d04273065e7e8755cc2c122ab26433c88228cfc8304a7711789e33f96970562e46eab198606f3d1223b7a70942be2adf979cb4573989263badce0ad6e0d03ecfd45b7785902358d0cab221b71f6ccc358d94447b6b5c2848d7f327fb557ee8dbf7b02e099b32fe522cfb0f0753aa902fa5ceff672f689255c2bff1a81e6a6e96302f5c806715780c6e77ae11e2f5c0de904ecbe01d019e3bb3d1a417cf30e6a8bcc7c45c03ff413c2fdbdd488fb11ee9d4c25556ce31e6e932efb91d29349ce532772e4983a2c998ccf0ea7601afab;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h78250cefc0f5230d93f596733c2c0c915cfec756450a6598da5b6214c8d1142928e1195b10c3e7877e6bc65d679ef4aff0801b82db357bc0120430294ed1137e80db2336156b76d9d78c89336e05f70a13c65c9674d57f9e2cc7e11979e130c82aafc565c9934acaed3f9c36088d0d35755778780307a2f09eca4ef12dafc45ff67fdb4a2d4805fc0b7b1241da51114aacdbf2a527311079286eace588987be85de222bff6c028f6f05e5c01f1de57ec02d0f4e795b146b13dc8d9daa04b705428a784ef8e3ea3255db2cd27c12ee7f0083f18df179cd7e53d37701d8534350b8631598405b27e5cb271035ba3ec21c6fe71a29161e0a788c0bccd7788a1e667e85715601f4a71db74ee3206a92b111eff3cf2c68935e53164944d7e333bd556221703b24330964b36f064170f9d5e7920f5d0998436d4cefcf8da1ca7766b56829d0e7aa2b22d17beb22766bd458a520d5c2a1e5f862ed7aecd439912486818e56b04ca88cac8c4ee8a3bc3162c1b1dc18b962ea492b5be7944f9c156c1cd0e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hf96bee2caa95b6337f473c985730279aded1b57ed40f0e74b307377fd6fb7dc4d01238ee4454fa8cfd8953d98fbddf9d1e67ae19d9e8c7773c0cb70f30e531a12fd0b78fdf77285a32fd5a3e45b890b6e123f5ca4e217326469987e1706d696d3b76ec32defc7104638b9a5c0846a8d16875c0c91187aa6aea4ea0b4bcae597f0d6d86d8908e1cee214fe23e6aed87beb70baff5d4324271224a51beb365e73a1e30be230179e81033a0a95c5fd7233af36a39b210834da315c46f2422372d27d1cf38176473da8ff55c4da407ce41f7e82d317b099922eb01d22cd033c0d718f66712eec6e0568f91e847c8af9290a3898ad46dbf231f44417a1607f7f6cab6536b18a8bbe3c3f482de9e3c4249c7d73c3071216ebce9b926a1978c24508158b1821739640593d67ad480308f4336c1fc450e0689c1fde63b0831bb70265e88481e61f2340e225c46f981e605113d7d68e3ebf5aedd60baa0326cb2fcb19987d5679851663cbb2b47d1dd3aaa3fe908c038c11fea9cdfb14ca30a11e9a02db;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'ha1efa792d270f038ac77650b3a0bcdd1ea112f34cff10a7ab984546f9c0b5ad0376957662da40288572bf387d1b52a3b094854fd10dd699c227ad4363bc166b5acc8c81770630a7b85521d5f0d8368bb1190452b148c9173f07225fc7de73fe8762fd15b4c63625c693716ef1234dd00e10bdbd33180e04b8d06dbc4fd04448f78f668fb9f64b5f8af7b62a3fd4a12e0e492331881c37b87332b5a0c6459b0472da14f202883a2fa14b254a0db7f271ee75b2ea8cdff310c6c4fb50090c02695439ffe1fb35c9e35ed8f171294f94efab91b8b7b7e36b1313d0c587ab297063a32cbee18b56efdfb4111081bee8decb33a9fb881252d4b84403e5ef8d46b37611077554aa11246bdad9c40b6023de9707d488a8ee9ba500bcafa6875c3ac596467ef4813f31b4be70ed15c5102cb463faa70656971ec5b1a3774ef7c2d6666cde0592d1fad030e8f21b5842924ef3ca06620cd08fe8e799611047c8268092c554b2c1d12b6a00d67c4e576ab33a47107224f19ce3547f23c1d99f5fd83ac2bf6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hd4f015be79519edf26f4523a22446fa91a9a3db9fcdc503bc9edc91aef77bc56d701b3598cb5b05314148e75099e7a96d643cd44d7f52aa3b18284ec7a27ba5b99bb1e00de74c35fd92c6b3890384e25ef976b7a4edbdaa50b4bd659f11b6108ff72275a568d8e265c35925deea51af492930bba0ab12f02d3d1faad337536886af592fc84bc23620005702f61fed8e2661e58393050af9ad5ff7d6f37ee6578686524b5f2c4b11db8e54fdc756482a9c8661d6ef071e40ab0c8c132ed78b23f61fc42b1230b04431ed1de7d99181e2979a4d1dddf548ebab185356bf1f40679d14a16fadfc0fc43528c8ab1f8b09c7cfc3d971ab59465fb4af55ec849c87556c5aeb5945717240f4eb3a9d25581cff75ac44c95f5a805a114ae40b1be0ea1ce31533370852eba55838ba7f5f4651259047bd510f24bb8a365dfd882a7bd47658d8edb10a4350f4c760db1042d469ff55486f9ae3068ea1508e37623ec4e75466edc6164a45a74494a71a1fc4115117c3636e5cbd9f5f596894dec2d1c25278a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h715766d5450bc596250befb7d5fefefb4d801c1c4e1497ba221d907c417ad80f231e3f6ef9366f21a70a64fb84855e11f55f73c23c277068c1455589e3def44b43f38af32815887a663a6f0536978287a23ba5a77bc1f7532d9ed2ab4edb0a4ea4e0929ff71262fe9aec09a3b9b319ae85f65140a8868028847bb5d8f8aaa7b9a8339c856a0f17722c180e7edd7d428ad4cc4d353405f82e3adbfcf0433e67b3303e09c1fb8cb4c626a77d2d6c323fe4655150af263b87ca972a29b060b8221c126ecb414af6cd3314b79d98dadd82688564c722cc24be2b6094d2e04f1deffc3395e6e4ef37668179a96a02271133dbce72e8044c391b4d62d11f5693e1b549e5e70b42c8524845539af113721c8aa3c855d4f26cd6ccd8a1aa4c0fc9ce60f24e3b953e27f88ed2868aae80adfd6d3c0b13667df5ae7e0c8dbdfe9c3f302cf339554e7f07b197043df1928aa10b323fa77e401f3e2c4e9946dc982d292c823c5b0a862b205628f08f91fdc8ea6d7d745ba7d0ed592aa43e5b9f8fce29b658c6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hac90c638fb77a72a67f561c1203b737e8d2e6b9dea95ee6337e0a7df9277ea2f6172f38856fecb432ffa3ebd28f6295100b7f4378737bf221c8b78d616c313bf87c1be2ebc680e409aa73dfed7c2011850cb29b734e3280ffef47e7b566322f2419fb35eb5c6edf8bfc769989fcbc3842d6f0f6a1f5e3d9027db3809e8b0d8e3b1c050b8adc938359a57c7fe64528549f920b2559f97efd99f4df3d1cb0f5eb78090642f24ec84722bf147fbc494ca9567f3818839d22a6fb3f67460db72f0134980852fe8ef608459ba4b640ccc971d7fb30d41074475c609edeac279712acb096e1dfdf260d3597b806b15278737376f42edfb9c60962ae15216e23ec1532c9f9e7bcb2bd8e828bcc7e25a5beadde1df58dacca42a82c7c20dc022cdd1021a30145cbf317f90940caefba624068cbecc6138e9db46360a8100c43736d66045df2c7e7b7ffee08132422d367559732bbff04fbc8975fc3e41c619e2f25763293b32a52f4b975cef10e11ef202e9f04675535a9b56c5dc649f08089bb09cdce4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hd37ea297c7ed31407129339972c1de4b79ed2379584f69555bb0c289d30c31a1086e27188b9059b56000503bb64191e23901f68e0b73db1813de3bbe2957efbf1b55f2551b0dbfbbf834f49a4ba33b4aee68315822619fff80e26d6b07f6feed4e1ed7279f2e4b99c86bc6c9a2552d5636994ba3189efa19533d2e2074a6d9a906286734bb4de7b3ae0c8d28c531a43ef2a1a857bb2950c998371a5fdd087cdb6bb1c9ddf4d752a765b08c68c1a8fc1d3cd0ded5e452a5e062c917cee99841c61059ac10e24b94db0ecbdc4d6194c9f39d603ab38fac061105722148dfaaed8bd28e0e722dce09c57966133b9aa0b01e41cf90aed4651b277de581e472e3d023845b0e81d36c69f6e3a0c9320bf4869be0c2c092fb0044ea1b350d2ba306b0bbd953192fddd7d5e845e6b7cc9e2d6cdfba41e42bbd450e18ee51fff5ec1eb6faf46a757dd22a8a1e4453c94ea2095f6f3a223629f963892edf114643973a70514b72a3982d90350edd4114ff52778c4f4dafbe0193987ed46b98c18a4127fc7b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h77dd7e98ae37363ed4bd769a7f04a240b91e9486e0f4cf6ebe2dfc054bb1d7a36e3d5b94b52a10f28035ce281aa4a4e89916042850ae92c69fdf542ee0f015a86033f4a55dbd704ed9530c4ec95b20ea1928f2c73de1db0f28955c0585886fed1719cd433163447674d52c532047bd4b81124df8c22d979b84d1fd001413afca32cd4d5b438aee44508920997183118ca1cf16a1579d7197b1c75e802bf2a23adfcf37423dd03a244d505d58742ee876445fa2c3dfeb7355a03ce7d499d8bfd4ad885f01009a420ee600cd2389e3f6bcc73c535a6b6776309da756847915fb995f1b3da0a581daeb2ca33776ff03cfe2104ff47911ff8bf3dd375a32ff31ffbb8bade8d141eb8842734c0ecdda9580feb553131e4a8278f636ef1c6f28c39c685dbefcf91e3816732e37b855f2f2464602d45b2c09b40cc98d0e34ed4249397c38ad90163241b5f9d6b34ba5f7571e581db73e8937e87a5880b2a5b0117e40fb2cba50461932a7977193b5ea72a6f408f3566c7ad38868379843fe5a0e758d50;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h3e779d69b6e45709aabdd87eef11fd2bb5bc4a748a039f85ec7f5709d5a1f3fd95ffcb21af1b7199259ae6fd8281dc89a504b6b6e6f2570ca73062b32c68aa39b60d45440dcc55e4963c49846e14a5950221d88086b7ab312876be10f334a376beb1000627fb1a1a412ca27bd9a3f9f8619a7015a7fc9abbf0f90000c4b3c10759a1518f2f74c39b432335723d668f0ff303dbac62f06e18e0990768bddbb93cfe670859a507fcabeae8f03ed95efc67a7f64350f1a1dec2d8a8663f0aa8cca39f5c42c5ffd772a3848f2dd065ddc2915bd8256e8acf03fb855d4466089ff0003f3a9ed4f2ec80f917a7814b70ffe645341a299c893e8c83f636e3f9261c6ceaabfa7bba6bda8e72ad9ac8440c27348339dc2f568efa86d75beab7d9875c1715fcef4ac6b3ea1d4af0d02676e61f9820ca3767ccf767b11d793c1eca1396cb611d800b6afedfdf047d0a437da07b311b77711058d9425e601dbb4c18f4ccbf001dc1e2f9edfeb2025038514a78a0abac5de4c96aa9efe602b954b4b231a3fc69;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h3caf24c04d0724f131229dc61f5d318165c559182cdd1d7737243c6d4f41cb3ec08f45564c7862d677ce411d4986f8da7b4ee3b2c74899db84e2a5f3c38fe6ebf7fd57095b7a7d9766e168b5a19148290404e119c294ba06394fa2739df9443bb64dd53ed8b1f9b287730fa233c81a6557376aee1828286e0b2a73d90f0b83123eaf458a5cc15c5deee9032f32caf42b172a6147f19007f5d2069df2755f2072a9ea39f5470872d3642be79aab408af8c128be36bf316f40e38de0f0cd4ce721f451af6bc19f04f4b00af0794eb63947cc3fea9572213412addac1e4392a944548fe802831f8ec52a293b319efb0871843df35a643aa6dc55f5a9d8919ad4ead51a6c36e5af0d510cec3012661fb67682edd149be013d3ad3ca85195cc956c6dc368081036aaa04941a48617be4f43e3433703563e90634cecae84b2f6e6654a1bf56f002acf3fffee804cc6642a18fdd7be38198ee1c3794aabdc0e8b3c9ad30886de9c776c0a6e692e57c0118906125f6ceef29b9586413a0acbf76bce8826;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hc8a489623139f9d93e2493964f0d92f7e1511c80778be82b2c2d492a9226283402c790f41d8687c29c65180407ab69baa2ae0e610eb65fbbc85892b5c794cba59a57235258102f53ef5307b4d5e41d8d785b20c2f2c6315707eba24794212a321563ef548667e90c9218e6b6838a496d807d451ef0c10cd9ad24237e1a114960d4557760579a2fb45993a59e78d6c8a0dff87055abda78e059adb9eec98a9da54047149407080cebaf204492956945e2d7513be16aaf667dd4785bb68f09f2066802139275405586972091acfc9190861d7464571159f8727ea080d247794f92bd85b75ea1e949bfb6114a3c336bc210a9f4cfe74ed6a7ff055a2b4ddeea2187de66a07a83e32749908ad4377c56cfed1ba2d02accb4480795af09c9195e14c0dfb14f3ef4c486801e37f76cd8c56b24ca4947045690fee5232354080eb55cc2e130ea3928ed90075ff6a8999ba284470a6792e7544ae364e9bd41423def938ee4d73e894ec9d42ee731fcc9a253df1f3d0cf2c317bfd600b803d8093c8c17;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hcdc810479394ac01851e72c9725fab2dcc2b2865cc2a2763636b4c69e2bfd866332e9249fd46f9264303eb9e8451765426487c827221e5a98f9203b4c98c6f5cda020fce673bc21499bc5c232d80793bce26ca4222f168057b8027d33a50e6931339f3ce189fd56bea5237044837ad71e0e36bd98b4e59268d73cdf45a4cc1294d7940ca322309620e9a00c207fea6f3c1ed47ab81be1279f242e9c5570a750d2093e014cd2c6318424d19d09604b44fb8faab98749ef348a2fa7674633eab903f5fe4be227d21dc508b03952415bf8f9c7c3f051a98f2480469f03d213b9bed1d6180dad3bc9195fda85c9823bbe8b8c0d9a94276b908d697b417c4e6ea4b20c72f32a932a7b75069ece995c7e2d09985ee9d320b97a1df2e38d8881d536178b8857215d55889547aa5e88c3ed7814977ece645c4863ba807a204b0768434b4c82379b605e662f363d39c97aba90a11e3e94b9f153ebe023c4c78accd5b81b02c769460a1782487cd72bcb3410736b24c50d4f5bda72f73cf1969580e14c6fb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hdbd6fb02b98854195ffd73872fd6faf0d213e59d8f1d424bb9713f5a3251511d5256d8df653fb8921883237ae3c212870eb2d483a7bd19f1b2a3654890a022e48a22616dac6ee7ed82f0fed182445bd0d724810cf1d72bec194d909414f5deb0a84fe80fbcfa63cf8788292bf42b104395b7d1aff528e59b8c7124379bd3b611002009cbb5722a58de92a0857785dbb87ef6ff043d21f4904494e3350b954ab5e641cebacac4ee44ac7b61680505d4a43ec7a97b71be18a99e9e6f39b521d09f60e51be3285435c0ae6521b10c1a91f48904ecd22cb4365c867cd5209be3e0cdd0c7b33c22e8bfe6c9bafdbae7729f34ebe360d9afa5f9cdde6d54edab5a5d26c2cd9d5af217227127234c6c12e4b3ecf6de8a186927ea38d6d7dda95f3345d39513b44b5e3c62b9ef6c47bc3584d260f0d35efe550992a6e920f1fad742dbe9fe0d5f51e10ace5926837fdd38faec87c98bf4806b97555b7a578caf5e9a264c00accc5dafd4c2f8f705b7048ea1055cdce9a79e77dd6ad0bbd7d742ef0f5c38;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h6700ca84c4d33528c0cd5d10f4811578846b9a4afd70e091b4b7936177e6dc032a7ad2144caccaf6e47dcd566e279d8bdfad81c37dd8af60bb7a28cb51e482b4e12531d379d0c415dfd9c3148f0198513f7963d5361968cfc09ffb5f0efb141f5aea0270ef51f8510a04298667fae9a16633392d294937949c2fde810c0c92e8a6e6c53ddff6bb15e7d762b924fc69c1fac3871b258b63bc0a05aa9b90ea433d8f48f0cdbeab1f4efe7ed64d6257ca9d8450dc954448cb8e9c27139ba1b0aa1cac930b774f2fd16a28f229d49a997b27f1e18bdeb1a6308fdac40472b54eca3933fa7756bcbc6acaadbfb0e795910d128b3eb4f9ef47d909345d5c3e9b7ef1ad05b578eba037d7f0c22bab05d8da06aff081b1639928989126ab9ae5e3d88d93d59431f68543f28685444869f3e9b6715a27b35ef7a08f5fcc2509f00a486f6a3ee45924b12564251f7ded29bd6b1053785731d163138a7444fbb7a1d726e5941d941446828f97a9241e02f10c7d6010fc399ebd209d45f635067b08d97d4be;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h228227544797c8eabddc7eca8017fc7aafe157ff4a0079ce3c56fb0782f26ce0abe7e75d2bdf517ef663d408a40ea41be400c2518836cb92b747c7ac1613a5476c3420c02bdd1223b980c0ccb1fa7b1dadf192a04b50548a8a55831b935b29d8087f6c3b217cc77cc1161028878a07df87546ac937990dfaa97ca6ae07b41e7b68403ef447407ad2f56d85921689a093d598dd3007b4b58007a510aa3da41280bdaa80d3d20f3927a6403d6dc3304029ff56c6a1299a751da6861a420358c34dcb44b6d8c8e9f9fef224d04adbe8a954869ecedfe77b22ac8c09a53ab5d54287739ac73a9ff6fff4b7c15d798715d9145ff76744fa9f12fb4d302f7dac5149974b0cd8cf57617c9e96ab46562e1e5697b82679f367ef9841fffb679982327e8ee3853c73f36b4a39f723bf835b890c46aca6be2aca7973965d6363be675577f6c9ac141c466edaea556f02a8d63556f43d3754792795f3f12e2a3ac6e37bf9d5f54e6e427d02a0b679be8a22273dfda2923fb02abc484d146629448a6cdc64b0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hbaae792647d2d2b34c989825a00e864a9a6faf9e3dcfe881a2d9923fd8a340dd985a53cf62b48995a2f483cb14f787330555a014bdae665ef8b15092cb7e97effd694264402438fe433c74788ec783acad7f509706489269ac953b7b52b6d744f1e4d6c593eb3b11d395a4616dd2a42240acc621808886717f79bfc68d45ee4a17c1d4e9d263655571a8c2db86a1dd1812d573ad4d711253d7883e76408e9729bd8827c348292e21d1591f2dd62214031556e5c0ae99d45985aad83ce443f2dd33df2e5bbfc9ad6fa064080d7fcfc58a2d5075d62e921c14724fd74b442addd7d6e68ba45a849d838b00073c5745dbd8efde60c6712b954f4e661475f885ea6bd97011b363fe1ec4ea21684362b48a7d84969ed72bd5bd7d90717245e702f197ff844f18b26dcef6cf1012870028381b089d6f423fb309c8dcb58d775aa71045f02b19b4f75609886dbe7da89fc3d0af6e85855b2b1ff49eca8a4a64ceeb6a3462c47fa1ff307b28dcffac4fae18da04ffc021411ee187e112b22f849f8f263a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hba7ea6e66519e5927aa829e8667333b136eb181a0c4df7f15a1859d802569168422f2a59beee6126665379414b80ad1f096a04a38d0b20b5c3f6786e72ab8ddd037e8ef7234d5906e876d6186e6d2dc151e24111864f43e867ff8c05db8972f45e20b58361752c3af8d2d19efd7dbf2cf4177775756af6ca69cee513160f4a43a3b28a7e3edabc1b267094a672c1e1154b61351f60bf934295f13f1f40d34cafa39a070a34851b99f4008d1139f6cbfbff8f7fc013328a7adeba5b641bb4d552e4b8a689ef8291b4c325eb286fef938ffb6c972d569056313ccb477b059c6cfda7d509dbf72b1408ec921120b029b13789c627802c631a44d6f8ad1cf602bb1047ac003dd3084e45a0098913d48816b046d106f9b672b914b8a49815f015cb59b4e10e99e4be3d665c9dbefdeb9b7aaa43b35df32eac83b2cffe8961ced4d6cb6970e10e874b7472c5d32f234e81776134dc2e2b70fd125dbbf4479ecc8b94fe6f83ebd3a6d7ec427abe9e2ea84e77cad9dcb343c82c108c82d8ef3b3bcda9d0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hf3da9c3e5033b26e3e61fed222fed274354bb4fe1f3276925fcac8d76ec90cc2d8c3a90149d787465884bf289b37b96d7186c450bd20de61c314a5ab2ac9ed6a3e95abdb372c3404dbba2cb4c3978dd8e8bf6ad313e90eacdebf01ceb434686a10c11e3aa556aa74464a2b5776cfa49926d502fb5a753a29ede6c531cb4e1cc1912b06a71884d990f957bef83e1fcf64702a0e0a7c0e53c4b148f2167f5da06571bdfe5b617cba659f020b3e4f9db177b4a5d91abc5a83034a05f659efe335a81a60122ae52254f69a56423d252063e8abbc711943e0a81ab4e110378939047d39aa991d8c0720f495190a7a681ce369bc93f8d0778b88d63cb146d8efae5abeed2bb8bac00f5117cfb868a69a7ececb59f6f0772fc4f4b6e5ba94c78acdeba6f012ef1e297d962ef19ebe775d3427d07aee3820c7727ba2bf28435a278fcbbd9b5ceaf6a0b702547bf33a1deb19015ec2ea237fd5627441387ef96d9068f3fbc44abbb853dba262ba037aeb29df43b022193294b9ad92e72d26f1c7ed3141e9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'ha7a967c9146a785d721eebb19617cc0288b11d19d2b68208904749988eaf1ab02583fc49404990884c9b2e9a5f013063dd7e29fb0f9e9b78e6ee10572138b32aa8ee938f45347131596741030a23b0569dd13132698af43ac9596068e653e367e3cc9e235dbd1ce33454f1ee9b84275d648d73b3c98f82568e24dc83dcd8152093217b61e7f93a74308df5fe9858027a0e3ea30df6fd9695df81a47d576a2060c0708b316e017d2013529e691ac8c2d935b771b218018b0826aa0a0fe68dc6b4a7e9815d10f6f96719be827f37a15f955352a00dd4221fac5a157d6f79614f4fa5c0eec38009739a212900942fa99d3bfd20689d02cba4e6851119915fc017250b76aa4b2cff5f411e4a3c66c93e058255a53c8e190bb9cc88b91f500ce8d723d36452381e4aa9b29d30f287770784b74e71fbdbce21420799a6f36640334253f9bef3f9eb130a9d49c25c202c00300c509c0b758239e7bf7be70345e2d9b9967dde5cf9646e55e5385866f1eb5828e20f16967178c2bc18ce9fbb8ba9276dbe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h1c413c6fd92c0979ae6db88ba6b552559b6a54dd52e3bd26e09daacc0fea36316e4fbb347dfbe8eafdf1b0ad0ab256d5f960f341a53c066d3575000e7507919bb4adc6953651622eae6cd82c71df2af7b14a9c92ec71f54b0d3d6c6c4e2129849df419ab0df8d796058ab37d00ce1a4fea9fa116976b41bf5af809104aad744d6ff8f2d8b62a84a28c3b7143edbc5cfe040928210a35cef1263ee6bc9245930a731b4401abdc842993632d934081d764b78a52a96bbe41f7dcb695ccf2b1119b966bc1160e768b7cc225e6c8fd171573f8d46843bcceaf93be4046461cbddd047c0647a359551e8dba10114eddc29d2540aa5e576b0804fc5c9f7650fb41a4a6a74c7657860c4c7709a5caec79e2c97b72d030e1dfa08ae1c153f9546b0d3f2bd52a2bdf1653a68c46f3e5353f3c0475d56f046f6847da8963233c04a72017e2ba62af5d6d6604cd85814ca0e1793a56631a41049ce626ffbaac4216ce8403cb81b925e2c2dfe2319fcf72638a88d76aaf1fe5cfb0a79f9f42e7c4d34a726b84;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'he891040f85598a9bc2d6f9905f6b1371fa163b6bd9dd87e2d91cc35ba1cd24bae8585732f5d755a9955c88cba48bd9acf2adefcb24f059c88985f9b65838fdfd2eb4caf4148989137a21e7ff1a1bff1a42595c183e68f7f955cb150cbd4c483c910d57663a0fef99b2f13880686b1baffdff40d5167672de1fe036ac7e7c4d2436227b1900b6275e9740c5434ccc19b6d5ca993fbbc8dcc52a16036920eae1bd04e79f424ab6ea53bf4e8b2caf5e11a410afcb37fb668ae1808d27bea0a8058caa6f207e81fcd634440bfef43932b2588dd5fc31f55e1e1da9fc5091348218727ac96101ae4cb569939c9a0ebc2a881d096a533c9781337b21bed6117143e7e5d048d3d85ea248e12d1d8c12bb0f1032793feb0feede5129e34a75d2e598604ff19e865a944d8d6a0a94bd12c4ec4c7cd80f7a530e7d16fd3dcd90e298a13ac7b011313c60d7dbbae553a4126fe155dfc1d34a4354263fd09b04534f03fe0dec525612c517c6cba2110afaa45fffa1d15fc36a0a946329db27199674e84fb288;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hfe504a6fc64433422a428fb6aabf37eb0926e1c4d371d06ad68aefdd1134d60e42e3ac468bf3a85e239f848e4ae0a0e4616e1dea46c27f84b5454d20fd4e06474606ae5e6a87cec066cf9a67ef39f42fcd00cddfa1df5c0daf9b5a97c730eb278e19530374ddada48d13c7c16bd139f9105b6aff5db4064bbc5f1fc32c90be330f08d866276d01c9a5bee4748e21963fe5d629ca9d3a59046c7a6d57d97606f18f89bfa1618672c8c11903ef7aa63ad1b5a2cd19a362268b7104267f7bc055b6473dda3fd658214491d0c2add266e008d9da63f8f86745cb6e2489e606f02a40d3de402401a28cea38b6b58be18abc46a3616a09093cbfe09a0cb4dcb58d06e5d42d23ea1ae7efc35a9417c6417e660ff650dfcbc76798b5caf43f66893af9647bc085ec29a7524fb5dad434d52528517f26ed93e6f0467b0d8eea4a12f91d8e00cdd4da169150ccb415d93cbc4aecf1b2a6242291b97add776185d8d74af9f76de7309a04c9923f68e7de0cc0185aa91fcd3b6a7af9e0d8a943cbe3deb9d2d9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h66c87fecdc702ca54aea10bb66c2d2cf347297464d3ebbd7d68ce7386289e6ac284be99d4d0d3ff9dd62cbf0e3b92147522c26aacda6c5881c831b50bab4b9ea66af5b3c73fbd13bd037cc58833177569f50f03d7486f201c293a644841039d0360191bdf86ef42894c1d0d47753220d454235213ffc52d88e7bff1995e9a71737c7c09d81140404f778a652457178d84ec75eda7a24258507d3df36c2bd6d652af2764607f50704425b902503153938fdb1252e20f1062bed9cdad6b09cfdbbdf5334d7aee2577bee479ed6856d30e17301d4407d1e6e71c9280725bc70d15087f749f1300603b5754345e9a30b46fe4ea186423e10f32890ff9b32b998a8d0a36f22b211975291f36c5f7a4bac03218f4071ed1f2cf6078488963fe0e916095502681b428970582de80668a96a01c86cb64c12200bf78e3ef2273b83a953894b16a8814b7472b11625d40a033ed7fd768ae121092c3d502af9e32c96e50f861db448e0afcd2150e2787ddbcf9414ea5692c9624c3d56f216e7489b433690d9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'ha03c0b9acdde6f254060ade628ec34d8be01b88bc0b10d85eabcea9622559d457ea1604b983eace659eb5317a3b496cda485944a75abe0f9f7bca9da9d78eb6196698d753c7055a407bad322390e16cbe73af5ace5fa7844ede90e187d61519e6f64f7aba55b1471cd95696bcdc76b55cf5e1b3f56b5954b9010f9a98dffd5064c180f808ee148b8487e580714fd0d31056a92f34e64f46ad543929a22f6c7a61fdda7730b6ae4afa50bc3633cf1cc991734fcf7c2771eb7864151492730aa02f4551516374e5ab1a865c629c834c8f0e1a83fd90d7f50a9b944e4772844d5f41779351ef04a506abbef4b4227519a87b62c34c8f79dea1e1ec8ec3ac050ff9b618a721ac9636358d74122b974eca7bcda4bdab4d45328c72d03a404249d21f4ae882009757f3876b21baf45f35d575596a34c5e43bef691e6fed081459205c20e7e6c9f3f6064960b30e55b86ddfc9776aecb0a446140794f02c5e4703de5ae0804e7ee56475dbe7b8d34177dfdb5331e9ebb539fa80272e00067b937115e92;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h371ff7d591dad77eaa1fba16d284a7df8632d7507d4e76ddd403db9a20dab1d6308c3dfafc8f1245e9d8af75c7e7d249ffba43959543e8da8b2104c1edfb1e3bf2ebaea47567177558dc121ead8e533d62b0f8394702b9db49fe2337b97d797d0ca51e90b033997577121633947a9abdb9347528a9522e011df685810a14f988242713937cf0df2bfc59ed320778b4b31e8b9768c8449cf1374677e02bbcfb7ee8941b633d41a2c8f41fa103e615eb01b9d4aed8c37c5283e76d5fc9b2dbf4ce8bb443a4cc118ab9417a2c930ce89cabae02ff9f169c2aed7aba2ac79852f4e553844a009f1c4742b6a03a9c1152efc188c28f4d73915b14dcdc73ca924f6583c510c81e56194fb0a11bdfd067aabf44d93abe65e828284c4115a429ff2e9c0df27494f599d906eb057b3680998bfd9868b21f26054892cf9922b0b6c0d9b97de39513644436e44a4cd675bf175657b1b61896865615c04c13549bcc226ac8de2982b497de0fb8cb961ca29a4f33ed28dfb35325fd31383d6a645ae18a174ecf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hf88819ad0caea0e080ff214e80d2534026fbf0ef13d36d20ed9fba30a1d0fe32caed7ab7995df9ef850951ed11174ea682dc837f8e7d3158d3697cefbe13a895d8f7a01480bca40499f15b901a1720cd805c2973af29ca8fe0e7eb21cda86211329865560a119d1bac7808ce64e5bb224f319b76edc099d249121779a3c58dd8db3f73152143c148036f376c9ba12a8545037c0361dff39dda38db1155cf703dd885da8bb084b9f4e91c98ada5af8826797699a9c5b215c11694b2c09721acc993ceaf41ace54f4f46a4dcb0e68ed8bb899e9b9ac025f2118d56d5c782274a55306fb5387861c95e61e99562596d20bac68655cc4a43182a31f31f7b89bd02b102051dda7e022ed2d5ec2cfcc1d39f65d16f6895815989bc3a125c8bf52d746e8af03945a9c01615fa6e021883744a3fbca074608e9cc7ed3e6d01f61dddfeb8b97ab7892443628ea6f1616240e7244e93261f1493c1762510a49e100236ec810356b7c783c9688cc10264c687d511631cb0e05f6c4889de74c0e0fc0ec4f51d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'haa51e57910e500856bfd7bbd5f89955902a9b7f027133481ac9543bc1d2fc649d1b7b993b88ed5d1155c4c250c2f8687efa3946480bd13801d1c2ae23769a96ef9be8095300ba5cbff571960a67e10dcd0f8100af246c96a44b594c71079e8c4b774928c613e0491fbb2ba1f2b6ec14b46d54840d4f5d60223066a1239e69bdff6f80e30acc9f439c24972040be966db4c59bf0cdd6076b0e8ee429529ce3cd843de6efec49f4d4b77816a2398f2d484fe35d31e65045608fe4c5364234dc39c421bdf7383a0970bb3d89b3336a4c969bb06fec466a725306da91887563a4b857e98b6a61dd185f962a7ca93fc0ee27a92c1ff062870c0da05f9b09f76c231ca7c6f732f6e72b1f690d701dbf5a7faa380c3c1d39be4be6c4155cc551d99a21263575d80cb842360409db28b65a2bd6b75b092a0ce77ab5e1891ba42696e37c0883f8c33e79e9a02d6cc8a3e7d6c7616302474a412d01b8d579e7265eaf27af2757628810cf6d8d41cec9f83fc20d9dda852623c17da805d0be1893b20ef8cbd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'haa33ff7734b9fb2a86e724a91552d89f58df10de62f30d990b7e91dbc79400dcf5ca53e2cc08b1191b2fabbe1772025872ea5f664da8942ddacdd444a5d636315f7618bd16575d49874085edc5c20bc6240053ba1e94a5b114eb6e5820df8708a410ca9d57593d328972ab850323423f84dff9683e67cdf61546397d1788f19805c29fef38537fd05303c43d87aca1255dae025cf6497e4b6e29ba67762135a288e02306378b264e5c6791c4f276348788681a1ee78823399b251c99fc4f376148eb1061fd4cc2e0385b13767bee19ed006d0de9caec391476d1efe2f9502734fe1530a6a39359f3e1fc297617036f21fecdba6b068a70e058ab2adc04bc36bc2ea21571ba0e8b0940c2880374c15a7b694e4dbb005f016db114e806e1df47e7ef2237fc7cd4fe29a3e100e0c99f05d933c8a6724be3cead4ae780355ad4c6e7de32db58a734ef02084f12f1936c08ec850d67a0bab94c846315962a5dc51e8b66154346dcc7c95d8f284176b896578de4be39de19e4b1f40809683411331f2b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'ha6e09136c6726941c17d49752c2d3b4e0254b01a289b1048781dd8904c93f880a20f103897975d007d80e65046466784f397e1c0fa1ea54d4b6f79e5dd741ad1c717b7240a85f3fe419ae42cb54f03e1c9d4045de76dd041c4165ecfd6f161d89915d11a667080a4689d68c07aaea9c8d425e76c215a7a81441bc856d677159d112cee663197c7e455a443ded55a96b084d26066288e7595b910ea1c54205094a4e1e6937e1eaeee1d0f463b7d0958478b6500bede9a75450c7d8aeff5a604a799a4c761c3607cd21b76a9e2de45ed183ecb3a3a54279bfe80b4138ff120ee16e5c5b61270d5be2444d801d57a4e510a9135dfea6d0c935d3f021a53d6788e2cd62a21187565459f7032e7739311e16f0157ba2da737879351da271664559200ca714fc5e07853af702bb4d53e503a37bce90d54d5ba6c4c2a55888a342a476441967054e13e3bc8bde816e99d8d7ca3fa43b0f7cfb9eef9e582df689be9728b6c6ce92a20d10161aa57f3b7f64692934c512331553a608898c5df8e41c430c3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hf07e86b5ec3a093d20c586409ec490fea804f29708367b6000ee9416e4a6cfd366cd7b536b800d46f8d5b4bc0662767f0b67a4792874e197df5c2a1fa595a69a4c88d66ca5efe5d4df5a2de83ece4452eed42fe933a5a05b50d61f5993a58a9da55f1adbe87fd690fb1a57951b1c0fc6f4d9ae747fdf741166a8ccc95811630e8241b00a3948e65f3e60f0ee867536f27f7a172676aca3a03512ca7ef287d082617778e4546dd8cddb17f0f06453e4a9aa0475cb62c06784d38a5248771f6cfc7d81ddd69da5b2cb58f130f18057b4a61e3a26a56283e6ec939923efb48a97416321ca6494e2ab49be1d9a27e7912d2aa1ef04d1f7dad7ce35f4c5d716afc091803ba34f34fe13f9ab6961d941f60f1eadb29ecba3e746b05a821834994b04b285b0b554d1b64389ad22486eb3a85580d0eeeebda9c2691277fcadb776188f6ab65d84b8b531f730c3a69b2e87810fb270616cde7c7add8f46dbe8226a50ea8834911bb8d92b6f5ffd388ee69febcf9ceed74feccc526a1288bc84ed832c89e5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h2e53bfed4a24f13ebff6615a012429bf0631bd94953eb7d606d0b6f5d460927aee19e4b73dc1c5c8668d68fddab65f4c10d24c033f97090a2a54245cf254170635d736b67b339189c993cdb3fde399e12946e8a60ced2df0aeca817e45f5a90bb15420c1564bc900703ba8b30e4693e80bb2b510cf6ca2db84ba6726ac97ef314c680e5905a10d78e0655355ac23bee32d5ff92dee77cc643db59540513c35dc0a589c19cc48aa905f0b86c27468ecaa08342b9457bc279a3389a470b33687eea5fcbb8e1514fbd325d93ce9a8d5d260268a4f31f0a25cb51a31bc5699c5c2b2da0e3d910dafb3e664080d9c36b4c80742161422c86580782689c0aec3fdedb8c48d2cabc14d3e1b0c80cb9d14c35d8da122b92398537190e839a08a4fb98acb9eccfc5ce926fd30bfccc47c8fcdd6c24fba93796134d72c653f0ab43873a2a43d7dc1460555af4c779a8c44dd41ec2f7e12c1719fd5b7befb9debbabd23c1f8e6f1cdc7d4670cadfe584e23fd65374c836634dd1ae82c513fcf30e5e0de2e59;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'he6d7c973fa4456ba86deb4d1f468d262bd4a144f4ab6d4e1f1dd855df3f1179e4eb0b8373ca44899c2c5524358e3109117a97b88b203bdf0f694c236bca45289068ff737253754161a7986b235f0fd03833f2873a39b31c724ffb2f5ab6eefac10ef53ba2900ab4ea19c3ea84c194455c81989131dfc49db7323cf0e4c04d0daeb8dd46cc376686c32667732cd4b02300a925b030fdb71345138248bb652b51172eda9653013577ae2bb230dc4440a37a5385fba7561055d8570a0d07e9ab957ea85728e81b478d86ca0948397e1e73507b95e6a9e519f1b98693cd9fa65852a3f5c88d5b21ff26c915c192a7feec66278d0bbf24fddc303073572e64f438729c1d45f21336ce7a93b53a1a41be50fdedab4e4cb53cbf70632b0672be0eef4dafeaf97cd19631401fa630642ddc878ca605275a862723dd1518fc2ffa313bf70faade36a74c40b6d6a51c8dd6a3825b8d63a36576c8b5c9ccd63b40934b35b717d1d893882d42759eecf9660d3021f994d2730e61ecd975a8de695879de4a48b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'haf00b517a87420befd444701976a5b2a980cebb48341c7ae15cccb85e41b48435f5aa61c8b65153ffaf131153789b0e00d8d3702a75c5c73c0c3f384fd88da42742d9f9a5279c8134aadfa4ffceb55c1c0d06be0253c3a55e371eeceb4fecf901fb8e62953c9fe10d3adb75c37b01c6c686e2fb84963fae968414790f3ed40326e143744987f35077949567a270d63a549b9bc20a004d63e86dfb5d2672f472cbe4d1a9bcfba2e17440a5d2aa1a8ac360216bfb5267a76f26fcf59feef7dd99d2d50bf62e8c3fd64d438d5ce037dcac94a51f40e0862a2c2ff2da2366b33d4ec818de71e55941d8abe72a42bb3681381de7909bac04d81c4def50157dbd26f566dba862540ae6c8644ee7ee82f2341fa2695d56f4ea077461b869854a1b3d529c90fd304615fe27942b54739f280e50d17e59f61902f14afc84c403c901eb88c8cee23bcb05ddba5245f726ab9bc6e0b23d93ad243474e471203322aaa902e05bbfdb096e27442a90c799c19f9111aa40df7b15046f332281cb7def215da7837;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h5adea7cc9f13d6dd72b5a6a7e08f23651b98a72bf9fe60158ec4e1064b02876052f8865eaf0e5b15c4d1b7e3733f45e1edc0298d1f3556d0edb35add380cfab0afe21e934d3bc7271e4c514fc2ddcfa0f856d8d92b7fb5cf9e10305c4bcfbcfb7fdc4a36fc943b9cb28a6a2aabb7f1d6e64c4888ffedc4c9f15daa1468169943d9d27a36cb6df1531a4a0f02fc2e9b4df9a9e0616c7d24b375b0f06ae6f76a1d9d0cdd398784e8a3e448fc3bf72a3a4e9513ae6a5f3353040cdbacb96bbaeb04839dc615efbccc8b261565fb9e9843c11cdeaeb7986c21612ad03307413367abf3c92e2ea56302d45dd2e8361cda3ea5f859a1fa417ce2beab942474c5feaad4c210039e4aab38c4ea685280305f13c11957622ae61836ae6d717132a400d5fe923a712e887f8d720b7d50dd432588449e5659722949f3b77135b857ad2efafeaeb0cb01cde02884c49fa2c85f3105347340640965b88364145e7e8adebb70ea7dc721306e49c551dc7bd580a241b5458a67126d8da1fcf60d058f043527b2cf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h36573598cdc327826a42bc5adc43e39d91948c9bd0b575e6cda2a332430ffa76d6d2648ca2488a2c0c874d83e85ed94757ff3f4135d58c956a6bdf90fcff511ff56861af138d1d1015889cd90a36dcd1a7201c00f2cc88c8e906ffcfacc41b41b5b439c30e1257eacc4bd29c8bb385f4d0035eaa4242a3a48c435684c3a84c2633fec8a04425f4d351bf61d4181060ebcc5234d49d58c61e570d401e02ebc0ecd163f8c1673c6f38636a97b7f4f63743e3b18b85d905942c306928e26164cea1e42959098e71e3601786e9b56d8b3fd99456a1117d2e946a78861da1b8c1269c03dce1cf168810e9429cec3038fb16daf1ea1eedbcee3ef852423b5087b8e199314313b79b504c74aec3c7a2e87d7dba02263cd982e34bcfbb262f2a7708192dbd708370492a30797fd6db70ac5f2b2f7d5608357cccb0098c1050c21050523f2e6c24f86c79efb66ff1480406f4825c05cc8bdd6ed9d2d238e835a15e10ebbb3dbfb23a2042ccba9320927b36dc328002563a2fed954af48839309f274ee975;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hd093599fc572b6d90471c54d65d259261c7edce53fc3e2b9fac7da9d110193acd524f5a3bce18a768d004241069429292b3c56fc8aee8c7e73342ced19315a1c5a7fce828f821e1b70b1720d603898825377ed152d63a95f07127cb7307eade8acb302e3c41aa4780dbb631f89f0a32387c39d36e8a705043f5d80e4e8c0297b56d83c96dc7e394d8275d3965a8842aeed86409c41f3ca0ebcae4339f873fa75be6b3c3fb4a3bcd401e4fd13366a2a210a30f27e8dc945aa704a740b2db844bde930ed19c2c99e997ce260dfc8b1d6808179d7c5246750a0bcec77435dade5af21d988454acb9ebf076e9a0460583cd9a3ef12f519412c2cb64d80aa9711acb8de2a9bcb4acd0d95864ab0e61b2d8ad6e2d0fdf3aaf2afce92ca0e2657cdc500eef9c79a1554fc7325ff462e0f5922efaab2ac09bc2a4a2b13d09d6dbd6a611b582ce8949d5b93e25596fca6389e1975fe6eeeb4b2fd151ea6de5919e089b8df3eb31a98c653db4b088b1740e217e31f9bf978409303cbad1ab8144ea69f8e77;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'he4137c6ce35fe741cfe8e2f95dd220806e0e990aeddd19ae00a77d0c7e34ae7b2785a880b1427abf096b3d21792507900dc7f3e94a9cee0d86e9144f36401ae73e61d142d906873ad11e81bc181483a5c30a9d037516b5c212deee81afeba800ec4cf14b09af4363c305a630af62514b20e7e61668993f05f95f49f2e8a8bb9f88bd467ac9d326dad9b3651fcc9b16b06e9690237119395b794771f5866f96a8935d699e87e845a553533dd64b22b6aa111087ea8b01377a6e20e7187cfd7d68c380beac03e2ca984febfff3cb970a841d88b0db78d5422400c3c4b3c93258c436f80a7e3d6f6fe2bf17eaec608a346b302353b9b459c0c0cd5fe0e834c35f2a20ccb5bd16db54d4b573207dbffb8cfec00d2e12c819c464cb666664218f79ac44940215d0abbde124c4edcd37fcd0652cb3a41c0a000beb8305091bb4d6a540e4663b283e4db534ac7ff07eb9017eb79c328f09ca057ee26793b55d93b4a6afec47a6f856470525ef788863a2ed17914a637688dcbc0266af13c76b3ca79e6a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hd3b858970d1bb32dd0937dcca385d23d8ce0a5609175a51cd27bb0850638e42b0b805e14288d28460ed83f352d1b78d29d9d44c0bb786c852826f8b58ea6db954b1884031528ec77b713bfb75f83aeaa310571215e479779883094f97c01bf629784d8e4d6393f4e92710ef9952e402049360df040a671d817576c002b53c10cbcd5caae16fa4887bd5b7bb6db587cd087abd014255cee21c8cb6d380aecfea81cdf587efbd1cbb8cd40dab85943412c3408dbb05ea2350936393b9573d92cbe70ab9e4743d9687ff8b3bd39019ec053e4344d6ae8451e4c06f4724fbdbc9534c02ba6023283335addf036411dfd37d780be7e5aa990f5ea9ffe7c14bdab5f9b40271ad5e71c803a23c5074d7ad8c18e44a3dec0b1e1ab1f57fa22d60c3c652dddf0f0783c9d8ee50841844eeab47c5c917eb816240d11691abf9126f28337c9dcebaa5555549c59c7535f52f98d2e55d6cabc35d9229942d2b86abbe0de3ea2fa764638e624081ffcc34cdda3ed8112c2799e1689376384107bebb9683a83d8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h18955bf6ea25955c306fba91bad0baa3ccdafd8bf5f8616d7d008b4b40257f22662f8699d6ef78fe245c99058c79c21bfa38a83f457192561267d54b75dc0398b5dcf8d407bf62ed6f804fdee6b32cf5daf4dd7709b0735f93082278b08263212ad14beed56e1e36e39f88057e6c9e37c846236eb6fbb860e3812bdc6fffee0f205038c569ac46cbc98d13fdbe547f7784d530f637db24ab44a2d833ed2409e6f716ad03c95a3b003955dc7cee4026df6a3542a5db7533ca78b959dfda04fda353d6184fee919f7ec1abec2fef92247c6d0add7d6d285a8d92aa6b8d0dfd0e143c3f6dc73f2493024d7fb17345307b151c8de2b4b7fde99f567e0bdcc93582907ef12b5b59037c70c9fcd3085784a9c42920ef88b5161065d80c434b21e0a339272eca9a448db01513536a192af2de567c08435f8ca68a45f86715336c8e31526c137cd48e73f626313e2f838eaf216f10d8e3f87eef66ca686a2f5bd3e0321ad591365b80e13b5960ff99cea563b4588bdf8e01a2fdaf42e7eeb3106429c776;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hc3df2efadda03cd890fa3c659fc7707747a8750ae0a09f4dd997348ef69895a487fbfb7ad3b0bfed1930461b4ee6b27750f769be72c37590dfb4fae8be1038540fed0f434b82598ef8bb7b7d4811f120c74a9bcc3a652b67d973ac8d95354ad8a035f622920beb7589836f58c45c8ad0becad655dbb11ed1beed4d0cc02488829b0d33a35da1086baff4954db2ab0197983ec742314724a0bc21a6f924d3dfbc92b1f9532e0e65c8d95906be06a143f28ef0572dcc0e594489a748b7928165d98a6bd99eee4b287f6d83826014067a10881dfa2e83bde330d4e5cae328e6745f35299f680aa96bfb00de23a5f94781b455de1b29a5c9431207eb4c2fe82787a6d67a7b37c1e5e2977a61b6937867838d6f6d2d75210041bed909235e665ed2ebdfaaf2da265c5d0ccfb6834f3bcdb69ae8379f4560ca634c407287f44db4c5334435db6cf399ea848b3c0fca227382f9f35740c888573f9e6a1cfd97213a03ea74783f00820a947aa3920a76149ba00990c9657b79b770c1a736d5f4da784cee;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h3d4c6820f62cac37462d4c8f5715031f6fa60206ee3d34ab320bed840df66abbd4d9c94aa56ba71c5f70e6c4bd0e3b038e0d9520c8299a60798c038e21bc0d8f4b1bde0b057737f9809ec81459b58e9e854d856033c0157bde16956a98edcfc669d515fb81877e323376aad0c47d49c41fd5b3341fb1196023ecb5d6a8d90cadd688ae847e81c7f241f37cbf4852cec20e48ecf3c1e5b20d7bdd3914fc95ce2a9efee3c1416af4bcd547ba47d736c3af39cebf4232cca08eeba003f912cdcad9ce477b52246d44a7129caa91f449b313298d3584e94c5dbaafce4f203333834e6a1193c7ba30671ff6f11833f59759fff819bd4253c64d2f4c8a8eb6253318c63154e4560a905da7253db5c164f6667d60efbdf9948e24990d4d146b80b5d6293a5759e7abb0b4a0f719f402a29807d6c3ee27cfd60b9dc4d2c3cfaa9195d9c1321ba7f573b7d775c1a7c933199cc1227f8e0d66b65f9fde1c39e895b25622fbd67f32525b41b2948677b5a7ba25786e1bfadf6d888a4cadb4f33315ab6beef6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hd80bd304946a1ee65fc1a91b3124e928baad8face2517077ca8cd65e3960305be3d675991cb6612b2edd3e7f684b581e03bf57cb77d7fa1edfedbfe656b8b732faa1fbf11c190dfb01ba54c7bd3b1440b637d4cba2bccd80d4999fdc5ce93cbcd2caaf6f38f110e6156627ce7d6e61f1c70af47dfee7630dde8be1feca2c98de980f0a3a77b5deb8f6107d9805ecb563384688432df1667b9bba44e540a5d268e9619a46736c7143c4a9ff6996b771f3f2bafdf829655726d2316d2b00ac47cd9969043d769da265cc25337842170d20882aa49370d8b3e00802f540b80f0274a2d9e0f40f2f29d74e228fe8db1b7bf37082fe356c4d15db57824cf4170ccb276fb6d81c98a843ef88e7469afdbea68ecf863485ccbb576e6d68206e04ee2329ff1a3d2f07be1c67bb58afba12ef1128ceaa1702a5dec04b118e2f59981f90c775174f0a4ae61b6f05a7fb09aed1c5dea87e09a56185fbc39613214b0e41c36bbf7f4643637834ac925e49c2eea03e36bc6575060e4576f1f483e4366201f0b2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h559fea244249462bf21ceb3d8a60f15224bd2ef28fcb26048ea8c2eb53578814f4c860d70683a468bcf5e7e42f4ebebe061e398f09e64d34d38e62658dce487a6e969e18a6fb5dfe8380e0744faea221d01d8bb20ccc28968041dc9c6d14a83381b780fb58d3f468f446d006ddf718b49f8ebce6adbfef9dd46e5ec2ae5ce646d52e806de80c73a4bb4b0f398997118b121b091effa3de43bf853f4851f735d5cf6c9d414213b0731fd4a5417b6e852fb0cce91fabfde1888a8a6b89404dbd02b170fc25e1b1753aa727b4d9d14f6cec19f10f03b127308fc5e9354423c0da7b7ddb1c64efdc0141ba47d0ca3178398abebf30d1f7a63b7f256e5ee5f0f3472416223cbb494f8144fdf8fbbabf08a8da02b65e5a477a4ab606f47cd23c73706d87f02ad8dd6c481cbbedf87c9d5c18b2a8a24ca74c2a3a70d9ebd103487f503f0bb0ef45e0c4b72a5c16ca8e0292b1819bb3f7a00760a73cc8d354455e9678a0c34ee63c377b55dd5552935f423f78a588489bbb4e5c39bcb75390b402223684;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h533f69040bf7fbb0fff72d377952ba810eae81366a7775f8c6d738ceeaa2f065d3ccef41046e9078fab44c965000b85d0e59560c7e395316ecfe73369981ac1d3f0a64c63cbe58a887094867d6d3263659b153ddc107130763efdef3d73ba0a8a5e103c4758ee3386896adda7e62c2d5385f80e70a4325b67d1070cbe5b838af5d154f8542efcc959736305a1221e75bac854585b17f8a6f8e3f4651d87e584ae5cef3f48e90bd052d184ced669157a76c19f9bc1bb65496e557ccb05d4089e9890e1c6ebbd44c232f8520f489fd9b09e0baab2cfc5458b9b036ffa03d2619c2355cd1e8721ed19c9a38840e452021c3c69e1dd151724129ea54ea8c0a43a2c99eabe850aa1c9e579f6f7e75bc5a44e4e1d30b8eb6630641f82566108a12311aa40160f24d2984a5e72d85bbf43a279dd9e48f3f2c61f1970e6dcaf2a686011485c1ee26b5e93c7ed3ec24c22874082923d203dc6e07538d85493c9fe03526790e1a758e3ad14804bb540e749256aa9c511fa01411dc6cd754ef28163a58eeeb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hc0eb9fa58219ef209dde259a7c557402767d95091203c349e6ddaec9b1c2451ec181487a8cc9e283a5c9ef6e9b117d684ecafac97c35655bf317be894c12fdc0e760b026660ced756219acfa1f0fd0f871a245a24cc60f91b4fc519b11c066ac56e47e630e08d5b9284be31a2ff1806fe767108fc45346b54415fe970d9fd10032cbb876f1dcf8b206d0f9f38b484159cad2d95974f41945e2eb2197d71027c4f6efe88e9353f57a8f6c6eed25eb1b9f40127aeb35d982b03120794951edeb8f845bb4f0b95a567061c9ca8181ea6e365c07729dddb6954aba3ce32b3d420e70fcff8131386a8c4f38ff8fe53f069996c7dc95b4d2b59db756f5fc501fdf45fd698ce3d6877b037858aae456993635ebd24542f0ceba45992aff693dff48234ac2b7c7b34103a484505b03a32cf7878b47177d0ba5ff54872a67ee7e3bbef276891242fac29ee1cf62c69ba7432d205d469363a4f69ef258520327561c12b3ab167962c81858fe05ad49afe322c325b8a71e8d0dd618bb1c002d68eebb1ae02c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h2a7e05f1175df0c5f700d7df4b71812ecb699400b22b621602414dac8bedf2f1e1de03d8aa2e9b600ebe3a10d9aac84381a69891fbae31d5dab7a483ed157c55f62830825ad0fce1de1b0f316cbd408a27be8f7c10acc49a4f1ba225a6360cee3bad4b7b835c236b19d60a562a17c7389a227dbd61faf999fba8be340ddfeafa1e882689afea502c2d87443767b0131547760360cbf967599e4f58dfb57479db0efea97ef36cfaaf1489d447f26a763ce486907fc6708c65129e73360c94ad316d6112fd9abbf43857157e84376da892c6b359320f0c4fa7bd7c2e4dc373ca0505d71060f1d12078c6e8c5420c61c77489b87efaedf9432f0745c7fa40e9a60f863cb0e43e3b19e700e793e9f77e10557a2d9f6ba7cf9bd8bed9a95271c7b8f91cb2069655a215ee7474b74d93e279a79ce34738b5ad74ab68329797c53bfdfa3caa57e4ded65a90888e2e53633266d9ac1951c475f9e4303dc3333671286bbe10f7a65645bf720d52369181f6a484219fc59b3bea46f63abbbfdb0b18a36098;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h9d5e752390148e8207adfd1dace5321bc9f0a2eeba25d75517ffce1e949f8f048dfbddcb4d6e35e9f34ddfc416c4a6dcf3f8f5fbb715183e5b623554e48d64f18e023f302f1303f69dcedf63c0855d5518f949e63581b2953495623e122c4a7e2ce5ae3c4b0a612857f1b1f910f34e101386aff4332f49020905db4e07d6b4218fba400a0809855ffa010a5d708ae058ede28c1403b7cd3cfbf76cd23b743300489e2b8f8acc5397b92ab789191daeb93b71286908eab412dc525bfe51d61ba6154cf8ad01eed1212db5a208df21b6cf05cf56e906a58101a2ce8234f26205b2aa2c9d7f186e07f17c8911fa7ad1f4245c2dbe4e902491e1f38e4108906c1908b4d3c7a7fe99e2c10069ad531d4d713aa1131a0cf5136f706be1512fa931860d32451ca4a8b857249e5303ddf715c29a537386f30505fb0d11fd4a1fd733f427c83ab9a4167504ab6baa038acc5882e19ade89260a5ca0f1f1f65ef5036211b1ee4e7d3f17c661f15e128c48389e9c0d76cf6f4b6b64a0c05336b78d56e78bc;
        #1
        $finish();
    end
endmodule
