module testbench();
    reg [12:0] src0;
    reg [12:0] src1;
    reg [12:0] src2;
    reg [12:0] src3;
    reg [12:0] src4;
    reg [12:0] src5;
    reg [12:0] src6;
    reg [12:0] src7;
    reg [12:0] src8;
    reg [12:0] src9;
    reg [12:0] src10;
    reg [12:0] src11;
    reg [12:0] src12;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [16:0] srcsum;
    wire [16:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6764c45cf875947cd442b7c4636b5e30622bf2d06b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h180f40942950dee6ebeb21e6e4627280f927a055f33;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dcb82def9fcc3c1889e786040303c138eac3e5ea03;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19b638f6366b41b3cc2d31f95eed2b03fbaad5ae13c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14b60f2592cab5e892eb1cb47ba7ad4c2e84c2b5583;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ce51794c2a7be99901358b09ff1b14cc0127b868f0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f830bb9515b00b6d4880a92ce003cf914bbcd3574b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h100cd26058e742b86c704675cd3af2f2531053d6376;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc45e69e89467d70db3b5a6b48f31d5429a903d5042;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc5ed622adb0d01877b16cc4dabd8a3e6f31eedd85;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fad6d2478624250991f1dd3f79e41aec30ddfd854e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ac5f07a0d8d74c8678cfb1ea21a0f28c5ace17540a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b6b5c45dbb514580002bea5f8261e41d30c2fd9f14;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h184172e03b608b23a6f154c7c4b01f43d3175bcd44a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4b7b88432678c7e78ea2c2a0eb37624b38700dcc3f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h27f85e7e268ef0b5e9e74c4726bcc93a0d9ec2b41c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha94cf5eed617784e7ade02fede914de1281c9a563f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4627bf82734afe8834935c043510961c48d9ddf84c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17a97786cd9fb15427a04073b17f48e8975eabb9505;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d11ac9956074ad58030ff54d42a4dcd22058737165;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17f1baad90ad79170d54840666433548224f8af64ec;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11f74ba0f5483f1e24bf45aeff864f986ee6d0af206;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h142cf15828d57879a64a10cb37b6f5e29add5fef78;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13b2511cb78818ee0c83cf92db47939a31c3bec5d14;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcb19eedb6bc8dc424715a06b0419f1664dc556ed2b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2a8c589bb753132bdcfb5c995247d1d2c86050ec7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b89ce4090f8c2120c8dc6befd21e798fa8f5532881;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18cd90bb4fb76763f07107307905d0d1cf771b29e1e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h100f7284d8d1fd0f728e667d48e2402d370b3ddd50f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h31126923eb4cd0c3c0149680c9e41bf69aabd3e580;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3e65f4374e1ce3350764b686df3680cf4ba6a48126;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd95f120febafd25e7c6692d4a7d9b85f856260872b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6a4a13b4e0d713e42ae92eb3ef3e62bb4e26197431;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he5e7c4aeb109a21a08886e609eb192151748c97573;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13938ca044fbe0a3a4cd70ffb99f9b33cb32fc29b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e5aaebedf24438662f8d1d8a450f6e11af2eca30b6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h69e9693d4cb0ddd701cafb9306c857672e4f8c5e1e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6434f6de832d3502f25223d259b618d8dc94532f67;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfe6c8e760260d65638d9b6619ab9665e4cd91c4d07;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cd10a9b9276540a3cff9b8748562a3243d39874c2e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aea4158a33551cbb008112d40df701472e9c7c9bc5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10e4e9809262a9a755ce4b78afa16f04db67e03552a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1348825cccc245dab054cd9a4d330bdfda1908543af;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6472bee7a8825e5782c2acba109ca08b8489816b1c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1005f911d61c72ca9124139dfb9b8b72282bdfac85;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hce43785c74c1f4f2c7f12ad291bb48083c594aff12;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10f08c2bf968a07f1cc70517ae16dfa7c5bcd2ea83;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1930694829a6b3b9988a5e5e4242b6ba2c35117118;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h192d4559bf576628e7221ea5713643ea00c5c73c278;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hce207e6cb5127a00d81706c8c28c4de0a1989a9809;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h156897cd9d29a72726fa66f02d930b2870bf7d1d901;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2851ae4c7eec34c67ff3ba221578f03d6a9465f2ae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1839ab8db8e6cd831485ac577a2e21e8a4e24f8c90f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1705a5ce91234df49f227d8cd18256eb04f64f98ddb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h615095be31dcc4a0e723ccf624f2d8c65ec686ff93;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11a2333d7ac3f8fe8d81f45323f2b08b1fda8b3b50;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1daa6367fa1ee042834e43c7cc81b3a86de6cf040b7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c1c8f2ba77a06bf0e70d21f588b9f04932d0fbc34f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11cc004baf85f344aa22de0e04fc0612f06149b8423;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1eecefc2d2242076ef45db3601a6c2bcfa466dc2da8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h125238d1b082e7906048e176f17f81d8fd3ac9e565e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h958925779eec43b291f9f4774600a6713b3d0e68a0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hac8b8416ae373508ced5140299aa733ab351c3f0e3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2828e037cda3bd7bea363cb181248790eb071cdfb3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14d089b5038622409c06f1432c5249f09e7ed95c43f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h249e6539f2294df578c72b5377270868b9587fd7a0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1635977bbc914458d6ae39a80b88b9ee76825907b9a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h53ea683352d799b5441010af5fd440ec2d262912eb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf5cc8703dd6bd2554295a5288663580a9f1c3e1386;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h84e5f9496cf4a920d071104b6119be567e82670c9e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2d6d60ce6a95ce57d21d612b65b2fa43ba76b001f0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ab4eed09e12c8c564a5877dd6e6bcf22a0cbcbaa5a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1536954d0560ac915211a6d3afdf36ba65d55dfc130;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1301dbd52f9999ef3f23a0f214ec7fc9213eeb895bf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h150b04e347c3ef61738c71f14da5f07ed97e48fca54;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12627bb088ebd220b9f2aee60871a5a60ff46045fa4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h87b472d41e3fac28f3d8f91ab19319a2e1d59792d9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbf289425b5de59d9b75f4a4702fd3582da4d25f75a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha1ef0085ea674baa2fe38abd27b4b13d9c5b2135d4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9342bd0653cc01ea29d7a0c881267b028beaf51186;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9242d225c537fb48a991acc95b64a90f2c254986c6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h62b8bdcb370ecf528e003a820bcc86b150ebe8bb6e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1283837e991e2f2b3c2f23c3024bed64ae49c21e308;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c1b3d542b33d4c3f02ef7debe6ca8b3391288b9114;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h389c01dcb2a1b2d41483a99c806ff1bf7605acae81;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17f8aeedb3e753f26f3c50c94ac4188749e9531fd4b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbefee6a1df26482570b69389c9b1426d520efe37d9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hac57f2c65c0b6b4083483dd15ac6aa56eb29535775;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h113f6f8dde76ff4dc3ab270ac9b49420403a07f77b8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7276bc63f9fee3e6cf171f110c2f53b9e2f726f352;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17d922d0279596842754d1a1285e093768c5f2c01d8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5cc61c2db3e9fa6529691d95b253162087b1ae6645;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2f7ae7c7892bc3df9667b68527e0a4a9a6e9e011fd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h24415dbaadf0cb078e39aa943e903e554de95915c6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc90b88f041e96826d63541e7da0b40bcd1aaf08146;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd14aeca74a683bc97b46611ffefd53834c9e295e7f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd280b8c86b53b3fe81b83ebffd002bc257d088dbde;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1018a3c569e7dfb58b61850aaec3bf8d5ea84640be4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d4c66039adba3742e6a3a2c14e016ba12ac6ced230;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cba70150f89c41e4ac27d6033c45ec36299b6d7e66;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h872dac97ee105b2b560ec2d27957400c66d38daef8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f32999dd16d5d9b97b55ca6c1c0e149e1709bcdd79;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1db891ec9cb02dffd29e8b08953e56b3791d94a8c92;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13c3118d811353e510ffacca35e0e7064746662efa6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h72d14c5d2551bebee88fb920b60c1acfd7f4ecb99c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ae8b96170b664d0fa9da7eebb2f11955881c5525c9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cdd940dda20f1d063d7fa519da23a508f391b37540;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h143ed660680e7959b29d6667388d8bcc3b3bd63c54d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1af1c28efcc3711f8630944162209170547fdd55c68;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1229dc3e98e9583f4acef81b4c68408ed14117b33e0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h114d961e15027eb90406d199cd38a1dca53b368e325;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13308f6efb3d7f77b4049cc055bc4abdbc8c52752c4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd9de219be817966768e476aed41c66faeaca69642b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf1032521aeebb5c20fc8c1489283c3b7491db797ba;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5cc2bc2544abadff573cf0756c362e801e49681dd9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bf0b7c559c4a439bf106d890b5d02b15722d25191b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1107224f78fa697d574294293eeae47d248af5f6b5e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf0557fe37ef9d4f440cfde7ee9221d497f82b43ac3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h29d98a560ccf592732238feedf0fcd47fb2dd0acc2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8553f689f2e0dc563fcc63487a4650e56274921682;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b736a6bdd0985acd67a60bf20373ddf21e3976ac55;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d7fbec6e8299a337af7d617eb76ad087da25c6f8f2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h147eacfe1680a8c6df31bac9e3b0759083a8c009256;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12f79c291a5a8603b0b72c3004216d18402c7d8168b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h153854a707e3049bec830ba699b2111008ffad4e6c5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h21e2a8dcc3de5c10d2da152cee71aa174f2e27c9a2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ca867022b31272ed70614a50b130f9a2a7bc60198;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc0980a815c4f3cc5c63cd4515f3a7ceed0752f8680;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cb5b9d3fdfae83c50b14f41c453e977237b495b44a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8197434aaa85996f037aabc765badefe98b0191214;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1555a89bf6873a6279c587e59ec0d3605b58bf3116a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbab563d496bc8d70842d736de552a08872faa80079;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11ed3624fb5248de3a920cb61567fde93555363263b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fab9291356b4b3b8f3c6bc5162902c94c88f5af986;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9313bb4d3528ec0bcba28a5a7be0b7971192c5b081;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3346a162036955f083aeae42164aeecaa6810d4f33;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h163bbd638fb4e28ebdc5417c25a388fd0168026041a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16f1b5c3263c13d584499578fdc217a236a184a23f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dbde68df325fc58f15510ae3d0532a44c8adb589d6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h157cc4346c12260a346bec24b2c1896e72afdb3a24c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1988aac325cbd9c3f31c7284f187161f32fd9fece15;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17fb48e76e6eeb4bd36ce791c9fb2a9f7907d4f718;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc5911441d12bc73825d8478d4ebdba4106d432e8a6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h965dfbd1dec9164a674680db000974123056b04275;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbec7cb5f24568aee61c30053edfe6f05a6310048a5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c3d0c4a8da21e86e21d1037df181ae28940c3a76ab;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hed965d1a8e1182f66182cb24162f65d67e68cf276e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1517f7636fd28d6a42fcffee9901a6ede8134c54c9d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4afdcfba7f294855845272407952a23d8b4ce81923;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d36b476bd9d725e0e2605a7848eee63f92761939e5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e2e6334024f178f99eebc5dec26ad5a6206d902efd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13f8b9b42a444c1997ab8f9b3ecc19a12eef0983b5c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6de1e6352bc4636fa09ba040bc3e8a73e212f31a7e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1673c4f6b743f0d8bc9d4e1017278eba74281d204dd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h20b5a6048fe8ee6b85927bb5254cf424f41196bdd8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12788f816e35726b47f8c68e9435c21a5604bdbe68a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb31fdb38d9c146027247de95b71f956a25b8e30bfa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bca96a2a7555c3da57ed77af059b2add6aee87da1a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h27f9b22e750521ca53af04bd3e75e78590d523074a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf6850f304cede42c82e3135064441feb5f66802e7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h462197b103ab48041d3b80689561f9a00da50aa560;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ce4a7a3972c071d828e3838caa6a10032bc4d0fc7a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heef0aa50f39ff9ad5d20d004cda183b0518a643f8b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c59baa73e91350557e9dc81b93357dd0214bb1782;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8b917f57f4a5dbcb50ac54385ad382fbdbc0a7f9bc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14b552e3112d57ac8496fce43eceebaa9d7c8fa2268;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18fb098e43cc21b5c65880ff039126ad0081b659bba;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb7ecb7035de6f9ee87620415c0491c6f8a87a5de09;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e36cc2a2355dc58f939c3addaf672409ec08601621;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h269ac7fc8ad50022d6debaffb36ba453b392e80865;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1083ea4539adcb013d1694d10b7ea45f7c116c262cd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1da7e424e7a3426ce1fb4df92ba0aaa7917eb045ca8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4799a3a83df3d36d59502f51f6e07febaccde3417e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h64bb0b5eeb6b5d6831988cc5096879708f00cba7bf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h170ae5c0207e140230376cb89b6f14e7ba20121e212;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd56b31ced45531c6a4539a725c159871ecb9915e56;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16aae00f64766497ce830afba84744166dc25882087;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e9eecf86b61562835a4a899660901ed82f8a9567da;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d6fc7fbdeb7a040c0475afbe05e577cab5f4176bfe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h502c746cf3caa6392b4ad0c1fb70adac4a71d487f8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h44eb41dfd2ccbb7cee623df7617d71419f6ecd33bf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h790dab84938673fa7f11e2dd433700652906a99cca;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3a2eb1c68cc1fac51a9829e1d09701b7b06166ace8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17a4ec2f13e2c582109629aa6303dea58f932c9f5be;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b5c07f6b761b517d7c1115bd702f70f1a0f2e55b44;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4b83405f77ca4b4e8bf54bb967917f9240c85ecd75;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14d3f19cc42cb2a375429d0584e3ccfd20ad83a7494;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b97c832d473253df8e9a462fd6ccc5c97916f81775;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h111986e5e0e7cee550638f358ad21d899c8b0252bc1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19ea00890d7a2ea60aa01bf8d2fde4d61e53f6383fa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cf601febba2b7a0f2b1bf4ad89f2c3bf8ba344a3d1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd92279686bb11cff11413bf9f302a19b009c8a2feb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h107c8181b6073ebc40de940d97d4c09668f33ef5fc7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2726e27522180d3a0fb40aadc0e6aae9f03f1e448d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h48c1cb79b95b94da03877a99105b149a90668ef7c6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h336fe95b6c38db83f8ecd8fbe14bf4a91e88e2a7e4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1285c21a6bced92dd5ee376e1a41ef3bcdc3ce0c024;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aab6d550a6eb5fe57c036d6d2c68e64ae5db4d2738;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7c62fe2a458c807d9fbc2de4681251990aea76cda6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h726267ec19a044bf5eaf8f24cd515dbcd00237ac57;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1808890354cd8fec9dd8ef4cf2740602c2acfb91146;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb2dec69bcc76717a1d58e5f593c57ea39789a186d6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h324701076b2669b8034cb82318c06503c1e2e5239;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16b87768bac33de405e80b51a16b1a8b801eba36377;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1df37c05a5c68a2bcbaeb69ff34f42b4f02a78beed1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf43403017cefea8fc1bde0028a513a9709dc4dac66;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h180aa5b0c613c5fde7a8e41716fea76661ec24d148b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haa103a45ca827103ab81c60fe5e3c03d7b9bb6f87f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10a415ad69dc896c241b4c6c428065e1bc6d0b38a0f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15cbcc85991c79b113adf9628a02e62fe9a26547407;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13a0dd21d735ce6709e626bbbe37f7efd4bde7a986d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13c92d861590e4b9122aca0a29dd5d6021759bce60b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h107a5e61c2642dff3ec6cdaaf37631a090fedea3eee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e65c92c193c828e7ace27835d1d3d1e8e0e488f1b9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha12c06a397e75c53c24c585e9aa2d3e86c2eb72bef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fdc2bb3fcb25388cd16cf3a67d79c5c80c51db1018;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hda251b02991b8e48ab339ccf746411d5c0b1ead5de;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9bb037bae63c6222713898d72a703faacbb7fb4892;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b4a3651477daa3869defb786ec9e5b3e147be68f71;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h123663d3ac8a556d8580dddadc617f281556ddb6e85;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a36a3f7f602ad5c42789af396d1c8cb0f9f4a0797;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18001709cc6e173b8062d9a2c1df9e2648b88f64983;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h245e3928523bb3d24e4c9b1a3aa4c4e281344862d5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fcba94229b1cf6940e2237a2181abab1cc758f0f29;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8093062860f18907c9ac65109add6b48cfd7c9fe1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1268a8b59d49574c55b245584bdbf58ca5a5a953721;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4d21b8747e283b56429685066ef93c54840b372dac;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdddd336d05b9c024e3fc8ce3869d91c5530b654529;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1529527afe59bcc61c5353e90c1aaa2ca26cecab678;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c38a252b9e25fd4df6b02e5227a16ed2c58b1ef5f3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h328caca78c37d792132ad04e22ac8484865fa80f5d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19d9244f84f3f9f1caa37b0219bcc1f5467ffa53cf8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1611af5fd995cb340860d9ec5003975bcf9c555634c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a4598e66186105ad427b96bc675b6ec1dc6b53f0d6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6bd7673953d945f44c439aec3bc9d358500ff9607b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6e40753d22a6e06caa3491edfa26f2ac9ab83ccd4b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5100c7afa373b8f4f11d6c23f6f0ee056303353c36;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc5eb417fff26786d305d5c43f99b8ba0d89e169cda;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9c157a2e7426b3ec8054e9d49db630823770d9fd8d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12bcc30a80c39904913e6787f50f078c33b5bffda45;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f543bb6929e1e4e73652215a6ff21c7993af6e2873;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6e72418d7c3c0cfe395dd23c6e65daa4838093cbbd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16ccdfe5bbaab63b75df7a1d47dc96f3c387d2aaeb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1302a7d1d04d657cad36a4a654570c05bdfd67ed36b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h632a471debacedebed22f75c40256f6dfbad87dc9c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha07ad7f4577d3024907d9c9604ca79bd07034ae230;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e520c3490aa9e140c60bd5ee98e1ebd9331f9a1c8a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h100e2883f06f27a8e1ba10fc531d67dcde0ca63b73;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hde37a5f6ba638a00f9c9ebfd9de49fa893ba010fcf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16123f2eb28fdac74488c4df6ba5492f41ac02de301;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h106755a0d932ed6e797f8808988f0734a5cbad02aee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4129a055cf1a93c4010371ff57e08146849db95e4b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h729c69bb84b5d5746033be7d8c671e955209a76038;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a496a9faeda6ec00cc67e52c3225e668d59a3332ae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10d15ec605e63caecc87c787ff05cfc92d3a9cb7822;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he427fdf3c3ed87c747d79a0fc1fbc79dd84f903825;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h82410065522b02f1d89bef649c0f66ce2231a4f337;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb2f16446627f0860ddc73ceb2fc7e1825734212324;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h965bf98dad2baa3d5a4fe5ba6b1738f4190ee7a387;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hede3e0d504935622d9f4c57399020cb143bb82629;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a80799af1a10fef57c9ab0a9cd2f120af13796a542;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hde7e9a3d0bbeaaa63afff21698e5ab2c5ec49f31f3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hac8ba126ba790f57afc05ab351152bde2482e0615;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15a737d35bf43ec9e92a4b051ac51357e0da9dfa49b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h135bcd4a9299cf1a2b17cb3a19d5741e6f3c254e7a8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h751c58d2fb54bc83d3eff90c6d90d1115c41f2dc86;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h111a2922e8695dd3bcde4a295255ca023e2200b17d8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1983d593b3c56be2afd73908dc7db07766ce617ca07;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a50f900e67fc29e0e7d24a3e0a0cf2a6ef6de106e0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8d5cc756a4723d8d2a73a0c71b84d6db2f7960fce6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15d9c11d46f7fdc735be02a31a26626fb1c2216d79;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5b0897fd18489194780e280fbf202305611722ca77;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha90fd9bf39b519d77cee589740eba75d3065de512f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5b9aba6231a26534e1465dfb5d7fc24f06e410b511;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5f323e62d6b7a26abd4c3f5bd3e8ab9573a506ecc7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7609ba236baa362e79be0d000ebbdb71c2866ece33;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11dc61add70acc9ee043f3c04b2cf9bc8b8ac1faeeb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdf064877d3545ebd291559c983f62fd14e0f21458c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he1484e257bdeebf0bfea4d9133a75714f7fd44210c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16eee724aff1f7f0a074d0bd3da60b8c3ff28bdb6bf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18e6210e957499489eb2daa5ee3d11fc0bb8fbf311c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c2ae2cdd324bcfdf1f88bbc1d1c0d1d97720d0edec;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h95abde34e07ca1a209bc1ef2107ecf39dc7d60af7c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6fe93d7ec62e7dcea953c021cb4ffc44383732e302;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h181619d366b17a3bf245b7f0422ed17819d88908939;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6f9c6a296e88d6be692d281636e61676e8320c308d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5c3f1a1a217d86ea66c31bb77f161951cf55751f15;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b4201df49a797904e70274921fc9450034fca128be;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a9de88cd60a2eb235fa08f8645f9e762f3a016485f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbc7a6cd9390cdfdd6a2004614b63e849afabbbfad7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1222a292913bf66cf880662291d795653dc60d14f1b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6688ded8c3db2a92483844fabce52361c8e0c83fd8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8531c1da02b49a572cd6ce33157adca36788d53554;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hff842ebf69660fc62cd1d0473c98183fd77bc1b213;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11cd5b998e6a43a2e9b382c21049d90874b98b97097;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h250b8be6e0e1273af62541f3bc7d5fadaf069d972d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5abf4312ac69ca2488151416bcbb58227e48cb590;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7b5f68b2fd6c34f38fd48fafd9f25b383840c38b98;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19628da283379225dc21bc4142360f0de296b328a0a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h106771081539d78088e104cabf8b8f1b9eda26d9635;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15834947f8ec4b8791b848c8fa661ef5633f0c5aa6e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d03649ae05c72261e1ca2e66d7f5c8f1aff6a4b830;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f2785cd148f7579400cf636f103a58402c15a0d22e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14847ad416ef55908921952d0f5013cb1df2a000dda;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17233e34b2261145d3245dbc25993b2a6f77b481395;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h360b8a843f6a551620fd7fbfb17efb4e0457232f61;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf2dd6446c97ab8c9df1d4c68bf325893400559fa47;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1de1b2e939ea342cfdd7aada4b5ebfe470a89782a89;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1af3221b5c23263361237e8809f36b419fb5dab16f1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8a5f432ddc4dea7be4bad56b6baa19726ed3b9c84e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd5facbc576762af3acf7fde39b3050be423768a1c1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13381994f727642ca019ab6bd9bc66ba397f595026a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h195c70c6cfb7a1deddf378430ce4246dfb6f3f745ff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc97ac38fccc5c83ea24c966a3acf0c9a793f39094e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2191c51fdff36ab990c64e81b278bad2762184133;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14338629d0ff59e582afcf7fe581d4d8cacfb156b0c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1edcb18a9b51b1d76530e3f8dc39e68bba2131778e4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5930d3f42e548fb2fac8b73707c9ac5cd84a9bbb45;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h41ab67502e507b0a24a52c5b9edf24745398b8e30;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h586016f2c5a24ffcc3a7df1379496f88e8cf0ae42a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8845ec6b18d404d0ab50096ba50050599f540365db;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heb106397faa4ac871ef6d83c9eafef6a35b42a909a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17bde719596d7a0a9519397207ef92294ed529bc55e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc0bf50a4b68b2ad0272635fc6ae80a5b5e654329a0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5ed251d7b8695c12b0fa929a61b890b31646281083;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h30e70b6692507547e7b3d69942959e2b73915936d2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb4bcd6dd35586727753c223e09ed668dad2d0261c3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hedff7145975a57de3dd0ca5a4a7c95909098845e67;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h553574cb216323955ae78ce015a6b22bbf4b81dd58;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h199a044c459f938ee166cd4921ea37aa8ccba584c05;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e4fb6115979405debcbc8e46dfb2166b46824d094d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h158da30572751bfbf466f32721f5ebe9d19253728d3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f5e28bbc73ae3e71176c928cbdfced65494f617caa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e6b079d21bb7f89e0bda18855af2d5c13dadc972d9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4349a240432def53e8ac0c26657e9f4ad3a5bf8f45;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19bf0e2cc2821ac83ba0d544baa9cc9de9ee2d38a22;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h52f3adf029108b66abba85c46b46407e6970563a28;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8e1607b9dd60abdc132958fcb940f123c75b7a8abf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haafeec7fa9516ea4a1d0b8e8bc0fcdc98e6adf2f04;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e13f8a79eaa487639dcfe255cec7b522de6e43e194;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf37a364c81d7e042bc7df5b8bb2b3df0339818f595;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1577eb47dccf222feca3f89aa82b8b422c59b33d672;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1683deb07b056fabc4e43eecb6396924675dabdcab3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc1af6d34fe999011931ea771492ea6da771dfb98dd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11bd8757a44edd83678b64bee3582d541d3037f20ee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd7afca1e1251c41f5fa0695af46d89012a1416450f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f5f509800f12731cbe5fe476354da8b05d51e15a8e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h205579ab12a3c8c50b9dd902b062e9f39ad2477bf6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb5aa178036b92a616d15f07de1b641465c1397c31c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15e7a71c6d179c27edb7e4b8e0c0b0ac9a76c0731a9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cf37e528a1fecbed4d1b3bd74c1af468d3b674b3b2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc76dabc9ffcf78a0c6c9304dc3af465391139f0af1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d3a2be9d9710d28d949c90e522a27b8c6a84381529;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h90f500da979af21387150b7267ce1b5a1d588956fb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1de2593b4e1fc88f10fad62b74d4f0bc9cbe1b9f96e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ee1c92d27c81d4b51c88f2eb6f4b400e28749aeb3d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1139f0b6630470ac0a6183fcf573f47a124bfec126f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h113ab74938f97a4b91a2c2a5356cd669a199b934d4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b65ad41154abebc98c4908afc60400f370f8bf2572;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6f8ff26e07f910b375eba6523434e74ed82be21804;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5bd3c91d0b5a4cabfafd38e131bda924e0386133b7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he9799c017473cef5bbf08414853e6975257fdc4ed;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1278aa5b0d38706386a27159444f1b3d770c860b06f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a1596bd28389c8e4313bbdb6fad472d48a2110873d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h24da87de9236b89f1ad68ae196c4d8bf5b60ca5e8a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e8318533bc311dc316f0d7094a53867090a82fe7f6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c793d53796a1f0d35083c4e669b95a621e82980a1f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfe5d7aaa1190a367255b8581960babca1b9741272b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a17c6364f9e6f79c720f3f0f7b48826b3140e9d8e8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf6d66c196e2d40180083d1cb2dd51d0a7994696579;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h26dd1d5286f4925ea2e8f8e71ccd80786872884473;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bed8f6598cde905e9825ab139b4eb01fefe2142287;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heda69c61c421ce625932866bb2719cc4fa519d6b3d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d0579f2e9e634a57ba959ebf393db2cdc2c1f6e4d3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d7a32c10a5a6ea8a66e6404c74b7f07af14499c36d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5e4343790a930ba683fcb8a5d25b3905a61b758952;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc4dd50a1bbcde5de9947eae9b8106c623b2f592366;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14cb6de512fa4c0b0bddc012b96c97879bb4253ed5e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hca4474612add2243f27151770ea21e5867aebf0c56;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3e0bdbe639ccaa4f0050614b946dfb033e3d76ad9c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5408ecf32834d7adcebee3793e28788c3f921af5f3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1585f7757642a35445701cb8c14ace6fa647b822e7f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2f30bd9adadd825b7d614118aed1bfe3116f469da2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1142ff837e6df038b0c4cad68bc9545282469f29331;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h188ecffdbde80ae060ca0d6b10ac92808ca546ca5a3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h917bf9d8a5b6db00c5adc7da490558e98a07b31736;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha21a5deb1d65ff48b051d1272caf0e9b1ce1f5e982;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7e5679036fd29b85fb349bc62968224d50cf5a8f64;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10e18a0e4cd96ace35b08d7afe8fa7e1dd100484cce;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he2d22414f742f497e2b23a31098a43f558a76a8ee1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1eff5ab044a09dabffb434448f594a4ceb0840337b4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14e0d1a81126f35d47be67f9a57c1e63b87796918b4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he87bbf2e3529d30202217f77af505e526e32cc7a73;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13d45754b14274644612b1186b3199f3fd72dc2e76f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc561024cd8415e4d7c237a32bd3c6dae257301975f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11dc453c85247830f883f69da405f548bb4092901c2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h76b1c435e26cb01660700ca4c8de3a682a3d78b6bd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8aa7048113f08a0e84916bd5b1fb388ec43efd6646;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7d7a5d1c1425e087e70dcf67156d5e745234a061e5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he9a9a2034ed21f5dfb4843db40356788cbe81c6655;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hed92cd941ca6741daac68560b19455f3cd696b0bdd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2feb24618e02a0a64d2f611435b1cbea825b66e3d6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14d13bf5d1f76bb6fa6de157887ace5a9c958c6c37e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19b75459e94e59e212375b4106a5704d6bc2b1d1909;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1555f77ca536324f8b940764b33e75ccf74f43cf097;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e1b29aaa1e0c5cf53b7bba0cdc73fe4f5221a637bf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bc2e64349a56ee99257e39938d7d1bf55f212ccc81;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he0249b8ce55a18fcf8b399d701a4366df20534ad33;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h198797dfd2616aef7aabe917500ad3e8f9d6ad05741;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha2cada7abe20fd0429da4ed7407a62212796c2d77d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ba16270982cd70f8da4879bee6fc0ec20b3cbdb8f9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17f21fbc9fcf5cf31de62aaae6ebfe8b3f095da4bb0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdb06147d7fa721ee8bef848d627e271e806c314f9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdadf0172db4444fac8e264be6fb3deab758f6a616;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d9fcc19d2fdd1bab7e949cb8183120b6462bfd13e8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'habe4cf532778969e54cbbf05e4933e337b9ec12ab7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he0df06ba03a1c7b7c0e54c8b9408036b3e4f89f0bf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h127c547261de0ccf9b0e4b2c316efa1a449cf728689;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15541564ed495ed3be4ba6b170b2426d14ebc4d9837;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b4c6e6b448ee7d04bdd2b8d435e2934a07f6946fb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h182cd811749cea7d06821d7fb38897932ab6234ab0c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h380b3c838ea957e99560294b8d5d338f81bbcc75ca;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10f14407e74d680c79285a61f1d6ddac621c9ac12b2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha932baeff71c9f4c6ae70180897a87d7a4aaec341c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cdd0b19d3669d5df3947add1353f403f0332049a6b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9c9accebd9b372360edae0c98267d4fae4ff9d50f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h31f2bd2573b6fe2d1a1c733de71c65c2cc61ae1178;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1018ff210160187fdfe1d9c2a96107e7f9816e651fc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16c18658d75e7ebb25be3bc7b115c5a44575961d704;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he113e6a168699f0c82abc056316a6a6de06d3f2bf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13e631ce73657028cce69d4b0f091f121c7b6c8ed82;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h379e08ce1121864a845977ad7560221b3db942d8fa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h24414ed3bb01f484533143e3b6d16804f4f341b703;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a7b0c48312eca3d143440260f377fbc86e6b1f7880;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb0634cbca1eb80a89a3e602314f9be6be2ed6f4686;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a6153755f6a93d5a57458c7e74fd09250b5f142ec2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h469db1669cec679e9be9e6a90efc7873d48dc59b1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16d95dcdcc33f51287e7c695ccf573fe632c78fb6e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e65c7be02fe5de204cd15f34953f08a9b05492e19d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcbe3dab6f9e4257e1bf42a3378a157d12d7af73bee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1636c70b177540e735bfac0a5d649796554c0f45f64;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14ed14fe7e58e2043d138cd4f35a8583158c208b08d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf6c4c4b1d66b8bbe6568ce8dc1934c7f04c17bb723;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12aeeb40f54e89acfb9aa762ec469a012177bb1b183;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd149107414c1a317a089814c6f5aff77e492a72ac2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h406ea2a24b1e2ffda20452001837b9bc31cb61e89f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha7517dd708fd01cf848d05ff5cab1b59e00b28fe3c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c1ce9885ed670179b8ffd0a6ea86f50df77ec6c518;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha34c3ecac5d7d7659c5a190e3b1f44b49742960bb2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2c0166f3051f90b01cb3c63710be0f1ceadd477438;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hab13409d2b05cbb8e67c0a3e858aa536fcb5c2784;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h63a60eb7b2a78d28ac0e0b66b89b2274b1b6eb63da;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1efcc5962e320bcaf01bec43085af9bc1bd3ddd5d44;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h146b6cc82fa95d7d20d3e411d2705b5f8dc49c986cc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e4b4f9943213930224a906d4be5f83bba00925bae0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h53ac52e8d552bacff995c4d3e664848b320291e5b3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h98c91f03cfccd728663b159f49d54f6439d26d3817;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he0f600af21dd68c1d9ebbff6d406880ad7023ccaa5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16b6589504476efa60a64727bf9fd69a9686cd74963;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5d516f05a35adfb61ee1d1aefc45217b3ce899cadf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h128314a0f78246a12c9281ba515d239f794f52f69f9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a26c3792d82ca159740bb857c7f2a22deb2add9899;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h73531a92759afa4057718a19845554c4df32d1b7bb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9483a96ffd62852ea54ffeb04bd8eeeac89f0cc9c1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c5dfed4d26ef978297755fdd1b1694bc27137584fa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb71f1cd32ea93c6e27e3bab64da566cdc23a6fd9f1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c5db4c60b23c1f037a27185769631e0ed19fa5e2bc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h47cde9e92d2f1a7b1bfd4a0b5fccf5a7b5fd3fe4b9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9ce0b58b52368b6ac7a972a99587dd46ed0378a6dc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16ba5ada033a1c1459989b2f3702e47c0b4d9e47b4c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf1bb1d5d96efa7998f55daa1aa60c98469b21a5cc7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf4cbffb43baafd332cdd5d0028de25ade9730b8e3d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha8e6270bf6792d28950768c6da20aa854c06ab169a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he27ae22e9260ee24c27084344a9977362224e4c7b4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h132635fd7fe7abcd46fdee06b86dc920497d4724473;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f4d0d2d0068dfd4fcc4620fb202e7e50243be13b78;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h31a949d600994df82cacece05500ec44a0d2b2309b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14a487ee5f126732698c5ad5bfd6694635034a74395;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h122a393c90e12960560fca3b961122d4f252bba43d8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11ba34919ff1876c50752fb9fffedb5588e7c3f9a56;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c2de9fad02d401c6d48eebbb7fedc868b832447be7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11136b1700b99e3d204fe36a0db0b4b92956a6ba5f2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17b05026bbd3c98456c0eda09308e173786ed505454;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h106ca7073dffe60d8916d2a63ad1d30c5c6162a74aa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1204581c266a7cc7c298ada4ff974264b8008c6d771;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb86d55409ec68f5d596cec615a4cc923fb9e511013;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dece501f90423956e62e42bf7961933907f6bb78fd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbfe64c5e550fdf600485887fb9e493a956bb4f46ca;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a06c6f0e1e47c272d94393374824a2925eb551a501;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf037f5ca6683c39c8998ace7a3e3e5026fea67a247;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aeed6293155b454cad5be100f90def2351493fa2a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8b6d084355e9860ba4e49b663c084727a35eb68bda;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5bad1579777bac60064c0c4ad1bd86ef3a528debb2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf488a46af4c96e2347d75b99513e02881e83c5f528;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf7e4d16756dd9e38014a8d6b52e0b142386b5e4ea5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h164fe7658376a258f63bc133bc0b5dd50f016b24602;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h22759f47d8a03fa0991e7d1c4a30873079ae0c15b0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h126dc1d600e5e6574a8d0971a89df847b9382dde409;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19653fc8f7cbae2fe7ec98d2bca9d2edb1a2b27b451;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f12584b63886973e759602dbf0d1e76b66fce5c7b3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d9cf7e8680ed1f76cdb563241dc0e4610657eb939b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15b403434aa62486d13108819ccab0667c6f97985e3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2e5fb2ea4c7bea917bbae2419e597c9411bf85caa7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12539f2dcf5bd644e9bfe885baa3d82c46189176f68;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aa0edb484d14e9bd9e38231bb4586b3b4dde30c1bb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14ef74cd24f0f20b509c31d434888fec3f059942b61;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18b69dc1faecc6538583dcde1e52bf70d757d8c2c32;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9ea3e56c4f2d13e8718e1473031be0d15d8926b6cf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ac19d799993f548ff3376754661647c8cb5cd2b999;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hafe8d7029247b406d2415dc5d58fb11bc909ef7bcf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19b74fb75394e4870181f875638aec356b1c7403114;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10dd901d25fd3024c6b8c49d3114f0be17dde437473;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8a9abad19f7770211df4a59a04c0e60fdd4f2afb7b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h119ffa33ba0ffa68d4d3f57259679a3e8aeb3ec0c4f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4c12a4281d518f5c804de53a3070b310c81df49793;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f6f12a40d0573f62fdc41d95b18b7945844e6f0abf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h199df43945537151bdc1216c97c32aee8dab7df197f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2144f19a78fb71a20060a0d06303732891bfb880bd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14d57f95f56ac0cc52fbf2721af43f4791399319e0e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h167aee944cf8b15392a01870c4e5d98851a90efd4f2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hac44c4cbf28624f3a3b228bdeddd9f3e48611dfd7f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9821aebff4c0474958872ae509fb5b3d18d76fd18e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha13d23b757735f149e425f51e1e0721b316e15417e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h23fea2895424855310e180fffa618dde5f8f401a8e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13f7cd71c326c7d4394857122865743f3b26a213954;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1abffb4aa2670121ff50285317b23ed04f46e640e74;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha1a286bd8b2cc75477362cb249fba9c84a44cefbf8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19f4961259a1686ebfbaf28d04ae874956b116e037b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13a462082461919ff38a935e07cebd918418b43cd56;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h195579354fd470b5e0d4b82d0d2255ba4016dc288d2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6b95daee11ab56c44e7401df273d6d6480e3cd23db;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4c6c6b6382c334fb9de40861c78301a15be07cd296;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1be7636360a0ddb76d1e928dc237e0f329dd14a02f2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h171444478d7666cd2878ee198c7d2a6da4bd43f6512;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb7b90811dde6355e2ea413d00aa0fe6606d3aaddcf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1158a195e853deac94bdfdf7821f67ba83fb49d2376;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbf36f4a553431adaf93efd662cde7a294c5c44b3fa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf00d451652dc1085da038f4f5998e836e13922b35c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha7609da45084dab0dcaa29c0389cb255b9a2ff725;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha945c94316eb588d0916850b61852edea739b81808;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h40d6d8ea5b38c590d9b79f7586d216d6f2d0bdb597;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf92986018b947557ddebaeb6ac6f11188da1340a66;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha1826013aa81e304566a7790d46b9d85ff78e40b9c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16292f8f96298adaad83bab2e57b74b7e0e8481ff1a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb1033034ae192d4a2276e8f8fbbe16fb45cab73a79;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18ad75f1484efe64aba01bd6fd115b0d33bd451bef4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13fa821115ce4150c90d1f60664ffdabadde017f2a6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5ee646dca672a1fdffd24bc8c9374eb8543fccab63;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h864c402314a75019676cb5b7147e44f83a85115640;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15e604cb8ef73c7014b8f8901616ca072ff48724062;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15727040b8b7dfa2ea10c087dcd1d81ebf017b260b5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h75e60a16155b9818c5c0131c62d2e7763fb5fb0865;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13e46238820bb820866ca6b1ede045bf6a2663e7ef9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h183b6aa78f1f7b87fc4d9990692e8c1373ee505c8a5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e150a07009f5a11dcb2cc1ccf73d3554075362179c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha4ac3880b8eed14b3684b67600f677f555e96bfb69;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hda998f5bd203ff7b75639ff198aefeb71066a81b43;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h746f8c324d96406cc1d7956cdd85f7bee9867acdc9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9e60c9f928cf6fd4a8c25c4d54ec39c33674b13834;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b995c467cb883ebf4c241d6ca1c817c841fe50e641;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h476acad068d892ea98d9a83c0f08a6505c84f5dbed;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1564fed26b1348f74faac8dad7792344be4d7f34eef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7aa908b2a09a610c3dd171045a68f268e69b44f453;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he433d508aed215065d2b12b2657a674cb22c2f7d76;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3256c055e4f3daa6274ea7ea535a9adb2dccffdc6f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h136521d2a7bc390d4a57e27122d7c4e861afbb05dad;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb451689768bed33e5b95e4c6687a60311039cfd7b8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2818a069af857a8fd76c20248243a2324763c8130;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19d3f39f5842ccbdc2e34618c9fea1ca182d2037839;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12982bbfd491f5436b1b537d25295c67ecd02eabd6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h167c76e3f16eb6218d2bf4b08ff1b12d168329eea95;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf505b02171894783cbc709239ddddb2ade45ce2327;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h45c03dbd6abe5e7dee327b1d31b0d3536bf9d78e6b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfa6707af8e4fd4dd7303b3fa3e0a8439da8c0551b0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h187c41020f22c5387ae3cab7010215c1e22e077bff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3799665b3943f0cdef3e79beaf53d6667ec8faecf7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ef9559913fe1f47feec80fb8562ef94020b56a7954;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14f492a673586a60f0ff2b3f2bae23b1f7e46cb6e42;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1083422ce25ea6078ba3af5ef8411efc908daf938db;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8c805bb1ddc81415f1dafe9e75dd1cf47a89b839c9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hffe35155a51a5d5d56e94fae9481709d8c3bdb5ba8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d92c7d20803f48e85da182162b55b09127f3c0e1dc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h883ff2de5ba9758e0941d4ad7a4421e353e0a9c1a2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17ab28b77648136610c64bfbceb3a9c8f622a0c801b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc9147efc0660fefa8df8ad3daa0a871c0cfe3272a8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9d9f7f3915e0925157fb19968f37cd25bfc3e7d695;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb1aa11811654d781ee411617a273ce89d75147d5af;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fe4d650fe5388e3f2fcf359f21bd423d4c8ac843d8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd32e70b37930c189665788b85bc6beaaba522c03d0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cca6655d6fcbf94389e74919b4a9665869351c948f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2b613aa68198be59fe926467fe2725ba1839caf3d0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h105c91393b072232bbee62b1485495f8b4f1e0702a8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ed8cbfd9e15becdff74ef2ffa05b195703d3ed1355;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16eee74227c4513d8e1e0a85d474865cd0bc3e93521;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heec4f25c9c8980eb0ab51e1c0f2cf522f240cecfdf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h774f88de57b210f0a171d5b49b61138b65750ce22a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3a8ab949bb7c64fd7f6bd413bcbcb4ba84bd61b4b6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9e149aa1b06b87aacbcfb98d3556eb0e13abb9e9ac;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1eaae97d74d783f743a993be13791f6d3161d7d92ef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf81e4a516da1f0cd050992c882c56507c6fdd8ac32;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h100cebde314870ee8bef1878185827a42fba0a922ba;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h183b09bd5f45d598bd27218d48ca829b62f46ebf31;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c45e8218f91db8f300b7f2eb32cc42fa40d3a6ae11;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h467011d1234398be80bb84af752d1f0cc698b03041;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1acec2e6a4834ff817cd255a842c33ebe572372da6f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd15ef7583f131c6b38c4053b844f911e62577fa0ed;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1142baed2d5b6ec28c29c452f1175514e8f2927ed33;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fbd81cd72e9ecd6dab5c8d76b9319e411ddab32fa8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19f28acd5e7c076f6691a339d550efa73c8040aa3e2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h154c9bf612a3a7830102dd2319b992711abf5e99b6e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he8ad192678bc354795edb72ae61ce51d7d8580e56b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9ded266374ecd8d3d39d1de4f46298979a0717fc5c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcc36b3fe6b8e03b058a411d92f18e8fdfcb11c4d19;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha8d30ca6c554108faad6ff6189891750f2a2368cf3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcf795eb36e9d907ef925e41a271408368246f78084;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf8136033987114b19a3605d2c7a61a6b01bd546ffb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfdc10c3b77dc01d1b52f625e649f510c9c6d83a956;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5a423c7cedddd335e38b1e2c6c4ae784512a6aa647;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7eb8c9c4f421473f4d29d20074839b2a389a78c378;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9f87154d042ed5b72389b459c1557a5ef05c81d853;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d275b0254bfc7756c91e36edb2cf986fba2da21310;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdb427ef0838dac5f86f19f24b8c657f8a22aeb781c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5d4f9830e01715a07e973b68ca451d6f111c1d795a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10213651b50c880b8c3ff23a7fa0ca4e4d001676ae9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8af89f90a14777338360ad0d9b60e9d6babbede498;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d5f63b54980597ab330035fb439dbcbf3a5b488581;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha935ecd49bcad20392619f2b8a4dd9f69ab16d0cab;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h25b3b279fbaa1f5b033a893cb15a2607358b656365;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1334d95b67f992afa6e8194fbcb5c8f7b704e8d86d2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19d5fd8959375e4b07ea9023b576d970b7c8197b0bc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h187549071e6a278e9ed63d818abbde32255e4193455;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h261441fece985bcbf171fe326a9f9c96efb6d607e6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17da8fa9b4b7709450bd45b2763a990349805f5cd28;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hca87cbcdf32b2fbb8005f7f1b705b905df273276a1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2fff6ecbab04234e915def710d67a9d100159938e1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c7ba43512b2e24ebdc7638ffa0f5d69f877234f69a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h774f17d648bd5907a7c000607f31fcddd3f92b836c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h108c67a2791bfd6cea720c95b36064a6b722e2bfe21;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd8d0b9ec08536c604e193fe78c146edebea2f43c56;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fbae243da4a95f1614921b548d051a37c3f913fec5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6911eb6818b446066ad0adcae29682a348f4494340;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3f5dee5636086f34be26cbbb075683690be5d42209;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12ba522ddbb3c9f3e1eaa328944da0daf1a88302e64;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14c6c71852647eab7afb4c20a1002b6d47b3ba54902;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6993e36ec4f7f33b33af40bda7511b694f907a3508;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h184f23118eaf36acf0efe49d104be17bbdd1637804;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hae0ac22b41c0f1dd51a1be3963d3d9b95e4c9abdb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19845d495585f139dbf0841f569e50a940aa5910799;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h87333f0aa550aed075f99e4e00386d4e2a79c7f9c0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2d4a0d42a91bbdaaffb45acd515cc9ca5b9ec9dd0f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9662772c88fa74d71b83ccaee425e7c6fe0eee5723;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1034bad73d9170cade6acbdcfda0a1671d6ba5ed218;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h926400e39e8b518dba23d69dc98a3492271fd01df5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c41939c06e5a6a81b7cc0a9620e1223f78fc94a720;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h720f41b005a7580fad088d242e8f022f4ca1bcb205;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c2daa177d017c5ea2207e953abaa9abe46b4585c39;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16857156cc3be041ba12bd034ca7cb068ad597d4469;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b991a0633f0acb4c27c1b2c1ff96f476dcf390445;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hae7b8939ddf2e1b4474c6e219e18fd5f04573e9b55;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h113b806c89cb9644f1d0df6440cc9e421286aefefe4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb2f845f1b681f65d8b1c1f3f968017abb1e2a6ba55;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b263b0410b81a228ff4861b7b852a5a0f2ab865978;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h476340fc21eb657369d1631f2fb4f4db403c840d1d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdfd6eb88670e6a1b1647bf7ec2769e2125455aa195;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc99072a0fc3c9b1a656931ab6846f402588140567d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1963b89ab416b194bb2b8caef10dd807a3e713d1ef1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d99216f69bb3307d19ed0a275bf51ba66aa9d41ff5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h126b713d4de33bbf00f31195a7988a18103b1bc9a98;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12c77c6f46c74d5c42fd041cc31b94f840665280183;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h50c4586ae80573fb3b93c741412cf6a97b0be75e87;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e1da406553a082c73a81d87d43f863a4144bd8da8b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1271c878b79e5f384f99756129f518310a102d8caaf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1856479c59a3a35277188a86d1068f9910e458e3bf1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17e9859c5afb71bf0f0a33c38d94dc09a07427275f0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16a60b2e88b24e1bfe4682c3a05bfaac4c045688a7d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h705a805df16c4a29c47d4c1eab1b633a5a63e9835d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc7f6822888e8077c16cc34551f1e07d7e140238fef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd579beedccc0a21ee04ea9d669e9a4dfc5fb9a0b2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cd7a226ab8b43beeeb839324f861eed55b37940929;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h97ae378eb66ee177b12e53b29f4488353581a37278;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6721539019549589a6177bae645fa8849fb834a175;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h168e4190f058fceaca3de0e4e71a120ebbb55ee6264;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h165ca40473980cd737b87cb28c805c0853a54093c78;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15820e23ac3960a684d776c38a24efb3904d8170038;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6fa9190ab8c7257ec69a05684f164fc7107e130b5d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h186c9b05f834c4079745144a94e0e51472bdaf65701;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1236099d94935c12c734d90d292cb6f56554a2ce45e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13df4e4b6aadd75618545279fdae05484119650dfcd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d2412eab1caf0999dc6b42f789e5f9e72a62cb08c9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c9f14363a7da3e34aa958b8d23a0a7744fe14fc183;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd5e28b5569a91f5eddb6ba43bc4575289c78fe4bcb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h152d9f2cc453c2a58a774c5f6c624bf19ccabbf6684;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h193dcbd5f73931bd9aa8870fee4eccb44fab7f211a0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18a4923dcfd899f6b9c9ff47f7e9f80e87361589ab2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13afeabb6c4ca812c92d8ba54a488782e96af016570;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1efbc43ce336feb2f82d1c827e1e6817a03e6ad5bbf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9de54a18b787793d7b7fe784c3435b5cb663697d2a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h153b564939f88b7ab6474285250f500f33003006530;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3d7afba88b10ca8d82c3781ec4d280d2a08b983e8c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h119b649849f6465d718606671a033f33c1fe7ef2a69;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h85dcc7aef931b5c783d9a95bb390e870e5025a8d8d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h130aee4f966619c84b762194224a8eeaa7776e48296;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c49706a264bb19b15c20e5197513bf2b4914bae97f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd865c7e19783a6133e89d0db199085f81017f1e4b6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f73feb14981fb3b65040a8facb50c3c8e002946cf5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18c5223a6cc58c71b4c679aed64cbe83ea3f2ebc41d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc38a943f4f5657a9781a7ac64eb51b2fa09ad1ce3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h130822e3aee88d31c2ca9ded1fd5b700c32d9877928;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19777866edcaaf6589123b18fcfb9eeb0087c15e79;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c36332d3774ccd003ddc81b2b94455fd5e6bdfa729;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h132a5d0b00bd2084146b29478cf78057bb087dfa81a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18da2850e54706e6f7b399e75222af0551ea2d1e8d6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d3869b920f9f56591231705dff60e083c1166db47f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h117b830749b66b74ff287c6059f67b9ec3d8377e64b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdd1eaf3fa487ceb033290e0cced22eb2e0924dfee7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h134ae6e57f6c6733a28e2d1a2847c5e246e3b5ec858;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f68ce4569c6d19a832aab80765a0ba38fc8cd91081;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b017846754bac9057f2f317212bb99a9397925fde9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b641a6013341939a14f1e4cc976cc9f3d8c2472d33;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h800b685220f26095f905236a15006e46c117b3325e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4a85cf02ffe9f5cdc876e17933bc0d7ae53f9f1a52;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1625bcdeb5b260e1d4e5fb19aeb14c3904f22918d5a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14894bbc402bb4e2a9fb6912bceb28e894afcff59ec;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h953e0c57de1e0ced2456df55c1a62962e33bbef32d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aa2a271e04b65a82120d42e1a1d3c73090eaa8451d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9b38b913e5555a405d09f5a2b6d682324817ba45c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h50a6a1f5ec6aa5aa7aaac86b10af010ed0127dd83a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h39341cd384b0d542aadf88d99f701bec241a21f743;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1118553517cab9949bb0037dca47cda2069b7f4da90;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h87316f4aedc215705d3db6f62dc3e9b52904502030;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e3571fb5dc15e1276b06ebc0307afb362c5d1f06f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f003c9a5d54560a6027cafce7f7a480815945b7f55;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1619d5a66a6820432eccbf823cb3ec2f22269d906e4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b2dd90c9c8ee77f4065c19375f904b64ebeb399146;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16be6d7bb0ebbd6f19d6cf349f28efd68cc04b8fe78;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h116c62958047a00a9774c62cf96b486e2eb21f823e3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc8495ee188aede2e4faade7686487f5afa39c7115e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h22c45176eaef90fb60b678a609d43846b34e254fbe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h85d0e6489907db26ca494b907d253fd0856284c107;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h83d7100d2b10f16b95e7cebde6dca370f4926f9401;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e166646dc424ea7a2db86a4e9c9fd98c588c8f5328;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14e2d062701c3d7c3af091edd6ceb5624d5371cbb4f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbfa5468cb29aeeaa67eab4c65cb95554e402ffedcf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfdf7ced9193054e096ef490f1fcedd65f9f217477d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fa914dff8c83431f23156e79e2df7d7bdf39cdce2b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he79dd13d073bc3a1452aba16b92c43d6ab4f6cfb0f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcceacdd40b41ed4131723a42c891a4e5e3e0a607e3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h199197dcf166dbd1d79ae8f3842c6001d5f0fd0b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd4d4cc624417924aca3c67495acb2316b33edf1246;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h73003c0770fd77b071a17672d21ad7e3ce2a012b1a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb224720a1a9a985d7ba464ed1c3ff7e941aff4518d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha94d1b1071c6daf61bf239a27abd64bb64d7239c93;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb75f900ecf177eb41e75508b7a6058712929b63e37;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf00d5fb76a4b9f2428c907aba17036b43a52e9f4ed;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h115a3e7def18110fc9d2343f9d2a2d49e154d9daa23;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e1ce042ad4622ae2733f7ed54d2b1a20b41f1becef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16ce5e61c1399efe9900a0e82bd4ca5e39d9d31c74f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h155177c741f15cbb8a69e87fa589b414ca3f12833f6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf62daf282f0ae97f548e4e167498cdf7077ac11b6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h856cde6ce43b9b9bf5613a8d64d7fc82149049d1aa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h60ca1e5eba0a954edae9649452637afc0a28c919f4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12132883d9ca82523568b81091d0d1b38fa8a61088f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf566c390fd59775d73cba8b04f22ba2982184c3a00;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h898c8f61d7ae2131a8eb0db5a5e8a36ebfa129b76a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1eebf443fd254242989df9e3116c112266da66ff598;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h117d52b5704e16078f28974fed67c9226934cf8307c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfe07645c3066db77e9f7f5217414174122f9d0398;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12c2d2095734ea409539fa0f480bd7fbc3ac4d3845a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h178f78072c21c2a95279d57751f1df22923d223e7c7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc4fc9c9f6eb8f01d02c63407ddde7aa55d529ee85d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dd7339ed42a7c13836ae4d86179f7795cbb06c3fa7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2b7dc2a8fa8525beebdafa4bdab3e5e6b9ee583bb3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1656d1e42b562d20c298b958e966191f6c0ed6cee0e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc8e5f13473924dd2afa607f4043a06c67d9a30cc5f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1994d60700eb6421ce44d9981e83ce0652356db01a1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9b286724cf49acbde9d68bb731f5f1e73b57ab47f9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12b89db4e45d17606ce678abe68be1ec884fec5a15a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d871b64f60f4c06295633f441c82cd1dfda06d064;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfefe09921b0f24125f18081c4c6ddccd96ff624d74;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h751554227556b46c4305eb04ec384a61166bf9173;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h190eadb9013bbb00706187c38f4a2119b9e1ebc3023;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h119e4fe9f19c0639612f49e72896ea92e52f1221f26;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12cbd2cb5a9d4f42dd5cce29c4d6286b373414ce4bc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b103d64a79b5661de4285db97e8de01f9003ad213b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ddbad58e25f23fa03c6c2d8fe38fc6c79642409418;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h132c86b62f2540d676f9ba464421fc2b1fdca66b679;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c77fe4246f9a8d43dfdfd3183bf3993f38ed4ce40c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15d103c499c7c7c8f45a65d1d9d548cf0185f66889e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4142ad8c43288dc39f6e93a2a2115b5613b480a534;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h178f23c813f1b5b14a6087afb5776cf0438c8aaf7c3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h107eedbfb12c0c879914586c39efd4ca0cbf6d329a2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6603a8e37c8694b13153affb78a634b7bc8263230f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3f869fc9a57922123bc4dea695621940a30860e6bd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h177ac1b5a72e8b8bde9301c6da1bb29ee1b47ef2ba;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdd25c4779b2ed50d1a8234bf8d1f48311bc0536888;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hca90cd50a6d802907fbcf021c4bcbeeb6f68377000;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfc86389b2f1b121f3308bd8ac9b27fbf5bd9da3a4f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h92a42d46ebe2a0a2058f7e82300e07366ff556d1c3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3b6a3cd0cb214307f80118a5499bf9cac961f06df0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9f2d024d5a7062980ce4d35195f7ea03442b8def5d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h887e457702c1af60b5e4f290ef40f816a89baf31d8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16aef323519be1aebb43719764f5a4e20bff822ab35;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6eeda728eb950ca0da6d6ee3b58c1dd8ca148f3234;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11b8fd30426c53e72c3930561d2e143eef96331195b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h111d0ee7ad8d6c70127ba1abbceb338cfda7b894c2b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcd8d0ebea6c49d33e74a1eea80d12767f9b361ec31;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e6b6251b7ccbe6ef0248326d76f1486ef4c90146bd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12be87b07884d30149c1efd6ecf5b0fed9f81e6ef8e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he7b3877afd053efee5ccdc56f56d965c59c7cffed;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h693e882af4529b0a416c7a7ca3c7241fcf95b8263c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h91457d07713ca19b4a646565980b730c96f09d1365;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h94603a58f650810a6561b5f2d5b3e1fbeaa39c47b8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h95b874a5ca67b82448b487db079f8a6260481a79cd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd7be7719fba8635c212cf7ef07a7b9531ad0e4a767;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haf2ba0c6ea534373b2fcc6ec3062a7b021be93977e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13455bd3ea26487cf0418a1df7e7b0e556744c5d323;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19ffda220f86e91fd77c2ebfb704eb8692442f5d30b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11ff617670dcff59a7c9e5c20411ef9ea41ace93fec;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dafec3fc22631efc8cee2e2a82e15b6cb629f6fd0a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a5b7395010e0d988042ac168bb92e57fc93047c570;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8e39d9961dc9644ecae8ea013c60ecd4445a18a965;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hac1eea2b41d44f110ffc3696b0e350f38c2c310458;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h81fe867a2f755b43fa3449136772a58dd96185f01f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7a7d206638519b35eaae808d6ee269babf1c99a595;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbc0e90b5a5b5a9bbda920df7fcde074f1c4bea00d7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd3448140294a775c6c5b88647f7dc4623a7910ddd6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b143e8c3403917981d02e21307eb886d8eb38ae60;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc7d8e41d1d40f7b15e0ea4e113c0dc423dda20f8c2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h47c15b268b8a7f57132634ec9908ca22fcf49352bd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he346815d10ee3c136f2f83242d2b76f0d1ff316828;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc56d42405905b962b1e1764d02093c817d08ee2d18;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a674311936c92fbd959f54702c7e4d5502615a36c9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hab373ab8486f7e2b1285bf2f850f03ef8e6c0463eb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h74bfc8b15ab7f9df8e07963a44ae9ea7bd683e6ed;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb7ca9c1ef63ab12c17e3bf8782d486fcfd8248c9df;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f960e0c7b6c4c6706ec0f7f107855d301a31892405;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2edde1237667ec73059fdc2c35dba7053e3db4a9bd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fa0ae0cb135f0de04930a64a169556e4a4a4dfe5ee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h162de2cdd511c61d68245ca64d472a0626fb08ae37b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fa56baa28af82ee8f91f16e6b8635b02fdd7121ec6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5f884b95d79d6af9781d7f58b4cdb73205bf55ca8f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h22c26b55e8b90ecbeac55179599428f808847f14c2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17207304c47eae81874492b5fd14ea8aac5cf032e0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10165ea05c3adbabca7c0e69c7093bad4c0fc00c2cf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e866bfbfade3f88ac50e2dd57f81ef9e3f8d264b22;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4d6d0611eaa3dc682934a2131e4ddde3273066d34f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h150d8c8b3b19c5a14b0c0d4ed872ef8177c752080cc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16eba809dabe5f3c0e46b63e465d30b0cb130c7a056;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1392a736986b1f4b8563a38531fbb9420f183640e36;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cc117a0a1d4170dc479a98d619445c5346ed6e4142;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h66d88af6c791b45a2e59e8051a81390cd5bd9d6d2c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13a3f0f150254984101b64cd55c8e3e9c5d1518b99f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc5efcb128dbe0fb28e35dfcb2408d1257f1b89a77;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bc5fb3ab5cac3f1933825da64fb73f104edba63831;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16841ba857c465bcb25526eaa7aef0c13578101f115;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1decd42a6672dd669aea11f027ddfe4c65c07987096;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1004f487b7c2051b4998313a4366a1b9fd9492ce4d1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1eede08c027910c53a2828738e87aa0f14b2874dd16;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc1ff973cd56f4468147adb1e3b9570e207585d14e2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8ab4509457c30987beaa4729715b19478447e461c0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11d9dcd1a8aff5053fe1a45a6cf4f768024ef0e410;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b26651d231b8c5fef21ee20faa8bb2f6b6d64daadf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bb445590524ef53a3fd57e94c29f95468f3b085739;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b29ba573121dd2521312ca0f4e7e94eab3179ed19a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15a02ef36edf383c5d9b94682568a6a355d1cde8773;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h191d25df779174d3ccc73138f7627b8b1f7458ca94f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fe84ce6b437118dd1c30eef601769050df35871f95;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1db09a73b408f626ee30f25c0b25654c68e98cd199b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hea783e93e9a9f5c8f2f2ff0dfbf2502bd00f0e3598;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aef9abc2c19115244ac91ef65d14f655bf18d56120;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha20994bc83860e2bda3b498632d1e0aa8c4b93731f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15438d16bc6646379a83d787c4ba5e5bb8030bfdeb7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1568dbc79454d52ef1fe52e0a374e51bfe92e25ec1d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h51feab1fb793ad5607ccfcd3726b97bf2114ad78b8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ffeaf8aee70664c9c6fdd34d61e2fba9f6761c2b64;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fb98ae981ace5de5e6dca95b72c4fe654bece560de;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h73ad310335dd15b81a26329502c770ad8d6003314a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hec0050c3d42901af4360bdc50401c844b2c9dd3c3d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2a1477dc10e48027b47751cc507878f8189b6a966e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8fad9b5a4b0dd40a1c8e59de80634b9bbaa83533d7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h98d4bfdee7d06d3f10ee52f50910723ec04b6bbd87;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha21f52b32df1d0f444ca7e520def78c9155612f20c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1244cd9c4087f96352dfa88bd4e34624d640aabe42f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fef52180eeb0eb71ea010ea53faf7892700a8637fe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8d353a93f5b1076c57ebd0001a5e495bdcdc1ac123;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1626f55147895f0fc10bec5ae8835c36865482ca62f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fab27ff6a259aed7c8c809706eab7aff9dbde9f40;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13b4f937dc563e540998ab0894a9da0d4f328e81152;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h156cbd81c0967ec023c72266c8f7d2a7f654ee5442e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1967a294392ede33f20db733934f6ada24b7ec0e718;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6a88d7656541d033f1930698d3e0559a5a46d68264;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1281d5193155895a56b4620302173d49d7b11394b1c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heeed697a89b4b1d5bc016e522950fcbbc1fc746db9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h152011c2a325ba7a59ddb1db4f008fb6578bcb38955;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h135b7788124d91108f9e44580b5b2c6df6d5116f298;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h133f88dc2c9bfb51aaa4c15934a908bae156520d216;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h103ce187c4179471731882cbe84aa4b91903f502060;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd0d187f58b3c58d41266080ef1f100ce89af8df094;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1769c730e267d373d581c5a89014ceedd2641a50c0e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d42919a4cafc9e1a416504a797b7ba596e29c041c5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h222dff0811730b8c70c3f4917200657dc775f8607a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h166addbfc180658cedabcf03de7d3f9de7b31f910aa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb205b7ba22337a23b1495eba4d665d5cb1640d7afa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1da89d15e87672bf451129e4963fed78667ad1308e2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdbec61f87e20872267a9ad19c04e3394060b95f718;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c81a7ecf451341d11004d7db7fb33ce128b19055f6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcd2fecd92b3ce223b3e53b5beaf61370527b6373ad;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16dcc7cc119adb7b62acaf21874ddfc5992411e2483;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d54cd03aac03f435a9743792b33402af7294b9d7c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d409c9fd3926ea2a34413399908a00a07c656be575;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdd6a6f2f2c3a1aff0c104e2da387c42e906e88faef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11d95ebed6276bd5f010cf43dc71567d561797d113e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hefb466ab4dd7fbaf5ae375290d9ed167a1fe5fd8a9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14c6d58849dceae4b950d2fce686049ea90aeee94a1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14d761482fb107bb61cd1c1ab022edff99095113a4e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1512d632939203445603abfd288dc0bab3504ee6d34;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hde0b237de1d76ff8f39a8e143f3815a0eb2068435;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf914323c7aa1404e2fff085c4672234a164f4513a9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b774addf97a13466d0737abafc61a3835a06d68dc9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b669e9520c7988d61df207288b4b2585262ac2d903;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4659b41c87978215c0bdb4a17b619d63e54a5d016f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18ad5f451710f20679e617aed004d77091e62a95a3d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16a7680de90eea4703aada69faa5b4cfa772fd570e4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17161494679df7a7d59174c618769f2a86cd937be32;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f8e7ce0dafa9d563b9b7681a9722b07b4e28159ab6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8c0d828a711f04e8d793f490f667eae9515752db45;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h705180fb75c9383de5092938a9564b2f33aba27149;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8ca3b4a2a108f8639852b47302051db4ca77257f0f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h119b80ce5895f6cb9e431f4524cbe74526f86687b82;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5620eb62e4ed19404f1149487ee252ddbc14881696;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h116cf5404e6d1878d7d19bf16f3f46b50a1a789f9d8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f2d5ef066163b59a265094273c0b2ea8102c4307f8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h57cbf8716b4e86a94272f7fac44a64b05006c1168;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d82d8805f4e085220e6f5553e76c99b40bd6583a33;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h630c0b6d9d8ba81dc2687228e46d601145be1f9de6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18b8c8c756df48ce3113a637903ef7222aa974f1ce;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h133eabf4a8ba7b1f0bf395931946aa26f0c30e5e975;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdf021ae964096bc0ea1068ac8e2ed31a3ab7e47a1a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13f9420e3c94f01be3fb9216f3cff66677758e9cc36;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h664610ab64bb95bd21ad776c7cd9cd5749705d9b9b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1647a7cee1b460f6dcc8b667475f38c3a1045864ef2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h933aa4e643a4cc8ebd1e8239ec194686d3fa9971f3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1074047e2a1f4676b9f7a168a8a23335c5ec1507108;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h603349055dfd68b9badb4bcb1b1951be82ff417ff5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h23b1a79c7cc4134c5ec7aff8626f98d7f1d8d1fcfb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11d39cd9d7c2db7f031b6c8fdd41379ddf32afb2df0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15083fb005910bedcdf1392bfe4b649f99c687119b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he5b8320839a9cee9b3b33e9cb80b2ffadaca63a194;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1288d7b939a343e6b44b7c04d5dc1a75a4c035469df;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13be6638d9fe41de9d71ed24b7a74b50d7317078890;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf0baca5e904ac396ba7b934903b3c77316691383a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1902e067ad29586892b2156a4da849d9fa89409b90;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h137f0f49c369ec5e894f6026b4b759f514784be10e3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h134484efa136c9871457150363b7dcba429f401919c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c8a66e833a2f7590b2f51d995cd8b4cb0b4c1b7e59;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdbfc6a232349f2e8470bf0f85c9b5a2a516f86687;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5da47d5d1519980864dd814c3628c4c6eacde3c87a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19667dafdb6e020be6a7c378d6d5b8443c84740ab7d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2f0d957a1162635baffc9f302238e2f3218b789c0a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9139af54a9236323c68eb70c4e1a447127566d0cdc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h43332c3dd523381e49686432e3103613a1f1256329;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9301dc19f846c07058915775a347a4ff076b43be66;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15e09efdaa880f109a28ef29524cc6cf62ea6efb587;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6217a3ffa1d3d164fdd5b304ae1df2c49186190834;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb4371cfef5159f61925377c3d7f5fd11a3710fd299;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9507e0ff843241c3d79c7ef72bc9b27433a3d9e2fe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5a8fa7f88974ad394a525d1dcc3f37ee5b3651f120;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12dc33834d67feabd78e053185382668c5d50392e50;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d45858ff5789e96d2c2c83de1ce33a908781a8ff0e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6c52a454a63c2736c677d3408e172503ed7d4ecd1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c8c2da2207ead47f1cf26460d7719347fda35ba7c5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'had713cf4df771d92b06e0656712f2b76344ccd8860;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16d853530a4dae4d3688d33b48495c67f9cfe6f90fe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h69e1bb03f7740e1b96262e3bbc83a4f000f7f913b4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcddfd3f347d1dbbd952698ec14c264333f8dc4a165;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1241a6f00c9d8524d2eba690894a09fdb4ef009a661;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1510375d87e6c3e7acb85cc415c01e0ac033edfe25b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e2b31d6a5998717be7068bde3f83fc381a8257e78b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb09bf6b1c7badf9103ade30d47c2597e9650423454;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19daac121c0c64495caccc84c07f77b0b180157ab4d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb036c440cb791ded0883a0f8c2fee11c1ad01407bc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6bb79dfa63de21f460559e74207ff224ec4c0369d6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12364af5be7e890c23fcf93fd389d70eb015ade765e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19be63aee8acf0067112c0bf7aed581cd8cbb3acbbf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a17a6234887cace41278177ed4b81d28221a79d7f1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9e6383c2d67081ec1e889f56507c711685db6ead96;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h163e106500e162983a15c4100c050a41c4c3fcf371;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d4c0c3d34ce172adfe06cf060172b4eebeedc6fbf9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1499772e1dcff34a887f688f16b846c746e0558f9f9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b5735373a7e10beb66dd37c289ec9c9af9d1f1410e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2e1d7ca9f97cd9fb7210ffecea1a9a715b4f394e55;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h174a36da49dea3db58a6d939dc2be297d427d4716f4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfcc1dfe13641de8b2b98117913c64d3b9213ddd647;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h961d59ba7afdb1ffbe827d83af9ddd802508bdcba2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1995067f76fe2ac14c6fd5b783fe0101df730ba4c1e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h196a6ffd5caa5fa34e64cdd3bbeb28f1f68215ebbfd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h869a358b1f005719e8993ba183b5240d89938464e3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc57a417c9c19dbb1e5f88be9b7c61d298fd2abe792;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h223fadb2e8e08de5c5b18e49a64fd733b4abd7a1e3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2d2abef9a288daa1af2edd2d3c9fbc56d6b4940962;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5100df67d2d6d5ed739fe271c738ce23ae982814dc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c258b0d1243bf240367c28de605d2cbf0472689980;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10e6e2a8380f5b1038a6c690e5eabd8a7ee45a2b62a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19e6172547e6c0d9342bc3f7b0ab1ee82dfb2eaf302;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf40be49688d6bcb931d751883735e37af8d59069b3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd431f96fccf4be568fe4057704d2a7163d1145dd2f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9241080371dcf8e3fffcb8aa96e0859637d6d171c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdb70e18ec28f8d38bebe6d200a25c81bb68b913c63;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8de04eb9ecf99d289e7501a6e75788c5c8b310a012;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h185dc04b77139a8386a9413dce1a2c9794e8a916974;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7e58d5c12179efae7b9c32bdb7a2e41dcef2e815eb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc453272758db0a17c92e3e5aed4ef8b74446d38da;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf773ebd8de68e6285a315dbe4dd55ae3164622520c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfda27531b96a96096635a3774acd3d5311c0502b84;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fd214ba1b9907fbd7e91abf1cc05e760767b64f19c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h21b08110424323776184c07d856b7524907778f98;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h507698df7c32500f7f89f5922d9eec0b74738aa878;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10b0300c80b913c18ec0bec62a2db111da83799c0b8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h81f001ab762df8d9f6eef9fbc9202b05d4b6368e1d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd3e94ada71d5473b147a8ddf0581827853fd05a76c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16080f313709e9a09cadd06273addbf176fe744e089;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c5476f49d7c4e16d488ac3fea9d2dcc2b23a7f63c4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h518e04422a475a41f7c06db9c62672cfdec0295d33;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbe947a2def7b88ad6f2d497aa3517dbbe483bfaa96;
        #1
        $finish();
    end
endmodule
