module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23);
    reg [255:0] src0;
    reg [255:0] src1;
    reg [255:0] src2;
    reg [255:0] src3;
    reg [255:0] src4;
    reg [255:0] src5;
    reg [255:0] src6;
    reg [255:0] src7;
    reg [255:0] src8;
    reg [255:0] src9;
    reg [255:0] src10;
    reg [255:0] src11;
    reg [255:0] src12;
    reg [255:0] src13;
    reg [255:0] src14;
    reg [255:0] src15;
    compressor_CLA256_16 compressor_CLA256_16(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23));
    initial begin
        src0 <= 256'h0;
        src1 <= 256'h0;
        src2 <= 256'h0;
        src3 <= 256'h0;
        src4 <= 256'h0;
        src5 <= 256'h0;
        src6 <= 256'h0;
        src7 <= 256'h0;
        src8 <= 256'h0;
        src9 <= 256'h0;
        src10 <= 256'h0;
        src11 <= 256'h0;
        src12 <= 256'h0;
        src13 <= 256'h0;
        src14 <= 256'h0;
        src15 <= 256'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
    end
endmodule
module compressor_CLA256_16(
    input [255:0]src0,
    input [255:0]src1,
    input [255:0]src2,
    input [255:0]src3,
    input [255:0]src4,
    input [255:0]src5,
    input [255:0]src6,
    input [255:0]src7,
    input [255:0]src8,
    input [255:0]src9,
    input [255:0]src10,
    input [255:0]src11,
    input [255:0]src12,
    input [255:0]src13,
    input [255:0]src14,
    input [255:0]src15,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [0:0] comp_out23;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [255:0] src0,
      input wire [255:0] src1,
      input wire [255:0] src2,
      input wire [255:0] src3,
      input wire [255:0] src4,
      input wire [255:0] src5,
      input wire [255:0] src6,
      input wire [255:0] src7,
      input wire [255:0] src8,
      input wire [255:0] src9,
      input wire [255:0] src10,
      input wire [255:0] src11,
      input wire [255:0] src12,
      input wire [255:0] src13,
      input wire [255:0] src14,
      input wire [255:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [0:0] dst23);

   wire [255:0] stage0_0;
   wire [255:0] stage0_1;
   wire [255:0] stage0_2;
   wire [255:0] stage0_3;
   wire [255:0] stage0_4;
   wire [255:0] stage0_5;
   wire [255:0] stage0_6;
   wire [255:0] stage0_7;
   wire [255:0] stage0_8;
   wire [255:0] stage0_9;
   wire [255:0] stage0_10;
   wire [255:0] stage0_11;
   wire [255:0] stage0_12;
   wire [255:0] stage0_13;
   wire [255:0] stage0_14;
   wire [255:0] stage0_15;
   wire [48:0] stage1_0;
   wire [97:0] stage1_1;
   wire [97:0] stage1_2;
   wire [113:0] stage1_3;
   wire [126:0] stage1_4;
   wire [104:0] stage1_5;
   wire [103:0] stage1_6;
   wire [114:0] stage1_7;
   wire [105:0] stage1_8;
   wire [115:0] stage1_9;
   wire [113:0] stage1_10;
   wire [114:0] stage1_11;
   wire [101:0] stage1_12;
   wire [132:0] stage1_13;
   wire [156:0] stage1_14;
   wire [75:0] stage1_15;
   wire [67:0] stage1_16;
   wire [41:0] stage1_17;
   wire [8:0] stage2_0;
   wire [25:0] stage2_1;
   wire [45:0] stage2_2;
   wire [33:0] stage2_3;
   wire [49:0] stage2_4;
   wire [54:0] stage2_5;
   wire [39:0] stage2_6;
   wire [58:0] stage2_7;
   wire [49:0] stage2_8;
   wire [47:0] stage2_9;
   wire [35:0] stage2_10;
   wire [47:0] stage2_11;
   wire [60:0] stage2_12;
   wire [44:0] stage2_13;
   wire [50:0] stage2_14;
   wire [50:0] stage2_15;
   wire [47:0] stage2_16;
   wire [33:0] stage2_17;
   wire [13:0] stage2_18;
   wire [4:0] stage2_19;
   wire [6:0] stage3_0;
   wire [5:0] stage3_1;
   wire [13:0] stage3_2;
   wire [13:0] stage3_3;
   wire [13:0] stage3_4;
   wire [19:0] stage3_5;
   wire [24:0] stage3_6;
   wire [22:0] stage3_7;
   wire [16:0] stage3_8;
   wire [20:0] stage3_9;
   wire [22:0] stage3_10;
   wire [16:0] stage3_11;
   wire [22:0] stage3_12;
   wire [20:0] stage3_13;
   wire [21:0] stage3_14;
   wire [24:0] stage3_15;
   wire [24:0] stage3_16;
   wire [18:0] stage3_17;
   wire [13:0] stage3_18;
   wire [11:0] stage3_19;
   wire [1:0] stage3_20;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [9:0] stage4_2;
   wire [5:0] stage4_3;
   wire [5:0] stage4_4;
   wire [5:0] stage4_5;
   wire [7:0] stage4_6;
   wire [16:0] stage4_7;
   wire [7:0] stage4_8;
   wire [8:0] stage4_9;
   wire [9:0] stage4_10;
   wire [9:0] stage4_11;
   wire [6:0] stage4_12;
   wire [7:0] stage4_13;
   wire [10:0] stage4_14;
   wire [8:0] stage4_15;
   wire [8:0] stage4_16;
   wire [9:0] stage4_17;
   wire [8:0] stage4_18;
   wire [9:0] stage4_19;
   wire [3:0] stage4_20;
   wire [1:0] stage4_21;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [5:0] stage5_2;
   wire [1:0] stage5_3;
   wire [6:0] stage5_4;
   wire [0:0] stage5_5;
   wire [4:0] stage5_6;
   wire [3:0] stage5_7;
   wire [3:0] stage5_8;
   wire [3:0] stage5_9;
   wire [5:0] stage5_10;
   wire [4:0] stage5_11;
   wire [2:0] stage5_12;
   wire [3:0] stage5_13;
   wire [3:0] stage5_14;
   wire [5:0] stage5_15;
   wire [4:0] stage5_16;
   wire [2:0] stage5_17;
   wire [3:0] stage5_18;
   wire [5:0] stage5_19;
   wire [5:0] stage5_20;
   wire [1:0] stage5_21;
   wire [0:0] stage5_22;
   wire [1:0] stage6_0;
   wire [1:0] stage6_1;
   wire [1:0] stage6_2;
   wire [1:0] stage6_3;
   wire [1:0] stage6_4;
   wire [1:0] stage6_5;
   wire [1:0] stage6_6;
   wire [1:0] stage6_7;
   wire [1:0] stage6_8;
   wire [1:0] stage6_9;
   wire [1:0] stage6_10;
   wire [1:0] stage6_11;
   wire [1:0] stage6_12;
   wire [1:0] stage6_13;
   wire [1:0] stage6_14;
   wire [1:0] stage6_15;
   wire [1:0] stage6_16;
   wire [1:0] stage6_17;
   wire [1:0] stage6_18;
   wire [1:0] stage6_19;
   wire [1:0] stage6_20;
   wire [1:0] stage6_21;
   wire [1:0] stage6_22;
   wire [0:0] stage6_23;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage6_0;
   assign dst1 = stage6_1;
   assign dst2 = stage6_2;
   assign dst3 = stage6_3;
   assign dst4 = stage6_4;
   assign dst5 = stage6_5;
   assign dst6 = stage6_6;
   assign dst7 = stage6_7;
   assign dst8 = stage6_8;
   assign dst9 = stage6_9;
   assign dst10 = stage6_10;
   assign dst11 = stage6_11;
   assign dst12 = stage6_12;
   assign dst13 = stage6_13;
   assign dst14 = stage6_14;
   assign dst15 = stage6_15;
   assign dst16 = stage6_16;
   assign dst17 = stage6_17;
   assign dst18 = stage6_18;
   assign dst19 = stage6_19;
   assign dst20 = stage6_20;
   assign dst21 = stage6_21;
   assign dst22 = stage6_22;
   assign dst23 = stage6_23;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc2135_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage0_3[4], stage0_3[5]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc2135_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[3]},
      {stage0_3[6], stage0_3[7]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc2135_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24]},
      {stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[4]},
      {stage0_3[8], stage0_3[9]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc2135_5 gpc5 (
      {stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[5]},
      {stage0_3[10], stage0_3[11]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc2135_5 gpc6 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_2[6]},
      {stage0_3[12], stage0_3[13]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc2135_5 gpc7 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39]},
      {stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[7]},
      {stage0_3[14], stage0_3[15]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc2135_5 gpc8 (
      {stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_1[24], stage0_1[25], stage0_1[26]},
      {stage0_2[8]},
      {stage0_3[16], stage0_3[17]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc2135_5 gpc9 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49]},
      {stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_2[9]},
      {stage0_3[18], stage0_3[19]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc2135_5 gpc10 (
      {stage0_0[50], stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54]},
      {stage0_1[30], stage0_1[31], stage0_1[32]},
      {stage0_2[10]},
      {stage0_3[20], stage0_3[21]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc2135_5 gpc11 (
      {stage0_0[55], stage0_0[56], stage0_0[57], stage0_0[58], stage0_0[59]},
      {stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_2[11]},
      {stage0_3[22], stage0_3[23]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc2135_5 gpc12 (
      {stage0_0[60], stage0_0[61], stage0_0[62], stage0_0[63], stage0_0[64]},
      {stage0_1[36], stage0_1[37], stage0_1[38]},
      {stage0_2[12]},
      {stage0_3[24], stage0_3[25]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc2135_5 gpc13 (
      {stage0_0[65], stage0_0[66], stage0_0[67], stage0_0[68], stage0_0[69]},
      {stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_2[13]},
      {stage0_3[26], stage0_3[27]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc2135_5 gpc14 (
      {stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74]},
      {stage0_1[42], stage0_1[43], stage0_1[44]},
      {stage0_2[14]},
      {stage0_3[28], stage0_3[29]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc2135_5 gpc15 (
      {stage0_0[75], stage0_0[76], stage0_0[77], stage0_0[78], stage0_0[79]},
      {stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_2[15]},
      {stage0_3[30], stage0_3[31]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc2135_5 gpc16 (
      {stage0_0[80], stage0_0[81], stage0_0[82], stage0_0[83], stage0_0[84]},
      {stage0_1[48], stage0_1[49], stage0_1[50]},
      {stage0_2[16]},
      {stage0_3[32], stage0_3[33]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc117_4 gpc17 (
      {stage0_0[85], stage0_0[86], stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91]},
      {stage0_1[51]},
      {stage0_2[17]},
      {stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc117_4 gpc18 (
      {stage0_0[92], stage0_0[93], stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97], stage0_0[98]},
      {stage0_1[52]},
      {stage0_2[18]},
      {stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc117_4 gpc19 (
      {stage0_0[99], stage0_0[100], stage0_0[101], stage0_0[102], stage0_0[103], stage0_0[104], stage0_0[105]},
      {stage0_1[53]},
      {stage0_2[19]},
      {stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc1163_5 gpc20 (
      {stage0_0[106], stage0_0[107], stage0_0[108]},
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59]},
      {stage0_2[20]},
      {stage0_3[34]},
      {stage1_4[17],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc1163_5 gpc21 (
      {stage0_0[109], stage0_0[110], stage0_0[111]},
      {stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65]},
      {stage0_2[21]},
      {stage0_3[35]},
      {stage1_4[18],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc1163_5 gpc22 (
      {stage0_0[112], stage0_0[113], stage0_0[114]},
      {stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71]},
      {stage0_2[22]},
      {stage0_3[36]},
      {stage1_4[19],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc1163_5 gpc23 (
      {stage0_0[115], stage0_0[116], stage0_0[117]},
      {stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77]},
      {stage0_2[23]},
      {stage0_3[37]},
      {stage1_4[20],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc1163_5 gpc24 (
      {stage0_0[118], stage0_0[119], stage0_0[120]},
      {stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83]},
      {stage0_2[24]},
      {stage0_3[38]},
      {stage1_4[21],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc1163_5 gpc25 (
      {stage0_0[121], stage0_0[122], stage0_0[123]},
      {stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89]},
      {stage0_2[25]},
      {stage0_3[39]},
      {stage1_4[22],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc1163_5 gpc26 (
      {stage0_0[124], stage0_0[125], stage0_0[126]},
      {stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95]},
      {stage0_2[26]},
      {stage0_3[40]},
      {stage1_4[23],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc1163_5 gpc27 (
      {stage0_0[127], stage0_0[128], stage0_0[129]},
      {stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101]},
      {stage0_2[27]},
      {stage0_3[41]},
      {stage1_4[24],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc606_5 gpc28 (
      {stage0_0[130], stage0_0[131], stage0_0[132], stage0_0[133], stage0_0[134], stage0_0[135]},
      {stage0_2[28], stage0_2[29], stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33]},
      {stage1_4[25],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc606_5 gpc29 (
      {stage0_0[136], stage0_0[137], stage0_0[138], stage0_0[139], stage0_0[140], stage0_0[141]},
      {stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39]},
      {stage1_4[26],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc606_5 gpc30 (
      {stage0_0[142], stage0_0[143], stage0_0[144], stage0_0[145], stage0_0[146], stage0_0[147]},
      {stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45]},
      {stage1_4[27],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc606_5 gpc31 (
      {stage0_0[148], stage0_0[149], stage0_0[150], stage0_0[151], stage0_0[152], stage0_0[153]},
      {stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49], stage0_2[50], stage0_2[51]},
      {stage1_4[28],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc606_5 gpc32 (
      {stage0_0[154], stage0_0[155], stage0_0[156], stage0_0[157], stage0_0[158], stage0_0[159]},
      {stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57]},
      {stage1_4[29],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc606_5 gpc33 (
      {stage0_0[160], stage0_0[161], stage0_0[162], stage0_0[163], stage0_0[164], stage0_0[165]},
      {stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61], stage0_2[62], stage0_2[63]},
      {stage1_4[30],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc606_5 gpc34 (
      {stage0_0[166], stage0_0[167], stage0_0[168], stage0_0[169], stage0_0[170], stage0_0[171]},
      {stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67], stage0_2[68], stage0_2[69]},
      {stage1_4[31],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc606_5 gpc35 (
      {stage0_0[172], stage0_0[173], stage0_0[174], stage0_0[175], stage0_0[176], stage0_0[177]},
      {stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73], stage0_2[74], stage0_2[75]},
      {stage1_4[32],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc606_5 gpc36 (
      {stage0_0[178], stage0_0[179], stage0_0[180], stage0_0[181], stage0_0[182], stage0_0[183]},
      {stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79], stage0_2[80], stage0_2[81]},
      {stage1_4[33],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc606_5 gpc37 (
      {stage0_0[184], stage0_0[185], stage0_0[186], stage0_0[187], stage0_0[188], stage0_0[189]},
      {stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85], stage0_2[86], stage0_2[87]},
      {stage1_4[34],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc606_5 gpc38 (
      {stage0_0[190], stage0_0[191], stage0_0[192], stage0_0[193], stage0_0[194], stage0_0[195]},
      {stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91], stage0_2[92], stage0_2[93]},
      {stage1_4[35],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc606_5 gpc39 (
      {stage0_0[196], stage0_0[197], stage0_0[198], stage0_0[199], stage0_0[200], stage0_0[201]},
      {stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97], stage0_2[98], stage0_2[99]},
      {stage1_4[36],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc606_5 gpc40 (
      {stage0_0[202], stage0_0[203], stage0_0[204], stage0_0[205], stage0_0[206], stage0_0[207]},
      {stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103], stage0_2[104], stage0_2[105]},
      {stage1_4[37],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc606_5 gpc41 (
      {stage0_0[208], stage0_0[209], stage0_0[210], stage0_0[211], stage0_0[212], stage0_0[213]},
      {stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109], stage0_2[110], stage0_2[111]},
      {stage1_4[38],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc606_5 gpc42 (
      {stage0_0[214], stage0_0[215], stage0_0[216], stage0_0[217], stage0_0[218], stage0_0[219]},
      {stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115], stage0_2[116], stage0_2[117]},
      {stage1_4[39],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc606_5 gpc43 (
      {stage0_0[220], stage0_0[221], stage0_0[222], stage0_0[223], stage0_0[224], stage0_0[225]},
      {stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121], stage0_2[122], stage0_2[123]},
      {stage1_4[40],stage1_3[43],stage1_2[43],stage1_1[43],stage1_0[43]}
   );
   gpc606_5 gpc44 (
      {stage0_0[226], stage0_0[227], stage0_0[228], stage0_0[229], stage0_0[230], stage0_0[231]},
      {stage0_2[124], stage0_2[125], stage0_2[126], stage0_2[127], stage0_2[128], stage0_2[129]},
      {stage1_4[41],stage1_3[44],stage1_2[44],stage1_1[44],stage1_0[44]}
   );
   gpc606_5 gpc45 (
      {stage0_0[232], stage0_0[233], stage0_0[234], stage0_0[235], stage0_0[236], stage0_0[237]},
      {stage0_2[130], stage0_2[131], stage0_2[132], stage0_2[133], stage0_2[134], stage0_2[135]},
      {stage1_4[42],stage1_3[45],stage1_2[45],stage1_1[45],stage1_0[45]}
   );
   gpc606_5 gpc46 (
      {stage0_0[238], stage0_0[239], stage0_0[240], stage0_0[241], stage0_0[242], stage0_0[243]},
      {stage0_2[136], stage0_2[137], stage0_2[138], stage0_2[139], stage0_2[140], stage0_2[141]},
      {stage1_4[43],stage1_3[46],stage1_2[46],stage1_1[46],stage1_0[46]}
   );
   gpc606_5 gpc47 (
      {stage0_0[244], stage0_0[245], stage0_0[246], stage0_0[247], stage0_0[248], stage0_0[249]},
      {stage0_2[142], stage0_2[143], stage0_2[144], stage0_2[145], stage0_2[146], stage0_2[147]},
      {stage1_4[44],stage1_3[47],stage1_2[47],stage1_1[47],stage1_0[47]}
   );
   gpc606_5 gpc48 (
      {stage0_0[250], stage0_0[251], stage0_0[252], stage0_0[253], stage0_0[254], stage0_0[255]},
      {stage0_2[148], stage0_2[149], stage0_2[150], stage0_2[151], stage0_2[152], stage0_2[153]},
      {stage1_4[45],stage1_3[48],stage1_2[48],stage1_1[48],stage1_0[48]}
   );
   gpc606_5 gpc49 (
      {stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107]},
      {stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47]},
      {stage1_5[0],stage1_4[46],stage1_3[49],stage1_2[49],stage1_1[49]}
   );
   gpc606_5 gpc50 (
      {stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113]},
      {stage0_3[48], stage0_3[49], stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53]},
      {stage1_5[1],stage1_4[47],stage1_3[50],stage1_2[50],stage1_1[50]}
   );
   gpc606_5 gpc51 (
      {stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119]},
      {stage0_3[54], stage0_3[55], stage0_3[56], stage0_3[57], stage0_3[58], stage0_3[59]},
      {stage1_5[2],stage1_4[48],stage1_3[51],stage1_2[51],stage1_1[51]}
   );
   gpc606_5 gpc52 (
      {stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125]},
      {stage0_3[60], stage0_3[61], stage0_3[62], stage0_3[63], stage0_3[64], stage0_3[65]},
      {stage1_5[3],stage1_4[49],stage1_3[52],stage1_2[52],stage1_1[52]}
   );
   gpc606_5 gpc53 (
      {stage0_1[126], stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131]},
      {stage0_3[66], stage0_3[67], stage0_3[68], stage0_3[69], stage0_3[70], stage0_3[71]},
      {stage1_5[4],stage1_4[50],stage1_3[53],stage1_2[53],stage1_1[53]}
   );
   gpc606_5 gpc54 (
      {stage0_1[132], stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137]},
      {stage0_3[72], stage0_3[73], stage0_3[74], stage0_3[75], stage0_3[76], stage0_3[77]},
      {stage1_5[5],stage1_4[51],stage1_3[54],stage1_2[54],stage1_1[54]}
   );
   gpc606_5 gpc55 (
      {stage0_1[138], stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143]},
      {stage0_3[78], stage0_3[79], stage0_3[80], stage0_3[81], stage0_3[82], stage0_3[83]},
      {stage1_5[6],stage1_4[52],stage1_3[55],stage1_2[55],stage1_1[55]}
   );
   gpc606_5 gpc56 (
      {stage0_1[144], stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149]},
      {stage0_3[84], stage0_3[85], stage0_3[86], stage0_3[87], stage0_3[88], stage0_3[89]},
      {stage1_5[7],stage1_4[53],stage1_3[56],stage1_2[56],stage1_1[56]}
   );
   gpc606_5 gpc57 (
      {stage0_1[150], stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155]},
      {stage0_3[90], stage0_3[91], stage0_3[92], stage0_3[93], stage0_3[94], stage0_3[95]},
      {stage1_5[8],stage1_4[54],stage1_3[57],stage1_2[57],stage1_1[57]}
   );
   gpc606_5 gpc58 (
      {stage0_1[156], stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161]},
      {stage0_3[96], stage0_3[97], stage0_3[98], stage0_3[99], stage0_3[100], stage0_3[101]},
      {stage1_5[9],stage1_4[55],stage1_3[58],stage1_2[58],stage1_1[58]}
   );
   gpc606_5 gpc59 (
      {stage0_1[162], stage0_1[163], stage0_1[164], stage0_1[165], stage0_1[166], stage0_1[167]},
      {stage0_3[102], stage0_3[103], stage0_3[104], stage0_3[105], stage0_3[106], stage0_3[107]},
      {stage1_5[10],stage1_4[56],stage1_3[59],stage1_2[59],stage1_1[59]}
   );
   gpc606_5 gpc60 (
      {stage0_1[168], stage0_1[169], stage0_1[170], stage0_1[171], stage0_1[172], stage0_1[173]},
      {stage0_3[108], stage0_3[109], stage0_3[110], stage0_3[111], stage0_3[112], stage0_3[113]},
      {stage1_5[11],stage1_4[57],stage1_3[60],stage1_2[60],stage1_1[60]}
   );
   gpc606_5 gpc61 (
      {stage0_1[174], stage0_1[175], stage0_1[176], stage0_1[177], stage0_1[178], stage0_1[179]},
      {stage0_3[114], stage0_3[115], stage0_3[116], stage0_3[117], stage0_3[118], stage0_3[119]},
      {stage1_5[12],stage1_4[58],stage1_3[61],stage1_2[61],stage1_1[61]}
   );
   gpc606_5 gpc62 (
      {stage0_1[180], stage0_1[181], stage0_1[182], stage0_1[183], stage0_1[184], stage0_1[185]},
      {stage0_3[120], stage0_3[121], stage0_3[122], stage0_3[123], stage0_3[124], stage0_3[125]},
      {stage1_5[13],stage1_4[59],stage1_3[62],stage1_2[62],stage1_1[62]}
   );
   gpc606_5 gpc63 (
      {stage0_1[186], stage0_1[187], stage0_1[188], stage0_1[189], stage0_1[190], stage0_1[191]},
      {stage0_3[126], stage0_3[127], stage0_3[128], stage0_3[129], stage0_3[130], stage0_3[131]},
      {stage1_5[14],stage1_4[60],stage1_3[63],stage1_2[63],stage1_1[63]}
   );
   gpc606_5 gpc64 (
      {stage0_1[192], stage0_1[193], stage0_1[194], stage0_1[195], stage0_1[196], stage0_1[197]},
      {stage0_3[132], stage0_3[133], stage0_3[134], stage0_3[135], stage0_3[136], stage0_3[137]},
      {stage1_5[15],stage1_4[61],stage1_3[64],stage1_2[64],stage1_1[64]}
   );
   gpc606_5 gpc65 (
      {stage0_1[198], stage0_1[199], stage0_1[200], stage0_1[201], stage0_1[202], stage0_1[203]},
      {stage0_3[138], stage0_3[139], stage0_3[140], stage0_3[141], stage0_3[142], stage0_3[143]},
      {stage1_5[16],stage1_4[62],stage1_3[65],stage1_2[65],stage1_1[65]}
   );
   gpc606_5 gpc66 (
      {stage0_1[204], stage0_1[205], stage0_1[206], stage0_1[207], stage0_1[208], stage0_1[209]},
      {stage0_3[144], stage0_3[145], stage0_3[146], stage0_3[147], stage0_3[148], stage0_3[149]},
      {stage1_5[17],stage1_4[63],stage1_3[66],stage1_2[66],stage1_1[66]}
   );
   gpc606_5 gpc67 (
      {stage0_1[210], stage0_1[211], stage0_1[212], stage0_1[213], stage0_1[214], stage0_1[215]},
      {stage0_3[150], stage0_3[151], stage0_3[152], stage0_3[153], stage0_3[154], stage0_3[155]},
      {stage1_5[18],stage1_4[64],stage1_3[67],stage1_2[67],stage1_1[67]}
   );
   gpc606_5 gpc68 (
      {stage0_1[216], stage0_1[217], stage0_1[218], stage0_1[219], stage0_1[220], stage0_1[221]},
      {stage0_3[156], stage0_3[157], stage0_3[158], stage0_3[159], stage0_3[160], stage0_3[161]},
      {stage1_5[19],stage1_4[65],stage1_3[68],stage1_2[68],stage1_1[68]}
   );
   gpc606_5 gpc69 (
      {stage0_1[222], stage0_1[223], stage0_1[224], stage0_1[225], stage0_1[226], stage0_1[227]},
      {stage0_3[162], stage0_3[163], stage0_3[164], stage0_3[165], stage0_3[166], stage0_3[167]},
      {stage1_5[20],stage1_4[66],stage1_3[69],stage1_2[69],stage1_1[69]}
   );
   gpc606_5 gpc70 (
      {stage0_2[154], stage0_2[155], stage0_2[156], stage0_2[157], stage0_2[158], stage0_2[159]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[21],stage1_4[67],stage1_3[70],stage1_2[70]}
   );
   gpc606_5 gpc71 (
      {stage0_2[160], stage0_2[161], stage0_2[162], stage0_2[163], stage0_2[164], stage0_2[165]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[22],stage1_4[68],stage1_3[71],stage1_2[71]}
   );
   gpc615_5 gpc72 (
      {stage0_2[166], stage0_2[167], stage0_2[168], stage0_2[169], stage0_2[170]},
      {stage0_3[168]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[23],stage1_4[69],stage1_3[72],stage1_2[72]}
   );
   gpc615_5 gpc73 (
      {stage0_2[171], stage0_2[172], stage0_2[173], stage0_2[174], stage0_2[175]},
      {stage0_3[169]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[24],stage1_4[70],stage1_3[73],stage1_2[73]}
   );
   gpc615_5 gpc74 (
      {stage0_2[176], stage0_2[177], stage0_2[178], stage0_2[179], stage0_2[180]},
      {stage0_3[170]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[25],stage1_4[71],stage1_3[74],stage1_2[74]}
   );
   gpc615_5 gpc75 (
      {stage0_2[181], stage0_2[182], stage0_2[183], stage0_2[184], stage0_2[185]},
      {stage0_3[171]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[26],stage1_4[72],stage1_3[75],stage1_2[75]}
   );
   gpc615_5 gpc76 (
      {stage0_2[186], stage0_2[187], stage0_2[188], stage0_2[189], stage0_2[190]},
      {stage0_3[172]},
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage1_6[6],stage1_5[27],stage1_4[73],stage1_3[76],stage1_2[76]}
   );
   gpc615_5 gpc77 (
      {stage0_2[191], stage0_2[192], stage0_2[193], stage0_2[194], stage0_2[195]},
      {stage0_3[173]},
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage1_6[7],stage1_5[28],stage1_4[74],stage1_3[77],stage1_2[77]}
   );
   gpc615_5 gpc78 (
      {stage0_2[196], stage0_2[197], stage0_2[198], stage0_2[199], stage0_2[200]},
      {stage0_3[174]},
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage1_6[8],stage1_5[29],stage1_4[75],stage1_3[78],stage1_2[78]}
   );
   gpc615_5 gpc79 (
      {stage0_2[201], stage0_2[202], stage0_2[203], stage0_2[204], stage0_2[205]},
      {stage0_3[175]},
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage1_6[9],stage1_5[30],stage1_4[76],stage1_3[79],stage1_2[79]}
   );
   gpc615_5 gpc80 (
      {stage0_2[206], stage0_2[207], stage0_2[208], stage0_2[209], stage0_2[210]},
      {stage0_3[176]},
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage1_6[10],stage1_5[31],stage1_4[77],stage1_3[80],stage1_2[80]}
   );
   gpc615_5 gpc81 (
      {stage0_2[211], stage0_2[212], stage0_2[213], stage0_2[214], stage0_2[215]},
      {stage0_3[177]},
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage1_6[11],stage1_5[32],stage1_4[78],stage1_3[81],stage1_2[81]}
   );
   gpc615_5 gpc82 (
      {stage0_2[216], stage0_2[217], stage0_2[218], stage0_2[219], stage0_2[220]},
      {stage0_3[178]},
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage1_6[12],stage1_5[33],stage1_4[79],stage1_3[82],stage1_2[82]}
   );
   gpc615_5 gpc83 (
      {stage0_2[221], stage0_2[222], stage0_2[223], stage0_2[224], stage0_2[225]},
      {stage0_3[179]},
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage1_6[13],stage1_5[34],stage1_4[80],stage1_3[83],stage1_2[83]}
   );
   gpc615_5 gpc84 (
      {stage0_2[226], stage0_2[227], stage0_2[228], stage0_2[229], stage0_2[230]},
      {stage0_3[180]},
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage1_6[14],stage1_5[35],stage1_4[81],stage1_3[84],stage1_2[84]}
   );
   gpc615_5 gpc85 (
      {stage0_2[231], stage0_2[232], stage0_2[233], stage0_2[234], stage0_2[235]},
      {stage0_3[181]},
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage1_6[15],stage1_5[36],stage1_4[82],stage1_3[85],stage1_2[85]}
   );
   gpc615_5 gpc86 (
      {stage0_2[236], stage0_2[237], stage0_2[238], stage0_2[239], stage0_2[240]},
      {stage0_3[182]},
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage1_6[16],stage1_5[37],stage1_4[83],stage1_3[86],stage1_2[86]}
   );
   gpc615_5 gpc87 (
      {stage0_2[241], stage0_2[242], stage0_2[243], stage0_2[244], stage0_2[245]},
      {stage0_3[183]},
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage1_6[17],stage1_5[38],stage1_4[84],stage1_3[87],stage1_2[87]}
   );
   gpc1343_5 gpc88 (
      {stage0_3[184], stage0_3[185], stage0_3[186]},
      {stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111]},
      {stage0_5[0], stage0_5[1], stage0_5[2]},
      {stage0_6[0]},
      {stage1_7[0],stage1_6[18],stage1_5[39],stage1_4[85],stage1_3[88]}
   );
   gpc615_5 gpc89 (
      {stage0_3[187], stage0_3[188], stage0_3[189], stage0_3[190], stage0_3[191]},
      {stage0_4[112]},
      {stage0_5[3], stage0_5[4], stage0_5[5], stage0_5[6], stage0_5[7], stage0_5[8]},
      {stage1_7[1],stage1_6[19],stage1_5[40],stage1_4[86],stage1_3[89]}
   );
   gpc615_5 gpc90 (
      {stage0_3[192], stage0_3[193], stage0_3[194], stage0_3[195], stage0_3[196]},
      {stage0_4[113]},
      {stage0_5[9], stage0_5[10], stage0_5[11], stage0_5[12], stage0_5[13], stage0_5[14]},
      {stage1_7[2],stage1_6[20],stage1_5[41],stage1_4[87],stage1_3[90]}
   );
   gpc615_5 gpc91 (
      {stage0_3[197], stage0_3[198], stage0_3[199], stage0_3[200], stage0_3[201]},
      {stage0_4[114]},
      {stage0_5[15], stage0_5[16], stage0_5[17], stage0_5[18], stage0_5[19], stage0_5[20]},
      {stage1_7[3],stage1_6[21],stage1_5[42],stage1_4[88],stage1_3[91]}
   );
   gpc615_5 gpc92 (
      {stage0_3[202], stage0_3[203], stage0_3[204], stage0_3[205], stage0_3[206]},
      {stage0_4[115]},
      {stage0_5[21], stage0_5[22], stage0_5[23], stage0_5[24], stage0_5[25], stage0_5[26]},
      {stage1_7[4],stage1_6[22],stage1_5[43],stage1_4[89],stage1_3[92]}
   );
   gpc615_5 gpc93 (
      {stage0_3[207], stage0_3[208], stage0_3[209], stage0_3[210], stage0_3[211]},
      {stage0_4[116]},
      {stage0_5[27], stage0_5[28], stage0_5[29], stage0_5[30], stage0_5[31], stage0_5[32]},
      {stage1_7[5],stage1_6[23],stage1_5[44],stage1_4[90],stage1_3[93]}
   );
   gpc615_5 gpc94 (
      {stage0_3[212], stage0_3[213], stage0_3[214], stage0_3[215], stage0_3[216]},
      {stage0_4[117]},
      {stage0_5[33], stage0_5[34], stage0_5[35], stage0_5[36], stage0_5[37], stage0_5[38]},
      {stage1_7[6],stage1_6[24],stage1_5[45],stage1_4[91],stage1_3[94]}
   );
   gpc615_5 gpc95 (
      {stage0_3[217], stage0_3[218], stage0_3[219], stage0_3[220], stage0_3[221]},
      {stage0_4[118]},
      {stage0_5[39], stage0_5[40], stage0_5[41], stage0_5[42], stage0_5[43], stage0_5[44]},
      {stage1_7[7],stage1_6[25],stage1_5[46],stage1_4[92],stage1_3[95]}
   );
   gpc615_5 gpc96 (
      {stage0_3[222], stage0_3[223], stage0_3[224], stage0_3[225], stage0_3[226]},
      {stage0_4[119]},
      {stage0_5[45], stage0_5[46], stage0_5[47], stage0_5[48], stage0_5[49], stage0_5[50]},
      {stage1_7[8],stage1_6[26],stage1_5[47],stage1_4[93],stage1_3[96]}
   );
   gpc615_5 gpc97 (
      {stage0_3[227], stage0_3[228], stage0_3[229], stage0_3[230], stage0_3[231]},
      {stage0_4[120]},
      {stage0_5[51], stage0_5[52], stage0_5[53], stage0_5[54], stage0_5[55], stage0_5[56]},
      {stage1_7[9],stage1_6[27],stage1_5[48],stage1_4[94],stage1_3[97]}
   );
   gpc615_5 gpc98 (
      {stage0_3[232], stage0_3[233], stage0_3[234], stage0_3[235], stage0_3[236]},
      {stage0_4[121]},
      {stage0_5[57], stage0_5[58], stage0_5[59], stage0_5[60], stage0_5[61], stage0_5[62]},
      {stage1_7[10],stage1_6[28],stage1_5[49],stage1_4[95],stage1_3[98]}
   );
   gpc615_5 gpc99 (
      {stage0_3[237], stage0_3[238], stage0_3[239], stage0_3[240], stage0_3[241]},
      {stage0_4[122]},
      {stage0_5[63], stage0_5[64], stage0_5[65], stage0_5[66], stage0_5[67], stage0_5[68]},
      {stage1_7[11],stage1_6[29],stage1_5[50],stage1_4[96],stage1_3[99]}
   );
   gpc606_5 gpc100 (
      {stage0_4[123], stage0_4[124], stage0_4[125], stage0_4[126], stage0_4[127], stage0_4[128]},
      {stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5], stage0_6[6]},
      {stage1_8[0],stage1_7[12],stage1_6[30],stage1_5[51],stage1_4[97]}
   );
   gpc606_5 gpc101 (
      {stage0_4[129], stage0_4[130], stage0_4[131], stage0_4[132], stage0_4[133], stage0_4[134]},
      {stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11], stage0_6[12]},
      {stage1_8[1],stage1_7[13],stage1_6[31],stage1_5[52],stage1_4[98]}
   );
   gpc606_5 gpc102 (
      {stage0_4[135], stage0_4[136], stage0_4[137], stage0_4[138], stage0_4[139], stage0_4[140]},
      {stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17], stage0_6[18]},
      {stage1_8[2],stage1_7[14],stage1_6[32],stage1_5[53],stage1_4[99]}
   );
   gpc606_5 gpc103 (
      {stage0_4[141], stage0_4[142], stage0_4[143], stage0_4[144], stage0_4[145], stage0_4[146]},
      {stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23], stage0_6[24]},
      {stage1_8[3],stage1_7[15],stage1_6[33],stage1_5[54],stage1_4[100]}
   );
   gpc606_5 gpc104 (
      {stage0_4[147], stage0_4[148], stage0_4[149], stage0_4[150], stage0_4[151], stage0_4[152]},
      {stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29], stage0_6[30]},
      {stage1_8[4],stage1_7[16],stage1_6[34],stage1_5[55],stage1_4[101]}
   );
   gpc606_5 gpc105 (
      {stage0_4[153], stage0_4[154], stage0_4[155], stage0_4[156], stage0_4[157], stage0_4[158]},
      {stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35], stage0_6[36]},
      {stage1_8[5],stage1_7[17],stage1_6[35],stage1_5[56],stage1_4[102]}
   );
   gpc606_5 gpc106 (
      {stage0_4[159], stage0_4[160], stage0_4[161], stage0_4[162], stage0_4[163], stage0_4[164]},
      {stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41], stage0_6[42]},
      {stage1_8[6],stage1_7[18],stage1_6[36],stage1_5[57],stage1_4[103]}
   );
   gpc606_5 gpc107 (
      {stage0_4[165], stage0_4[166], stage0_4[167], stage0_4[168], stage0_4[169], stage0_4[170]},
      {stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47], stage0_6[48]},
      {stage1_8[7],stage1_7[19],stage1_6[37],stage1_5[58],stage1_4[104]}
   );
   gpc606_5 gpc108 (
      {stage0_4[171], stage0_4[172], stage0_4[173], stage0_4[174], stage0_4[175], stage0_4[176]},
      {stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53], stage0_6[54]},
      {stage1_8[8],stage1_7[20],stage1_6[38],stage1_5[59],stage1_4[105]}
   );
   gpc606_5 gpc109 (
      {stage0_4[177], stage0_4[178], stage0_4[179], stage0_4[180], stage0_4[181], stage0_4[182]},
      {stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59], stage0_6[60]},
      {stage1_8[9],stage1_7[21],stage1_6[39],stage1_5[60],stage1_4[106]}
   );
   gpc606_5 gpc110 (
      {stage0_4[183], stage0_4[184], stage0_4[185], stage0_4[186], stage0_4[187], stage0_4[188]},
      {stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65], stage0_6[66]},
      {stage1_8[10],stage1_7[22],stage1_6[40],stage1_5[61],stage1_4[107]}
   );
   gpc615_5 gpc111 (
      {stage0_4[189], stage0_4[190], stage0_4[191], stage0_4[192], stage0_4[193]},
      {stage0_5[69]},
      {stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71], stage0_6[72]},
      {stage1_8[11],stage1_7[23],stage1_6[41],stage1_5[62],stage1_4[108]}
   );
   gpc615_5 gpc112 (
      {stage0_4[194], stage0_4[195], stage0_4[196], stage0_4[197], stage0_4[198]},
      {stage0_5[70]},
      {stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77], stage0_6[78]},
      {stage1_8[12],stage1_7[24],stage1_6[42],stage1_5[63],stage1_4[109]}
   );
   gpc615_5 gpc113 (
      {stage0_4[199], stage0_4[200], stage0_4[201], stage0_4[202], stage0_4[203]},
      {stage0_5[71]},
      {stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83], stage0_6[84]},
      {stage1_8[13],stage1_7[25],stage1_6[43],stage1_5[64],stage1_4[110]}
   );
   gpc615_5 gpc114 (
      {stage0_4[204], stage0_4[205], stage0_4[206], stage0_4[207], stage0_4[208]},
      {stage0_5[72]},
      {stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89], stage0_6[90]},
      {stage1_8[14],stage1_7[26],stage1_6[44],stage1_5[65],stage1_4[111]}
   );
   gpc615_5 gpc115 (
      {stage0_4[209], stage0_4[210], stage0_4[211], stage0_4[212], stage0_4[213]},
      {stage0_5[73]},
      {stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95], stage0_6[96]},
      {stage1_8[15],stage1_7[27],stage1_6[45],stage1_5[66],stage1_4[112]}
   );
   gpc615_5 gpc116 (
      {stage0_4[214], stage0_4[215], stage0_4[216], stage0_4[217], stage0_4[218]},
      {stage0_5[74]},
      {stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101], stage0_6[102]},
      {stage1_8[16],stage1_7[28],stage1_6[46],stage1_5[67],stage1_4[113]}
   );
   gpc615_5 gpc117 (
      {stage0_4[219], stage0_4[220], stage0_4[221], stage0_4[222], stage0_4[223]},
      {stage0_5[75]},
      {stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107], stage0_6[108]},
      {stage1_8[17],stage1_7[29],stage1_6[47],stage1_5[68],stage1_4[114]}
   );
   gpc615_5 gpc118 (
      {stage0_4[224], stage0_4[225], stage0_4[226], stage0_4[227], stage0_4[228]},
      {stage0_5[76]},
      {stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113], stage0_6[114]},
      {stage1_8[18],stage1_7[30],stage1_6[48],stage1_5[69],stage1_4[115]}
   );
   gpc615_5 gpc119 (
      {stage0_4[229], stage0_4[230], stage0_4[231], stage0_4[232], stage0_4[233]},
      {stage0_5[77]},
      {stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119], stage0_6[120]},
      {stage1_8[19],stage1_7[31],stage1_6[49],stage1_5[70],stage1_4[116]}
   );
   gpc615_5 gpc120 (
      {stage0_4[234], stage0_4[235], stage0_4[236], stage0_4[237], stage0_4[238]},
      {stage0_5[78]},
      {stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125], stage0_6[126]},
      {stage1_8[20],stage1_7[32],stage1_6[50],stage1_5[71],stage1_4[117]}
   );
   gpc615_5 gpc121 (
      {stage0_4[239], stage0_4[240], stage0_4[241], stage0_4[242], stage0_4[243]},
      {stage0_5[79]},
      {stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131], stage0_6[132]},
      {stage1_8[21],stage1_7[33],stage1_6[51],stage1_5[72],stage1_4[118]}
   );
   gpc615_5 gpc122 (
      {stage0_4[244], stage0_4[245], stage0_4[246], stage0_4[247], stage0_4[248]},
      {stage0_5[80]},
      {stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137], stage0_6[138]},
      {stage1_8[22],stage1_7[34],stage1_6[52],stage1_5[73],stage1_4[119]}
   );
   gpc606_5 gpc123 (
      {stage0_5[81], stage0_5[82], stage0_5[83], stage0_5[84], stage0_5[85], stage0_5[86]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[23],stage1_7[35],stage1_6[53],stage1_5[74]}
   );
   gpc606_5 gpc124 (
      {stage0_5[87], stage0_5[88], stage0_5[89], stage0_5[90], stage0_5[91], stage0_5[92]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[24],stage1_7[36],stage1_6[54],stage1_5[75]}
   );
   gpc606_5 gpc125 (
      {stage0_5[93], stage0_5[94], stage0_5[95], stage0_5[96], stage0_5[97], stage0_5[98]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[25],stage1_7[37],stage1_6[55],stage1_5[76]}
   );
   gpc606_5 gpc126 (
      {stage0_5[99], stage0_5[100], stage0_5[101], stage0_5[102], stage0_5[103], stage0_5[104]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[26],stage1_7[38],stage1_6[56],stage1_5[77]}
   );
   gpc606_5 gpc127 (
      {stage0_5[105], stage0_5[106], stage0_5[107], stage0_5[108], stage0_5[109], stage0_5[110]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[27],stage1_7[39],stage1_6[57],stage1_5[78]}
   );
   gpc606_5 gpc128 (
      {stage0_5[111], stage0_5[112], stage0_5[113], stage0_5[114], stage0_5[115], stage0_5[116]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[28],stage1_7[40],stage1_6[58],stage1_5[79]}
   );
   gpc606_5 gpc129 (
      {stage0_5[117], stage0_5[118], stage0_5[119], stage0_5[120], stage0_5[121], stage0_5[122]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[29],stage1_7[41],stage1_6[59],stage1_5[80]}
   );
   gpc606_5 gpc130 (
      {stage0_5[123], stage0_5[124], stage0_5[125], stage0_5[126], stage0_5[127], stage0_5[128]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[30],stage1_7[42],stage1_6[60],stage1_5[81]}
   );
   gpc606_5 gpc131 (
      {stage0_5[129], stage0_5[130], stage0_5[131], stage0_5[132], stage0_5[133], stage0_5[134]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[31],stage1_7[43],stage1_6[61],stage1_5[82]}
   );
   gpc606_5 gpc132 (
      {stage0_5[135], stage0_5[136], stage0_5[137], stage0_5[138], stage0_5[139], stage0_5[140]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[32],stage1_7[44],stage1_6[62],stage1_5[83]}
   );
   gpc606_5 gpc133 (
      {stage0_5[141], stage0_5[142], stage0_5[143], stage0_5[144], stage0_5[145], stage0_5[146]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[33],stage1_7[45],stage1_6[63],stage1_5[84]}
   );
   gpc606_5 gpc134 (
      {stage0_5[147], stage0_5[148], stage0_5[149], stage0_5[150], stage0_5[151], stage0_5[152]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[34],stage1_7[46],stage1_6[64],stage1_5[85]}
   );
   gpc606_5 gpc135 (
      {stage0_5[153], stage0_5[154], stage0_5[155], stage0_5[156], stage0_5[157], stage0_5[158]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[35],stage1_7[47],stage1_6[65],stage1_5[86]}
   );
   gpc606_5 gpc136 (
      {stage0_5[159], stage0_5[160], stage0_5[161], stage0_5[162], stage0_5[163], stage0_5[164]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[36],stage1_7[48],stage1_6[66],stage1_5[87]}
   );
   gpc606_5 gpc137 (
      {stage0_5[165], stage0_5[166], stage0_5[167], stage0_5[168], stage0_5[169], stage0_5[170]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[37],stage1_7[49],stage1_6[67],stage1_5[88]}
   );
   gpc606_5 gpc138 (
      {stage0_5[171], stage0_5[172], stage0_5[173], stage0_5[174], stage0_5[175], stage0_5[176]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[38],stage1_7[50],stage1_6[68],stage1_5[89]}
   );
   gpc606_5 gpc139 (
      {stage0_5[177], stage0_5[178], stage0_5[179], stage0_5[180], stage0_5[181], stage0_5[182]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[39],stage1_7[51],stage1_6[69],stage1_5[90]}
   );
   gpc606_5 gpc140 (
      {stage0_5[183], stage0_5[184], stage0_5[185], stage0_5[186], stage0_5[187], stage0_5[188]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[40],stage1_7[52],stage1_6[70],stage1_5[91]}
   );
   gpc606_5 gpc141 (
      {stage0_5[189], stage0_5[190], stage0_5[191], stage0_5[192], stage0_5[193], stage0_5[194]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[41],stage1_7[53],stage1_6[71],stage1_5[92]}
   );
   gpc606_5 gpc142 (
      {stage0_5[195], stage0_5[196], stage0_5[197], stage0_5[198], stage0_5[199], stage0_5[200]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[42],stage1_7[54],stage1_6[72],stage1_5[93]}
   );
   gpc606_5 gpc143 (
      {stage0_5[201], stage0_5[202], stage0_5[203], stage0_5[204], stage0_5[205], stage0_5[206]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[43],stage1_7[55],stage1_6[73],stage1_5[94]}
   );
   gpc606_5 gpc144 (
      {stage0_5[207], stage0_5[208], stage0_5[209], stage0_5[210], stage0_5[211], stage0_5[212]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[44],stage1_7[56],stage1_6[74],stage1_5[95]}
   );
   gpc606_5 gpc145 (
      {stage0_5[213], stage0_5[214], stage0_5[215], stage0_5[216], stage0_5[217], stage0_5[218]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[45],stage1_7[57],stage1_6[75],stage1_5[96]}
   );
   gpc606_5 gpc146 (
      {stage0_5[219], stage0_5[220], stage0_5[221], stage0_5[222], stage0_5[223], stage0_5[224]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[46],stage1_7[58],stage1_6[76],stage1_5[97]}
   );
   gpc606_5 gpc147 (
      {stage0_5[225], stage0_5[226], stage0_5[227], stage0_5[228], stage0_5[229], stage0_5[230]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[47],stage1_7[59],stage1_6[77],stage1_5[98]}
   );
   gpc606_5 gpc148 (
      {stage0_5[231], stage0_5[232], stage0_5[233], stage0_5[234], stage0_5[235], stage0_5[236]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[48],stage1_7[60],stage1_6[78],stage1_5[99]}
   );
   gpc606_5 gpc149 (
      {stage0_5[237], stage0_5[238], stage0_5[239], stage0_5[240], stage0_5[241], stage0_5[242]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[49],stage1_7[61],stage1_6[79],stage1_5[100]}
   );
   gpc606_5 gpc150 (
      {stage0_5[243], stage0_5[244], stage0_5[245], stage0_5[246], stage0_5[247], stage0_5[248]},
      {stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167]},
      {stage1_9[27],stage1_8[50],stage1_7[62],stage1_6[80],stage1_5[101]}
   );
   gpc615_5 gpc151 (
      {stage0_5[249], stage0_5[250], stage0_5[251], stage0_5[252], stage0_5[253]},
      {stage0_6[139]},
      {stage0_7[168], stage0_7[169], stage0_7[170], stage0_7[171], stage0_7[172], stage0_7[173]},
      {stage1_9[28],stage1_8[51],stage1_7[63],stage1_6[81],stage1_5[102]}
   );
   gpc606_5 gpc152 (
      {stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143], stage0_6[144], stage0_6[145]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[29],stage1_8[52],stage1_7[64],stage1_6[82]}
   );
   gpc606_5 gpc153 (
      {stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149], stage0_6[150], stage0_6[151]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[30],stage1_8[53],stage1_7[65],stage1_6[83]}
   );
   gpc606_5 gpc154 (
      {stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155], stage0_6[156], stage0_6[157]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[31],stage1_8[54],stage1_7[66],stage1_6[84]}
   );
   gpc606_5 gpc155 (
      {stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161], stage0_6[162], stage0_6[163]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[32],stage1_8[55],stage1_7[67],stage1_6[85]}
   );
   gpc606_5 gpc156 (
      {stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167], stage0_6[168], stage0_6[169]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[33],stage1_8[56],stage1_7[68],stage1_6[86]}
   );
   gpc606_5 gpc157 (
      {stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173], stage0_6[174], stage0_6[175]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[34],stage1_8[57],stage1_7[69],stage1_6[87]}
   );
   gpc606_5 gpc158 (
      {stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179], stage0_6[180], stage0_6[181]},
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage1_10[6],stage1_9[35],stage1_8[58],stage1_7[70],stage1_6[88]}
   );
   gpc606_5 gpc159 (
      {stage0_6[182], stage0_6[183], stage0_6[184], stage0_6[185], stage0_6[186], stage0_6[187]},
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage1_10[7],stage1_9[36],stage1_8[59],stage1_7[71],stage1_6[89]}
   );
   gpc606_5 gpc160 (
      {stage0_6[188], stage0_6[189], stage0_6[190], stage0_6[191], stage0_6[192], stage0_6[193]},
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage1_10[8],stage1_9[37],stage1_8[60],stage1_7[72],stage1_6[90]}
   );
   gpc606_5 gpc161 (
      {stage0_6[194], stage0_6[195], stage0_6[196], stage0_6[197], stage0_6[198], stage0_6[199]},
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage1_10[9],stage1_9[38],stage1_8[61],stage1_7[73],stage1_6[91]}
   );
   gpc615_5 gpc162 (
      {stage0_6[200], stage0_6[201], stage0_6[202], stage0_6[203], stage0_6[204]},
      {stage0_7[174]},
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage1_10[10],stage1_9[39],stage1_8[62],stage1_7[74],stage1_6[92]}
   );
   gpc615_5 gpc163 (
      {stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208], stage0_6[209]},
      {stage0_7[175]},
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage1_10[11],stage1_9[40],stage1_8[63],stage1_7[75],stage1_6[93]}
   );
   gpc615_5 gpc164 (
      {stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214]},
      {stage0_7[176]},
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77]},
      {stage1_10[12],stage1_9[41],stage1_8[64],stage1_7[76],stage1_6[94]}
   );
   gpc615_5 gpc165 (
      {stage0_6[215], stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219]},
      {stage0_7[177]},
      {stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83]},
      {stage1_10[13],stage1_9[42],stage1_8[65],stage1_7[77],stage1_6[95]}
   );
   gpc615_5 gpc166 (
      {stage0_6[220], stage0_6[221], stage0_6[222], stage0_6[223], stage0_6[224]},
      {stage0_7[178]},
      {stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89]},
      {stage1_10[14],stage1_9[43],stage1_8[66],stage1_7[78],stage1_6[96]}
   );
   gpc615_5 gpc167 (
      {stage0_6[225], stage0_6[226], stage0_6[227], stage0_6[228], stage0_6[229]},
      {stage0_7[179]},
      {stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95]},
      {stage1_10[15],stage1_9[44],stage1_8[67],stage1_7[79],stage1_6[97]}
   );
   gpc615_5 gpc168 (
      {stage0_6[230], stage0_6[231], stage0_6[232], stage0_6[233], stage0_6[234]},
      {stage0_7[180]},
      {stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101]},
      {stage1_10[16],stage1_9[45],stage1_8[68],stage1_7[80],stage1_6[98]}
   );
   gpc615_5 gpc169 (
      {stage0_6[235], stage0_6[236], stage0_6[237], stage0_6[238], stage0_6[239]},
      {stage0_7[181]},
      {stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107]},
      {stage1_10[17],stage1_9[46],stage1_8[69],stage1_7[81],stage1_6[99]}
   );
   gpc615_5 gpc170 (
      {stage0_6[240], stage0_6[241], stage0_6[242], stage0_6[243], stage0_6[244]},
      {stage0_7[182]},
      {stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113]},
      {stage1_10[18],stage1_9[47],stage1_8[70],stage1_7[82],stage1_6[100]}
   );
   gpc615_5 gpc171 (
      {stage0_6[245], stage0_6[246], stage0_6[247], stage0_6[248], stage0_6[249]},
      {stage0_7[183]},
      {stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119]},
      {stage1_10[19],stage1_9[48],stage1_8[71],stage1_7[83],stage1_6[101]}
   );
   gpc615_5 gpc172 (
      {stage0_6[250], stage0_6[251], stage0_6[252], stage0_6[253], stage0_6[254]},
      {stage0_7[184]},
      {stage0_8[120], stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125]},
      {stage1_10[20],stage1_9[49],stage1_8[72],stage1_7[84],stage1_6[102]}
   );
   gpc606_5 gpc173 (
      {stage0_7[185], stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189], stage0_7[190]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[21],stage1_9[50],stage1_8[73],stage1_7[85]}
   );
   gpc615_5 gpc174 (
      {stage0_7[191], stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195]},
      {stage0_8[126]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[22],stage1_9[51],stage1_8[74],stage1_7[86]}
   );
   gpc615_5 gpc175 (
      {stage0_7[196], stage0_7[197], stage0_7[198], stage0_7[199], stage0_7[200]},
      {stage0_8[127]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[23],stage1_9[52],stage1_8[75],stage1_7[87]}
   );
   gpc615_5 gpc176 (
      {stage0_7[201], stage0_7[202], stage0_7[203], stage0_7[204], stage0_7[205]},
      {stage0_8[128]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[24],stage1_9[53],stage1_8[76],stage1_7[88]}
   );
   gpc615_5 gpc177 (
      {stage0_7[206], stage0_7[207], stage0_7[208], stage0_7[209], stage0_7[210]},
      {stage0_8[129]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[25],stage1_9[54],stage1_8[77],stage1_7[89]}
   );
   gpc615_5 gpc178 (
      {stage0_7[211], stage0_7[212], stage0_7[213], stage0_7[214], stage0_7[215]},
      {stage0_8[130]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[26],stage1_9[55],stage1_8[78],stage1_7[90]}
   );
   gpc615_5 gpc179 (
      {stage0_7[216], stage0_7[217], stage0_7[218], stage0_7[219], stage0_7[220]},
      {stage0_8[131]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[27],stage1_9[56],stage1_8[79],stage1_7[91]}
   );
   gpc615_5 gpc180 (
      {stage0_7[221], stage0_7[222], stage0_7[223], stage0_7[224], stage0_7[225]},
      {stage0_8[132]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[28],stage1_9[57],stage1_8[80],stage1_7[92]}
   );
   gpc615_5 gpc181 (
      {stage0_7[226], stage0_7[227], stage0_7[228], stage0_7[229], stage0_7[230]},
      {stage0_8[133]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[29],stage1_9[58],stage1_8[81],stage1_7[93]}
   );
   gpc615_5 gpc182 (
      {stage0_7[231], stage0_7[232], stage0_7[233], stage0_7[234], stage0_7[235]},
      {stage0_8[134]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[30],stage1_9[59],stage1_8[82],stage1_7[94]}
   );
   gpc606_5 gpc183 (
      {stage0_8[135], stage0_8[136], stage0_8[137], stage0_8[138], stage0_8[139], stage0_8[140]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[10],stage1_10[31],stage1_9[60],stage1_8[83]}
   );
   gpc606_5 gpc184 (
      {stage0_8[141], stage0_8[142], stage0_8[143], stage0_8[144], stage0_8[145], stage0_8[146]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[11],stage1_10[32],stage1_9[61],stage1_8[84]}
   );
   gpc606_5 gpc185 (
      {stage0_8[147], stage0_8[148], stage0_8[149], stage0_8[150], stage0_8[151], stage0_8[152]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[12],stage1_10[33],stage1_9[62],stage1_8[85]}
   );
   gpc606_5 gpc186 (
      {stage0_8[153], stage0_8[154], stage0_8[155], stage0_8[156], stage0_8[157], stage0_8[158]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[13],stage1_10[34],stage1_9[63],stage1_8[86]}
   );
   gpc606_5 gpc187 (
      {stage0_8[159], stage0_8[160], stage0_8[161], stage0_8[162], stage0_8[163], stage0_8[164]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[14],stage1_10[35],stage1_9[64],stage1_8[87]}
   );
   gpc606_5 gpc188 (
      {stage0_8[165], stage0_8[166], stage0_8[167], stage0_8[168], stage0_8[169], stage0_8[170]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[15],stage1_10[36],stage1_9[65],stage1_8[88]}
   );
   gpc606_5 gpc189 (
      {stage0_8[171], stage0_8[172], stage0_8[173], stage0_8[174], stage0_8[175], stage0_8[176]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[16],stage1_10[37],stage1_9[66],stage1_8[89]}
   );
   gpc606_5 gpc190 (
      {stage0_8[177], stage0_8[178], stage0_8[179], stage0_8[180], stage0_8[181], stage0_8[182]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[17],stage1_10[38],stage1_9[67],stage1_8[90]}
   );
   gpc606_5 gpc191 (
      {stage0_8[183], stage0_8[184], stage0_8[185], stage0_8[186], stage0_8[187], stage0_8[188]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[18],stage1_10[39],stage1_9[68],stage1_8[91]}
   );
   gpc606_5 gpc192 (
      {stage0_8[189], stage0_8[190], stage0_8[191], stage0_8[192], stage0_8[193], stage0_8[194]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[19],stage1_10[40],stage1_9[69],stage1_8[92]}
   );
   gpc615_5 gpc193 (
      {stage0_8[195], stage0_8[196], stage0_8[197], stage0_8[198], stage0_8[199]},
      {stage0_9[60]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[20],stage1_10[41],stage1_9[70],stage1_8[93]}
   );
   gpc615_5 gpc194 (
      {stage0_8[200], stage0_8[201], stage0_8[202], stage0_8[203], stage0_8[204]},
      {stage0_9[61]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[21],stage1_10[42],stage1_9[71],stage1_8[94]}
   );
   gpc615_5 gpc195 (
      {stage0_8[205], stage0_8[206], stage0_8[207], stage0_8[208], stage0_8[209]},
      {stage0_9[62]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[22],stage1_10[43],stage1_9[72],stage1_8[95]}
   );
   gpc615_5 gpc196 (
      {stage0_8[210], stage0_8[211], stage0_8[212], stage0_8[213], stage0_8[214]},
      {stage0_9[63]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[23],stage1_10[44],stage1_9[73],stage1_8[96]}
   );
   gpc615_5 gpc197 (
      {stage0_8[215], stage0_8[216], stage0_8[217], stage0_8[218], stage0_8[219]},
      {stage0_9[64]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[24],stage1_10[45],stage1_9[74],stage1_8[97]}
   );
   gpc615_5 gpc198 (
      {stage0_8[220], stage0_8[221], stage0_8[222], stage0_8[223], stage0_8[224]},
      {stage0_9[65]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[25],stage1_10[46],stage1_9[75],stage1_8[98]}
   );
   gpc615_5 gpc199 (
      {stage0_8[225], stage0_8[226], stage0_8[227], stage0_8[228], stage0_8[229]},
      {stage0_9[66]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[26],stage1_10[47],stage1_9[76],stage1_8[99]}
   );
   gpc615_5 gpc200 (
      {stage0_8[230], stage0_8[231], stage0_8[232], stage0_8[233], stage0_8[234]},
      {stage0_9[67]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[27],stage1_10[48],stage1_9[77],stage1_8[100]}
   );
   gpc615_5 gpc201 (
      {stage0_8[235], stage0_8[236], stage0_8[237], stage0_8[238], stage0_8[239]},
      {stage0_9[68]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[28],stage1_10[49],stage1_9[78],stage1_8[101]}
   );
   gpc615_5 gpc202 (
      {stage0_8[240], stage0_8[241], stage0_8[242], stage0_8[243], stage0_8[244]},
      {stage0_9[69]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[29],stage1_10[50],stage1_9[79],stage1_8[102]}
   );
   gpc615_5 gpc203 (
      {stage0_8[245], stage0_8[246], stage0_8[247], stage0_8[248], stage0_8[249]},
      {stage0_9[70]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[30],stage1_10[51],stage1_9[80],stage1_8[103]}
   );
   gpc615_5 gpc204 (
      {stage0_8[250], stage0_8[251], stage0_8[252], stage0_8[253], stage0_8[254]},
      {stage0_9[71]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[31],stage1_10[52],stage1_9[81],stage1_8[104]}
   );
   gpc606_5 gpc205 (
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[22],stage1_11[32],stage1_10[53],stage1_9[82]}
   );
   gpc606_5 gpc206 (
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[23],stage1_11[33],stage1_10[54],stage1_9[83]}
   );
   gpc606_5 gpc207 (
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[24],stage1_11[34],stage1_10[55],stage1_9[84]}
   );
   gpc606_5 gpc208 (
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[25],stage1_11[35],stage1_10[56],stage1_9[85]}
   );
   gpc606_5 gpc209 (
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[26],stage1_11[36],stage1_10[57],stage1_9[86]}
   );
   gpc606_5 gpc210 (
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[27],stage1_11[37],stage1_10[58],stage1_9[87]}
   );
   gpc606_5 gpc211 (
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[28],stage1_11[38],stage1_10[59],stage1_9[88]}
   );
   gpc606_5 gpc212 (
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[29],stage1_11[39],stage1_10[60],stage1_9[89]}
   );
   gpc606_5 gpc213 (
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[30],stage1_11[40],stage1_10[61],stage1_9[90]}
   );
   gpc606_5 gpc214 (
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[31],stage1_11[41],stage1_10[62],stage1_9[91]}
   );
   gpc606_5 gpc215 (
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[32],stage1_11[42],stage1_10[63],stage1_9[92]}
   );
   gpc606_5 gpc216 (
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[33],stage1_11[43],stage1_10[64],stage1_9[93]}
   );
   gpc606_5 gpc217 (
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[34],stage1_11[44],stage1_10[65],stage1_9[94]}
   );
   gpc606_5 gpc218 (
      {stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[35],stage1_11[45],stage1_10[66],stage1_9[95]}
   );
   gpc615_5 gpc219 (
      {stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160]},
      {stage0_10[132]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[36],stage1_11[46],stage1_10[67],stage1_9[96]}
   );
   gpc615_5 gpc220 (
      {stage0_9[161], stage0_9[162], stage0_9[163], stage0_9[164], stage0_9[165]},
      {stage0_10[133]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[37],stage1_11[47],stage1_10[68],stage1_9[97]}
   );
   gpc615_5 gpc221 (
      {stage0_9[166], stage0_9[167], stage0_9[168], stage0_9[169], stage0_9[170]},
      {stage0_10[134]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[38],stage1_11[48],stage1_10[69],stage1_9[98]}
   );
   gpc615_5 gpc222 (
      {stage0_9[171], stage0_9[172], stage0_9[173], stage0_9[174], stage0_9[175]},
      {stage0_10[135]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[39],stage1_11[49],stage1_10[70],stage1_9[99]}
   );
   gpc615_5 gpc223 (
      {stage0_9[176], stage0_9[177], stage0_9[178], stage0_9[179], stage0_9[180]},
      {stage0_10[136]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[40],stage1_11[50],stage1_10[71],stage1_9[100]}
   );
   gpc615_5 gpc224 (
      {stage0_9[181], stage0_9[182], stage0_9[183], stage0_9[184], stage0_9[185]},
      {stage0_10[137]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[41],stage1_11[51],stage1_10[72],stage1_9[101]}
   );
   gpc615_5 gpc225 (
      {stage0_9[186], stage0_9[187], stage0_9[188], stage0_9[189], stage0_9[190]},
      {stage0_10[138]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[42],stage1_11[52],stage1_10[73],stage1_9[102]}
   );
   gpc615_5 gpc226 (
      {stage0_9[191], stage0_9[192], stage0_9[193], stage0_9[194], stage0_9[195]},
      {stage0_10[139]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[43],stage1_11[53],stage1_10[74],stage1_9[103]}
   );
   gpc615_5 gpc227 (
      {stage0_9[196], stage0_9[197], stage0_9[198], stage0_9[199], stage0_9[200]},
      {stage0_10[140]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[44],stage1_11[54],stage1_10[75],stage1_9[104]}
   );
   gpc615_5 gpc228 (
      {stage0_9[201], stage0_9[202], stage0_9[203], stage0_9[204], stage0_9[205]},
      {stage0_10[141]},
      {stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage1_13[23],stage1_12[45],stage1_11[55],stage1_10[76],stage1_9[105]}
   );
   gpc615_5 gpc229 (
      {stage0_9[206], stage0_9[207], stage0_9[208], stage0_9[209], stage0_9[210]},
      {stage0_10[142]},
      {stage0_11[144], stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage1_13[24],stage1_12[46],stage1_11[56],stage1_10[77],stage1_9[106]}
   );
   gpc615_5 gpc230 (
      {stage0_9[211], stage0_9[212], stage0_9[213], stage0_9[214], stage0_9[215]},
      {stage0_10[143]},
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154], stage0_11[155]},
      {stage1_13[25],stage1_12[47],stage1_11[57],stage1_10[78],stage1_9[107]}
   );
   gpc615_5 gpc231 (
      {stage0_9[216], stage0_9[217], stage0_9[218], stage0_9[219], stage0_9[220]},
      {stage0_10[144]},
      {stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159], stage0_11[160], stage0_11[161]},
      {stage1_13[26],stage1_12[48],stage1_11[58],stage1_10[79],stage1_9[108]}
   );
   gpc615_5 gpc232 (
      {stage0_9[221], stage0_9[222], stage0_9[223], stage0_9[224], stage0_9[225]},
      {stage0_10[145]},
      {stage0_11[162], stage0_11[163], stage0_11[164], stage0_11[165], stage0_11[166], stage0_11[167]},
      {stage1_13[27],stage1_12[49],stage1_11[59],stage1_10[80],stage1_9[109]}
   );
   gpc615_5 gpc233 (
      {stage0_9[226], stage0_9[227], stage0_9[228], stage0_9[229], stage0_9[230]},
      {stage0_10[146]},
      {stage0_11[168], stage0_11[169], stage0_11[170], stage0_11[171], stage0_11[172], stage0_11[173]},
      {stage1_13[28],stage1_12[50],stage1_11[60],stage1_10[81],stage1_9[110]}
   );
   gpc615_5 gpc234 (
      {stage0_9[231], stage0_9[232], stage0_9[233], stage0_9[234], stage0_9[235]},
      {stage0_10[147]},
      {stage0_11[174], stage0_11[175], stage0_11[176], stage0_11[177], stage0_11[178], stage0_11[179]},
      {stage1_13[29],stage1_12[51],stage1_11[61],stage1_10[82],stage1_9[111]}
   );
   gpc615_5 gpc235 (
      {stage0_9[236], stage0_9[237], stage0_9[238], stage0_9[239], stage0_9[240]},
      {stage0_10[148]},
      {stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183], stage0_11[184], stage0_11[185]},
      {stage1_13[30],stage1_12[52],stage1_11[62],stage1_10[83],stage1_9[112]}
   );
   gpc615_5 gpc236 (
      {stage0_9[241], stage0_9[242], stage0_9[243], stage0_9[244], stage0_9[245]},
      {stage0_10[149]},
      {stage0_11[186], stage0_11[187], stage0_11[188], stage0_11[189], stage0_11[190], stage0_11[191]},
      {stage1_13[31],stage1_12[53],stage1_11[63],stage1_10[84],stage1_9[113]}
   );
   gpc615_5 gpc237 (
      {stage0_9[246], stage0_9[247], stage0_9[248], stage0_9[249], stage0_9[250]},
      {stage0_10[150]},
      {stage0_11[192], stage0_11[193], stage0_11[194], stage0_11[195], stage0_11[196], stage0_11[197]},
      {stage1_13[32],stage1_12[54],stage1_11[64],stage1_10[85],stage1_9[114]}
   );
   gpc615_5 gpc238 (
      {stage0_9[251], stage0_9[252], stage0_9[253], stage0_9[254], stage0_9[255]},
      {stage0_10[151]},
      {stage0_11[198], stage0_11[199], stage0_11[200], stage0_11[201], stage0_11[202], stage0_11[203]},
      {stage1_13[33],stage1_12[55],stage1_11[65],stage1_10[86],stage1_9[115]}
   );
   gpc606_5 gpc239 (
      {stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155], stage0_10[156], stage0_10[157]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[34],stage1_12[56],stage1_11[66],stage1_10[87]}
   );
   gpc606_5 gpc240 (
      {stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161], stage0_10[162], stage0_10[163]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[35],stage1_12[57],stage1_11[67],stage1_10[88]}
   );
   gpc606_5 gpc241 (
      {stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167], stage0_10[168], stage0_10[169]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[36],stage1_12[58],stage1_11[68],stage1_10[89]}
   );
   gpc606_5 gpc242 (
      {stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173], stage0_10[174], stage0_10[175]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[37],stage1_12[59],stage1_11[69],stage1_10[90]}
   );
   gpc606_5 gpc243 (
      {stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179], stage0_10[180], stage0_10[181]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[38],stage1_12[60],stage1_11[70],stage1_10[91]}
   );
   gpc606_5 gpc244 (
      {stage0_10[182], stage0_10[183], stage0_10[184], stage0_10[185], stage0_10[186], stage0_10[187]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[39],stage1_12[61],stage1_11[71],stage1_10[92]}
   );
   gpc606_5 gpc245 (
      {stage0_10[188], stage0_10[189], stage0_10[190], stage0_10[191], stage0_10[192], stage0_10[193]},
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage1_14[6],stage1_13[40],stage1_12[62],stage1_11[72],stage1_10[93]}
   );
   gpc606_5 gpc246 (
      {stage0_10[194], stage0_10[195], stage0_10[196], stage0_10[197], stage0_10[198], stage0_10[199]},
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage1_14[7],stage1_13[41],stage1_12[63],stage1_11[73],stage1_10[94]}
   );
   gpc606_5 gpc247 (
      {stage0_10[200], stage0_10[201], stage0_10[202], stage0_10[203], stage0_10[204], stage0_10[205]},
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage1_14[8],stage1_13[42],stage1_12[64],stage1_11[74],stage1_10[95]}
   );
   gpc606_5 gpc248 (
      {stage0_10[206], stage0_10[207], stage0_10[208], stage0_10[209], stage0_10[210], stage0_10[211]},
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage1_14[9],stage1_13[43],stage1_12[65],stage1_11[75],stage1_10[96]}
   );
   gpc606_5 gpc249 (
      {stage0_10[212], stage0_10[213], stage0_10[214], stage0_10[215], stage0_10[216], stage0_10[217]},
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage1_14[10],stage1_13[44],stage1_12[66],stage1_11[76],stage1_10[97]}
   );
   gpc606_5 gpc250 (
      {stage0_10[218], stage0_10[219], stage0_10[220], stage0_10[221], stage0_10[222], stage0_10[223]},
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage1_14[11],stage1_13[45],stage1_12[67],stage1_11[77],stage1_10[98]}
   );
   gpc606_5 gpc251 (
      {stage0_10[224], stage0_10[225], stage0_10[226], stage0_10[227], stage0_10[228], stage0_10[229]},
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage1_14[12],stage1_13[46],stage1_12[68],stage1_11[78],stage1_10[99]}
   );
   gpc615_5 gpc252 (
      {stage0_10[230], stage0_10[231], stage0_10[232], stage0_10[233], stage0_10[234]},
      {stage0_11[204]},
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage1_14[13],stage1_13[47],stage1_12[69],stage1_11[79],stage1_10[100]}
   );
   gpc615_5 gpc253 (
      {stage0_10[235], stage0_10[236], stage0_10[237], stage0_10[238], stage0_10[239]},
      {stage0_11[205]},
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89]},
      {stage1_14[14],stage1_13[48],stage1_12[70],stage1_11[80],stage1_10[101]}
   );
   gpc615_5 gpc254 (
      {stage0_10[240], stage0_10[241], stage0_10[242], stage0_10[243], stage0_10[244]},
      {stage0_11[206]},
      {stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95]},
      {stage1_14[15],stage1_13[49],stage1_12[71],stage1_11[81],stage1_10[102]}
   );
   gpc615_5 gpc255 (
      {stage0_11[207], stage0_11[208], stage0_11[209], stage0_11[210], stage0_11[211]},
      {stage0_12[96]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[16],stage1_13[50],stage1_12[72],stage1_11[82]}
   );
   gpc615_5 gpc256 (
      {stage0_11[212], stage0_11[213], stage0_11[214], stage0_11[215], stage0_11[216]},
      {stage0_12[97]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[17],stage1_13[51],stage1_12[73],stage1_11[83]}
   );
   gpc615_5 gpc257 (
      {stage0_11[217], stage0_11[218], stage0_11[219], stage0_11[220], stage0_11[221]},
      {stage0_12[98]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[18],stage1_13[52],stage1_12[74],stage1_11[84]}
   );
   gpc615_5 gpc258 (
      {stage0_11[222], stage0_11[223], stage0_11[224], stage0_11[225], stage0_11[226]},
      {stage0_12[99]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[19],stage1_13[53],stage1_12[75],stage1_11[85]}
   );
   gpc606_5 gpc259 (
      {stage0_12[100], stage0_12[101], stage0_12[102], stage0_12[103], stage0_12[104], stage0_12[105]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[4],stage1_14[20],stage1_13[54],stage1_12[76]}
   );
   gpc606_5 gpc260 (
      {stage0_12[106], stage0_12[107], stage0_12[108], stage0_12[109], stage0_12[110], stage0_12[111]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[5],stage1_14[21],stage1_13[55],stage1_12[77]}
   );
   gpc606_5 gpc261 (
      {stage0_12[112], stage0_12[113], stage0_12[114], stage0_12[115], stage0_12[116], stage0_12[117]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[6],stage1_14[22],stage1_13[56],stage1_12[78]}
   );
   gpc606_5 gpc262 (
      {stage0_12[118], stage0_12[119], stage0_12[120], stage0_12[121], stage0_12[122], stage0_12[123]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[7],stage1_14[23],stage1_13[57],stage1_12[79]}
   );
   gpc606_5 gpc263 (
      {stage0_12[124], stage0_12[125], stage0_12[126], stage0_12[127], stage0_12[128], stage0_12[129]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[8],stage1_14[24],stage1_13[58],stage1_12[80]}
   );
   gpc606_5 gpc264 (
      {stage0_12[130], stage0_12[131], stage0_12[132], stage0_12[133], stage0_12[134], stage0_12[135]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[9],stage1_14[25],stage1_13[59],stage1_12[81]}
   );
   gpc606_5 gpc265 (
      {stage0_12[136], stage0_12[137], stage0_12[138], stage0_12[139], stage0_12[140], stage0_12[141]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[10],stage1_14[26],stage1_13[60],stage1_12[82]}
   );
   gpc606_5 gpc266 (
      {stage0_12[142], stage0_12[143], stage0_12[144], stage0_12[145], stage0_12[146], stage0_12[147]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[11],stage1_14[27],stage1_13[61],stage1_12[83]}
   );
   gpc606_5 gpc267 (
      {stage0_12[148], stage0_12[149], stage0_12[150], stage0_12[151], stage0_12[152], stage0_12[153]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[12],stage1_14[28],stage1_13[62],stage1_12[84]}
   );
   gpc606_5 gpc268 (
      {stage0_12[154], stage0_12[155], stage0_12[156], stage0_12[157], stage0_12[158], stage0_12[159]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[13],stage1_14[29],stage1_13[63],stage1_12[85]}
   );
   gpc606_5 gpc269 (
      {stage0_12[160], stage0_12[161], stage0_12[162], stage0_12[163], stage0_12[164], stage0_12[165]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[14],stage1_14[30],stage1_13[64],stage1_12[86]}
   );
   gpc606_5 gpc270 (
      {stage0_12[166], stage0_12[167], stage0_12[168], stage0_12[169], stage0_12[170], stage0_12[171]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[15],stage1_14[31],stage1_13[65],stage1_12[87]}
   );
   gpc606_5 gpc271 (
      {stage0_12[172], stage0_12[173], stage0_12[174], stage0_12[175], stage0_12[176], stage0_12[177]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[16],stage1_14[32],stage1_13[66],stage1_12[88]}
   );
   gpc606_5 gpc272 (
      {stage0_12[178], stage0_12[179], stage0_12[180], stage0_12[181], stage0_12[182], stage0_12[183]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[17],stage1_14[33],stage1_13[67],stage1_12[89]}
   );
   gpc606_5 gpc273 (
      {stage0_12[184], stage0_12[185], stage0_12[186], stage0_12[187], stage0_12[188], stage0_12[189]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[18],stage1_14[34],stage1_13[68],stage1_12[90]}
   );
   gpc606_5 gpc274 (
      {stage0_12[190], stage0_12[191], stage0_12[192], stage0_12[193], stage0_12[194], stage0_12[195]},
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage1_16[15],stage1_15[19],stage1_14[35],stage1_13[69],stage1_12[91]}
   );
   gpc606_5 gpc275 (
      {stage0_12[196], stage0_12[197], stage0_12[198], stage0_12[199], stage0_12[200], stage0_12[201]},
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage1_16[16],stage1_15[20],stage1_14[36],stage1_13[70],stage1_12[92]}
   );
   gpc606_5 gpc276 (
      {stage0_12[202], stage0_12[203], stage0_12[204], stage0_12[205], stage0_12[206], stage0_12[207]},
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage1_16[17],stage1_15[21],stage1_14[37],stage1_13[71],stage1_12[93]}
   );
   gpc606_5 gpc277 (
      {stage0_12[208], stage0_12[209], stage0_12[210], stage0_12[211], stage0_12[212], stage0_12[213]},
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113]},
      {stage1_16[18],stage1_15[22],stage1_14[38],stage1_13[72],stage1_12[94]}
   );
   gpc606_5 gpc278 (
      {stage0_12[214], stage0_12[215], stage0_12[216], stage0_12[217], stage0_12[218], stage0_12[219]},
      {stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119]},
      {stage1_16[19],stage1_15[23],stage1_14[39],stage1_13[73],stage1_12[95]}
   );
   gpc606_5 gpc279 (
      {stage0_12[220], stage0_12[221], stage0_12[222], stage0_12[223], stage0_12[224], stage0_12[225]},
      {stage0_14[120], stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125]},
      {stage1_16[20],stage1_15[24],stage1_14[40],stage1_13[74],stage1_12[96]}
   );
   gpc606_5 gpc280 (
      {stage0_12[226], stage0_12[227], stage0_12[228], stage0_12[229], stage0_12[230], stage0_12[231]},
      {stage0_14[126], stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131]},
      {stage1_16[21],stage1_15[25],stage1_14[41],stage1_13[75],stage1_12[97]}
   );
   gpc606_5 gpc281 (
      {stage0_12[232], stage0_12[233], stage0_12[234], stage0_12[235], stage0_12[236], stage0_12[237]},
      {stage0_14[132], stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137]},
      {stage1_16[22],stage1_15[26],stage1_14[42],stage1_13[76],stage1_12[98]}
   );
   gpc606_5 gpc282 (
      {stage0_12[238], stage0_12[239], stage0_12[240], stage0_12[241], stage0_12[242], stage0_12[243]},
      {stage0_14[138], stage0_14[139], stage0_14[140], stage0_14[141], stage0_14[142], stage0_14[143]},
      {stage1_16[23],stage1_15[27],stage1_14[43],stage1_13[77],stage1_12[99]}
   );
   gpc606_5 gpc283 (
      {stage0_12[244], stage0_12[245], stage0_12[246], stage0_12[247], stage0_12[248], stage0_12[249]},
      {stage0_14[144], stage0_14[145], stage0_14[146], stage0_14[147], stage0_14[148], stage0_14[149]},
      {stage1_16[24],stage1_15[28],stage1_14[44],stage1_13[78],stage1_12[100]}
   );
   gpc606_5 gpc284 (
      {stage0_12[250], stage0_12[251], stage0_12[252], stage0_12[253], stage0_12[254], stage0_12[255]},
      {stage0_14[150], stage0_14[151], stage0_14[152], stage0_14[153], stage0_14[154], stage0_14[155]},
      {stage1_16[25],stage1_15[29],stage1_14[45],stage1_13[79],stage1_12[101]}
   );
   gpc606_5 gpc285 (
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[26],stage1_15[30],stage1_14[46],stage1_13[80]}
   );
   gpc606_5 gpc286 (
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[27],stage1_15[31],stage1_14[47],stage1_13[81]}
   );
   gpc606_5 gpc287 (
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[28],stage1_15[32],stage1_14[48],stage1_13[82]}
   );
   gpc606_5 gpc288 (
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[29],stage1_15[33],stage1_14[49],stage1_13[83]}
   );
   gpc606_5 gpc289 (
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[30],stage1_15[34],stage1_14[50],stage1_13[84]}
   );
   gpc606_5 gpc290 (
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[31],stage1_15[35],stage1_14[51],stage1_13[85]}
   );
   gpc606_5 gpc291 (
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[32],stage1_15[36],stage1_14[52],stage1_13[86]}
   );
   gpc606_5 gpc292 (
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[33],stage1_15[37],stage1_14[53],stage1_13[87]}
   );
   gpc606_5 gpc293 (
      {stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[34],stage1_15[38],stage1_14[54],stage1_13[88]}
   );
   gpc606_5 gpc294 (
      {stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[35],stage1_15[39],stage1_14[55],stage1_13[89]}
   );
   gpc606_5 gpc295 (
      {stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87], stage0_13[88], stage0_13[89]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[36],stage1_15[40],stage1_14[56],stage1_13[90]}
   );
   gpc615_5 gpc296 (
      {stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93], stage0_13[94]},
      {stage0_14[156]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[37],stage1_15[41],stage1_14[57],stage1_13[91]}
   );
   gpc615_5 gpc297 (
      {stage0_13[95], stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99]},
      {stage0_14[157]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[38],stage1_15[42],stage1_14[58],stage1_13[92]}
   );
   gpc615_5 gpc298 (
      {stage0_13[100], stage0_13[101], stage0_13[102], stage0_13[103], stage0_13[104]},
      {stage0_14[158]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[39],stage1_15[43],stage1_14[59],stage1_13[93]}
   );
   gpc615_5 gpc299 (
      {stage0_13[105], stage0_13[106], stage0_13[107], stage0_13[108], stage0_13[109]},
      {stage0_14[159]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[40],stage1_15[44],stage1_14[60],stage1_13[94]}
   );
   gpc615_5 gpc300 (
      {stage0_13[110], stage0_13[111], stage0_13[112], stage0_13[113], stage0_13[114]},
      {stage0_14[160]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[41],stage1_15[45],stage1_14[61],stage1_13[95]}
   );
   gpc615_5 gpc301 (
      {stage0_13[115], stage0_13[116], stage0_13[117], stage0_13[118], stage0_13[119]},
      {stage0_14[161]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[42],stage1_15[46],stage1_14[62],stage1_13[96]}
   );
   gpc615_5 gpc302 (
      {stage0_13[120], stage0_13[121], stage0_13[122], stage0_13[123], stage0_13[124]},
      {stage0_14[162]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[43],stage1_15[47],stage1_14[63],stage1_13[97]}
   );
   gpc615_5 gpc303 (
      {stage0_13[125], stage0_13[126], stage0_13[127], stage0_13[128], stage0_13[129]},
      {stage0_14[163]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[44],stage1_15[48],stage1_14[64],stage1_13[98]}
   );
   gpc615_5 gpc304 (
      {stage0_13[130], stage0_13[131], stage0_13[132], stage0_13[133], stage0_13[134]},
      {stage0_14[164]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[45],stage1_15[49],stage1_14[65],stage1_13[99]}
   );
   gpc615_5 gpc305 (
      {stage0_13[135], stage0_13[136], stage0_13[137], stage0_13[138], stage0_13[139]},
      {stage0_14[165]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[46],stage1_15[50],stage1_14[66],stage1_13[100]}
   );
   gpc615_5 gpc306 (
      {stage0_13[140], stage0_13[141], stage0_13[142], stage0_13[143], stage0_13[144]},
      {stage0_14[166]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[47],stage1_15[51],stage1_14[67],stage1_13[101]}
   );
   gpc615_5 gpc307 (
      {stage0_13[145], stage0_13[146], stage0_13[147], stage0_13[148], stage0_13[149]},
      {stage0_14[167]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[48],stage1_15[52],stage1_14[68],stage1_13[102]}
   );
   gpc615_5 gpc308 (
      {stage0_13[150], stage0_13[151], stage0_13[152], stage0_13[153], stage0_13[154]},
      {stage0_14[168]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[49],stage1_15[53],stage1_14[69],stage1_13[103]}
   );
   gpc615_5 gpc309 (
      {stage0_13[155], stage0_13[156], stage0_13[157], stage0_13[158], stage0_13[159]},
      {stage0_14[169]},
      {stage0_15[144], stage0_15[145], stage0_15[146], stage0_15[147], stage0_15[148], stage0_15[149]},
      {stage1_17[24],stage1_16[50],stage1_15[54],stage1_14[70],stage1_13[104]}
   );
   gpc615_5 gpc310 (
      {stage0_13[160], stage0_13[161], stage0_13[162], stage0_13[163], stage0_13[164]},
      {stage0_14[170]},
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155]},
      {stage1_17[25],stage1_16[51],stage1_15[55],stage1_14[71],stage1_13[105]}
   );
   gpc615_5 gpc311 (
      {stage0_13[165], stage0_13[166], stage0_13[167], stage0_13[168], stage0_13[169]},
      {stage0_14[171]},
      {stage0_15[156], stage0_15[157], stage0_15[158], stage0_15[159], stage0_15[160], stage0_15[161]},
      {stage1_17[26],stage1_16[52],stage1_15[56],stage1_14[72],stage1_13[106]}
   );
   gpc615_5 gpc312 (
      {stage0_13[170], stage0_13[171], stage0_13[172], stage0_13[173], stage0_13[174]},
      {stage0_14[172]},
      {stage0_15[162], stage0_15[163], stage0_15[164], stage0_15[165], stage0_15[166], stage0_15[167]},
      {stage1_17[27],stage1_16[53],stage1_15[57],stage1_14[73],stage1_13[107]}
   );
   gpc615_5 gpc313 (
      {stage0_13[175], stage0_13[176], stage0_13[177], stage0_13[178], stage0_13[179]},
      {stage0_14[173]},
      {stage0_15[168], stage0_15[169], stage0_15[170], stage0_15[171], stage0_15[172], stage0_15[173]},
      {stage1_17[28],stage1_16[54],stage1_15[58],stage1_14[74],stage1_13[108]}
   );
   gpc615_5 gpc314 (
      {stage0_13[180], stage0_13[181], stage0_13[182], stage0_13[183], stage0_13[184]},
      {stage0_14[174]},
      {stage0_15[174], stage0_15[175], stage0_15[176], stage0_15[177], stage0_15[178], stage0_15[179]},
      {stage1_17[29],stage1_16[55],stage1_15[59],stage1_14[75],stage1_13[109]}
   );
   gpc615_5 gpc315 (
      {stage0_13[185], stage0_13[186], stage0_13[187], stage0_13[188], stage0_13[189]},
      {stage0_14[175]},
      {stage0_15[180], stage0_15[181], stage0_15[182], stage0_15[183], stage0_15[184], stage0_15[185]},
      {stage1_17[30],stage1_16[56],stage1_15[60],stage1_14[76],stage1_13[110]}
   );
   gpc615_5 gpc316 (
      {stage0_13[190], stage0_13[191], stage0_13[192], stage0_13[193], stage0_13[194]},
      {stage0_14[176]},
      {stage0_15[186], stage0_15[187], stage0_15[188], stage0_15[189], stage0_15[190], stage0_15[191]},
      {stage1_17[31],stage1_16[57],stage1_15[61],stage1_14[77],stage1_13[111]}
   );
   gpc615_5 gpc317 (
      {stage0_13[195], stage0_13[196], stage0_13[197], stage0_13[198], stage0_13[199]},
      {stage0_14[177]},
      {stage0_15[192], stage0_15[193], stage0_15[194], stage0_15[195], stage0_15[196], stage0_15[197]},
      {stage1_17[32],stage1_16[58],stage1_15[62],stage1_14[78],stage1_13[112]}
   );
   gpc615_5 gpc318 (
      {stage0_13[200], stage0_13[201], stage0_13[202], stage0_13[203], stage0_13[204]},
      {stage0_14[178]},
      {stage0_15[198], stage0_15[199], stage0_15[200], stage0_15[201], stage0_15[202], stage0_15[203]},
      {stage1_17[33],stage1_16[59],stage1_15[63],stage1_14[79],stage1_13[113]}
   );
   gpc615_5 gpc319 (
      {stage0_13[205], stage0_13[206], stage0_13[207], stage0_13[208], stage0_13[209]},
      {stage0_14[179]},
      {stage0_15[204], stage0_15[205], stage0_15[206], stage0_15[207], stage0_15[208], stage0_15[209]},
      {stage1_17[34],stage1_16[60],stage1_15[64],stage1_14[80],stage1_13[114]}
   );
   gpc615_5 gpc320 (
      {stage0_13[210], stage0_13[211], stage0_13[212], stage0_13[213], stage0_13[214]},
      {stage0_14[180]},
      {stage0_15[210], stage0_15[211], stage0_15[212], stage0_15[213], stage0_15[214], stage0_15[215]},
      {stage1_17[35],stage1_16[61],stage1_15[65],stage1_14[81],stage1_13[115]}
   );
   gpc615_5 gpc321 (
      {stage0_13[215], stage0_13[216], stage0_13[217], stage0_13[218], stage0_13[219]},
      {stage0_14[181]},
      {stage0_15[216], stage0_15[217], stage0_15[218], stage0_15[219], stage0_15[220], stage0_15[221]},
      {stage1_17[36],stage1_16[62],stage1_15[66],stage1_14[82],stage1_13[116]}
   );
   gpc615_5 gpc322 (
      {stage0_13[220], stage0_13[221], stage0_13[222], stage0_13[223], stage0_13[224]},
      {stage0_14[182]},
      {stage0_15[222], stage0_15[223], stage0_15[224], stage0_15[225], stage0_15[226], stage0_15[227]},
      {stage1_17[37],stage1_16[63],stage1_15[67],stage1_14[83],stage1_13[117]}
   );
   gpc615_5 gpc323 (
      {stage0_13[225], stage0_13[226], stage0_13[227], stage0_13[228], stage0_13[229]},
      {stage0_14[183]},
      {stage0_15[228], stage0_15[229], stage0_15[230], stage0_15[231], stage0_15[232], stage0_15[233]},
      {stage1_17[38],stage1_16[64],stage1_15[68],stage1_14[84],stage1_13[118]}
   );
   gpc615_5 gpc324 (
      {stage0_13[230], stage0_13[231], stage0_13[232], stage0_13[233], stage0_13[234]},
      {stage0_14[184]},
      {stage0_15[234], stage0_15[235], stage0_15[236], stage0_15[237], stage0_15[238], stage0_15[239]},
      {stage1_17[39],stage1_16[65],stage1_15[69],stage1_14[85],stage1_13[119]}
   );
   gpc615_5 gpc325 (
      {stage0_13[235], stage0_13[236], stage0_13[237], stage0_13[238], stage0_13[239]},
      {stage0_14[185]},
      {stage0_15[240], stage0_15[241], stage0_15[242], stage0_15[243], stage0_15[244], stage0_15[245]},
      {stage1_17[40],stage1_16[66],stage1_15[70],stage1_14[86],stage1_13[120]}
   );
   gpc615_5 gpc326 (
      {stage0_13[240], stage0_13[241], stage0_13[242], stage0_13[243], stage0_13[244]},
      {stage0_14[186]},
      {stage0_15[246], stage0_15[247], stage0_15[248], stage0_15[249], stage0_15[250], stage0_15[251]},
      {stage1_17[41],stage1_16[67],stage1_15[71],stage1_14[87],stage1_13[121]}
   );
   gpc1_1 gpc327 (
      {stage0_1[228]},
      {stage1_1[70]}
   );
   gpc1_1 gpc328 (
      {stage0_1[229]},
      {stage1_1[71]}
   );
   gpc1_1 gpc329 (
      {stage0_1[230]},
      {stage1_1[72]}
   );
   gpc1_1 gpc330 (
      {stage0_1[231]},
      {stage1_1[73]}
   );
   gpc1_1 gpc331 (
      {stage0_1[232]},
      {stage1_1[74]}
   );
   gpc1_1 gpc332 (
      {stage0_1[233]},
      {stage1_1[75]}
   );
   gpc1_1 gpc333 (
      {stage0_1[234]},
      {stage1_1[76]}
   );
   gpc1_1 gpc334 (
      {stage0_1[235]},
      {stage1_1[77]}
   );
   gpc1_1 gpc335 (
      {stage0_1[236]},
      {stage1_1[78]}
   );
   gpc1_1 gpc336 (
      {stage0_1[237]},
      {stage1_1[79]}
   );
   gpc1_1 gpc337 (
      {stage0_1[238]},
      {stage1_1[80]}
   );
   gpc1_1 gpc338 (
      {stage0_1[239]},
      {stage1_1[81]}
   );
   gpc1_1 gpc339 (
      {stage0_1[240]},
      {stage1_1[82]}
   );
   gpc1_1 gpc340 (
      {stage0_1[241]},
      {stage1_1[83]}
   );
   gpc1_1 gpc341 (
      {stage0_1[242]},
      {stage1_1[84]}
   );
   gpc1_1 gpc342 (
      {stage0_1[243]},
      {stage1_1[85]}
   );
   gpc1_1 gpc343 (
      {stage0_1[244]},
      {stage1_1[86]}
   );
   gpc1_1 gpc344 (
      {stage0_1[245]},
      {stage1_1[87]}
   );
   gpc1_1 gpc345 (
      {stage0_1[246]},
      {stage1_1[88]}
   );
   gpc1_1 gpc346 (
      {stage0_1[247]},
      {stage1_1[89]}
   );
   gpc1_1 gpc347 (
      {stage0_1[248]},
      {stage1_1[90]}
   );
   gpc1_1 gpc348 (
      {stage0_1[249]},
      {stage1_1[91]}
   );
   gpc1_1 gpc349 (
      {stage0_1[250]},
      {stage1_1[92]}
   );
   gpc1_1 gpc350 (
      {stage0_1[251]},
      {stage1_1[93]}
   );
   gpc1_1 gpc351 (
      {stage0_1[252]},
      {stage1_1[94]}
   );
   gpc1_1 gpc352 (
      {stage0_1[253]},
      {stage1_1[95]}
   );
   gpc1_1 gpc353 (
      {stage0_1[254]},
      {stage1_1[96]}
   );
   gpc1_1 gpc354 (
      {stage0_1[255]},
      {stage1_1[97]}
   );
   gpc1_1 gpc355 (
      {stage0_2[246]},
      {stage1_2[88]}
   );
   gpc1_1 gpc356 (
      {stage0_2[247]},
      {stage1_2[89]}
   );
   gpc1_1 gpc357 (
      {stage0_2[248]},
      {stage1_2[90]}
   );
   gpc1_1 gpc358 (
      {stage0_2[249]},
      {stage1_2[91]}
   );
   gpc1_1 gpc359 (
      {stage0_2[250]},
      {stage1_2[92]}
   );
   gpc1_1 gpc360 (
      {stage0_2[251]},
      {stage1_2[93]}
   );
   gpc1_1 gpc361 (
      {stage0_2[252]},
      {stage1_2[94]}
   );
   gpc1_1 gpc362 (
      {stage0_2[253]},
      {stage1_2[95]}
   );
   gpc1_1 gpc363 (
      {stage0_2[254]},
      {stage1_2[96]}
   );
   gpc1_1 gpc364 (
      {stage0_2[255]},
      {stage1_2[97]}
   );
   gpc1_1 gpc365 (
      {stage0_3[242]},
      {stage1_3[100]}
   );
   gpc1_1 gpc366 (
      {stage0_3[243]},
      {stage1_3[101]}
   );
   gpc1_1 gpc367 (
      {stage0_3[244]},
      {stage1_3[102]}
   );
   gpc1_1 gpc368 (
      {stage0_3[245]},
      {stage1_3[103]}
   );
   gpc1_1 gpc369 (
      {stage0_3[246]},
      {stage1_3[104]}
   );
   gpc1_1 gpc370 (
      {stage0_3[247]},
      {stage1_3[105]}
   );
   gpc1_1 gpc371 (
      {stage0_3[248]},
      {stage1_3[106]}
   );
   gpc1_1 gpc372 (
      {stage0_3[249]},
      {stage1_3[107]}
   );
   gpc1_1 gpc373 (
      {stage0_3[250]},
      {stage1_3[108]}
   );
   gpc1_1 gpc374 (
      {stage0_3[251]},
      {stage1_3[109]}
   );
   gpc1_1 gpc375 (
      {stage0_3[252]},
      {stage1_3[110]}
   );
   gpc1_1 gpc376 (
      {stage0_3[253]},
      {stage1_3[111]}
   );
   gpc1_1 gpc377 (
      {stage0_3[254]},
      {stage1_3[112]}
   );
   gpc1_1 gpc378 (
      {stage0_3[255]},
      {stage1_3[113]}
   );
   gpc1_1 gpc379 (
      {stage0_4[249]},
      {stage1_4[120]}
   );
   gpc1_1 gpc380 (
      {stage0_4[250]},
      {stage1_4[121]}
   );
   gpc1_1 gpc381 (
      {stage0_4[251]},
      {stage1_4[122]}
   );
   gpc1_1 gpc382 (
      {stage0_4[252]},
      {stage1_4[123]}
   );
   gpc1_1 gpc383 (
      {stage0_4[253]},
      {stage1_4[124]}
   );
   gpc1_1 gpc384 (
      {stage0_4[254]},
      {stage1_4[125]}
   );
   gpc1_1 gpc385 (
      {stage0_4[255]},
      {stage1_4[126]}
   );
   gpc1_1 gpc386 (
      {stage0_5[254]},
      {stage1_5[103]}
   );
   gpc1_1 gpc387 (
      {stage0_5[255]},
      {stage1_5[104]}
   );
   gpc1_1 gpc388 (
      {stage0_6[255]},
      {stage1_6[103]}
   );
   gpc1_1 gpc389 (
      {stage0_7[236]},
      {stage1_7[95]}
   );
   gpc1_1 gpc390 (
      {stage0_7[237]},
      {stage1_7[96]}
   );
   gpc1_1 gpc391 (
      {stage0_7[238]},
      {stage1_7[97]}
   );
   gpc1_1 gpc392 (
      {stage0_7[239]},
      {stage1_7[98]}
   );
   gpc1_1 gpc393 (
      {stage0_7[240]},
      {stage1_7[99]}
   );
   gpc1_1 gpc394 (
      {stage0_7[241]},
      {stage1_7[100]}
   );
   gpc1_1 gpc395 (
      {stage0_7[242]},
      {stage1_7[101]}
   );
   gpc1_1 gpc396 (
      {stage0_7[243]},
      {stage1_7[102]}
   );
   gpc1_1 gpc397 (
      {stage0_7[244]},
      {stage1_7[103]}
   );
   gpc1_1 gpc398 (
      {stage0_7[245]},
      {stage1_7[104]}
   );
   gpc1_1 gpc399 (
      {stage0_7[246]},
      {stage1_7[105]}
   );
   gpc1_1 gpc400 (
      {stage0_7[247]},
      {stage1_7[106]}
   );
   gpc1_1 gpc401 (
      {stage0_7[248]},
      {stage1_7[107]}
   );
   gpc1_1 gpc402 (
      {stage0_7[249]},
      {stage1_7[108]}
   );
   gpc1_1 gpc403 (
      {stage0_7[250]},
      {stage1_7[109]}
   );
   gpc1_1 gpc404 (
      {stage0_7[251]},
      {stage1_7[110]}
   );
   gpc1_1 gpc405 (
      {stage0_7[252]},
      {stage1_7[111]}
   );
   gpc1_1 gpc406 (
      {stage0_7[253]},
      {stage1_7[112]}
   );
   gpc1_1 gpc407 (
      {stage0_7[254]},
      {stage1_7[113]}
   );
   gpc1_1 gpc408 (
      {stage0_7[255]},
      {stage1_7[114]}
   );
   gpc1_1 gpc409 (
      {stage0_8[255]},
      {stage1_8[105]}
   );
   gpc1_1 gpc410 (
      {stage0_10[245]},
      {stage1_10[103]}
   );
   gpc1_1 gpc411 (
      {stage0_10[246]},
      {stage1_10[104]}
   );
   gpc1_1 gpc412 (
      {stage0_10[247]},
      {stage1_10[105]}
   );
   gpc1_1 gpc413 (
      {stage0_10[248]},
      {stage1_10[106]}
   );
   gpc1_1 gpc414 (
      {stage0_10[249]},
      {stage1_10[107]}
   );
   gpc1_1 gpc415 (
      {stage0_10[250]},
      {stage1_10[108]}
   );
   gpc1_1 gpc416 (
      {stage0_10[251]},
      {stage1_10[109]}
   );
   gpc1_1 gpc417 (
      {stage0_10[252]},
      {stage1_10[110]}
   );
   gpc1_1 gpc418 (
      {stage0_10[253]},
      {stage1_10[111]}
   );
   gpc1_1 gpc419 (
      {stage0_10[254]},
      {stage1_10[112]}
   );
   gpc1_1 gpc420 (
      {stage0_10[255]},
      {stage1_10[113]}
   );
   gpc1_1 gpc421 (
      {stage0_11[227]},
      {stage1_11[86]}
   );
   gpc1_1 gpc422 (
      {stage0_11[228]},
      {stage1_11[87]}
   );
   gpc1_1 gpc423 (
      {stage0_11[229]},
      {stage1_11[88]}
   );
   gpc1_1 gpc424 (
      {stage0_11[230]},
      {stage1_11[89]}
   );
   gpc1_1 gpc425 (
      {stage0_11[231]},
      {stage1_11[90]}
   );
   gpc1_1 gpc426 (
      {stage0_11[232]},
      {stage1_11[91]}
   );
   gpc1_1 gpc427 (
      {stage0_11[233]},
      {stage1_11[92]}
   );
   gpc1_1 gpc428 (
      {stage0_11[234]},
      {stage1_11[93]}
   );
   gpc1_1 gpc429 (
      {stage0_11[235]},
      {stage1_11[94]}
   );
   gpc1_1 gpc430 (
      {stage0_11[236]},
      {stage1_11[95]}
   );
   gpc1_1 gpc431 (
      {stage0_11[237]},
      {stage1_11[96]}
   );
   gpc1_1 gpc432 (
      {stage0_11[238]},
      {stage1_11[97]}
   );
   gpc1_1 gpc433 (
      {stage0_11[239]},
      {stage1_11[98]}
   );
   gpc1_1 gpc434 (
      {stage0_11[240]},
      {stage1_11[99]}
   );
   gpc1_1 gpc435 (
      {stage0_11[241]},
      {stage1_11[100]}
   );
   gpc1_1 gpc436 (
      {stage0_11[242]},
      {stage1_11[101]}
   );
   gpc1_1 gpc437 (
      {stage0_11[243]},
      {stage1_11[102]}
   );
   gpc1_1 gpc438 (
      {stage0_11[244]},
      {stage1_11[103]}
   );
   gpc1_1 gpc439 (
      {stage0_11[245]},
      {stage1_11[104]}
   );
   gpc1_1 gpc440 (
      {stage0_11[246]},
      {stage1_11[105]}
   );
   gpc1_1 gpc441 (
      {stage0_11[247]},
      {stage1_11[106]}
   );
   gpc1_1 gpc442 (
      {stage0_11[248]},
      {stage1_11[107]}
   );
   gpc1_1 gpc443 (
      {stage0_11[249]},
      {stage1_11[108]}
   );
   gpc1_1 gpc444 (
      {stage0_11[250]},
      {stage1_11[109]}
   );
   gpc1_1 gpc445 (
      {stage0_11[251]},
      {stage1_11[110]}
   );
   gpc1_1 gpc446 (
      {stage0_11[252]},
      {stage1_11[111]}
   );
   gpc1_1 gpc447 (
      {stage0_11[253]},
      {stage1_11[112]}
   );
   gpc1_1 gpc448 (
      {stage0_11[254]},
      {stage1_11[113]}
   );
   gpc1_1 gpc449 (
      {stage0_11[255]},
      {stage1_11[114]}
   );
   gpc1_1 gpc450 (
      {stage0_13[245]},
      {stage1_13[122]}
   );
   gpc1_1 gpc451 (
      {stage0_13[246]},
      {stage1_13[123]}
   );
   gpc1_1 gpc452 (
      {stage0_13[247]},
      {stage1_13[124]}
   );
   gpc1_1 gpc453 (
      {stage0_13[248]},
      {stage1_13[125]}
   );
   gpc1_1 gpc454 (
      {stage0_13[249]},
      {stage1_13[126]}
   );
   gpc1_1 gpc455 (
      {stage0_13[250]},
      {stage1_13[127]}
   );
   gpc1_1 gpc456 (
      {stage0_13[251]},
      {stage1_13[128]}
   );
   gpc1_1 gpc457 (
      {stage0_13[252]},
      {stage1_13[129]}
   );
   gpc1_1 gpc458 (
      {stage0_13[253]},
      {stage1_13[130]}
   );
   gpc1_1 gpc459 (
      {stage0_13[254]},
      {stage1_13[131]}
   );
   gpc1_1 gpc460 (
      {stage0_13[255]},
      {stage1_13[132]}
   );
   gpc1_1 gpc461 (
      {stage0_14[187]},
      {stage1_14[88]}
   );
   gpc1_1 gpc462 (
      {stage0_14[188]},
      {stage1_14[89]}
   );
   gpc1_1 gpc463 (
      {stage0_14[189]},
      {stage1_14[90]}
   );
   gpc1_1 gpc464 (
      {stage0_14[190]},
      {stage1_14[91]}
   );
   gpc1_1 gpc465 (
      {stage0_14[191]},
      {stage1_14[92]}
   );
   gpc1_1 gpc466 (
      {stage0_14[192]},
      {stage1_14[93]}
   );
   gpc1_1 gpc467 (
      {stage0_14[193]},
      {stage1_14[94]}
   );
   gpc1_1 gpc468 (
      {stage0_14[194]},
      {stage1_14[95]}
   );
   gpc1_1 gpc469 (
      {stage0_14[195]},
      {stage1_14[96]}
   );
   gpc1_1 gpc470 (
      {stage0_14[196]},
      {stage1_14[97]}
   );
   gpc1_1 gpc471 (
      {stage0_14[197]},
      {stage1_14[98]}
   );
   gpc1_1 gpc472 (
      {stage0_14[198]},
      {stage1_14[99]}
   );
   gpc1_1 gpc473 (
      {stage0_14[199]},
      {stage1_14[100]}
   );
   gpc1_1 gpc474 (
      {stage0_14[200]},
      {stage1_14[101]}
   );
   gpc1_1 gpc475 (
      {stage0_14[201]},
      {stage1_14[102]}
   );
   gpc1_1 gpc476 (
      {stage0_14[202]},
      {stage1_14[103]}
   );
   gpc1_1 gpc477 (
      {stage0_14[203]},
      {stage1_14[104]}
   );
   gpc1_1 gpc478 (
      {stage0_14[204]},
      {stage1_14[105]}
   );
   gpc1_1 gpc479 (
      {stage0_14[205]},
      {stage1_14[106]}
   );
   gpc1_1 gpc480 (
      {stage0_14[206]},
      {stage1_14[107]}
   );
   gpc1_1 gpc481 (
      {stage0_14[207]},
      {stage1_14[108]}
   );
   gpc1_1 gpc482 (
      {stage0_14[208]},
      {stage1_14[109]}
   );
   gpc1_1 gpc483 (
      {stage0_14[209]},
      {stage1_14[110]}
   );
   gpc1_1 gpc484 (
      {stage0_14[210]},
      {stage1_14[111]}
   );
   gpc1_1 gpc485 (
      {stage0_14[211]},
      {stage1_14[112]}
   );
   gpc1_1 gpc486 (
      {stage0_14[212]},
      {stage1_14[113]}
   );
   gpc1_1 gpc487 (
      {stage0_14[213]},
      {stage1_14[114]}
   );
   gpc1_1 gpc488 (
      {stage0_14[214]},
      {stage1_14[115]}
   );
   gpc1_1 gpc489 (
      {stage0_14[215]},
      {stage1_14[116]}
   );
   gpc1_1 gpc490 (
      {stage0_14[216]},
      {stage1_14[117]}
   );
   gpc1_1 gpc491 (
      {stage0_14[217]},
      {stage1_14[118]}
   );
   gpc1_1 gpc492 (
      {stage0_14[218]},
      {stage1_14[119]}
   );
   gpc1_1 gpc493 (
      {stage0_14[219]},
      {stage1_14[120]}
   );
   gpc1_1 gpc494 (
      {stage0_14[220]},
      {stage1_14[121]}
   );
   gpc1_1 gpc495 (
      {stage0_14[221]},
      {stage1_14[122]}
   );
   gpc1_1 gpc496 (
      {stage0_14[222]},
      {stage1_14[123]}
   );
   gpc1_1 gpc497 (
      {stage0_14[223]},
      {stage1_14[124]}
   );
   gpc1_1 gpc498 (
      {stage0_14[224]},
      {stage1_14[125]}
   );
   gpc1_1 gpc499 (
      {stage0_14[225]},
      {stage1_14[126]}
   );
   gpc1_1 gpc500 (
      {stage0_14[226]},
      {stage1_14[127]}
   );
   gpc1_1 gpc501 (
      {stage0_14[227]},
      {stage1_14[128]}
   );
   gpc1_1 gpc502 (
      {stage0_14[228]},
      {stage1_14[129]}
   );
   gpc1_1 gpc503 (
      {stage0_14[229]},
      {stage1_14[130]}
   );
   gpc1_1 gpc504 (
      {stage0_14[230]},
      {stage1_14[131]}
   );
   gpc1_1 gpc505 (
      {stage0_14[231]},
      {stage1_14[132]}
   );
   gpc1_1 gpc506 (
      {stage0_14[232]},
      {stage1_14[133]}
   );
   gpc1_1 gpc507 (
      {stage0_14[233]},
      {stage1_14[134]}
   );
   gpc1_1 gpc508 (
      {stage0_14[234]},
      {stage1_14[135]}
   );
   gpc1_1 gpc509 (
      {stage0_14[235]},
      {stage1_14[136]}
   );
   gpc1_1 gpc510 (
      {stage0_14[236]},
      {stage1_14[137]}
   );
   gpc1_1 gpc511 (
      {stage0_14[237]},
      {stage1_14[138]}
   );
   gpc1_1 gpc512 (
      {stage0_14[238]},
      {stage1_14[139]}
   );
   gpc1_1 gpc513 (
      {stage0_14[239]},
      {stage1_14[140]}
   );
   gpc1_1 gpc514 (
      {stage0_14[240]},
      {stage1_14[141]}
   );
   gpc1_1 gpc515 (
      {stage0_14[241]},
      {stage1_14[142]}
   );
   gpc1_1 gpc516 (
      {stage0_14[242]},
      {stage1_14[143]}
   );
   gpc1_1 gpc517 (
      {stage0_14[243]},
      {stage1_14[144]}
   );
   gpc1_1 gpc518 (
      {stage0_14[244]},
      {stage1_14[145]}
   );
   gpc1_1 gpc519 (
      {stage0_14[245]},
      {stage1_14[146]}
   );
   gpc1_1 gpc520 (
      {stage0_14[246]},
      {stage1_14[147]}
   );
   gpc1_1 gpc521 (
      {stage0_14[247]},
      {stage1_14[148]}
   );
   gpc1_1 gpc522 (
      {stage0_14[248]},
      {stage1_14[149]}
   );
   gpc1_1 gpc523 (
      {stage0_14[249]},
      {stage1_14[150]}
   );
   gpc1_1 gpc524 (
      {stage0_14[250]},
      {stage1_14[151]}
   );
   gpc1_1 gpc525 (
      {stage0_14[251]},
      {stage1_14[152]}
   );
   gpc1_1 gpc526 (
      {stage0_14[252]},
      {stage1_14[153]}
   );
   gpc1_1 gpc527 (
      {stage0_14[253]},
      {stage1_14[154]}
   );
   gpc1_1 gpc528 (
      {stage0_14[254]},
      {stage1_14[155]}
   );
   gpc1_1 gpc529 (
      {stage0_14[255]},
      {stage1_14[156]}
   );
   gpc1_1 gpc530 (
      {stage0_15[252]},
      {stage1_15[72]}
   );
   gpc1_1 gpc531 (
      {stage0_15[253]},
      {stage1_15[73]}
   );
   gpc1_1 gpc532 (
      {stage0_15[254]},
      {stage1_15[74]}
   );
   gpc1_1 gpc533 (
      {stage0_15[255]},
      {stage1_15[75]}
   );
   gpc606_5 gpc534 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc535 (
      {stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc606_5 gpc536 (
      {stage1_0[12], stage1_0[13], stage1_0[14], stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc606_5 gpc537 (
      {stage1_0[18], stage1_0[19], stage1_0[20], stage1_0[21], stage1_0[22], stage1_0[23]},
      {stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc606_5 gpc538 (
      {stage1_0[24], stage1_0[25], stage1_0[26], stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27], stage1_2[28], stage1_2[29]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc606_5 gpc539 (
      {stage1_0[30], stage1_0[31], stage1_0[32], stage1_0[33], stage1_0[34], stage1_0[35]},
      {stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33], stage1_2[34], stage1_2[35]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc606_5 gpc540 (
      {stage1_0[36], stage1_0[37], stage1_0[38], stage1_0[39], stage1_0[40], stage1_0[41]},
      {stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39], stage1_2[40], stage1_2[41]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc606_5 gpc541 (
      {stage1_0[42], stage1_0[43], stage1_0[44], stage1_0[45], stage1_0[46], stage1_0[47]},
      {stage1_2[42], stage1_2[43], stage1_2[44], stage1_2[45], stage1_2[46], stage1_2[47]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc606_5 gpc542 (
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage2_5[0],stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8]}
   );
   gpc606_5 gpc543 (
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage2_5[1],stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9]}
   );
   gpc606_5 gpc544 (
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage2_5[2],stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10]}
   );
   gpc606_5 gpc545 (
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23]},
      {stage2_5[3],stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11]}
   );
   gpc606_5 gpc546 (
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27], stage1_3[28], stage1_3[29]},
      {stage2_5[4],stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12]}
   );
   gpc606_5 gpc547 (
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_3[30], stage1_3[31], stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35]},
      {stage2_5[5],stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13]}
   );
   gpc606_5 gpc548 (
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_3[36], stage1_3[37], stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41]},
      {stage2_5[6],stage2_4[14],stage2_3[14],stage2_2[14],stage2_1[14]}
   );
   gpc606_5 gpc549 (
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_3[42], stage1_3[43], stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47]},
      {stage2_5[7],stage2_4[15],stage2_3[15],stage2_2[15],stage2_1[15]}
   );
   gpc606_5 gpc550 (
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_3[48], stage1_3[49], stage1_3[50], stage1_3[51], stage1_3[52], stage1_3[53]},
      {stage2_5[8],stage2_4[16],stage2_3[16],stage2_2[16],stage2_1[16]}
   );
   gpc606_5 gpc551 (
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59]},
      {stage1_3[54], stage1_3[55], stage1_3[56], stage1_3[57], stage1_3[58], stage1_3[59]},
      {stage2_5[9],stage2_4[17],stage2_3[17],stage2_2[17],stage2_1[17]}
   );
   gpc606_5 gpc552 (
      {stage1_1[60], stage1_1[61], stage1_1[62], stage1_1[63], stage1_1[64], stage1_1[65]},
      {stage1_3[60], stage1_3[61], stage1_3[62], stage1_3[63], stage1_3[64], stage1_3[65]},
      {stage2_5[10],stage2_4[18],stage2_3[18],stage2_2[18],stage2_1[18]}
   );
   gpc606_5 gpc553 (
      {stage1_1[66], stage1_1[67], stage1_1[68], stage1_1[69], stage1_1[70], stage1_1[71]},
      {stage1_3[66], stage1_3[67], stage1_3[68], stage1_3[69], stage1_3[70], stage1_3[71]},
      {stage2_5[11],stage2_4[19],stage2_3[19],stage2_2[19],stage2_1[19]}
   );
   gpc606_5 gpc554 (
      {stage1_1[72], stage1_1[73], stage1_1[74], stage1_1[75], stage1_1[76], stage1_1[77]},
      {stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75], stage1_3[76], stage1_3[77]},
      {stage2_5[12],stage2_4[20],stage2_3[20],stage2_2[20],stage2_1[20]}
   );
   gpc606_5 gpc555 (
      {stage1_1[78], stage1_1[79], stage1_1[80], stage1_1[81], stage1_1[82], stage1_1[83]},
      {stage1_3[78], stage1_3[79], stage1_3[80], stage1_3[81], stage1_3[82], stage1_3[83]},
      {stage2_5[13],stage2_4[21],stage2_3[21],stage2_2[21],stage2_1[21]}
   );
   gpc606_5 gpc556 (
      {stage1_1[84], stage1_1[85], stage1_1[86], stage1_1[87], stage1_1[88], stage1_1[89]},
      {stage1_3[84], stage1_3[85], stage1_3[86], stage1_3[87], stage1_3[88], stage1_3[89]},
      {stage2_5[14],stage2_4[22],stage2_3[22],stage2_2[22],stage2_1[22]}
   );
   gpc606_5 gpc557 (
      {stage1_1[90], stage1_1[91], stage1_1[92], stage1_1[93], stage1_1[94], stage1_1[95]},
      {stage1_3[90], stage1_3[91], stage1_3[92], stage1_3[93], stage1_3[94], stage1_3[95]},
      {stage2_5[15],stage2_4[23],stage2_3[23],stage2_2[23],stage2_1[23]}
   );
   gpc606_5 gpc558 (
      {stage1_2[48], stage1_2[49], stage1_2[50], stage1_2[51], stage1_2[52], stage1_2[53]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[16],stage2_4[24],stage2_3[24],stage2_2[24]}
   );
   gpc606_5 gpc559 (
      {stage1_2[54], stage1_2[55], stage1_2[56], stage1_2[57], stage1_2[58], stage1_2[59]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[17],stage2_4[25],stage2_3[25],stage2_2[25]}
   );
   gpc606_5 gpc560 (
      {stage1_2[60], stage1_2[61], stage1_2[62], stage1_2[63], stage1_2[64], stage1_2[65]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[18],stage2_4[26],stage2_3[26],stage2_2[26]}
   );
   gpc606_5 gpc561 (
      {stage1_2[66], stage1_2[67], stage1_2[68], stage1_2[69], stage1_2[70], stage1_2[71]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[19],stage2_4[27],stage2_3[27],stage2_2[27]}
   );
   gpc615_5 gpc562 (
      {stage1_2[72], stage1_2[73], stage1_2[74], stage1_2[75], stage1_2[76]},
      {stage1_3[96]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[20],stage2_4[28],stage2_3[28],stage2_2[28]}
   );
   gpc615_5 gpc563 (
      {stage1_2[77], stage1_2[78], stage1_2[79], stage1_2[80], stage1_2[81]},
      {stage1_3[97]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[21],stage2_4[29],stage2_3[29],stage2_2[29]}
   );
   gpc615_5 gpc564 (
      {stage1_3[98], stage1_3[99], stage1_3[100], stage1_3[101], stage1_3[102]},
      {stage1_4[36]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[6],stage2_5[22],stage2_4[30],stage2_3[30]}
   );
   gpc615_5 gpc565 (
      {stage1_3[103], stage1_3[104], stage1_3[105], stage1_3[106], stage1_3[107]},
      {stage1_4[37]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[7],stage2_5[23],stage2_4[31],stage2_3[31]}
   );
   gpc615_5 gpc566 (
      {stage1_3[108], stage1_3[109], stage1_3[110], stage1_3[111], stage1_3[112]},
      {stage1_4[38]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[8],stage2_5[24],stage2_4[32],stage2_3[32]}
   );
   gpc606_5 gpc567 (
      {stage1_4[39], stage1_4[40], stage1_4[41], stage1_4[42], stage1_4[43], stage1_4[44]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[3],stage2_6[9],stage2_5[25],stage2_4[33]}
   );
   gpc606_5 gpc568 (
      {stage1_4[45], stage1_4[46], stage1_4[47], stage1_4[48], stage1_4[49], stage1_4[50]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[4],stage2_6[10],stage2_5[26],stage2_4[34]}
   );
   gpc606_5 gpc569 (
      {stage1_4[51], stage1_4[52], stage1_4[53], stage1_4[54], stage1_4[55], stage1_4[56]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[5],stage2_6[11],stage2_5[27],stage2_4[35]}
   );
   gpc615_5 gpc570 (
      {stage1_4[57], stage1_4[58], stage1_4[59], stage1_4[60], stage1_4[61]},
      {stage1_5[18]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[6],stage2_6[12],stage2_5[28],stage2_4[36]}
   );
   gpc615_5 gpc571 (
      {stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65], stage1_4[66]},
      {stage1_5[19]},
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage2_8[4],stage2_7[7],stage2_6[13],stage2_5[29],stage2_4[37]}
   );
   gpc615_5 gpc572 (
      {stage1_4[67], stage1_4[68], stage1_4[69], stage1_4[70], stage1_4[71]},
      {stage1_5[20]},
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage2_8[5],stage2_7[8],stage2_6[14],stage2_5[30],stage2_4[38]}
   );
   gpc615_5 gpc573 (
      {stage1_4[72], stage1_4[73], stage1_4[74], stage1_4[75], stage1_4[76]},
      {stage1_5[21]},
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage2_8[6],stage2_7[9],stage2_6[15],stage2_5[31],stage2_4[39]}
   );
   gpc615_5 gpc574 (
      {stage1_4[77], stage1_4[78], stage1_4[79], stage1_4[80], stage1_4[81]},
      {stage1_5[22]},
      {stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47]},
      {stage2_8[7],stage2_7[10],stage2_6[16],stage2_5[32],stage2_4[40]}
   );
   gpc615_5 gpc575 (
      {stage1_4[82], stage1_4[83], stage1_4[84], stage1_4[85], stage1_4[86]},
      {stage1_5[23]},
      {stage1_6[48], stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53]},
      {stage2_8[8],stage2_7[11],stage2_6[17],stage2_5[33],stage2_4[41]}
   );
   gpc615_5 gpc576 (
      {stage1_4[87], stage1_4[88], stage1_4[89], stage1_4[90], stage1_4[91]},
      {stage1_5[24]},
      {stage1_6[54], stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59]},
      {stage2_8[9],stage2_7[12],stage2_6[18],stage2_5[34],stage2_4[42]}
   );
   gpc615_5 gpc577 (
      {stage1_4[92], stage1_4[93], stage1_4[94], stage1_4[95], stage1_4[96]},
      {stage1_5[25]},
      {stage1_6[60], stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65]},
      {stage2_8[10],stage2_7[13],stage2_6[19],stage2_5[35],stage2_4[43]}
   );
   gpc615_5 gpc578 (
      {stage1_4[97], stage1_4[98], stage1_4[99], stage1_4[100], stage1_4[101]},
      {stage1_5[26]},
      {stage1_6[66], stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71]},
      {stage2_8[11],stage2_7[14],stage2_6[20],stage2_5[36],stage2_4[44]}
   );
   gpc615_5 gpc579 (
      {stage1_4[102], stage1_4[103], stage1_4[104], stage1_4[105], stage1_4[106]},
      {stage1_5[27]},
      {stage1_6[72], stage1_6[73], stage1_6[74], stage1_6[75], stage1_6[76], stage1_6[77]},
      {stage2_8[12],stage2_7[15],stage2_6[21],stage2_5[37],stage2_4[45]}
   );
   gpc615_5 gpc580 (
      {stage1_4[107], stage1_4[108], stage1_4[109], stage1_4[110], stage1_4[111]},
      {stage1_5[28]},
      {stage1_6[78], stage1_6[79], stage1_6[80], stage1_6[81], stage1_6[82], stage1_6[83]},
      {stage2_8[13],stage2_7[16],stage2_6[22],stage2_5[38],stage2_4[46]}
   );
   gpc615_5 gpc581 (
      {stage1_4[112], stage1_4[113], stage1_4[114], stage1_4[115], stage1_4[116]},
      {stage1_5[29]},
      {stage1_6[84], stage1_6[85], stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89]},
      {stage2_8[14],stage2_7[17],stage2_6[23],stage2_5[39],stage2_4[47]}
   );
   gpc615_5 gpc582 (
      {stage1_4[117], stage1_4[118], stage1_4[119], stage1_4[120], stage1_4[121]},
      {stage1_5[30]},
      {stage1_6[90], stage1_6[91], stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95]},
      {stage2_8[15],stage2_7[18],stage2_6[24],stage2_5[40],stage2_4[48]}
   );
   gpc615_5 gpc583 (
      {stage1_4[122], stage1_4[123], stage1_4[124], stage1_4[125], stage1_4[126]},
      {stage1_5[31]},
      {stage1_6[96], stage1_6[97], stage1_6[98], stage1_6[99], stage1_6[100], stage1_6[101]},
      {stage2_8[16],stage2_7[19],stage2_6[25],stage2_5[41],stage2_4[49]}
   );
   gpc606_5 gpc584 (
      {stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35], stage1_5[36], stage1_5[37]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[17],stage2_7[20],stage2_6[26],stage2_5[42]}
   );
   gpc606_5 gpc585 (
      {stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41], stage1_5[42], stage1_5[43]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[18],stage2_7[21],stage2_6[27],stage2_5[43]}
   );
   gpc606_5 gpc586 (
      {stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47], stage1_5[48], stage1_5[49]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[19],stage2_7[22],stage2_6[28],stage2_5[44]}
   );
   gpc606_5 gpc587 (
      {stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53], stage1_5[54], stage1_5[55]},
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage2_9[3],stage2_8[20],stage2_7[23],stage2_6[29],stage2_5[45]}
   );
   gpc606_5 gpc588 (
      {stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59], stage1_5[60], stage1_5[61]},
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29]},
      {stage2_9[4],stage2_8[21],stage2_7[24],stage2_6[30],stage2_5[46]}
   );
   gpc606_5 gpc589 (
      {stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65], stage1_5[66], stage1_5[67]},
      {stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35]},
      {stage2_9[5],stage2_8[22],stage2_7[25],stage2_6[31],stage2_5[47]}
   );
   gpc606_5 gpc590 (
      {stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71], stage1_5[72], stage1_5[73]},
      {stage1_7[36], stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage2_9[6],stage2_8[23],stage2_7[26],stage2_6[32],stage2_5[48]}
   );
   gpc606_5 gpc591 (
      {stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77], stage1_5[78], stage1_5[79]},
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47]},
      {stage2_9[7],stage2_8[24],stage2_7[27],stage2_6[33],stage2_5[49]}
   );
   gpc606_5 gpc592 (
      {stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83], stage1_5[84], stage1_5[85]},
      {stage1_7[48], stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53]},
      {stage2_9[8],stage2_8[25],stage2_7[28],stage2_6[34],stage2_5[50]}
   );
   gpc606_5 gpc593 (
      {stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89], stage1_5[90], stage1_5[91]},
      {stage1_7[54], stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58], stage1_7[59]},
      {stage2_9[9],stage2_8[26],stage2_7[29],stage2_6[35],stage2_5[51]}
   );
   gpc606_5 gpc594 (
      {stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95], stage1_5[96], stage1_5[97]},
      {stage1_7[60], stage1_7[61], stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65]},
      {stage2_9[10],stage2_8[27],stage2_7[30],stage2_6[36],stage2_5[52]}
   );
   gpc606_5 gpc595 (
      {stage1_5[98], stage1_5[99], stage1_5[100], stage1_5[101], stage1_5[102], stage1_5[103]},
      {stage1_7[66], stage1_7[67], stage1_7[68], stage1_7[69], stage1_7[70], stage1_7[71]},
      {stage2_9[11],stage2_8[28],stage2_7[31],stage2_6[37],stage2_5[53]}
   );
   gpc615_5 gpc596 (
      {stage1_7[72], stage1_7[73], stage1_7[74], stage1_7[75], stage1_7[76]},
      {stage1_8[0]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[0],stage2_9[12],stage2_8[29],stage2_7[32]}
   );
   gpc615_5 gpc597 (
      {stage1_7[77], stage1_7[78], stage1_7[79], stage1_7[80], stage1_7[81]},
      {stage1_8[1]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[1],stage2_9[13],stage2_8[30],stage2_7[33]}
   );
   gpc615_5 gpc598 (
      {stage1_7[82], stage1_7[83], stage1_7[84], stage1_7[85], stage1_7[86]},
      {stage1_8[2]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[2],stage2_9[14],stage2_8[31],stage2_7[34]}
   );
   gpc615_5 gpc599 (
      {stage1_7[87], stage1_7[88], stage1_7[89], stage1_7[90], stage1_7[91]},
      {stage1_8[3]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[3],stage2_9[15],stage2_8[32],stage2_7[35]}
   );
   gpc606_5 gpc600 (
      {stage1_8[4], stage1_8[5], stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[4],stage2_10[4],stage2_9[16],stage2_8[33]}
   );
   gpc606_5 gpc601 (
      {stage1_8[10], stage1_8[11], stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[5],stage2_10[5],stage2_9[17],stage2_8[34]}
   );
   gpc606_5 gpc602 (
      {stage1_8[16], stage1_8[17], stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[6],stage2_10[6],stage2_9[18],stage2_8[35]}
   );
   gpc606_5 gpc603 (
      {stage1_8[22], stage1_8[23], stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[7],stage2_10[7],stage2_9[19],stage2_8[36]}
   );
   gpc606_5 gpc604 (
      {stage1_8[28], stage1_8[29], stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[8],stage2_10[8],stage2_9[20],stage2_8[37]}
   );
   gpc606_5 gpc605 (
      {stage1_8[34], stage1_8[35], stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[9],stage2_10[9],stage2_9[21],stage2_8[38]}
   );
   gpc606_5 gpc606 (
      {stage1_8[40], stage1_8[41], stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45]},
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage2_12[6],stage2_11[10],stage2_10[10],stage2_9[22],stage2_8[39]}
   );
   gpc606_5 gpc607 (
      {stage1_8[46], stage1_8[47], stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51]},
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage2_12[7],stage2_11[11],stage2_10[11],stage2_9[23],stage2_8[40]}
   );
   gpc606_5 gpc608 (
      {stage1_8[52], stage1_8[53], stage1_8[54], stage1_8[55], stage1_8[56], stage1_8[57]},
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage2_12[8],stage2_11[12],stage2_10[12],stage2_9[24],stage2_8[41]}
   );
   gpc606_5 gpc609 (
      {stage1_8[58], stage1_8[59], stage1_8[60], stage1_8[61], stage1_8[62], stage1_8[63]},
      {stage1_10[54], stage1_10[55], stage1_10[56], stage1_10[57], stage1_10[58], stage1_10[59]},
      {stage2_12[9],stage2_11[13],stage2_10[13],stage2_9[25],stage2_8[42]}
   );
   gpc606_5 gpc610 (
      {stage1_8[64], stage1_8[65], stage1_8[66], stage1_8[67], stage1_8[68], stage1_8[69]},
      {stage1_10[60], stage1_10[61], stage1_10[62], stage1_10[63], stage1_10[64], stage1_10[65]},
      {stage2_12[10],stage2_11[14],stage2_10[14],stage2_9[26],stage2_8[43]}
   );
   gpc606_5 gpc611 (
      {stage1_8[70], stage1_8[71], stage1_8[72], stage1_8[73], stage1_8[74], stage1_8[75]},
      {stage1_10[66], stage1_10[67], stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71]},
      {stage2_12[11],stage2_11[15],stage2_10[15],stage2_9[27],stage2_8[44]}
   );
   gpc606_5 gpc612 (
      {stage1_8[76], stage1_8[77], stage1_8[78], stage1_8[79], stage1_8[80], stage1_8[81]},
      {stage1_10[72], stage1_10[73], stage1_10[74], stage1_10[75], stage1_10[76], stage1_10[77]},
      {stage2_12[12],stage2_11[16],stage2_10[16],stage2_9[28],stage2_8[45]}
   );
   gpc606_5 gpc613 (
      {stage1_8[82], stage1_8[83], stage1_8[84], stage1_8[85], stage1_8[86], stage1_8[87]},
      {stage1_10[78], stage1_10[79], stage1_10[80], stage1_10[81], stage1_10[82], stage1_10[83]},
      {stage2_12[13],stage2_11[17],stage2_10[17],stage2_9[29],stage2_8[46]}
   );
   gpc606_5 gpc614 (
      {stage1_8[88], stage1_8[89], stage1_8[90], stage1_8[91], stage1_8[92], stage1_8[93]},
      {stage1_10[84], stage1_10[85], stage1_10[86], stage1_10[87], stage1_10[88], stage1_10[89]},
      {stage2_12[14],stage2_11[18],stage2_10[18],stage2_9[30],stage2_8[47]}
   );
   gpc606_5 gpc615 (
      {stage1_8[94], stage1_8[95], stage1_8[96], stage1_8[97], stage1_8[98], stage1_8[99]},
      {stage1_10[90], stage1_10[91], stage1_10[92], stage1_10[93], stage1_10[94], stage1_10[95]},
      {stage2_12[15],stage2_11[19],stage2_10[19],stage2_9[31],stage2_8[48]}
   );
   gpc606_5 gpc616 (
      {stage1_8[100], stage1_8[101], stage1_8[102], stage1_8[103], stage1_8[104], stage1_8[105]},
      {stage1_10[96], stage1_10[97], stage1_10[98], stage1_10[99], stage1_10[100], stage1_10[101]},
      {stage2_12[16],stage2_11[20],stage2_10[20],stage2_9[32],stage2_8[49]}
   );
   gpc117_4 gpc617 (
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29], stage1_9[30]},
      {stage1_10[102]},
      {stage1_11[0]},
      {stage2_12[17],stage2_11[21],stage2_10[21],stage2_9[33]}
   );
   gpc117_4 gpc618 (
      {stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35], stage1_9[36], stage1_9[37]},
      {stage1_10[103]},
      {stage1_11[1]},
      {stage2_12[18],stage2_11[22],stage2_10[22],stage2_9[34]}
   );
   gpc117_4 gpc619 (
      {stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41], stage1_9[42], stage1_9[43], stage1_9[44]},
      {stage1_10[104]},
      {stage1_11[2]},
      {stage2_12[19],stage2_11[23],stage2_10[23],stage2_9[35]}
   );
   gpc117_4 gpc620 (
      {stage1_9[45], stage1_9[46], stage1_9[47], stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51]},
      {stage1_10[105]},
      {stage1_11[3]},
      {stage2_12[20],stage2_11[24],stage2_10[24],stage2_9[36]}
   );
   gpc117_4 gpc621 (
      {stage1_9[52], stage1_9[53], stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58]},
      {stage1_10[106]},
      {stage1_11[4]},
      {stage2_12[21],stage2_11[25],stage2_10[25],stage2_9[37]}
   );
   gpc117_4 gpc622 (
      {stage1_9[59], stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage1_10[107]},
      {stage1_11[5]},
      {stage2_12[22],stage2_11[26],stage2_10[26],stage2_9[38]}
   );
   gpc117_4 gpc623 (
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71], stage1_9[72]},
      {stage1_10[108]},
      {stage1_11[6]},
      {stage2_12[23],stage2_11[27],stage2_10[27],stage2_9[39]}
   );
   gpc606_5 gpc624 (
      {stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77], stage1_9[78]},
      {stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11], stage1_11[12]},
      {stage2_13[0],stage2_12[24],stage2_11[28],stage2_10[28],stage2_9[40]}
   );
   gpc606_5 gpc625 (
      {stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83], stage1_9[84]},
      {stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17], stage1_11[18]},
      {stage2_13[1],stage2_12[25],stage2_11[29],stage2_10[29],stage2_9[41]}
   );
   gpc606_5 gpc626 (
      {stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89], stage1_9[90]},
      {stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23], stage1_11[24]},
      {stage2_13[2],stage2_12[26],stage2_11[30],stage2_10[30],stage2_9[42]}
   );
   gpc606_5 gpc627 (
      {stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95], stage1_9[96]},
      {stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29], stage1_11[30]},
      {stage2_13[3],stage2_12[27],stage2_11[31],stage2_10[31],stage2_9[43]}
   );
   gpc606_5 gpc628 (
      {stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100], stage1_9[101], stage1_9[102]},
      {stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35], stage1_11[36]},
      {stage2_13[4],stage2_12[28],stage2_11[32],stage2_10[32],stage2_9[44]}
   );
   gpc606_5 gpc629 (
      {stage1_9[103], stage1_9[104], stage1_9[105], stage1_9[106], stage1_9[107], stage1_9[108]},
      {stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41], stage1_11[42]},
      {stage2_13[5],stage2_12[29],stage2_11[33],stage2_10[33],stage2_9[45]}
   );
   gpc606_5 gpc630 (
      {stage1_9[109], stage1_9[110], stage1_9[111], stage1_9[112], stage1_9[113], stage1_9[114]},
      {stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47], stage1_11[48]},
      {stage2_13[6],stage2_12[30],stage2_11[34],stage2_10[34],stage2_9[46]}
   );
   gpc615_5 gpc631 (
      {stage1_10[109], stage1_10[110], stage1_10[111], stage1_10[112], stage1_10[113]},
      {stage1_11[49]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[7],stage2_12[31],stage2_11[35],stage2_10[35]}
   );
   gpc606_5 gpc632 (
      {stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53], stage1_11[54], stage1_11[55]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[1],stage2_13[8],stage2_12[32],stage2_11[36]}
   );
   gpc606_5 gpc633 (
      {stage1_11[56], stage1_11[57], stage1_11[58], stage1_11[59], stage1_11[60], stage1_11[61]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[2],stage2_13[9],stage2_12[33],stage2_11[37]}
   );
   gpc606_5 gpc634 (
      {stage1_11[62], stage1_11[63], stage1_11[64], stage1_11[65], stage1_11[66], stage1_11[67]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[3],stage2_13[10],stage2_12[34],stage2_11[38]}
   );
   gpc606_5 gpc635 (
      {stage1_11[68], stage1_11[69], stage1_11[70], stage1_11[71], stage1_11[72], stage1_11[73]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[4],stage2_13[11],stage2_12[35],stage2_11[39]}
   );
   gpc606_5 gpc636 (
      {stage1_11[74], stage1_11[75], stage1_11[76], stage1_11[77], stage1_11[78], stage1_11[79]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[5],stage2_13[12],stage2_12[36],stage2_11[40]}
   );
   gpc615_5 gpc637 (
      {stage1_11[80], stage1_11[81], stage1_11[82], stage1_11[83], stage1_11[84]},
      {stage1_12[6]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[6],stage2_13[13],stage2_12[37],stage2_11[41]}
   );
   gpc615_5 gpc638 (
      {stage1_11[85], stage1_11[86], stage1_11[87], stage1_11[88], stage1_11[89]},
      {stage1_12[7]},
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage2_15[6],stage2_14[7],stage2_13[14],stage2_12[38],stage2_11[42]}
   );
   gpc615_5 gpc639 (
      {stage1_11[90], stage1_11[91], stage1_11[92], stage1_11[93], stage1_11[94]},
      {stage1_12[8]},
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage2_15[7],stage2_14[8],stage2_13[15],stage2_12[39],stage2_11[43]}
   );
   gpc615_5 gpc640 (
      {stage1_11[95], stage1_11[96], stage1_11[97], stage1_11[98], stage1_11[99]},
      {stage1_12[9]},
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage2_15[8],stage2_14[9],stage2_13[16],stage2_12[40],stage2_11[44]}
   );
   gpc615_5 gpc641 (
      {stage1_11[100], stage1_11[101], stage1_11[102], stage1_11[103], stage1_11[104]},
      {stage1_12[10]},
      {stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59]},
      {stage2_15[9],stage2_14[10],stage2_13[17],stage2_12[41],stage2_11[45]}
   );
   gpc615_5 gpc642 (
      {stage1_11[105], stage1_11[106], stage1_11[107], stage1_11[108], stage1_11[109]},
      {stage1_12[11]},
      {stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage2_15[10],stage2_14[11],stage2_13[18],stage2_12[42],stage2_11[46]}
   );
   gpc615_5 gpc643 (
      {stage1_11[110], stage1_11[111], stage1_11[112], stage1_11[113], stage1_11[114]},
      {stage1_12[12]},
      {stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69], stage1_13[70], stage1_13[71]},
      {stage2_15[11],stage2_14[12],stage2_13[19],stage2_12[43],stage2_11[47]}
   );
   gpc606_5 gpc644 (
      {stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17], stage1_12[18]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[12],stage2_14[13],stage2_13[20],stage2_12[44]}
   );
   gpc606_5 gpc645 (
      {stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23], stage1_12[24]},
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage2_16[1],stage2_15[13],stage2_14[14],stage2_13[21],stage2_12[45]}
   );
   gpc606_5 gpc646 (
      {stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29], stage1_12[30]},
      {stage1_14[12], stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17]},
      {stage2_16[2],stage2_15[14],stage2_14[15],stage2_13[22],stage2_12[46]}
   );
   gpc606_5 gpc647 (
      {stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35], stage1_12[36]},
      {stage1_14[18], stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23]},
      {stage2_16[3],stage2_15[15],stage2_14[16],stage2_13[23],stage2_12[47]}
   );
   gpc615_5 gpc648 (
      {stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage1_13[72]},
      {stage1_14[24], stage1_14[25], stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29]},
      {stage2_16[4],stage2_15[16],stage2_14[17],stage2_13[24],stage2_12[48]}
   );
   gpc615_5 gpc649 (
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46]},
      {stage1_13[73]},
      {stage1_14[30], stage1_14[31], stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35]},
      {stage2_16[5],stage2_15[17],stage2_14[18],stage2_13[25],stage2_12[49]}
   );
   gpc615_5 gpc650 (
      {stage1_12[47], stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51]},
      {stage1_13[74]},
      {stage1_14[36], stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41]},
      {stage2_16[6],stage2_15[18],stage2_14[19],stage2_13[26],stage2_12[50]}
   );
   gpc615_5 gpc651 (
      {stage1_12[52], stage1_12[53], stage1_12[54], stage1_12[55], stage1_12[56]},
      {stage1_13[75]},
      {stage1_14[42], stage1_14[43], stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47]},
      {stage2_16[7],stage2_15[19],stage2_14[20],stage2_13[27],stage2_12[51]}
   );
   gpc615_5 gpc652 (
      {stage1_12[57], stage1_12[58], stage1_12[59], stage1_12[60], stage1_12[61]},
      {stage1_13[76]},
      {stage1_14[48], stage1_14[49], stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53]},
      {stage2_16[8],stage2_15[20],stage2_14[21],stage2_13[28],stage2_12[52]}
   );
   gpc615_5 gpc653 (
      {stage1_12[62], stage1_12[63], stage1_12[64], stage1_12[65], stage1_12[66]},
      {stage1_13[77]},
      {stage1_14[54], stage1_14[55], stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59]},
      {stage2_16[9],stage2_15[21],stage2_14[22],stage2_13[29],stage2_12[53]}
   );
   gpc615_5 gpc654 (
      {stage1_12[67], stage1_12[68], stage1_12[69], stage1_12[70], stage1_12[71]},
      {stage1_13[78]},
      {stage1_14[60], stage1_14[61], stage1_14[62], stage1_14[63], stage1_14[64], stage1_14[65]},
      {stage2_16[10],stage2_15[22],stage2_14[23],stage2_13[30],stage2_12[54]}
   );
   gpc615_5 gpc655 (
      {stage1_12[72], stage1_12[73], stage1_12[74], stage1_12[75], stage1_12[76]},
      {stage1_13[79]},
      {stage1_14[66], stage1_14[67], stage1_14[68], stage1_14[69], stage1_14[70], stage1_14[71]},
      {stage2_16[11],stage2_15[23],stage2_14[24],stage2_13[31],stage2_12[55]}
   );
   gpc615_5 gpc656 (
      {stage1_12[77], stage1_12[78], stage1_12[79], stage1_12[80], stage1_12[81]},
      {stage1_13[80]},
      {stage1_14[72], stage1_14[73], stage1_14[74], stage1_14[75], stage1_14[76], stage1_14[77]},
      {stage2_16[12],stage2_15[24],stage2_14[25],stage2_13[32],stage2_12[56]}
   );
   gpc615_5 gpc657 (
      {stage1_12[82], stage1_12[83], stage1_12[84], stage1_12[85], stage1_12[86]},
      {stage1_13[81]},
      {stage1_14[78], stage1_14[79], stage1_14[80], stage1_14[81], stage1_14[82], stage1_14[83]},
      {stage2_16[13],stage2_15[25],stage2_14[26],stage2_13[33],stage2_12[57]}
   );
   gpc615_5 gpc658 (
      {stage1_12[87], stage1_12[88], stage1_12[89], stage1_12[90], stage1_12[91]},
      {stage1_13[82]},
      {stage1_14[84], stage1_14[85], stage1_14[86], stage1_14[87], stage1_14[88], stage1_14[89]},
      {stage2_16[14],stage2_15[26],stage2_14[27],stage2_13[34],stage2_12[58]}
   );
   gpc615_5 gpc659 (
      {stage1_12[92], stage1_12[93], stage1_12[94], stage1_12[95], stage1_12[96]},
      {stage1_13[83]},
      {stage1_14[90], stage1_14[91], stage1_14[92], stage1_14[93], stage1_14[94], stage1_14[95]},
      {stage2_16[15],stage2_15[27],stage2_14[28],stage2_13[35],stage2_12[59]}
   );
   gpc615_5 gpc660 (
      {stage1_12[97], stage1_12[98], stage1_12[99], stage1_12[100], stage1_12[101]},
      {stage1_13[84]},
      {stage1_14[96], stage1_14[97], stage1_14[98], stage1_14[99], stage1_14[100], stage1_14[101]},
      {stage2_16[16],stage2_15[28],stage2_14[29],stage2_13[36],stage2_12[60]}
   );
   gpc606_5 gpc661 (
      {stage1_13[85], stage1_13[86], stage1_13[87], stage1_13[88], stage1_13[89], stage1_13[90]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[17],stage2_15[29],stage2_14[30],stage2_13[37]}
   );
   gpc606_5 gpc662 (
      {stage1_13[91], stage1_13[92], stage1_13[93], stage1_13[94], stage1_13[95], stage1_13[96]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[18],stage2_15[30],stage2_14[31],stage2_13[38]}
   );
   gpc606_5 gpc663 (
      {stage1_13[97], stage1_13[98], stage1_13[99], stage1_13[100], stage1_13[101], stage1_13[102]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[19],stage2_15[31],stage2_14[32],stage2_13[39]}
   );
   gpc606_5 gpc664 (
      {stage1_13[103], stage1_13[104], stage1_13[105], stage1_13[106], stage1_13[107], stage1_13[108]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[20],stage2_15[32],stage2_14[33],stage2_13[40]}
   );
   gpc606_5 gpc665 (
      {stage1_13[109], stage1_13[110], stage1_13[111], stage1_13[112], stage1_13[113], stage1_13[114]},
      {stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29]},
      {stage2_17[4],stage2_16[21],stage2_15[33],stage2_14[34],stage2_13[41]}
   );
   gpc606_5 gpc666 (
      {stage1_13[115], stage1_13[116], stage1_13[117], stage1_13[118], stage1_13[119], stage1_13[120]},
      {stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35]},
      {stage2_17[5],stage2_16[22],stage2_15[34],stage2_14[35],stage2_13[42]}
   );
   gpc606_5 gpc667 (
      {stage1_13[121], stage1_13[122], stage1_13[123], stage1_13[124], stage1_13[125], stage1_13[126]},
      {stage1_15[36], stage1_15[37], stage1_15[38], stage1_15[39], stage1_15[40], stage1_15[41]},
      {stage2_17[6],stage2_16[23],stage2_15[35],stage2_14[36],stage2_13[43]}
   );
   gpc606_5 gpc668 (
      {stage1_13[127], stage1_13[128], stage1_13[129], stage1_13[130], stage1_13[131], stage1_13[132]},
      {stage1_15[42], stage1_15[43], stage1_15[44], stage1_15[45], stage1_15[46], stage1_15[47]},
      {stage2_17[7],stage2_16[24],stage2_15[36],stage2_14[37],stage2_13[44]}
   );
   gpc606_5 gpc669 (
      {stage1_14[102], stage1_14[103], stage1_14[104], stage1_14[105], stage1_14[106], stage1_14[107]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[8],stage2_16[25],stage2_15[37],stage2_14[38]}
   );
   gpc606_5 gpc670 (
      {stage1_14[108], stage1_14[109], stage1_14[110], stage1_14[111], stage1_14[112], stage1_14[113]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[9],stage2_16[26],stage2_15[38],stage2_14[39]}
   );
   gpc606_5 gpc671 (
      {stage1_14[114], stage1_14[115], stage1_14[116], stage1_14[117], stage1_14[118], stage1_14[119]},
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage2_18[2],stage2_17[10],stage2_16[27],stage2_15[39],stage2_14[40]}
   );
   gpc606_5 gpc672 (
      {stage1_14[120], stage1_14[121], stage1_14[122], stage1_14[123], stage1_14[124], stage1_14[125]},
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage2_18[3],stage2_17[11],stage2_16[28],stage2_15[40],stage2_14[41]}
   );
   gpc606_5 gpc673 (
      {stage1_14[126], stage1_14[127], stage1_14[128], stage1_14[129], stage1_14[130], stage1_14[131]},
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage2_18[4],stage2_17[12],stage2_16[29],stage2_15[41],stage2_14[42]}
   );
   gpc606_5 gpc674 (
      {stage1_14[132], stage1_14[133], stage1_14[134], stage1_14[135], stage1_14[136], stage1_14[137]},
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage2_18[5],stage2_17[13],stage2_16[30],stage2_15[42],stage2_14[43]}
   );
   gpc615_5 gpc675 (
      {stage1_14[138], stage1_14[139], stage1_14[140], stage1_14[141], stage1_14[142]},
      {stage1_15[48]},
      {stage1_16[36], stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41]},
      {stage2_18[6],stage2_17[14],stage2_16[31],stage2_15[43],stage2_14[44]}
   );
   gpc615_5 gpc676 (
      {stage1_14[143], stage1_14[144], stage1_14[145], stage1_14[146], stage1_14[147]},
      {stage1_15[49]},
      {stage1_16[42], stage1_16[43], stage1_16[44], stage1_16[45], stage1_16[46], stage1_16[47]},
      {stage2_18[7],stage2_17[15],stage2_16[32],stage2_15[44],stage2_14[45]}
   );
   gpc615_5 gpc677 (
      {stage1_14[148], stage1_14[149], stage1_14[150], stage1_14[151], stage1_14[152]},
      {stage1_15[50]},
      {stage1_16[48], stage1_16[49], stage1_16[50], stage1_16[51], stage1_16[52], stage1_16[53]},
      {stage2_18[8],stage2_17[16],stage2_16[33],stage2_15[45],stage2_14[46]}
   );
   gpc615_5 gpc678 (
      {stage1_15[51], stage1_15[52], stage1_15[53], stage1_15[54], stage1_15[55]},
      {stage1_16[54]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[9],stage2_17[17],stage2_16[34],stage2_15[46]}
   );
   gpc615_5 gpc679 (
      {stage1_15[56], stage1_15[57], stage1_15[58], stage1_15[59], stage1_15[60]},
      {stage1_16[55]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[10],stage2_17[18],stage2_16[35],stage2_15[47]}
   );
   gpc615_5 gpc680 (
      {stage1_15[61], stage1_15[62], stage1_15[63], stage1_15[64], stage1_15[65]},
      {stage1_16[56]},
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage2_19[2],stage2_18[11],stage2_17[19],stage2_16[36],stage2_15[48]}
   );
   gpc615_5 gpc681 (
      {stage1_15[66], stage1_15[67], stage1_15[68], stage1_15[69], stage1_15[70]},
      {stage1_16[57]},
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage2_19[3],stage2_18[12],stage2_17[20],stage2_16[37],stage2_15[49]}
   );
   gpc615_5 gpc682 (
      {stage1_15[71], stage1_15[72], stage1_15[73], stage1_15[74], stage1_15[75]},
      {stage1_16[58]},
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage2_19[4],stage2_18[13],stage2_17[21],stage2_16[38],stage2_15[50]}
   );
   gpc1_1 gpc683 (
      {stage1_0[48]},
      {stage2_0[8]}
   );
   gpc1_1 gpc684 (
      {stage1_1[96]},
      {stage2_1[24]}
   );
   gpc1_1 gpc685 (
      {stage1_1[97]},
      {stage2_1[25]}
   );
   gpc1_1 gpc686 (
      {stage1_2[82]},
      {stage2_2[30]}
   );
   gpc1_1 gpc687 (
      {stage1_2[83]},
      {stage2_2[31]}
   );
   gpc1_1 gpc688 (
      {stage1_2[84]},
      {stage2_2[32]}
   );
   gpc1_1 gpc689 (
      {stage1_2[85]},
      {stage2_2[33]}
   );
   gpc1_1 gpc690 (
      {stage1_2[86]},
      {stage2_2[34]}
   );
   gpc1_1 gpc691 (
      {stage1_2[87]},
      {stage2_2[35]}
   );
   gpc1_1 gpc692 (
      {stage1_2[88]},
      {stage2_2[36]}
   );
   gpc1_1 gpc693 (
      {stage1_2[89]},
      {stage2_2[37]}
   );
   gpc1_1 gpc694 (
      {stage1_2[90]},
      {stage2_2[38]}
   );
   gpc1_1 gpc695 (
      {stage1_2[91]},
      {stage2_2[39]}
   );
   gpc1_1 gpc696 (
      {stage1_2[92]},
      {stage2_2[40]}
   );
   gpc1_1 gpc697 (
      {stage1_2[93]},
      {stage2_2[41]}
   );
   gpc1_1 gpc698 (
      {stage1_2[94]},
      {stage2_2[42]}
   );
   gpc1_1 gpc699 (
      {stage1_2[95]},
      {stage2_2[43]}
   );
   gpc1_1 gpc700 (
      {stage1_2[96]},
      {stage2_2[44]}
   );
   gpc1_1 gpc701 (
      {stage1_2[97]},
      {stage2_2[45]}
   );
   gpc1_1 gpc702 (
      {stage1_3[113]},
      {stage2_3[33]}
   );
   gpc1_1 gpc703 (
      {stage1_5[104]},
      {stage2_5[54]}
   );
   gpc1_1 gpc704 (
      {stage1_6[102]},
      {stage2_6[38]}
   );
   gpc1_1 gpc705 (
      {stage1_6[103]},
      {stage2_6[39]}
   );
   gpc1_1 gpc706 (
      {stage1_7[92]},
      {stage2_7[36]}
   );
   gpc1_1 gpc707 (
      {stage1_7[93]},
      {stage2_7[37]}
   );
   gpc1_1 gpc708 (
      {stage1_7[94]},
      {stage2_7[38]}
   );
   gpc1_1 gpc709 (
      {stage1_7[95]},
      {stage2_7[39]}
   );
   gpc1_1 gpc710 (
      {stage1_7[96]},
      {stage2_7[40]}
   );
   gpc1_1 gpc711 (
      {stage1_7[97]},
      {stage2_7[41]}
   );
   gpc1_1 gpc712 (
      {stage1_7[98]},
      {stage2_7[42]}
   );
   gpc1_1 gpc713 (
      {stage1_7[99]},
      {stage2_7[43]}
   );
   gpc1_1 gpc714 (
      {stage1_7[100]},
      {stage2_7[44]}
   );
   gpc1_1 gpc715 (
      {stage1_7[101]},
      {stage2_7[45]}
   );
   gpc1_1 gpc716 (
      {stage1_7[102]},
      {stage2_7[46]}
   );
   gpc1_1 gpc717 (
      {stage1_7[103]},
      {stage2_7[47]}
   );
   gpc1_1 gpc718 (
      {stage1_7[104]},
      {stage2_7[48]}
   );
   gpc1_1 gpc719 (
      {stage1_7[105]},
      {stage2_7[49]}
   );
   gpc1_1 gpc720 (
      {stage1_7[106]},
      {stage2_7[50]}
   );
   gpc1_1 gpc721 (
      {stage1_7[107]},
      {stage2_7[51]}
   );
   gpc1_1 gpc722 (
      {stage1_7[108]},
      {stage2_7[52]}
   );
   gpc1_1 gpc723 (
      {stage1_7[109]},
      {stage2_7[53]}
   );
   gpc1_1 gpc724 (
      {stage1_7[110]},
      {stage2_7[54]}
   );
   gpc1_1 gpc725 (
      {stage1_7[111]},
      {stage2_7[55]}
   );
   gpc1_1 gpc726 (
      {stage1_7[112]},
      {stage2_7[56]}
   );
   gpc1_1 gpc727 (
      {stage1_7[113]},
      {stage2_7[57]}
   );
   gpc1_1 gpc728 (
      {stage1_7[114]},
      {stage2_7[58]}
   );
   gpc1_1 gpc729 (
      {stage1_9[115]},
      {stage2_9[47]}
   );
   gpc1_1 gpc730 (
      {stage1_14[153]},
      {stage2_14[47]}
   );
   gpc1_1 gpc731 (
      {stage1_14[154]},
      {stage2_14[48]}
   );
   gpc1_1 gpc732 (
      {stage1_14[155]},
      {stage2_14[49]}
   );
   gpc1_1 gpc733 (
      {stage1_14[156]},
      {stage2_14[50]}
   );
   gpc1_1 gpc734 (
      {stage1_16[59]},
      {stage2_16[39]}
   );
   gpc1_1 gpc735 (
      {stage1_16[60]},
      {stage2_16[40]}
   );
   gpc1_1 gpc736 (
      {stage1_16[61]},
      {stage2_16[41]}
   );
   gpc1_1 gpc737 (
      {stage1_16[62]},
      {stage2_16[42]}
   );
   gpc1_1 gpc738 (
      {stage1_16[63]},
      {stage2_16[43]}
   );
   gpc1_1 gpc739 (
      {stage1_16[64]},
      {stage2_16[44]}
   );
   gpc1_1 gpc740 (
      {stage1_16[65]},
      {stage2_16[45]}
   );
   gpc1_1 gpc741 (
      {stage1_16[66]},
      {stage2_16[46]}
   );
   gpc1_1 gpc742 (
      {stage1_16[67]},
      {stage2_16[47]}
   );
   gpc1_1 gpc743 (
      {stage1_17[30]},
      {stage2_17[22]}
   );
   gpc1_1 gpc744 (
      {stage1_17[31]},
      {stage2_17[23]}
   );
   gpc1_1 gpc745 (
      {stage1_17[32]},
      {stage2_17[24]}
   );
   gpc1_1 gpc746 (
      {stage1_17[33]},
      {stage2_17[25]}
   );
   gpc1_1 gpc747 (
      {stage1_17[34]},
      {stage2_17[26]}
   );
   gpc1_1 gpc748 (
      {stage1_17[35]},
      {stage2_17[27]}
   );
   gpc1_1 gpc749 (
      {stage1_17[36]},
      {stage2_17[28]}
   );
   gpc1_1 gpc750 (
      {stage1_17[37]},
      {stage2_17[29]}
   );
   gpc1_1 gpc751 (
      {stage1_17[38]},
      {stage2_17[30]}
   );
   gpc1_1 gpc752 (
      {stage1_17[39]},
      {stage2_17[31]}
   );
   gpc1_1 gpc753 (
      {stage1_17[40]},
      {stage2_17[32]}
   );
   gpc1_1 gpc754 (
      {stage1_17[41]},
      {stage2_17[33]}
   );
   gpc1163_5 gpc755 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc756 (
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5], stage2_3[6]},
      {stage3_5[0],stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1]}
   );
   gpc606_5 gpc757 (
      {stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15], stage2_1[16], stage2_1[17]},
      {stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11], stage2_3[12]},
      {stage3_5[1],stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2]}
   );
   gpc606_5 gpc758 (
      {stage2_1[18], stage2_1[19], stage2_1[20], stage2_1[21], stage2_1[22], stage2_1[23]},
      {stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17], stage2_3[18]},
      {stage3_5[2],stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3]}
   );
   gpc606_5 gpc759 (
      {stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[3],stage3_4[4],stage3_3[4],stage3_2[4]}
   );
   gpc606_5 gpc760 (
      {stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11], stage2_2[12]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[4],stage3_4[5],stage3_3[5],stage3_2[5]}
   );
   gpc606_5 gpc761 (
      {stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17], stage2_2[18]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage3_6[2],stage3_5[5],stage3_4[6],stage3_3[6],stage3_2[6]}
   );
   gpc615_5 gpc762 (
      {stage2_2[19], stage2_2[20], stage2_2[21], stage2_2[22], stage2_2[23]},
      {stage2_3[19]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage3_6[3],stage3_5[6],stage3_4[7],stage3_3[7],stage3_2[7]}
   );
   gpc615_5 gpc763 (
      {stage2_2[24], stage2_2[25], stage2_2[26], stage2_2[27], stage2_2[28]},
      {stage2_3[20]},
      {stage2_4[24], stage2_4[25], stage2_4[26], stage2_4[27], stage2_4[28], stage2_4[29]},
      {stage3_6[4],stage3_5[7],stage3_4[8],stage3_3[8],stage3_2[8]}
   );
   gpc615_5 gpc764 (
      {stage2_2[29], stage2_2[30], stage2_2[31], stage2_2[32], stage2_2[33]},
      {stage2_3[21]},
      {stage2_4[30], stage2_4[31], stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35]},
      {stage3_6[5],stage3_5[8],stage3_4[9],stage3_3[9],stage3_2[9]}
   );
   gpc615_5 gpc765 (
      {stage2_2[34], stage2_2[35], stage2_2[36], stage2_2[37], stage2_2[38]},
      {stage2_3[22]},
      {stage2_4[36], stage2_4[37], stage2_4[38], stage2_4[39], stage2_4[40], stage2_4[41]},
      {stage3_6[6],stage3_5[9],stage3_4[10],stage3_3[10],stage3_2[10]}
   );
   gpc615_5 gpc766 (
      {stage2_2[39], stage2_2[40], stage2_2[41], stage2_2[42], stage2_2[43]},
      {stage2_3[23]},
      {stage2_4[42], stage2_4[43], stage2_4[44], stage2_4[45], stage2_4[46], stage2_4[47]},
      {stage3_6[7],stage3_5[10],stage3_4[11],stage3_3[11],stage3_2[11]}
   );
   gpc615_5 gpc767 (
      {stage2_3[24], stage2_3[25], stage2_3[26], stage2_3[27], stage2_3[28]},
      {stage2_4[48]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[8],stage3_5[11],stage3_4[12],stage3_3[12]}
   );
   gpc615_5 gpc768 (
      {stage2_3[29], stage2_3[30], stage2_3[31], stage2_3[32], stage2_3[33]},
      {stage2_4[49]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[9],stage3_5[12],stage3_4[13],stage3_3[13]}
   );
   gpc7_3 gpc769 (
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17], stage2_5[18]},
      {stage3_7[2],stage3_6[10],stage3_5[13]}
   );
   gpc207_4 gpc770 (
      {stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23], stage2_5[24], stage2_5[25]},
      {stage2_7[0], stage2_7[1]},
      {stage3_8[0],stage3_7[3],stage3_6[11],stage3_5[14]}
   );
   gpc606_5 gpc771 (
      {stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29], stage2_5[30], stage2_5[31]},
      {stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5], stage2_7[6], stage2_7[7]},
      {stage3_9[0],stage3_8[1],stage3_7[4],stage3_6[12],stage3_5[15]}
   );
   gpc606_5 gpc772 (
      {stage2_5[32], stage2_5[33], stage2_5[34], stage2_5[35], stage2_5[36], stage2_5[37]},
      {stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11], stage2_7[12], stage2_7[13]},
      {stage3_9[1],stage3_8[2],stage3_7[5],stage3_6[13],stage3_5[16]}
   );
   gpc606_5 gpc773 (
      {stage2_5[38], stage2_5[39], stage2_5[40], stage2_5[41], stage2_5[42], stage2_5[43]},
      {stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17], stage2_7[18], stage2_7[19]},
      {stage3_9[2],stage3_8[3],stage3_7[6],stage3_6[14],stage3_5[17]}
   );
   gpc606_5 gpc774 (
      {stage2_5[44], stage2_5[45], stage2_5[46], stage2_5[47], stage2_5[48], stage2_5[49]},
      {stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23], stage2_7[24], stage2_7[25]},
      {stage3_9[3],stage3_8[4],stage3_7[7],stage3_6[15],stage3_5[18]}
   );
   gpc606_5 gpc775 (
      {stage2_5[50], stage2_5[51], stage2_5[52], stage2_5[53], stage2_5[54], 1'b0},
      {stage2_7[26], stage2_7[27], stage2_7[28], stage2_7[29], stage2_7[30], stage2_7[31]},
      {stage3_9[4],stage3_8[5],stage3_7[8],stage3_6[16],stage3_5[19]}
   );
   gpc615_5 gpc776 (
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4]},
      {stage2_7[32]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[5],stage3_8[6],stage3_7[9],stage3_6[17]}
   );
   gpc615_5 gpc777 (
      {stage2_6[5], stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9]},
      {stage2_7[33]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[6],stage3_8[7],stage3_7[10],stage3_6[18]}
   );
   gpc615_5 gpc778 (
      {stage2_6[10], stage2_6[11], stage2_6[12], stage2_6[13], stage2_6[14]},
      {stage2_7[34]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[7],stage3_8[8],stage3_7[11],stage3_6[19]}
   );
   gpc615_5 gpc779 (
      {stage2_6[15], stage2_6[16], stage2_6[17], stage2_6[18], stage2_6[19]},
      {stage2_7[35]},
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23]},
      {stage3_10[3],stage3_9[8],stage3_8[9],stage3_7[12],stage3_6[20]}
   );
   gpc615_5 gpc780 (
      {stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23], stage2_6[24]},
      {stage2_7[36]},
      {stage2_8[24], stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29]},
      {stage3_10[4],stage3_9[9],stage3_8[10],stage3_7[13],stage3_6[21]}
   );
   gpc615_5 gpc781 (
      {stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29]},
      {stage2_7[37]},
      {stage2_8[30], stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35]},
      {stage3_10[5],stage3_9[10],stage3_8[11],stage3_7[14],stage3_6[22]}
   );
   gpc615_5 gpc782 (
      {stage2_6[30], stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34]},
      {stage2_7[38]},
      {stage2_8[36], stage2_8[37], stage2_8[38], stage2_8[39], stage2_8[40], stage2_8[41]},
      {stage3_10[6],stage3_9[11],stage3_8[12],stage3_7[15],stage3_6[23]}
   );
   gpc615_5 gpc783 (
      {stage2_6[35], stage2_6[36], stage2_6[37], stage2_6[38], stage2_6[39]},
      {stage2_7[39]},
      {stage2_8[42], stage2_8[43], stage2_8[44], stage2_8[45], stage2_8[46], stage2_8[47]},
      {stage3_10[7],stage3_9[12],stage3_8[13],stage3_7[16],stage3_6[24]}
   );
   gpc606_5 gpc784 (
      {stage2_7[40], stage2_7[41], stage2_7[42], stage2_7[43], stage2_7[44], stage2_7[45]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[8],stage3_9[13],stage3_8[14],stage3_7[17]}
   );
   gpc615_5 gpc785 (
      {stage2_7[46], stage2_7[47], stage2_7[48], stage2_7[49], stage2_7[50]},
      {stage2_8[48]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[9],stage3_9[14],stage3_8[15],stage3_7[18]}
   );
   gpc615_5 gpc786 (
      {stage2_7[51], stage2_7[52], stage2_7[53], stage2_7[54], stage2_7[55]},
      {stage2_8[49]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[10],stage3_9[15],stage3_8[16],stage3_7[19]}
   );
   gpc606_5 gpc787 (
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[0],stage3_11[3],stage3_10[11],stage3_9[16]}
   );
   gpc606_5 gpc788 (
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage3_13[1],stage3_12[1],stage3_11[4],stage3_10[12],stage3_9[17]}
   );
   gpc606_5 gpc789 (
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17]},
      {stage3_13[2],stage3_12[2],stage3_11[5],stage3_10[13],stage3_9[18]}
   );
   gpc606_5 gpc790 (
      {stage2_9[36], stage2_9[37], stage2_9[38], stage2_9[39], stage2_9[40], stage2_9[41]},
      {stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23]},
      {stage3_13[3],stage3_12[3],stage3_11[6],stage3_10[14],stage3_9[19]}
   );
   gpc606_5 gpc791 (
      {stage2_9[42], stage2_9[43], stage2_9[44], stage2_9[45], stage2_9[46], stage2_9[47]},
      {stage2_11[24], stage2_11[25], stage2_11[26], stage2_11[27], stage2_11[28], stage2_11[29]},
      {stage3_13[4],stage3_12[4],stage3_11[7],stage3_10[15],stage3_9[20]}
   );
   gpc606_5 gpc792 (
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[5],stage3_12[5],stage3_11[8],stage3_10[16]}
   );
   gpc615_5 gpc793 (
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10]},
      {stage2_11[30]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[6],stage3_12[6],stage3_11[9],stage3_10[17]}
   );
   gpc615_5 gpc794 (
      {stage2_10[11], stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15]},
      {stage2_11[31]},
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage3_14[2],stage3_13[7],stage3_12[7],stage3_11[10],stage3_10[18]}
   );
   gpc615_5 gpc795 (
      {stage2_10[16], stage2_10[17], stage2_10[18], stage2_10[19], stage2_10[20]},
      {stage2_11[32]},
      {stage2_12[18], stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23]},
      {stage3_14[3],stage3_13[8],stage3_12[8],stage3_11[11],stage3_10[19]}
   );
   gpc615_5 gpc796 (
      {stage2_10[21], stage2_10[22], stage2_10[23], stage2_10[24], stage2_10[25]},
      {stage2_11[33]},
      {stage2_12[24], stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29]},
      {stage3_14[4],stage3_13[9],stage3_12[9],stage3_11[12],stage3_10[20]}
   );
   gpc615_5 gpc797 (
      {stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29], stage2_10[30]},
      {stage2_11[34]},
      {stage2_12[30], stage2_12[31], stage2_12[32], stage2_12[33], stage2_12[34], stage2_12[35]},
      {stage3_14[5],stage3_13[10],stage3_12[10],stage3_11[13],stage3_10[21]}
   );
   gpc615_5 gpc798 (
      {stage2_10[31], stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35]},
      {stage2_11[35]},
      {stage2_12[36], stage2_12[37], stage2_12[38], stage2_12[39], stage2_12[40], stage2_12[41]},
      {stage3_14[6],stage3_13[11],stage3_12[11],stage3_11[14],stage3_10[22]}
   );
   gpc606_5 gpc799 (
      {stage2_11[36], stage2_11[37], stage2_11[38], stage2_11[39], stage2_11[40], stage2_11[41]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[7],stage3_13[12],stage3_12[12],stage3_11[15]}
   );
   gpc606_5 gpc800 (
      {stage2_11[42], stage2_11[43], stage2_11[44], stage2_11[45], stage2_11[46], stage2_11[47]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[8],stage3_13[13],stage3_12[13],stage3_11[16]}
   );
   gpc606_5 gpc801 (
      {stage2_12[42], stage2_12[43], stage2_12[44], stage2_12[45], stage2_12[46], stage2_12[47]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[2],stage3_14[9],stage3_13[14],stage3_12[14]}
   );
   gpc606_5 gpc802 (
      {stage2_12[48], stage2_12[49], stage2_12[50], stage2_12[51], stage2_12[52], stage2_12[53]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[3],stage3_14[10],stage3_13[15],stage3_12[15]}
   );
   gpc117_4 gpc803 (
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17], stage2_13[18]},
      {stage2_14[12]},
      {stage2_15[0]},
      {stage3_16[2],stage3_15[4],stage3_14[11],stage3_13[16]}
   );
   gpc117_4 gpc804 (
      {stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23], stage2_13[24], stage2_13[25]},
      {stage2_14[13]},
      {stage2_15[1]},
      {stage3_16[3],stage3_15[5],stage3_14[12],stage3_13[17]}
   );
   gpc117_4 gpc805 (
      {stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29], stage2_13[30], stage2_13[31], stage2_13[32]},
      {stage2_14[14]},
      {stage2_15[2]},
      {stage3_16[4],stage3_15[6],stage3_14[13],stage3_13[18]}
   );
   gpc606_5 gpc806 (
      {stage2_13[33], stage2_13[34], stage2_13[35], stage2_13[36], stage2_13[37], stage2_13[38]},
      {stage2_15[3], stage2_15[4], stage2_15[5], stage2_15[6], stage2_15[7], stage2_15[8]},
      {stage3_17[0],stage3_16[5],stage3_15[7],stage3_14[14],stage3_13[19]}
   );
   gpc606_5 gpc807 (
      {stage2_13[39], stage2_13[40], stage2_13[41], stage2_13[42], stage2_13[43], stage2_13[44]},
      {stage2_15[9], stage2_15[10], stage2_15[11], stage2_15[12], stage2_15[13], stage2_15[14]},
      {stage3_17[1],stage3_16[6],stage3_15[8],stage3_14[15],stage3_13[20]}
   );
   gpc117_4 gpc808 (
      {stage2_14[15], stage2_14[16], stage2_14[17], stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21]},
      {stage2_15[15]},
      {stage2_16[0]},
      {stage3_17[2],stage3_16[7],stage3_15[9],stage3_14[16]}
   );
   gpc606_5 gpc809 (
      {stage2_14[22], stage2_14[23], stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27]},
      {stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5], stage2_16[6]},
      {stage3_18[0],stage3_17[3],stage3_16[8],stage3_15[10],stage3_14[17]}
   );
   gpc606_5 gpc810 (
      {stage2_14[28], stage2_14[29], stage2_14[30], stage2_14[31], stage2_14[32], stage2_14[33]},
      {stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11], stage2_16[12]},
      {stage3_18[1],stage3_17[4],stage3_16[9],stage3_15[11],stage3_14[18]}
   );
   gpc606_5 gpc811 (
      {stage2_14[34], stage2_14[35], stage2_14[36], stage2_14[37], stage2_14[38], stage2_14[39]},
      {stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17], stage2_16[18]},
      {stage3_18[2],stage3_17[5],stage3_16[10],stage3_15[12],stage3_14[19]}
   );
   gpc606_5 gpc812 (
      {stage2_14[40], stage2_14[41], stage2_14[42], stage2_14[43], stage2_14[44], stage2_14[45]},
      {stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23], stage2_16[24]},
      {stage3_18[3],stage3_17[6],stage3_16[11],stage3_15[13],stage3_14[20]}
   );
   gpc606_5 gpc813 (
      {stage2_14[46], stage2_14[47], stage2_14[48], stage2_14[49], stage2_14[50], 1'b0},
      {stage2_16[25], stage2_16[26], stage2_16[27], stage2_16[28], stage2_16[29], stage2_16[30]},
      {stage3_18[4],stage3_17[7],stage3_16[12],stage3_15[14],stage3_14[21]}
   );
   gpc606_5 gpc814 (
      {stage2_15[16], stage2_15[17], stage2_15[18], stage2_15[19], stage2_15[20], stage2_15[21]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[5],stage3_17[8],stage3_16[13],stage3_15[15]}
   );
   gpc606_5 gpc815 (
      {stage2_15[22], stage2_15[23], stage2_15[24], stage2_15[25], stage2_15[26], stage2_15[27]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[6],stage3_17[9],stage3_16[14],stage3_15[16]}
   );
   gpc606_5 gpc816 (
      {stage2_15[28], stage2_15[29], stage2_15[30], stage2_15[31], stage2_15[32], stage2_15[33]},
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage3_19[2],stage3_18[7],stage3_17[10],stage3_16[15],stage3_15[17]}
   );
   gpc606_5 gpc817 (
      {stage2_15[34], stage2_15[35], stage2_15[36], stage2_15[37], stage2_15[38], stage2_15[39]},
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23]},
      {stage3_19[3],stage3_18[8],stage3_17[11],stage3_16[16],stage3_15[18]}
   );
   gpc606_5 gpc818 (
      {stage2_15[40], stage2_15[41], stage2_15[42], stage2_15[43], stage2_15[44], stage2_15[45]},
      {stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29]},
      {stage3_19[4],stage3_18[9],stage3_17[12],stage3_16[17],stage3_15[19]}
   );
   gpc606_5 gpc819 (
      {stage2_16[31], stage2_16[32], stage2_16[33], stage2_16[34], stage2_16[35], stage2_16[36]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[5],stage3_18[10],stage3_17[13],stage3_16[18]}
   );
   gpc606_5 gpc820 (
      {stage2_16[37], stage2_16[38], stage2_16[39], stage2_16[40], stage2_16[41], stage2_16[42]},
      {stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10], stage2_18[11]},
      {stage3_20[1],stage3_19[6],stage3_18[11],stage3_17[14],stage3_16[19]}
   );
   gpc1_1 gpc821 (
      {stage2_0[3]},
      {stage3_0[1]}
   );
   gpc1_1 gpc822 (
      {stage2_0[4]},
      {stage3_0[2]}
   );
   gpc1_1 gpc823 (
      {stage2_0[5]},
      {stage3_0[3]}
   );
   gpc1_1 gpc824 (
      {stage2_0[6]},
      {stage3_0[4]}
   );
   gpc1_1 gpc825 (
      {stage2_0[7]},
      {stage3_0[5]}
   );
   gpc1_1 gpc826 (
      {stage2_0[8]},
      {stage3_0[6]}
   );
   gpc1_1 gpc827 (
      {stage2_1[24]},
      {stage3_1[4]}
   );
   gpc1_1 gpc828 (
      {stage2_1[25]},
      {stage3_1[5]}
   );
   gpc1_1 gpc829 (
      {stage2_2[44]},
      {stage3_2[12]}
   );
   gpc1_1 gpc830 (
      {stage2_2[45]},
      {stage3_2[13]}
   );
   gpc1_1 gpc831 (
      {stage2_7[56]},
      {stage3_7[20]}
   );
   gpc1_1 gpc832 (
      {stage2_7[57]},
      {stage3_7[21]}
   );
   gpc1_1 gpc833 (
      {stage2_7[58]},
      {stage3_7[22]}
   );
   gpc1_1 gpc834 (
      {stage2_12[54]},
      {stage3_12[16]}
   );
   gpc1_1 gpc835 (
      {stage2_12[55]},
      {stage3_12[17]}
   );
   gpc1_1 gpc836 (
      {stage2_12[56]},
      {stage3_12[18]}
   );
   gpc1_1 gpc837 (
      {stage2_12[57]},
      {stage3_12[19]}
   );
   gpc1_1 gpc838 (
      {stage2_12[58]},
      {stage3_12[20]}
   );
   gpc1_1 gpc839 (
      {stage2_12[59]},
      {stage3_12[21]}
   );
   gpc1_1 gpc840 (
      {stage2_12[60]},
      {stage3_12[22]}
   );
   gpc1_1 gpc841 (
      {stage2_15[46]},
      {stage3_15[20]}
   );
   gpc1_1 gpc842 (
      {stage2_15[47]},
      {stage3_15[21]}
   );
   gpc1_1 gpc843 (
      {stage2_15[48]},
      {stage3_15[22]}
   );
   gpc1_1 gpc844 (
      {stage2_15[49]},
      {stage3_15[23]}
   );
   gpc1_1 gpc845 (
      {stage2_15[50]},
      {stage3_15[24]}
   );
   gpc1_1 gpc846 (
      {stage2_16[43]},
      {stage3_16[20]}
   );
   gpc1_1 gpc847 (
      {stage2_16[44]},
      {stage3_16[21]}
   );
   gpc1_1 gpc848 (
      {stage2_16[45]},
      {stage3_16[22]}
   );
   gpc1_1 gpc849 (
      {stage2_16[46]},
      {stage3_16[23]}
   );
   gpc1_1 gpc850 (
      {stage2_16[47]},
      {stage3_16[24]}
   );
   gpc1_1 gpc851 (
      {stage2_17[30]},
      {stage3_17[15]}
   );
   gpc1_1 gpc852 (
      {stage2_17[31]},
      {stage3_17[16]}
   );
   gpc1_1 gpc853 (
      {stage2_17[32]},
      {stage3_17[17]}
   );
   gpc1_1 gpc854 (
      {stage2_17[33]},
      {stage3_17[18]}
   );
   gpc1_1 gpc855 (
      {stage2_18[12]},
      {stage3_18[12]}
   );
   gpc1_1 gpc856 (
      {stage2_18[13]},
      {stage3_18[13]}
   );
   gpc1_1 gpc857 (
      {stage2_19[0]},
      {stage3_19[7]}
   );
   gpc1_1 gpc858 (
      {stage2_19[1]},
      {stage3_19[8]}
   );
   gpc1_1 gpc859 (
      {stage2_19[2]},
      {stage3_19[9]}
   );
   gpc1_1 gpc860 (
      {stage2_19[3]},
      {stage3_19[10]}
   );
   gpc1_1 gpc861 (
      {stage2_19[4]},
      {stage3_19[11]}
   );
   gpc606_5 gpc862 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc606_5 gpc863 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc615_5 gpc864 (
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10]},
      {stage3_4[0]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[0],stage4_5[1],stage4_4[2],stage4_3[2]}
   );
   gpc606_5 gpc865 (
      {stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5], stage3_4[6]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[1],stage4_6[1],stage4_5[2],stage4_4[3]}
   );
   gpc606_5 gpc866 (
      {stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11], stage3_4[12]},
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10], stage3_6[11]},
      {stage4_8[1],stage4_7[2],stage4_6[2],stage4_5[3],stage4_4[4]}
   );
   gpc7_3 gpc867 (
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11], stage3_5[12]},
      {stage4_7[3],stage4_6[3],stage4_5[4]}
   );
   gpc7_3 gpc868 (
      {stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17], stage3_5[18], stage3_5[19]},
      {stage4_7[4],stage4_6[4],stage4_5[5]}
   );
   gpc207_4 gpc869 (
      {stage3_6[12], stage3_6[13], stage3_6[14], stage3_6[15], stage3_6[16], stage3_6[17], stage3_6[18]},
      {stage3_8[0], stage3_8[1]},
      {stage4_9[0],stage4_8[2],stage4_7[5],stage4_6[5]}
   );
   gpc615_5 gpc870 (
      {stage3_6[19], stage3_6[20], stage3_6[21], stage3_6[22], stage3_6[23]},
      {stage3_7[0]},
      {stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5], stage3_8[6], stage3_8[7]},
      {stage4_10[0],stage4_9[1],stage4_8[3],stage4_7[6],stage4_6[6]}
   );
   gpc615_5 gpc871 (
      {stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage3_8[8]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[1],stage4_9[2],stage4_8[4],stage4_7[7]}
   );
   gpc615_5 gpc872 (
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10]},
      {stage3_8[9]},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage4_11[1],stage4_10[2],stage4_9[3],stage4_8[5],stage4_7[8]}
   );
   gpc615_5 gpc873 (
      {stage3_7[11], stage3_7[12], stage3_7[13], stage3_7[14], stage3_7[15]},
      {stage3_8[10]},
      {stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15], stage3_9[16], stage3_9[17]},
      {stage4_11[2],stage4_10[3],stage4_9[4],stage4_8[6],stage4_7[9]}
   );
   gpc606_5 gpc874 (
      {stage3_8[11], stage3_8[12], stage3_8[13], stage3_8[14], stage3_8[15], stage3_8[16]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage4_12[0],stage4_11[3],stage4_10[4],stage4_9[5],stage4_8[7]}
   );
   gpc615_5 gpc875 (
      {stage3_10[6], stage3_10[7], stage3_10[8], stage3_10[9], stage3_10[10]},
      {stage3_11[0]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[0],stage4_12[1],stage4_11[4],stage4_10[5]}
   );
   gpc615_5 gpc876 (
      {stage3_10[11], stage3_10[12], stage3_10[13], stage3_10[14], stage3_10[15]},
      {stage3_11[1]},
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage4_14[1],stage4_13[1],stage4_12[2],stage4_11[5],stage4_10[6]}
   );
   gpc615_5 gpc877 (
      {stage3_10[16], stage3_10[17], stage3_10[18], stage3_10[19], stage3_10[20]},
      {stage3_11[2]},
      {stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15], stage3_12[16], stage3_12[17]},
      {stage4_14[2],stage4_13[2],stage4_12[3],stage4_11[6],stage4_10[7]}
   );
   gpc207_4 gpc878 (
      {stage3_11[3], stage3_11[4], stage3_11[5], stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9]},
      {stage3_13[0], stage3_13[1]},
      {stage4_14[3],stage4_13[3],stage4_12[4],stage4_11[7]}
   );
   gpc606_5 gpc879 (
      {stage3_11[10], stage3_11[11], stage3_11[12], stage3_11[13], stage3_11[14], stage3_11[15]},
      {stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5], stage3_13[6], stage3_13[7]},
      {stage4_15[0],stage4_14[4],stage4_13[4],stage4_12[5],stage4_11[8]}
   );
   gpc615_5 gpc880 (
      {stage3_12[18], stage3_12[19], stage3_12[20], stage3_12[21], stage3_12[22]},
      {stage3_13[8]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[1],stage4_14[5],stage4_13[5],stage4_12[6]}
   );
   gpc606_5 gpc881 (
      {stage3_13[9], stage3_13[10], stage3_13[11], stage3_13[12], stage3_13[13], stage3_13[14]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[1],stage4_15[2],stage4_14[6],stage4_13[6]}
   );
   gpc606_5 gpc882 (
      {stage3_13[15], stage3_13[16], stage3_13[17], stage3_13[18], stage3_13[19], stage3_13[20]},
      {stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11]},
      {stage4_17[1],stage4_16[2],stage4_15[3],stage4_14[7],stage4_13[7]}
   );
   gpc606_5 gpc883 (
      {stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10], stage3_14[11]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[2],stage4_16[3],stage4_15[4],stage4_14[8]}
   );
   gpc615_5 gpc884 (
      {stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15], stage3_14[16]},
      {stage3_15[12]},
      {stage3_16[6], stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11]},
      {stage4_18[1],stage4_17[3],stage4_16[4],stage4_15[5],stage4_14[9]}
   );
   gpc615_5 gpc885 (
      {stage3_14[17], stage3_14[18], stage3_14[19], stage3_14[20], stage3_14[21]},
      {stage3_15[13]},
      {stage3_16[12], stage3_16[13], stage3_16[14], stage3_16[15], stage3_16[16], stage3_16[17]},
      {stage4_18[2],stage4_17[4],stage4_16[5],stage4_15[6],stage4_14[10]}
   );
   gpc606_5 gpc886 (
      {stage3_15[14], stage3_15[15], stage3_15[16], stage3_15[17], stage3_15[18], stage3_15[19]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage4_19[0],stage4_18[3],stage4_17[5],stage4_16[6],stage4_15[7]}
   );
   gpc615_5 gpc887 (
      {stage3_15[20], stage3_15[21], stage3_15[22], stage3_15[23], stage3_15[24]},
      {stage3_16[18]},
      {stage3_17[6], stage3_17[7], stage3_17[8], stage3_17[9], stage3_17[10], stage3_17[11]},
      {stage4_19[1],stage4_18[4],stage4_17[6],stage4_16[7],stage4_15[8]}
   );
   gpc606_5 gpc888 (
      {stage3_16[19], stage3_16[20], stage3_16[21], stage3_16[22], stage3_16[23], stage3_16[24]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[2],stage4_18[5],stage4_17[7],stage4_16[8]}
   );
   gpc606_5 gpc889 (
      {stage3_17[12], stage3_17[13], stage3_17[14], stage3_17[15], stage3_17[16], stage3_17[17]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[1],stage4_19[3],stage4_18[6],stage4_17[8]}
   );
   gpc117_4 gpc890 (
      {stage3_18[6], stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11], stage3_18[12]},
      {stage3_19[6]},
      {stage3_20[0]},
      {stage4_21[1],stage4_20[2],stage4_19[4],stage4_18[7]}
   );
   gpc1_1 gpc891 (
      {stage3_0[6]},
      {stage4_0[1]}
   );
   gpc1_1 gpc892 (
      {stage3_2[6]},
      {stage4_2[2]}
   );
   gpc1_1 gpc893 (
      {stage3_2[7]},
      {stage4_2[3]}
   );
   gpc1_1 gpc894 (
      {stage3_2[8]},
      {stage4_2[4]}
   );
   gpc1_1 gpc895 (
      {stage3_2[9]},
      {stage4_2[5]}
   );
   gpc1_1 gpc896 (
      {stage3_2[10]},
      {stage4_2[6]}
   );
   gpc1_1 gpc897 (
      {stage3_2[11]},
      {stage4_2[7]}
   );
   gpc1_1 gpc898 (
      {stage3_2[12]},
      {stage4_2[8]}
   );
   gpc1_1 gpc899 (
      {stage3_2[13]},
      {stage4_2[9]}
   );
   gpc1_1 gpc900 (
      {stage3_3[11]},
      {stage4_3[3]}
   );
   gpc1_1 gpc901 (
      {stage3_3[12]},
      {stage4_3[4]}
   );
   gpc1_1 gpc902 (
      {stage3_3[13]},
      {stage4_3[5]}
   );
   gpc1_1 gpc903 (
      {stage3_4[13]},
      {stage4_4[5]}
   );
   gpc1_1 gpc904 (
      {stage3_6[24]},
      {stage4_6[7]}
   );
   gpc1_1 gpc905 (
      {stage3_7[16]},
      {stage4_7[10]}
   );
   gpc1_1 gpc906 (
      {stage3_7[17]},
      {stage4_7[11]}
   );
   gpc1_1 gpc907 (
      {stage3_7[18]},
      {stage4_7[12]}
   );
   gpc1_1 gpc908 (
      {stage3_7[19]},
      {stage4_7[13]}
   );
   gpc1_1 gpc909 (
      {stage3_7[20]},
      {stage4_7[14]}
   );
   gpc1_1 gpc910 (
      {stage3_7[21]},
      {stage4_7[15]}
   );
   gpc1_1 gpc911 (
      {stage3_7[22]},
      {stage4_7[16]}
   );
   gpc1_1 gpc912 (
      {stage3_9[18]},
      {stage4_9[6]}
   );
   gpc1_1 gpc913 (
      {stage3_9[19]},
      {stage4_9[7]}
   );
   gpc1_1 gpc914 (
      {stage3_9[20]},
      {stage4_9[8]}
   );
   gpc1_1 gpc915 (
      {stage3_10[21]},
      {stage4_10[8]}
   );
   gpc1_1 gpc916 (
      {stage3_10[22]},
      {stage4_10[9]}
   );
   gpc1_1 gpc917 (
      {stage3_11[16]},
      {stage4_11[9]}
   );
   gpc1_1 gpc918 (
      {stage3_17[18]},
      {stage4_17[9]}
   );
   gpc1_1 gpc919 (
      {stage3_18[13]},
      {stage4_18[8]}
   );
   gpc1_1 gpc920 (
      {stage3_19[7]},
      {stage4_19[5]}
   );
   gpc1_1 gpc921 (
      {stage3_19[8]},
      {stage4_19[6]}
   );
   gpc1_1 gpc922 (
      {stage3_19[9]},
      {stage4_19[7]}
   );
   gpc1_1 gpc923 (
      {stage3_19[10]},
      {stage4_19[8]}
   );
   gpc1_1 gpc924 (
      {stage3_19[11]},
      {stage4_19[9]}
   );
   gpc1_1 gpc925 (
      {stage3_20[1]},
      {stage4_20[3]}
   );
   gpc15_3 gpc926 (
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4]},
      {stage4_3[0]},
      {stage5_4[0],stage5_3[0],stage5_2[0]}
   );
   gpc615_5 gpc927 (
      {stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5]},
      {stage4_4[0]},
      {stage4_5[0], stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5]},
      {stage5_7[0],stage5_6[0],stage5_5[0],stage5_4[1],stage5_3[1]}
   );
   gpc1163_5 gpc928 (
      {stage4_6[0], stage4_6[1], stage4_6[2]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5]},
      {stage4_8[0]},
      {stage4_9[0]},
      {stage5_10[0],stage5_9[0],stage5_8[0],stage5_7[1],stage5_6[1]}
   );
   gpc1163_5 gpc929 (
      {stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage4_7[6], stage4_7[7], stage4_7[8], stage4_7[9], stage4_7[10], stage4_7[11]},
      {stage4_8[1]},
      {stage4_9[1]},
      {stage5_10[1],stage5_9[1],stage5_8[1],stage5_7[2],stage5_6[2]}
   );
   gpc615_5 gpc930 (
      {stage4_7[12], stage4_7[13], stage4_7[14], stage4_7[15], stage4_7[16]},
      {stage4_8[2]},
      {stage4_9[2], stage4_9[3], stage4_9[4], stage4_9[5], stage4_9[6], stage4_9[7]},
      {stage5_11[0],stage5_10[2],stage5_9[2],stage5_8[2],stage5_7[3]}
   );
   gpc615_5 gpc931 (
      {stage4_8[3], stage4_8[4], stage4_8[5], stage4_8[6], stage4_8[7]},
      {stage4_9[8]},
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5]},
      {stage5_12[0],stage5_11[1],stage5_10[3],stage5_9[3],stage5_8[3]}
   );
   gpc1163_5 gpc932 (
      {stage4_10[6], stage4_10[7], stage4_10[8]},
      {stage4_11[0], stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5]},
      {stage4_12[0]},
      {stage4_13[0]},
      {stage5_14[0],stage5_13[0],stage5_12[1],stage5_11[2],stage5_10[4]}
   );
   gpc1163_5 gpc933 (
      {stage4_11[6], stage4_11[7], stage4_11[8]},
      {stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5], stage4_12[6]},
      {stage4_13[1]},
      {stage4_14[0]},
      {stage5_15[0],stage5_14[1],stage5_13[1],stage5_12[2],stage5_11[3]}
   );
   gpc135_4 gpc934 (
      {stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5], stage4_13[6]},
      {stage4_14[1], stage4_14[2], stage4_14[3]},
      {stage4_15[0]},
      {stage5_16[0],stage5_15[1],stage5_14[2],stage5_13[2]}
   );
   gpc7_3 gpc935 (
      {stage4_14[4], stage4_14[5], stage4_14[6], stage4_14[7], stage4_14[8], stage4_14[9], stage4_14[10]},
      {stage5_16[1],stage5_15[2],stage5_14[3]}
   );
   gpc606_5 gpc936 (
      {stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5], stage4_15[6]},
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage5_19[0],stage5_18[0],stage5_17[0],stage5_16[2],stage5_15[3]}
   );
   gpc2135_5 gpc937 (
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4]},
      {stage4_17[6], stage4_17[7], stage4_17[8]},
      {stage4_18[0]},
      {stage4_19[0], stage4_19[1]},
      {stage5_20[0],stage5_19[1],stage5_18[1],stage5_17[1],stage5_16[3]}
   );
   gpc615_5 gpc938 (
      {stage4_16[5], stage4_16[6], stage4_16[7], stage4_16[8], 1'b0},
      {stage4_17[9]},
      {stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5], stage4_18[6]},
      {stage5_20[1],stage5_19[2],stage5_18[2],stage5_17[2],stage5_16[4]}
   );
   gpc1163_5 gpc939 (
      {stage4_18[7], stage4_18[8], 1'b0},
      {stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5], stage4_19[6], stage4_19[7]},
      {stage4_20[0]},
      {stage4_21[0]},
      {stage5_22[0],stage5_21[0],stage5_20[2],stage5_19[3],stage5_18[3]}
   );
   gpc1_1 gpc940 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc941 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc942 (
      {stage4_1[0]},
      {stage5_1[0]}
   );
   gpc1_1 gpc943 (
      {stage4_1[1]},
      {stage5_1[1]}
   );
   gpc1_1 gpc944 (
      {stage4_2[5]},
      {stage5_2[1]}
   );
   gpc1_1 gpc945 (
      {stage4_2[6]},
      {stage5_2[2]}
   );
   gpc1_1 gpc946 (
      {stage4_2[7]},
      {stage5_2[3]}
   );
   gpc1_1 gpc947 (
      {stage4_2[8]},
      {stage5_2[4]}
   );
   gpc1_1 gpc948 (
      {stage4_2[9]},
      {stage5_2[5]}
   );
   gpc1_1 gpc949 (
      {stage4_4[1]},
      {stage5_4[2]}
   );
   gpc1_1 gpc950 (
      {stage4_4[2]},
      {stage5_4[3]}
   );
   gpc1_1 gpc951 (
      {stage4_4[3]},
      {stage5_4[4]}
   );
   gpc1_1 gpc952 (
      {stage4_4[4]},
      {stage5_4[5]}
   );
   gpc1_1 gpc953 (
      {stage4_4[5]},
      {stage5_4[6]}
   );
   gpc1_1 gpc954 (
      {stage4_6[6]},
      {stage5_6[3]}
   );
   gpc1_1 gpc955 (
      {stage4_6[7]},
      {stage5_6[4]}
   );
   gpc1_1 gpc956 (
      {stage4_10[9]},
      {stage5_10[5]}
   );
   gpc1_1 gpc957 (
      {stage4_11[9]},
      {stage5_11[4]}
   );
   gpc1_1 gpc958 (
      {stage4_13[7]},
      {stage5_13[3]}
   );
   gpc1_1 gpc959 (
      {stage4_15[7]},
      {stage5_15[4]}
   );
   gpc1_1 gpc960 (
      {stage4_15[8]},
      {stage5_15[5]}
   );
   gpc1_1 gpc961 (
      {stage4_19[8]},
      {stage5_19[4]}
   );
   gpc1_1 gpc962 (
      {stage4_19[9]},
      {stage5_19[5]}
   );
   gpc1_1 gpc963 (
      {stage4_20[1]},
      {stage5_20[3]}
   );
   gpc1_1 gpc964 (
      {stage4_20[2]},
      {stage5_20[4]}
   );
   gpc1_1 gpc965 (
      {stage4_20[3]},
      {stage5_20[5]}
   );
   gpc1_1 gpc966 (
      {stage4_21[1]},
      {stage5_21[1]}
   );
   gpc615_5 gpc967 (
      {stage5_2[0], stage5_2[1], stage5_2[2], stage5_2[3], stage5_2[4]},
      {stage5_3[0]},
      {stage5_4[0], stage5_4[1], stage5_4[2], stage5_4[3], stage5_4[4], stage5_4[5]},
      {stage6_6[0],stage6_5[0],stage6_4[0],stage6_3[0],stage6_2[0]}
   );
   gpc135_4 gpc968 (
      {stage5_6[0], stage5_6[1], stage5_6[2], stage5_6[3], stage5_6[4]},
      {stage5_7[0], stage5_7[1], stage5_7[2]},
      {stage5_8[0]},
      {stage6_9[0],stage6_8[0],stage6_7[0],stage6_6[1]}
   );
   gpc1343_5 gpc969 (
      {stage5_8[1], stage5_8[2], stage5_8[3]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3]},
      {stage5_10[0], stage5_10[1], stage5_10[2]},
      {stage5_11[0]},
      {stage6_12[0],stage6_11[0],stage6_10[0],stage6_9[1],stage6_8[1]}
   );
   gpc1343_5 gpc970 (
      {stage5_10[3], stage5_10[4], stage5_10[5]},
      {stage5_11[1], stage5_11[2], stage5_11[3], stage5_11[4]},
      {stage5_12[0], stage5_12[1], stage5_12[2]},
      {stage5_13[0]},
      {stage6_14[0],stage6_13[0],stage6_12[1],stage6_11[1],stage6_10[1]}
   );
   gpc1343_5 gpc971 (
      {stage5_13[1], stage5_13[2], stage5_13[3]},
      {stage5_14[0], stage5_14[1], stage5_14[2], stage5_14[3]},
      {stage5_15[0], stage5_15[1], stage5_15[2]},
      {stage5_16[0]},
      {stage6_17[0],stage6_16[0],stage6_15[0],stage6_14[1],stage6_13[1]}
   );
   gpc1343_5 gpc972 (
      {stage5_15[3], stage5_15[4], stage5_15[5]},
      {stage5_16[1], stage5_16[2], stage5_16[3], stage5_16[4]},
      {stage5_17[0], stage5_17[1], stage5_17[2]},
      {stage5_18[0]},
      {stage6_19[0],stage6_18[0],stage6_17[1],stage6_16[1],stage6_15[1]}
   );
   gpc1163_5 gpc973 (
      {stage5_18[1], stage5_18[2], stage5_18[3]},
      {stage5_19[0], stage5_19[1], stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5]},
      {stage5_20[0]},
      {stage5_21[0]},
      {stage6_22[0],stage6_21[0],stage6_20[0],stage6_19[1],stage6_18[1]}
   );
   gpc135_4 gpc974 (
      {stage5_20[1], stage5_20[2], stage5_20[3], stage5_20[4], stage5_20[5]},
      {stage5_21[1], 1'b0, 1'b0},
      {stage5_22[0]},
      {stage6_23[0],stage6_22[1],stage6_21[1],stage6_20[1]}
   );
   gpc1_1 gpc975 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc976 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc977 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc978 (
      {stage5_1[1]},
      {stage6_1[1]}
   );
   gpc1_1 gpc979 (
      {stage5_2[5]},
      {stage6_2[1]}
   );
   gpc1_1 gpc980 (
      {stage5_3[1]},
      {stage6_3[1]}
   );
   gpc1_1 gpc981 (
      {stage5_4[6]},
      {stage6_4[1]}
   );
   gpc1_1 gpc982 (
      {stage5_5[0]},
      {stage6_5[1]}
   );
   gpc1_1 gpc983 (
      {stage5_7[3]},
      {stage6_7[1]}
   );
endmodule

module testbench();
    reg [255:0] src0;
    reg [255:0] src1;
    reg [255:0] src2;
    reg [255:0] src3;
    reg [255:0] src4;
    reg [255:0] src5;
    reg [255:0] src6;
    reg [255:0] src7;
    reg [255:0] src8;
    reg [255:0] src9;
    reg [255:0] src10;
    reg [255:0] src11;
    reg [255:0] src12;
    reg [255:0] src13;
    reg [255:0] src14;
    reg [255:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [23:0] srcsum;
    wire [23:0] dstsum;
    wire test;
    compressor_CLA256_16 compressor_CLA256_16(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161] + src12[162] + src12[163] + src12[164] + src12[165] + src12[166] + src12[167] + src12[168] + src12[169] + src12[170] + src12[171] + src12[172] + src12[173] + src12[174] + src12[175] + src12[176] + src12[177] + src12[178] + src12[179] + src12[180] + src12[181] + src12[182] + src12[183] + src12[184] + src12[185] + src12[186] + src12[187] + src12[188] + src12[189] + src12[190] + src12[191] + src12[192] + src12[193] + src12[194] + src12[195] + src12[196] + src12[197] + src12[198] + src12[199] + src12[200] + src12[201] + src12[202] + src12[203] + src12[204] + src12[205] + src12[206] + src12[207] + src12[208] + src12[209] + src12[210] + src12[211] + src12[212] + src12[213] + src12[214] + src12[215] + src12[216] + src12[217] + src12[218] + src12[219] + src12[220] + src12[221] + src12[222] + src12[223] + src12[224] + src12[225] + src12[226] + src12[227] + src12[228] + src12[229] + src12[230] + src12[231] + src12[232] + src12[233] + src12[234] + src12[235] + src12[236] + src12[237] + src12[238] + src12[239] + src12[240] + src12[241] + src12[242] + src12[243] + src12[244] + src12[245] + src12[246] + src12[247] + src12[248] + src12[249] + src12[250] + src12[251] + src12[252] + src12[253] + src12[254] + src12[255])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161] + src13[162] + src13[163] + src13[164] + src13[165] + src13[166] + src13[167] + src13[168] + src13[169] + src13[170] + src13[171] + src13[172] + src13[173] + src13[174] + src13[175] + src13[176] + src13[177] + src13[178] + src13[179] + src13[180] + src13[181] + src13[182] + src13[183] + src13[184] + src13[185] + src13[186] + src13[187] + src13[188] + src13[189] + src13[190] + src13[191] + src13[192] + src13[193] + src13[194] + src13[195] + src13[196] + src13[197] + src13[198] + src13[199] + src13[200] + src13[201] + src13[202] + src13[203] + src13[204] + src13[205] + src13[206] + src13[207] + src13[208] + src13[209] + src13[210] + src13[211] + src13[212] + src13[213] + src13[214] + src13[215] + src13[216] + src13[217] + src13[218] + src13[219] + src13[220] + src13[221] + src13[222] + src13[223] + src13[224] + src13[225] + src13[226] + src13[227] + src13[228] + src13[229] + src13[230] + src13[231] + src13[232] + src13[233] + src13[234] + src13[235] + src13[236] + src13[237] + src13[238] + src13[239] + src13[240] + src13[241] + src13[242] + src13[243] + src13[244] + src13[245] + src13[246] + src13[247] + src13[248] + src13[249] + src13[250] + src13[251] + src13[252] + src13[253] + src13[254] + src13[255])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161] + src14[162] + src14[163] + src14[164] + src14[165] + src14[166] + src14[167] + src14[168] + src14[169] + src14[170] + src14[171] + src14[172] + src14[173] + src14[174] + src14[175] + src14[176] + src14[177] + src14[178] + src14[179] + src14[180] + src14[181] + src14[182] + src14[183] + src14[184] + src14[185] + src14[186] + src14[187] + src14[188] + src14[189] + src14[190] + src14[191] + src14[192] + src14[193] + src14[194] + src14[195] + src14[196] + src14[197] + src14[198] + src14[199] + src14[200] + src14[201] + src14[202] + src14[203] + src14[204] + src14[205] + src14[206] + src14[207] + src14[208] + src14[209] + src14[210] + src14[211] + src14[212] + src14[213] + src14[214] + src14[215] + src14[216] + src14[217] + src14[218] + src14[219] + src14[220] + src14[221] + src14[222] + src14[223] + src14[224] + src14[225] + src14[226] + src14[227] + src14[228] + src14[229] + src14[230] + src14[231] + src14[232] + src14[233] + src14[234] + src14[235] + src14[236] + src14[237] + src14[238] + src14[239] + src14[240] + src14[241] + src14[242] + src14[243] + src14[244] + src14[245] + src14[246] + src14[247] + src14[248] + src14[249] + src14[250] + src14[251] + src14[252] + src14[253] + src14[254] + src14[255])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161] + src15[162] + src15[163] + src15[164] + src15[165] + src15[166] + src15[167] + src15[168] + src15[169] + src15[170] + src15[171] + src15[172] + src15[173] + src15[174] + src15[175] + src15[176] + src15[177] + src15[178] + src15[179] + src15[180] + src15[181] + src15[182] + src15[183] + src15[184] + src15[185] + src15[186] + src15[187] + src15[188] + src15[189] + src15[190] + src15[191] + src15[192] + src15[193] + src15[194] + src15[195] + src15[196] + src15[197] + src15[198] + src15[199] + src15[200] + src15[201] + src15[202] + src15[203] + src15[204] + src15[205] + src15[206] + src15[207] + src15[208] + src15[209] + src15[210] + src15[211] + src15[212] + src15[213] + src15[214] + src15[215] + src15[216] + src15[217] + src15[218] + src15[219] + src15[220] + src15[221] + src15[222] + src15[223] + src15[224] + src15[225] + src15[226] + src15[227] + src15[228] + src15[229] + src15[230] + src15[231] + src15[232] + src15[233] + src15[234] + src15[235] + src15[236] + src15[237] + src15[238] + src15[239] + src15[240] + src15[241] + src15[242] + src15[243] + src15[244] + src15[245] + src15[246] + src15[247] + src15[248] + src15[249] + src15[250] + src15[251] + src15[252] + src15[253] + src15[254] + src15[255])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hafae780abcb47fe4bba49a6f898593ad17cc69dd09f5b8be323b9023d1cf47c8ce9be86b409c57e3b6a5615e59e0568b0ffb9f47c6e146789908349f1e3538c988199ef1e63ea911e9d37cae2aa5c8b1c923e9b3474fef0a570898b928026c5e89cca94c21cfdc49347394cbeef657d2585d8ca1198c3644d8bd33ac9b9a52b6f6863888b00c45549acce9fcb5c4d12e99644707eaf695d5143643c8857b9b052379c4466b2e0b590554f693a7f5f59489f2fb2685f51ebf9f40f9a5378ed84072116a000d98ad7019759b7886b7eb279bb9f2fa5d0164754d87df712946a62fa65a306eada53e74b0242a6e0030c7f31acda66500c10bf849d07721d24aa538f0682bc904e90c1bb7f2330119bd70accff0d7d641f20b0872ac9b5c5d04fb0cd3a60181e3ca131959ba9252067551c54abf0f2f8f44bfe2ab9fe80acde77165bc6cdcde1b92ec283da963027fb2f500b79c995808983ee48f4a81cee5feffe4444cdd047d083eb8ae510d15d168d8141341dc851b75138cc9e54657e42025122dee93bfd618600c8f21d44cc0b91d76aaf13d315b3a9c8f0b0fa7a1342dd7316bd6299fe6d85315968a9d8fc967ce0b18707aea587ba4233e302286bf33c87a6ee44bbf8e69e0d90fce9a82d59c414c1fed4cde2569b4a6f4c28aade426b54fb160fac883da213f8758196281b91577f614035e40311c7db92b17db06c88c87;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h4f160a3d1d81230520ff6e8f3510cf8d9ccd7907cff4f255d5aaeaa522a424695c83e29e996528f9b22f51cc73cbe5a9e307625268db2b961666e6a6641943b92bc0cbfc74c2ce3083a80e88aae214a2228d06bea4c0602cb51a2a274a8330554fb592d86ff6efbb0b1e3bd12fde61dcf96b00c975a16eeb0b39d3f54c062f10957c1d4709939ee4aba0ae3432480224de003e31992e6b7f98d639301d3eec0f595b804b345f52272cc4b8cc48168cff531169e6e790483797c5e76e05dd9e93a6d57712cfa73bf6b16756f194cdc0fd04e48fd3330b69eab318e144c64dee17e12187aef17264099cb6c9bf72a03f85e92948db9956504770f7d5682c78d53b26a922072193b1b624c341e0f94ae8ee85c0f869fd6b5b843282c2118211e90a2c9fc708743c15df4c1207c9d53145ee3965101aff739e1f4fa273140510e28a71a6d20a88f33c9f235c82f7ba4ac9b3443a874f831fc302ffd9f874a68c093def812d540912742e25a50ee8b7dbeecbea982e902ff2c21f179e2cd8f7a6ef85a06b2b159ff1e0627dd1b64864ba861333c21fde8ae83229e548be972a3073007df3737aea54dd072fa9401280016ff0b19e6d10b50e3df12dcde68316c68471a6d3ac5e1b0a1f7934fafbe9a5876f81263aa7df21662493ad92e677456e487bc11362c51c76ae42947341e93e5c60eeafd4875a2ef57f1d850903a52f06abb9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hfb3cbad6081c4d92ec430625a2438ab73db8624f88fd601b92487608d34e30ecaa1b74631f5eb5f6d23809a64c6c2b1311892cebde6d44fa2373416bc74b39fadd5e44b9697b0650287d77cc3a6108038f5e461de6e56eeb7fba5a65c86ff1c15416bed5b819234acbec07dec32e2a29c404644ddfa57cd9dbe7a5165d56dc3185ffe77dc85e5391f0f15aff8202018073b82f114a779da2add0ff37cc03e631ff0f2dd4f1882cf179013b6e93c81034c48999593a60a50f029f85601c05fa24246765631edec608fd8b5552047a5ac836e55d53821d839a8da7b014b5c188035bd671a0d289d9e16bfa90202709731b20204feef66f0740d79c0ad10c347d3f5025d647dee6e48b09c191af64fda601f6f2979288d512517e1ee0b602027563434a1e27ffb130b3831ee0f9282a96149c332e9f1474dc20071a082b870fc92d8776b2b23030febafd336c339495de6c2b994748989a1d2edb410a3705b065ceabb1a0c1bdd44d9772921e2cf49603db9694592d09d7e150fa4d58a2417dd6c4e71cbc0abbb40ccf1b9634fac5a0b82406552c559a1d7b2002e0069b06b78e7f4694511d26f4f6e6a5b043d7e8dc3e4eebe6c219ad260b89838a6e03454712d2f2d551c55597600924c693a6cff3b5159bc81ac563beef9a680c55e464d00ba1b7e30439606813957d38af4e4de8be52329c9cad3462a76baf26bec6512df01c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3bd3d642246856e477d5c46b53d8ca1dcb2b7ffb8c035018afc8fa2be3322226efa196cf39b6138f67d297a38455ca1287ededf08df36fb7660ff11ee593a81b3599bc745f084fcf72ce9afc3e1af53262c8a9c60050d83c59553ce374a785e360ca09b77e2c21f23f04d309ccacd2650bb946c96957a1e6cb2dab693da10f235a21776125842bfd51fa72f878b9266e09bef3a878513561d937b279de592df0226163e80e826b125bdfc9272e4490676b0755a8243669edbbb2f89b3e26c9e236b388b8e4eae8e4785a4336a414d379846ec9ed67abf3fd563b9100721007b9abeaba218d57183c9969b0744bac1c93020c221455fdd7ca430726c6591c0c3896dbf945541557cc154f5e5f45b8fa038322279ed9936a3e0ee23305e213705cc173ed75452f039f90c14b6e6de8f953f7d5421124586c2906390b214f6f8f572ed3ea1d8564ab05414364090a5f144973ac05d6c7cf6a264f563bf51737bc62c76bda5aef4393d8e13433bcffdd3bdac05d84d5a7a971a313b48ec20542a8f5296e9e69b68b6003ccf3c2afe540098f57ed0f5f0c1c25e0c04ebb0bd1ed8f339b8ee416f4ca5ee7e24edc1a7a8b2e7de5a1459ae4d0f06cad922cd00def535bd2e9b452664e27907cab9abe4adee4f9c709a4823e822e526477c09fce09a77f76435cf72504c8ec1521f116170ef77d175d3d66c274451c808b3ee6f61141f4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf4fddad5efba5fe0847a1be09da88424dcb71477c6fb4fcbe17cb66d591aa5263c40c5192cd99a4ccea67076e3333a74666021fadfd13f335b45faee72ee35fc55119fc0d2d44dab523d904eef553aeff0c42fab3ed603d80a2c325c716ee5d2693540991f4289c1d5e8325cc4c48911718210fb9c9d7b0333d3b7aa4acc110161ae390c6250cc512138687568e8bcfb5b5448dfc1ce79023c9a1debb546cb32745b38da5156cc717cb44351a5b8eacb9b9f6ffba0a74731ce45c6af37da4dcc5a859384a65a8efb28873928f256bdc57dd38a27e4e3529bab2b568db857c4aea08be6406ef6b03ed3569e5106d55b4d1c0f7e11f13b9305e27be4ff39037142b9bd458a10be61d12a0513ac6daf12bc3467051555cfe32181b5ba574e3b865b739e7eef3b98ee0d4c21c8c4ae9b824ef082a0f687dbef8edd096fd2e83f6cf2f30212c5d0c6603e4841ac2da020584f84f8c5c9835293fc9d0e08501227584587d7de88a25409eaf11ee9423f5e188b707c38ffac3d535f85671ddf01228f33359e914b3870f4a6b1107dba19b11bd2518bdc30a0e7a64f57b29de4ce087911cbe846d87e4493d9aba1e1694d0d343170e344429fae9cc21bd9789a3019265dd1a7809697fc11272e8dfcc95f37a48b4aae4f7dd780d6c3a543e5d91f4a12f3aad207dd4c570678b8500f25f0bb35c6edb052780fb25109bac17c570d02bb1c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h506ddc646947bab64607b76261e54becda328224de85c43fad2c2d5ebf71a374c5fc52e80e3ca9379a9188ef1e07f8947f4ed38ed178c60fcb6a10028eb7ddac895f76843a6d7dce2b3ca8aa824e16304b095cb21ab836a7bfede782145c3bbd270a60e601599fe6fbd7b730884472e2ba3e240268a7323461d3d4d3416d538c0fdee2bcd63c6bdd963150b2e72d4b6408b81c184d37b16e5cf4004a3d782854b1e99188b19cdfefef7c953e55a258a2e4bf8962d3be08c925d14adf40e30a4d65956346ab9215505fa870c80f334ac8d4f6a5d8df01e520e22c80fa9bc334c198dfff0c7844c86fbab5b6628a33760c16807c660f58804b70cc6878ccc9808648183b7dd1a00ed4cc633f660a01bd93143b7d58a830e31f27f2b8b6df60613558a628eb0cc816b37c78da40bd6159ed6cf24db7d581046a7f22a2428ea5e64857c54e720c4957d4bc0fd11333c568dbf4745808c50fe039acdd6d1a4d2a8e58da1022b6728a35a51a49e2f112728cd703228b288a735f0ce59ba804af1547d470daeddfbd79f393fdbe1ef71f8720090310286caee451464639f850f745f5c621be5918d9d5e183674bcb844339813d9ede95123ad6a8a27384156e8dc403d1367a1ff967018ece67458ca3c77682b94e02900b409deed1fe58ca4d5dcec2081e4c8209d7de6a6c640d96e5801c3bae56b94d04e37305ad1dcf20c41d51c86f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h2b26e0fcdc01150656ad5f746ff8491fdc9cec3b7f307a48ae7b32a0474bcaae5f81ccf565de8119b78eb48bd283bc300cd15b14634ad61236bdf5972e64241d7063a0d6925dd563256aac9dfd9525cb204fa65a8d0ff41b17302ef5610ad8fd2e17445300eb17eff4068ffc28b817591cf57777626518bc370e3e397d77bc456b364d75448f30b6dbf4852aaf94086b9fab6c3e7661b5a6289e22d2d3f016e1481c24e5105b4834ba1ca941dd826b76df6c474c7a0cca70b84a22b05090f0c4c7b5824dd5d352dc72359b05f07f17bdd2924554d9c12aa6d5c9a0d1de470aaceedcfb378adbb67471d4cfa26ad07268943c54da23ff9d232a723530cddcf52516a80e8da4d20cf497ae14c31dfd500f8e3c5c7599e37312f1a952e40de6e4e3607a619343b9ed303365c6ca5b6c9a7593ef42ad67f323900e208d117dec99a5b61a07d96b80e5470abb54513e7e738190ce9c39d59935fbbb766a3e5167205db468dc94f3783e91f33ab5d1c8dc3ed93e6f982fee6ac1eb2e70cdcad0227cf4d2ad5c7f0172a10e10082e9f158bd04c6428812efa91fa4a119053f3a656c388e62f09434924b2fcb643b316c4241cb9abe11494d39fb3a300d5d5e63450c1cc6441a6a4f7414eca4f5e7879029f2d829a48e41f1f118200f107c2e281cb6ff495d9bb3d16abce442cfc28a8ae23c5de69026d14df66d40c4c4bc73ed9e9f362;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hcdd08dd02ff25b8966b6f7420ca757895c4278d727b2d30236ceb77cbf7dcc1adace7dce96ed090e8fe0df6f2570757c02d6c31b1b22ec5db850faadbd1ce22ec2edcbc8eba9931ae6f0cc80408c9eb5e15698e23c7b942d41f418177fb8abc728eb3689a67ebc4accdfb3d41c7d337cd630bed92e42c74e4d6eac24514c571c80aa2db2f066ee24fb5ba4de03aa243a572b81a593bd2ed64d13eba5cdc38a28e298ad9572f93f2936ce0020899254ee421884157ed948c11e8dc1df9573eecfa21d73ec2fdccd8430a09cb0e0c95f9a8428895943822b2acc9609d54b9cdef65ac7bcc62cd82268f38d4df0efaad32f921293cfbb34d76157fc559d078b3967772d235ace2c3867f1bacdcd0d4d433b4dc528d90254948abb63802688359b44bf7b55c60d00767d98c115522806ca891f01db35ce9c95c7bc272de7b01a025ac2bac85dfab4f205d0e49a306d1146c5be7aeeefcfbdde08b31e18e18f6ea41331c239c2e3afc0dd5e1ae913d5707761412204f1ae1754b09ea111c2a5f0f93f6f313bc8858622cda5261f2d7d43d60fc5273dcb274080e3f3fdef17300578fbfee19a44c9c5f22d93d483911653fedadba65198abd35ca90944d00833fc0acd560d8c6312815b59f28184e083f56f452d7867fb197e01d0ef9591d198b6dbf91d961043c1230b4332847991b229942cbfb87e5e1a7c91627ba32fc11c94d722;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hbcb67593cc00d7bd5c3cb029d04d79272a1861678387dff48be35fa43e4a303651e2d9015a3df55c51cc76e9627132bf0d2877150b2fe96264d54b828ac81615af14f5c96f5d8d29ea6680bb184f8515b840322d56a935ec6b7b12d091bfa401f8009c506d4169073176661ac73816a92c0ba2267ae669e30a98ad8d6006cf7db2d15f3ea04ece15b9868483b83685db9b208bc7647ff3ccc42d66eddbae2da3f1a9a9dd24545b63812e15695ee8016ebff8dbdc8d22c4ffb02ec84a62460fa548ee6181553610999c4bc35a9bbee1dded2748c0e48f5ad2162a08fabe221555c52d044cc88bc7676f2f0f9cbd362bf436dc2a0e6a900d4bffe1ae84629716d311e9f1e780b2fada5d7c073ba5ebf91ba4df1d548465c91d5a7e25051c3db622b1841477d19ff82dfae4763858f3bcb1fc4e9ef5cc5319dcfe317ea5a8580a7c320bb6be4068fdc0127ecd308af02b405f6a8c480b93243c4dcc72fadd6c106907e08ec067ce6e353c502d4b49e942752cf261c2cc57f51c798309ea76eed211d98f67b5dbaaf8aef9bd33a59ec037bebca23e9a4965f9265f260b770f7a264e4f063227f3e8db24580bb0bc493255e3aa42a77c99e10fb1a004405af12a75ead675bdb65df566c619533df2948a2294568da6a81cc9b7f13908dc01f20110ff55270ef9de319d7d69918b45836a0fa88d5701d969f4d7856c1f98d3c50b5713;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h27917ef65b3380f4bac4ada14ac492ae659782fea8da6835636d1179d3335a0c75df441be990c884e34cd39417270ed8ad955034dd23544431e318245879e6e7a722258c549e7c3b74345fe543ca966e0e57a213437624bfb5a282a7cc3b52584add666b00bd49a44aa2e35c870a66221e590e04edd28a2a1868a963de8f7ed7da5af2c453322305b0f139431043a3044437548ce3cdf22250f02b2806fb45b96603607aafbc41a00fab4daa979f2a26b21d92d0448b230c2e2c00e6525f5886c1695f7571d68344b28c04380b582408183499b77bbe9bcf7cb5ccd3725b485372e9bb4770ed61d0ecb525222d337da67250da69a3069524cc87f0114da0b36ebe8b1d942141b300509aa587e93b8e6ac5cb90edeed431e46ed4f87fc10f4d973a145ca19bfa7aba7e5816704867d95d09703718dc5e3a00b69b99218ada8b8febf8da2fdf7448cb7faf4c83d7e76884043676808018b75cb068fd8e38a34544d5345951dacd2b8d99df609ca2b58d6aac95bad91954b3f972b12d5e5275740ba4e9daf45996a2b835c4278f5c3bbc093aa8a3f487fc910a25e68fe90eeadcb463ad09507fcced598e731a6206a70d6c26fce8b897a52bc6bbf69935ddab8ea7bac69687eaba0c1a0817eaa98970608f7ebbaaecf940881ef213cd5e29e3d7a218c708a1789f0f838bdc32e94904d40bad79dd31b5212ddf0145237f19a64e11;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hdc16b1dc3af33f0a6ecc38838b7acf4791c37830dff65c03fa4c09dd7b31f50f043826650d20309f323d7ac652d717c9132ab8e832a9f7747485585288ec62174a500febcc1fe045651f6ff2179e963495a7483930eeeee291fb72b4dadeb790136271205a5734a6ca9f390fdc07b11da6b7cb9cd2bccc693446326bd1ba3b6746f234fc66eb5ed4d337dde93ea8e662bf78f59e8e75fd4a7a371b876dc153f354d6208cfa75f8d09f7b3fd07513d6b7e8a1a85d578d2acbf724db05bb53fb3b07dbd336936ded82aef2d5569a6b93f5834db0a115f34db7bc173dfea7e25e229f618cede052f75d214affdf4b54626e86918a8d7c75847829ef2bbfbb26f3d2fc8e3e0fbc0f7b2376625e8cab72f16a833f318494faede1bff3502da0e0665b93c90009ab7c37e5af9aac8360f082bcbb199e295a0dd455862876fec553b80f6a1ef6314193200b329da63fd245f8f6639ad888432fbf5b90257287b3f47b1aadd48ea4765a2b309f466015ed623b9d582f9723c7d6b7c42e197876927a5a6ca1f9e6080b0ea839575eb65403adb0be2fe475b868d55f40c3e7a13bd380efac99375cb8ee04488fc97ec45743af3403b487e811f39c33850b253be410e68ee2d902fad5c5f4126cb45a8230976e2a782c418e2a297a72a9b01d8a5f4b224c900972b0dd856ca0134249d0c6606c7c5be0e2903a5b98846befde8970241805ca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h1453fd54268009b07873bd574b8d26a3c62cb57f069b244a3e3cd092ceb8209b3bd962584dc330427eab1cc6a5c722ba019874f9206a2dc101f0cc587e7d353012a114f027a81cfbbd6bf40019fdeea9cbacbaa4d2fa67f781834fa9e3cb3df4a307c563d461b0970e8ec4e43729692d3a96628ac260a735fe5f20b5dbc9c7d4c8d2ebfcc44b4044a523b58490659751cc0851d2755c1f33a2dbd3913f3755ccd2a4c200ac8035862b3c23e1d76ee991eb287d95abd5f577634587fdf4d599b83a51afc06fb31ee46831604aca963bb11e0dda787a4face4f89b05304d547eae7021e5d878b043bec22cfbaa8087bcafe7f1e93db97e471ac5d059970d28b09bca341ed31b1c097cd73b60bc05eb2a216d7e73e75ce89796b90ec16b5cd5781ecaa31c1c936dd2962df499625552638583581e5aa3360653dd5b7715a0fcb6034073601ee2145c865e845928bc2a082377f9e268428c77cb2b5f16568a4617fdd5823db9beae0868dc90c067b21e858425dcb8f465d5c3e445113b06946c4bb80b4056cf28b2daefb6a8ac99a176916bbc33176039973956901d8c472d4916e08cf1c86f5f2a383d41db2d2feb42338acb1f0ab1556b5a88d25247314828ef730114b7b5d69dc2f1414081268cf69bfac6cb263b98cd834a6aac925659d97313672743f80cd54ace1b755a4f0fbcb0116a079d3de5ffa238ce64e164f1032458;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h53cfd7abd9619e2d74ba8b95c2fc2c6870d4ec9aaacd669a1f8e0fa354aae78ba588f4db34f78e465e49b00ab3393a3800f23cbdb86aa562f47dbe743ba9217ab9baccbdd92b4c7a0e3e918d98b18e0b057e64d7cc0634f57e9b454827c83f175c0a5183018d580720ae376ed89b37abeb0a03913b02b5433b50df29192d845d218df966a75c96eb5a212df1a8bb6cf6f0bc0cd39bba15a80c7d12292db9c5d5642edc6d05e827dc7f265a000672c30fba9dd5d7aa8b0cd1fc936dc0a272301423ddfbb8d79486c60657e45e85e09e9af154b50056a8328eba1863f1e91fe62713195a6e11fcea356561e865d39b2b6f01c07e6dff72cf48ee595085a27c24de4e31f49d5c27a12bf21da587773dd28235e98d055485bc026f8ebf2aa4fb9baa645fa7f66efdb76520eafeff33689edba59415d534c3b2379457cdb82bdd30b82b8f80580dd2bb1e32fba14be288a9c18d0f9c1c3bcb429ab93574086624cdfd6a74dc3385a49047912e26743a5f7bb28dec79e32f98d51d5fce1e2125195f6ae80fc5f047f92c65c8e888b36aba5e6c9b18a5461744495f55b43639728a18cc3e0bb7014725d25617da2ac4d8945756bd85c3897a39e57d109c21bb4bcdcea17520a157ba8b7f9790ac73f14104bbddade28ec1995ee6cfd179e7776a11f415df38b2d93aca840bb135346f7fbdc08ad3c378fbf7825222577c19446f47b296;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h7723c267b92edeb3c15585426a97afa81a611a1383d7a920b3639c73d46f210ab743d3a5905516037edbd05164fbd17c48c9170109367fd6cbb22835bd2777a97d3882ef9d9fed0b82dd83055bad755c543f09904ef62859af23a6916efaade5874fd66724931a5833c90f0b421c89f462262d59c8bb478c6a384047e13ab73d6ee0ede05fc388bcfe1ca0884bcf6a33975462cc2576fd42354a59c53e7f6b078bc517906a4aa02335e32c6f32868045a9773ac068ebb002c1bc5903cd456c5bcddea493e6906da828d1aa022c6b2371e1eb7cb330dc311d4ea6b2a5b83147f32c323bb3d9f80ddf4a1d6e2a3467cee1e6d9403018ca734ee775381e909e07447c2a2db173e94bf3e8415dfb4eef219a9abe82c6969a52ee32dc1b6c3a298e497cc4ab2b41e2f6c66427da6a6c9e54f26a64a9571a861b286e6a6e81c1c90190c4376de1031604da28920812c9c2da9e65eedfbd566d52a1b3d9b9001a8efa1b36cf523a3d802b4f004b32b7536a1b68153d1e73cbf49356166b522f2ac1afbcd9cc6fea3be82ff379f01086ef3dba12ef8ce47a4946d3bc9f3bce81ffd8f5a9eaa5673f793ce2309b5ccd617c9d905f8027c080ce4b7c4524a4e0875e5baffe3fd8e57ef27c55012a3f13783b50ded3727440449b71aa2979af30a4382da1583b547bb3295a304ad1309b40d483b04265bb7ff4b2aacc97d5a21637e15cbfa3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hd978d44b03e328851a717b928b94c67d7fab02230c7f8683bfeb605135617114baa3d3c5e8926fdf0a7b4e9e5034b2af865dcf8314de39c3bf4f5cced3898a09dbec5ae0e974b4d4dc1903beb0c807cfa23d37493ab266acea78e72f0462f00672fe630dad4c8f0c03c131915174ab199f53f102b8e188fd6cd1b6a45399c3192ff223b23e5c6fa5252e83c9d127bba6c014d6c281360c71543b9d3338144bf12416823e1cfddc7a0a5ebf3208345edad7da7a80720910110666c72888dee9d81fae0aad59381e4f1d257b292a91c1e4871bdd331229ed890e867c577d28d09cac91c73eb34c73c7deab7ef87b1ee66ccca207902721de418078dc7969dbcafddd8920705851f7be3989f5840e6b1e8ba5ff5bf6bdb67db5ebe50e821d9cf082339ecfbc0cb8b6faaa49c10205a5f50f81fe8705126807cb9053f3f650e0c99573a44535bf4960233f1c0ac52148dc30054e10c87a3eb22be0f38725e84d94f80eb1ce3446a1592127e9071749b402bdc760ae799cca2ceda870b325f5b5c5b0b566169f28cb97b87de7c65794d2b39236ffea16338d59266a57f79eea114916d10520b2ad3546b316b2057b3f3ad7b48f8bb06be157dbb1cf39c7496c8004ed61a1c25f5f6f21ac4cf3369a47123e0acf30241e2595a302da63c5efe8461d397a3fc3b02e1f2839f76f621698bd1f037f47af135f26776cb548dc7e7b29d821;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h5f1be8351041a9c82c121e74bf0137c7a9aa0a890638b122e89919e5bd4656195541a0086b02d215f0c787d97425120fee29a59eece3f16bad49fec92a2662986bc7bdcfbe775a3bbcce19b0f2aeac481315c5b15b80d6ebb11bdf2c31e3b4996e1d9d1e3a014eeffe78bc5dc096591d45622e68042432ae6c15c4c5e39c89d0066695d19d63ca58e66998a2868539ddf717d8d03e00e22b8c5c0004d84e4d5a4d7757a5e3d128c2e6f7e573e184a538ecb827bc4d7dcffb46867f38a80f5dfc3eecbf2bd6a2476e0780d48ce4f8b62060c7f325c5e0305652f8cf082dff2f9870b53e57a7c87056fb5499b31b1a3bbd359f2af715315b7b2aaec49558b17cfd4512d6a9476ffbea7b0465d23ce14897e62419a43feca975b72205687ad17fc80569a3431c3d2b6a5ef7323587ac9c58564b16a6610b8fff1c432113be925c871fc8f488eb3d9b1a5abfc2b8011248097b8fe6a23221c66891e7e017d63660444cc6d9ee0af933980a44dc35463c2c10f780a093d5ec32bba3c2e4f32448d943736c1521f5595fb4b8fd2f63cd67c147946b83ce10786053eace5be1ec44686a8dbf1361317ed04073d1f43d327d744aa6d312e0b37619392c85aa1a6dc97ca76999f43f9f4ddf992c413c084a298dc3d8626a85765a98b0486df677917a7b38652fcf3f0d62c5ea5093aa6e3a85606c3d17bf282d176a64906b4c4fa233a1a5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h303129eda02a73c68f520310ba6551af090bf2f0488230efb3dd12ca181f90a16f596518001f35fb4d2c4a62eb8cda8bf1b1e8f2209efd8316ddef34720ff76ecf8a2abe411cbd862c443bc897c9776e5ca065c32261e872e94e0a64ea46fa45274907136161ab4166995eba19e7bb06c8a6318b9bbf171df28818dc0db75e4843dd9a6480d185fb7b26f8ea1eddf9cbe0a6d2e908a092c925869dedc7d5a2fec7edacf697a90348f725fdc55ecd67babe74f19cdf128176118824a7c84eb43a2220547f94c52d73839694f8d5b341174cbaf6b3d073d86e0c550cd989467eab618a8ae8220363fa7d00d389e14ba476aa0e212157863f2ce26cd99be56f56008cc7bd1d7c99a5f62add0a2b9c24861c7a8fb3c3c992b7454a9e0c94dc24e711c77078be53301a2526b3726b514d4afba72354314c589e217ceb41587fa9a3d0729fd015bac7b72d7266aa17e2e2d6e6d80b7aab44daa85d82b092d7881b373990a0e514d21b0e9555781a7bd9d53c64c13a9508ed0a501d5be2e03d9a54ca6b1e966e9f8257c8ad637912a6ca73410c46454c39718761ac625c121b4c8cd98db8f7b5baf5f36ba755acf1a22492290029c740dad1c436737f6a22f026b5a44962d855521d368835cef29bd1932cc3759a2a59260a325ed0654d3478d0532488dc09cff4ae465c1d1aad22af5766769b045beffa736b9069c9958c87032472ea;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h39e3150d235301f2e999ea867ccce2692d1f0bb891f1e582a0d353ce075a3393a091099ecddaa2992020aad32c276ac99ae9b1164358df1fc4bab2c9256269d5537c788826b5f9b6d5e2552dbb98d2b431e97bd6f82cb92a25fab8373d7f4798a7f1d3f2b8c804fb89844bd548ca3e3df3c870f2b460568d25fdce089ce6bbf85cf732f85743dd52663e83d9c244557560706b1857fb756294fcba93fb06548a3925531ba8102ef15ae4472c3bea96d240af5b99963503258fda5dc515ce18ceb7403690d5b05a280141937e72115dbd0764d904650e608742e3970655e84ade874f015afb87487fbbee9a9ee70e16266741b00091e6837b11cb1050175cf937e601142c2ff33459d0ab418510ef9b9fe6df652a845d2b90c17b84d4abacb55117daa970a6547ba3b0a1a47aa8478630c6b8592d6f72401896a6bc0d4bdc3c15be6ad933eca99353700f9901b8e204d52ec06335f91c06805eac9b160e2d40466658a59ebc0c328051b7eaa99bb5cfffff787866765936f78b9071f151047f09d9b222e5277f039abde697286c1c14a93ee3fbbbe16dd3896bb553d527986e34f799ab13685856338f94f935938f9292d153c0aa5e251042c49b66cd9971258e344a54f654c0fb819e56735a2f2504edb55eeb41f51f841d3b80878b49bac0481f6216ca1e4c7970cd2d774bd6b288f00ecbb47fa501af6e2dfb81a003808db6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb3d835ee1ff87b5107bf413f67d59cc9184eab1c84a23ccb686794e74c385927703c3a4ac98be3e6afe207199f34381f78f1550adcc7cfaffeb19ad7886370d89e8fd656c819240e7cbaae26f241feb1ed9b9abb575b57a8663f4c7969ac1bef53a91d2bf946cbed72b2d2ecb7b2eafe8e284aa6d16b2e6f3715bd7a4ee54460ccdf4e34788c39c5e3ae6b4fe760773464902e62f4b9a6dae0a8ca545bfeb1140e70051ad7a248190c5b6f355446746e0d9e5464bb5ba267d88ac2284dcb6eddcf2f4c30679aa2d197611b17740b2e60b5263c94a6b87f9819135d645fc8930807db7574ed07400db490814f34535b3363ed32d8eaff75e2b6004f4a3e9f2be73cbb2bc95908676c2c1f2e24adfaf1ba9e9473fffbe2152df69e9924fd319f4334acf345085dc1c42d01346ef68e10a5a3e646c4cdf2d1857d88c4a5f79c94dbc5152a52559e6f7f9f9bea39d59999f9b36d26fbe0fc2cc45ad3233f52a5f25bb6d3e3541f19e1545cc56d4497c9b5b66337079d8cf19d41d1f471f0d8a57edcc549dd22108ad9a69aac2cb46c71e8275f283e297e967e3b395a3c4deb0c4415eb09b434495693b11f174982ab732467b2e3f8ad1b2a504f31260941a9ee3e651acddd43db1eb259ec50042743e6d1b62f2d8b1368168a3374e3c076a1d76cfaba89809d516d118a05244ed9a2bf515e35733e4b2e0cb1be0d340af08b0932b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h7a0dc1488ebdcfc3882374c42c431f57b068bbfc396236fd31099a944916c25d05196e4cbd9408f8338d3cecda8d9d41a791a5f6b4e0d5ccb4698331e7442a15361c9d9ce0460c2575c8d8494ef2d747778e3ac0a05f958d626827ba245460b906f00a3c8fcb9fac6b6ab7cdb98dfbd98d1cb72d62c9c1ba4b3a1fc35fc0fb4a3e722b49b38ac8ae6d1229b54637850d28bc7686ae782fca957d313e13dee8e73d00265cf4acf4e27f80130a36015f2f92bf2dc95c02dd3abac5988de7f499b88cb6f34ca47328546a03d4ff8e6fd83a229a496a3164186befe2516134d945eb8e0e26c220285d64719863291069c49379106ad3059e7f9655e71febcabce2e2566d4e1fb38613e5503d17263c900ba3c9a7b05e28129a6ef5736dcba4dcc10c473f2eee9bdfe725ab15eed4149dbe79263445b5f8c4438a82a6f6458cd325ba8ec77e068ba0eea98f8bb84da6f1e833c4f553a856a5ede51f0ae208b749f1cee255971161b1350547f7ef3dd6216de1ed263e2aba79eec22b560f5d3f4726d36a6fd4adef5202ea9ed2c7130bacfcbae1305c864ade6e396dfa70e127e9ddefcd3121801542cbfbc1ac4447bb6b8be956cf665ed5eddfba6da4160962def7361a75bd6ea397c0121e15ab9f82f532b1db3ace9e6be308ec6c8a8a7ff8af61fd3c05b3b877ac96c136087b2630e3b0bdf7d136fa7556a07d9e07f087ddebbcb7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h2286281fc8984499c813645e58c836006b1d686d2f52b8ae653c7e56c5799731e30024aed62471d5bd156fa6b10729998d53c351b73c44ff3d0a31d3077762d55244f23b01fce56c8a98e57b982f12a56377c01f27768f7a8c971b14981ed7017394b3070e9939ca351555233a86cee68dbdc7de98c79c6414a77a38aa64b25bdd96e2efbdee6bd5947cc1aa2159b986c3e050e48a8903da69933d182af64e2f5637511d636e5fff0a0df2e964b7e718d6cd4a77c54a1c55c89bedf32797db9676ad707483c6f3907a20ea9eff9bff8745ef36edf84aec9b18c9bb5d3a75342e8c8a8fb7406a7fb3916730283105f60809b9eaaf181d29a36aea1cfb4befc399af34477437a520a9d3d8fc17a161fcb4a8833a35cac9f3e39dffd2e0d2da672f76b61c0ea6c5bd087c20a85047038511e15cd84bf011fd2fb32e8b768d8fdf1c62b5d8a56f704ad55f84fc00fe14cdb351ed740200e67b6f897bbd953c6cbe271aa96baed3d5796e0606caae6b2e22b575d3a7b776b7aab671b4d800adf10b29e93c093c16233e7c7e50e8fa3ae243b9232d926e32929a334faec180bf0c56aab4c6fcf66d37410722d4eb1f96fe16bde9139534e7f4887ad5a2f1e085dd22f64f04917c5c3ec0df404f328e455d198e2bbe51160a4f283c61e99bcab09d90a4fb7f3b09aaa5b8ea130a06926132e7409beddf6ed69a07256f07f6924d501a89;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h76a92cb315f4a75906e7d8117e29691b93334053f37ecfbad76a6e483d7ba21ede759534cfa60ded52f9de97dd97376aad310185e32eb1ab2a64583cab617df9b3ed69c321c6a6ea53c38a5e472c92c09827f667053843915e9772c507ebb9f94520460c2e1c80aef71c83abf47c710a00928655ac29c1aa678b00d73e772498af4b1b708502950483e88e1ad91834ad38cfc6c505654fdd0787583717ef9188d6c0718f8e937ff190c308bdff1ba891613305bc5a105fe585669bbb71b236574e525cc93b1154122146c7dc7b3110c31b0278ed64ae9a2a643572702038f2c65fe3d41c7ef2ebabbe767e1735c1425245ebbfd5b1836d63e58ef849a37ea0e39dbceb6bc2dfe75d1797b7223a52f33223ea83dbc08416cd8bd100e29fc3380b0114557578b84d8aa1f3d123767789bfcf06563c7f139d5653ed624ff32ffb9d5e5e0246ffc1c5c85170578124966da97f1e5c8e9145df769e28c55189394bf95e9d58dd8e8bcea43062e4653f4e56d7db0502b7e4dbfc5fe4b44e3b9049c4c451785d108c65d7a6e944d1586ac190f873e43c12623b9da3affcd2428798decd9d4f6db8aabcc8dd560e99482587581d2ef852e03cf6c425e3bd13e7a46a0dde3035d2faa9772ece0bde589a22cc676784d88de41d8e007fe9a8563d5619efcad05816722424630bea2289487e7e1c747b6ec9fa1bd2a5f660f05cf6a6e43480;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf0b294daa7a47d966603beed3abb7689fef57fd76354ba0bcce3e2d28c86a1be0c6b38f4c51d88d3630781a8250f286a95f6a8ba57bd934d45b982058a83f7a517cb6a5dfa9e71502d23bf414e0d01493a4a4b010b30c6074ea64030650b983d0b64aef90c52e5a56ecf0737a16852866221440db283473f096b6bd116466206fafcf0159ffb5327d4185457a4d3d998cfafea12cff9108e1e9e1363cf4c5329122634d056c3746df51f935068575fd8ad10f5b439f2d446b7bcca47a6e7a72e931b6c5f51ded9cd8bcaf34c09717eb64236359497a6cf1de4e8535a0b5436b78a31ac9df900bf25918f8b2b3534495f7d8f47b3e6da528b3067a3db0098d169e4b0b39dd9913813c2133a157caf6b097cb552fe214c30e7368b1ce8c7e6702be775bf77e96ea346ff682c22145acb36775f65ba473d1a0367ba947c2117342f7396085480fddaff0bcc3377e7ecb1a7723ceb0ee3d5dfa7c5bad22d96346da28863ea92b4577f1cee784d2e9c02d91a6558209702114c3a6e7b6472ad9f730a3ae6ca520429eeab86c12343a4fed00377c9bc21484192c1ee57c7751de6042933210e323945834071a7e90849f84fec2dc95ecc8a7ebf25d48991ff889cd902f027dc18e26aef338342eb64d188574c605681f6fd490988faf9bd9293f33a99e5a478b5279aaaf3702992a21916f8bdaed19ed27565a505d377b9240d0b2599;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hcbcb93fea2a3305316c5c8b6ef8b691ce76b6490733c1233bb4abee7b59443dc0ae00896dd83853b1d32c37411720cc2077b5f14326d0a64d0f3f808365ac2d4073a16462cbe658c43d392c9b50da60be38d0a4f3c49b13185a4c439807f934f5860bb47c23b22975fe21ec4378f52e5ce5c896dfa9cae9443894866148dc90435bdcc1dd0b528defb6a151d6b214869742bc6e31f36d24a3c15c7db36d978ddae2fb60ce1212696f885bb3ba87719cae6b795f1f447c048b17d3dfb9d38820ad1bb08638f867e4780fb559ece7fd060deac80317817431087a470fb014c44b529d121c9d4c5662d3dcad93b4a32ac922d95a76e8a9bfb80fe4da29587bde13542a0b906518e9350325bdef3ab9f11f19f89b1c20a0dfddaa0b2236e2e35f7793885f142c12549520038d3b9c7a671cd85651c6c846b524986cf59ba68f6887c2e7d94322c16c8cb73c3f0a5d90621d9f382c890e725bca70f3d4c472564cfa9c8a2e7044bcc5241e79be5c690d7f853e2b13603a987f9fa23997ce62ad7c22919f668c2b1b689d708e3381c433771afc4ecced220bd3bac779069d11f555fc4e28436b8df7379ac6c315f133991f5103ea4062a6e8c5d520e2864c691d54a11d1482d6ba1c24d16f1d91061ec890e835e198f7823fe4758bf85d0e28c0ab96bf375b1019bd721b4487147ab0b82f7a2766cae7f4b1e437cf8e9d756a799f443;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h29f13753e0d746b5a358e152ea12ab9ae1390c95c7bf7d090710027959ca26aebe9dc2e0ae657f428d81281e97d21aa3c6f08ee4d5f8c495e4cca197fb08497ceb412d3801762577960300229d5769688b728c3b369d68a39ef3c39becdffec0a656039dcd1c53d63dd9d16e38e93b6e275070cdb31fb5ed5712cb98e97041cc5265635990e79890f70a67cf69769c5db4c226922ee8e1593ec13ccfb6ff03b8126ac01e79f4f49f66ba6853fb1c912890523c84eeb270a6ad280ca44dea9af70559c70bc5a877ae7801beb212ee95e5a9648256cc3b0237d4964e0c4e0bf336d9a9a2f5103f383b7cd5cb2f53a8d6a52bfded3a524d35c61462eed22cd48aba3748fc698969407c53eb2502bdf927bc7d4c1c174723f9ee1926c4ea4e6f0ca173f67a42c722187045f3c6e6a195dea678ed4844de864ba96006c19da4119b1145565a994e9ff8d20ff77d60c5964cbb0dccf99a104ced665415f3734e4f24791674b9933207da8a61cf6364f7ecccaf15782ed54d382a86375e7a6eeafdb7503313cd8c7faee1ef47e9ad66432b06405129b1bd0e971033b3ea68ba52b94c829f63d2caa03301cd285a56d64afc9789f3e9494feadd7b8248d1975a4894edc83e1ca4c90dcbb6f3a198b3b6151077e5b4ff88cb811e340159987bec98d29d4996e847e7fe8063c2cfdd7bdb05c3f08a87f3ecf637496ec3f4809965d4866ec2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h5262ccdc086f5fb4b30b8c765d688623d2141ad642acccd3a72c5cda0a62422329872667a065cefc58f275de0367926b40ba604cb62244848d00cd147f04963e4d6fa59447a5bb6e59fc50a00e882a2b397ff74033b55f943769c503fa4ffd39a71ddd22d7e9debf1ab5ad77add53916cdf8f6b92ebaa00fadadbe8f695da8a1c02e66e8222801fc2e2d151691b532ca0534f6ef020618fa45ba2600dafab9718b786c7060a744eb191dc802243e9d3d688142236d917690ba92a729846d214074f95d9f1f7f1258d0735cba14fddd8a20f968a6bd0bb77ce26b8dd46ca37178bdf4219e51212ff23b1c75436e51a1eb952b1745df26865eecf93dc9091cdb0dd5e795a8697f55c9424460be36a0ca78d48579b7bf49393e645fc2efe7cef7f0eed0f0d59e9253e0e6ca7c4773ef61572e8e1026eb5cb577a24edb51fbf2294468f59a954dcafd5ebe52a96d74213e4ba1c4b63976bd39024c1e1366924aff3c3f499515dde1e67f0f529d15f01f021dca25a0b8c7460a9289a21fd8566d7a805365c69373af30357af7dbe3facdcecb13041889e33fe63caeb43840dd2031278590ebaf395c8ca9d9226592cd97f8108b069f1e0b611c87af6e6ea65dccdbf73d65851759a9612fc14a760e78b1cb5433aad6bc37e684dac68e0e4013d2cfaa452dbd3e9140b92ab9d2cc9bb14edf37a949ae61c9d8ff93e0329158bc736789;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h27000de33fb46e9f7897ebdf46bc9ea3d3976f73e2d4a3066916603dc3b057bf187c79c27ea987308038a9bf039d2ef537b26330ebdd7cd1ffb2e839feba476a977f449354033911a0a928dc682bbfd2b47340a7fa2a4947ce2eb34db9b9e6590a163a2e1137c4dd31423b2deb481b3234d8b0739663f3aacec772005bacceb8e0c2855625d223f96e43017a0981fe221429d9185f8c1e81067a1a0e51eb998a5a37d0129c25440977b24ce473b261859d6a34ef33901c2d21048798c02696c5107c1344d2fbf797cda6165c417a62a9f5ba6b4e1eceddce55ddeae1c67d7a4608454eb2073e77187453d21e63b58ab84593e213db79048df1d2ac04d987e49e7dd868a794e4515b4dae44a7a10bae9ef9ed65b62a71c06e939da0e60030120cf73c72aaa17b812d0d7024c4c268a626293041678ea4b714563d71e91ae4f33b6dfac5c7d2ad6effab434dca7602052ecea3b984ef40c68612cd0e60eba8038dc85d96c1706dca239e7007d49df6ded0388c163cb6a772b05c66c163f0e19201d59024fcd59885f6d549323837e47e9f505da8635f52851dc4c274075fae8cb608d588891087949565b9763a4bae433081b5307cc8ac1294f2d7cc5388a30eea54e4474579affa5bb4ad938dea5199e9e928172932bb4c4ec288247fd3bc870ff95e94647c684298544560423f64095baa7940f74d780b8f3d936f77930e6ac1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h807a4c5af4f47bbd6c7751a3a4bca3a0992884e38ed114d0457784ea6aa56b6ddf985cc98ffd441b03506a8ddd0f92ba53041a6ae32c2647d505993e2639828ebe66688efe35d387219ec8f1b0e02683a15ba3a108dbafd85241784a117d49d80c13e0eae0db3502ab5d412186f6adcc121fcf52dc6c5c1f83234f25c87d81edf519d6cfd0386101c8cb598a4e5ae92cdc983670b05401780bf393d41f84b66abddc15ab2c527115e94b337c488edffae6d542ee5e2a39c02e5a6bfe5eea7721377a18a420b5d71ce79507d563123812d4524a97c2247b91c70ceea310e038fc5fb9b6f5bfc996672d38c63291312bbfa85016b7ffc95782cfb9e8d672e33ac9ee79d3807764939c1d04d3fcf76857aaaecd9236cb9fbda32d5a45779c5f62c0c7ce80ac47ea7a48591ab508108015cd429f31e5a97afc4ce4f1bd2e5c1d6ef56ea50d298eb77dda124cea79c7bb82412acef161127121e2a37d97293999f1b9fd4a64986bb2fd4ccf16ecb84f04305539a0da200402f72a3f1fdcd7fbae04c7cf1d5d0e6af1ce32b75415058c0c7723e72cce7673f9fcd8531f04c91cb96c95d2a4376c8e70242d69258185b3337bc70f7d3762d3b5936633c0463099a3cdfc44bfb2bd28107d874d9d677ef6ac1ac59dfd4ce688e29ee9544c53ebe82f2d425dffb414acfc05b42bc94299336d928ff9799c71c81cf41fb7fc8436964bb4e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hfa39480f9d0b4890f049c1204f738ae523c78f760057a2399cf3eedfb787de047a8e442f15e7af7e4fbc6fbbecf53db9f2972887a15a8e1117d0ea6a087c56d8a9556c1513da0efe7e9c4d26e5863e11970113ee68723dd0c13515aec1659a83a87b5a04c1c4e4f856bb0bacea6b052b2b8a1ad1bf8b9493d991b512212694e41c56f4394c0e7a66c61773e65c91f62ef37e802aeafabf05b081eb058ff5dd9a39b76391d7994b5713a448c94180110130c47d0f7da3dbfe176a91105d7dee7328587fad29044cb2fd6aacb6a63535db89db94644b00cf84ee2c68c5d6ec9229791eb56c48e03fc510695f1b2b56e4e1f1b0a2e20e6388f7852c186a230d5347b921ebc78179f5b45fd50641af1288349cfb0491879f06ede362a34e7820ca01f4b561adfc3b94a2f8ddb31dae8909092aed1a6fc37d75838bf29bd5c3b91fe8623b9311c4b0b280ee7b2caa85ef3839b6e0e7018975855e10632d5b6c95eb75fb015933bbb2bf4a41de2eda18cdddac89f9dd73761fe38c2be1614ff2cfc2254c2e2ee1fb8ba3d221462ebd905863673278eb69bfd63506b0995f5b81a0d86b955a6d8a66ba9ad3f2e1c468f6247b92117b89186e213a6d2e8672c27a25ee444a7bcb8b3af82370ed7a4f08a855ce34c1f65034fb3ef8956727869dceb84a23229c81df81a840eac2bc8fb4dd982ec862874fee32b3521cb527c1c65f08d7d9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h2ccead2edb267ff7ae8e13de1a94a1ed0c739d3723a000a6a36fbe619801a0cc668d33d4f67eb8b5b00a9b8d3ad5ffc668d2e3fe9890f8869a1343e082c52077bd0ba4832423b4e9c0c3fbcaf4e5f5bffeeb8feb99975d84796fb2ec6aafc882f3f5b507789c39558070190d715ff53a19f4fda3eb939bfb96507e64ab59cccca4ceb5f3a23cdcfb31426cae2126d1f26b6c59cd5f1670ffe61e43f1ebae4a0b1699ab5322d7b8e687f8c5baa711bed7ab72f87c4be1648d2c9d3117e5d91fa1e4cb503bb6237738f785f1a6857c89578a47f2849d220c2d356cdc9397f0434d4fb63931ed43366476b5c2cd5e3977da4921e26b81c3890f768f5237ca005da3642198c4d7cc0550eafc922f30b4ab0af0cad314fb02bf66c0ad433efdedc1640aa04a9bae50eadc16ddcd64bb98bb467743b54933b15d7e67d826d0b54dd9b686683aab3982ff1694fb37012a695bbd6b203a252ac8246580e1b1501b76662f4d688534fb11a9751a35301e4323a084f574ad5c3f247bebdd51740728168e2a830fc363db6a938fed44a94b3dd76a7dff61626328b1a6b41f9120cc5057a4aeda13d4843fdbe9c766b02a92ca2668f7463bddce41b3017cbfa47f2660684ad7701e277e15e658924af6a3f4c98cfa6bd531b264d53bf1d87c773d6243fac47d91942494f464a69392177eeb3dacb7ae1ef10042736fdaa218122c7fc8b50d3a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h2544c5238d21eb159d739b965e7f8aa335bcfa8cc9aa499976f516805642ff3f8a540b8a301d703daf4cb9870e5583604f89176cee10c51b5f96362a8c315db866ebbb972c699a6c111dd21af6ccb9d25e2f02843a34645c5e0139558be2bb9a6e539fc898f2cf71a6d72fbbf249d1f7bfc01451ee841e04b76bb9aa8cd0e41f9ef8dbbad32a51fba6c83b8aede4afa786046a7bcd6178e5147096e0a16239032c7b66e51e02044b96de060b8a8eeac5e681df0a4c2f7d20154df696b18dbb3512f63353c141a6cc5c493168dc77d422bdb1434d2f9c1a08b6703d57ac24700cb610aea90c0cc3c08163c7924bd0455371068af943a98e0ec8585c10bd7dd5986986f1a2713ec6acb0fb130f7d88a293a1f35db4692fee9c28b64392b9ce04b886d0390116081c49ee119844fdb1939a67b91c6fcb848ddba26ca4e0562f5569ecacdd6c69428c15cd504ba9574c602691b3c7014177a56caa33aeb147e1b1141492ec392b45ce47df3359ff313b3a0d9041a02203b56b983e61d042d0fe4cc40546db5bccca55ff7f78b181b02ec8e32ea4e757a0eceb439851a2c1dc4ad1e9398083db93b8999f16cab6501a677c6c0c4cfa2e46ca1353e54d91a77a43ca0a0307b68930dedb9e6a41dcf84011c4836347c92a2010ed5fe8769cffc969b320e069a3d926fbf0f4fa57ab53104f95e17727a9a67c6d15dc26ebdca3ad01cf84;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h8198c6bb6f049430cfe396bd75d6cbdd5dcc1b6b4e6ed6be57cd4fa8a662f6cf94261cf793379b4775047cf3e178d84457144553f91035e24ab866c7bea62fffe8b71a04a909eb1107145389a4e01a18c648d984f11cd6797858c859d890fc5320de22ffabfa15e0514bd70aa565048fd053bb7f95633fe910048a8e7ad99bad854c2778146e9c416fec7baa0d1a118113148e0fade58b1058bc8e3e168cae67e50105ce61bd1653a223193c28a6133dd51018f3aa1577580f7ce5fba68ad64253d466573ca0979d69b23fb1554ab75629ec923f673ff5611d64547aadd2708357b54f2cd9560c8a9c668493f933de6d0f83b1be96a2f7b9010abad12b3e514f093b9d0222ffc71efb06fa8a5b2a4bb49c6ad91672bbbe8216275082cd2a8aee2688a1ec98212e7bc8f5982cd9cb7b1677d9ffa601d2e65371165838344152130d6fa2aa7a71bec52d0b636c119f64ccdd3abf02f3c0bba167076887925cd095a4964723fad1c181de8fb2e2c54e64018611fb33eff153eb8ce03beb6d05969606d33b2449c0b832f3cb73cd345b961d872e447670a09f70614cf2a8dd525f69306a54db78087771df7b39f2d033ccda2cf7d8cdf362b244da5c8d1e39ee9b5b3c6fa8de234ebae720d57a282d7e21ff3ee36b574c550520d52883eacb245ba14aa695cb01605a73579b4849730c01bc33031a0bde32139a46dc2b3e8075b9bf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h649107e7c62729c3b1b656f1e2ae88414d111ab12f34b3253382df34be7559a4776d71aa46c43e5c68308d4d206b893a05642f39c50b7c0b4d38ef729da899dbfdcf8e8c8cf5ceb0f556bfe52779cf36ecf07918885e579c7e690077254ce678310b56edb0b92718788100f0322bc484e52dbb465278740fb898a5cdf4b5a3b43b9e47e9a51ecaa66fbb65ace67a53bd7dc17a92f56c73cf577ba12f551f7fe80f05fe040c69e2953e3b8720f1430dac9e85213ed30af7886ef3e36b661da29101abc03cf5c74189533a0fd4f424d96eade64c4405c143a10433034bd58b75442b871ce6ea136651cdd0d3a8cd99dd9f23aec699ff60e78f2e675ebb67bd3a06ab60ba4e140181951c3a6531fcef3ac6a61dea70df56ff27932dcd787d093d8826497a32e70363edf1052ac82b359992a6cff71523765ab495b8bdf9ced026e5672c3ef09119f3bfea825fe66ba35ce1082d89bd3adc127a5a794b7848eb49fa3a8ec97cc44e5d1945a610a41e340f8b78c426c215c3f423e506469bc145416972451ec1cfad9824e04695a80f6f06145068188da23caace4435de339f7d9dfba0924b205171aebcce0fa6dd9dff7f4ed2e55b8aeccc67b3d36a907d5ed2e845c138e189ecdaa8dce6cd848ae5e39f3eaddadb558eb80d775e6da634009072350f0e37c3d02029fa62b62c1e06196f869205c81d5700a8f9c846c094a8a5099f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h2de11148ae157ed49a291d8210044cd97bb94b727fb0b917e6f147b9bee8f6130c8b560027bbb41767f0c3ba766c716ae56cf02611a47ab031841b580a0af6bc9a8923a233b0564ae468f9e87241a6dd58e39c259c46e2aead80b25aa327c010d1fae48385f50fffb6fbe7c4ed7a809405e59f35e3f15619261c63c39a2bebdd3ed46990826ee41396031e9001e201e7ad9cce795cd90603ed567e426f8f696d3ea140c240898e05a3bc3084c279eb6d02cce2c7af3769a1ce6429d2f3623824658acf3eb1131b069d5f3d69f2a4c09482169f30d9eca8412f0068f97b3fd129121b48dd17853ed34a13e6561dd648027baf41b96347558472898407d5eda9a8465be428962324e39c85a2a2ecf524018006a2a7f9f9aefe53628126f02c20cd130e0e0d941c6c741770be4502e0c880c9f6384ea95e5b977f21676aeda9dab7a03e7195b9665bd1c4bf413d89c36e7d394ec39203590b7c9f06bc33cfb8fbfc711379447f9fa16d5f71770320ebd645ce9961c8e980f0e3a3c537f71e6576307a0197d5b40c223594b5d31ef72cd30fcbe0e436058f8c33adfdb80031c1b197e0c22153eb229caed29442571f3b0984f1a05545e634f08180870efaa8682443da43132b85c95b1c6b03c68c805edcbc66b7a7d8dc91182541d917d2d3e3e85c5918e5db4afb01ed48ee0db928f740664916cea4477eb4231081b72bf0d8e158;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h92d512b7854d4def49958c58c5d2e9a199959d259c01b5247b8d117a94812f9a9f245ef13c8226c7365944462908b05476164afb5e48a2ea63c11abaa54a0506c65b3a2f3a445093ac9c6e4079f82eda9c5ee383d415a6ef503cbf9283488e68a830358c15fb1feeea04b88dc2eb635db6b7493ff866e7b36abe60639fa0829d4364cc985d7e8d93c47ca145f04205dff77b4c1832676737fabc8a1bdefc23bd3a288b55b71f73585c370a77bc0a4ba960e13c0684a36eea23400cc3b1b373630c36394e6a32ec5c9e05f7f091fc2f7a3f985997a198171175d1de78202bc0da3707272ba897f8fc39aac04541276671cd9935cb1f414976f2d04e24b79a14949355c0ce1848a1c1a892a5e9ef36f03468c9a45c5d9155839f05449e0961d961c3f5e9746d2786694eac957a7c982285c0cd330ea77a43aeac1d479208cedcc013f002fbc5f1265b74882db027742e69fc302df65a3d387629968e6cb7f6ce360c71bf82a1ce7ad79b5817a78f5ba49264034b592f8fa6943e5d03aa43155d8256f030d61df37d4dedba14334a0ecaf6a768736d109f8bd1af806ed7f902d0e264dd389ad74f36df9c416f47ce2a0e512d0c93a085e8f61099ae247cc8e62c30c30622e03753d6a6330b751dff66b69a4c4f00106d54c6c57ff0bbef449931879a2287144f310b1f49c9b393d9e571bbce7890a03b7cddce9bea6b73714bdd7e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h434b352d3fdb984042f92a4ee92d86b62b39fe2f396b04e4f8571e6bbc53b13eaa11f6c502619f94d55a44ae8ff00120542c63839d91a60efe8b6da4c0768d6763d622c7733d125e8d099da95c3f6f90b5f9e0aa6ec1a1ad29ca87756a396331934eafd12bf8ab678c048d6ed577680b96e3a50d263553358b76014fda29bcc13045b80fab38ab4d05588766cbd56dd693ef3f82964876d312801c94638f7fcedde0300f3c0485ab4bce9e8721c33d5587d7bc958331720f5ec9f2d75280fd61e1283083aca5941e824a0999e458afbfda55b906690941769db92bf61809c18b60ade0a2c5f0b13eabacfc7045458adee4a11e4a579d62f10bd7be95820e4f60379ecd00c0e9f013fa71f52840c6e7c26ffb285f00907574965c31e5e250dfd25950b33fa57ea5a10aeb7681c08141ef529c2b6035176358c1ad4189ead945f0cf34cec94af378c35d2d3288ac7d9587c83187c46d98f63e324d26f8b22e77051d32ea710c7a0f70acff7513518aa78ab554184c318e4579ee933ce626ec98e70c8d9034938f8fb9f7b55a0f557ab159ec8e42d77ccdfcc1d3e016378ac4245ccd8827ece50bc83149bc6bf763f84b70a8f846dbcf82c32f46bbbb313391f43d7ec3362bb035862a4b929ae986ce0ca3b88aff933d2ea7a01d9fd957f759b6066f9a922267604722c7b4e7e5b75d95859c5336727a8e3a91a8988633db921f73;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h65ba5ade30347fd9c5c027a0f54bb996ea6193ebb5c46a0ccd51abfcfc5b53d42bb3e4d21c9923b5ddd9cca4682128cd9b8a0b72ed31698c2622a0f6b8e3c2ae1971d3b3038fb8ba8628a4281eba6397cfaf93d69b16ec0c2a640245b3f179a7d835e8c8f0719422b83525ec501a7f89ea74dd8376fc10bcc4ec5c3003c01b348db2bf812c2ab3158e1780ab04e3787b89cb49365beea646dfa501214fdd229abe202edea936c7f52439d2a416d21968b9a1dcbb8ae787033089723a0e06e62da7d895315b8679948b2631f506b3a8c7a0d9aa9ebd65574609144928cf02c82b9ce5d98636c3323b974fa5b94a487362f5132c7f49ac81f4a2b773bf595b6510cadf3a52cd711d81d8f61d0c7bdeea9ab9edd8b6a3fc7ddf60174f466c5acddb954bb1ce44acd03befcbc44b4a5c92d43566baf7c7dd966a6b9d3a6bb85af6206d4099c0245e812fad2792d48af9120f82fb1e375a8b1a032d5b328a37c3500e41c85d9e024a0e7c79b8bea8dcdb6429ba586ef9dd5b67140e322331e3a1686900a287a1faceec87b4caa5f1452b233d21388d41296979debc257f988fdea96b2aeb8295796a6b2672fcf9c3738dcaa1094417cb5dbc1e3856a3d967de6d7c2585e5eaaac7d40575d0d89b9a6edfacffd3201b7a31ee90f77b80cb7744ba77db950025dbd10e93785617969f9f13d0612cf77a2acc3ddd42d94948f4935d53d7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'he96373e3633003e9f3692558a0fde06426f1d8ef45ea601d2e21e81ca4610f1b2af949fb248947ab183da12d93488e16f900fdcc830ad429de038a0b165d3a0a9898641ae3d9b732a131c6545f96b4789e44cbc1ec0d5ed3bf16c5f3dfa37acfad96fc7f37e2f15ad26993c38c886d61377e9970588d6d4e1f06d8b27b10d8b90fbcaf080573d3ba89d87182109d8165db0c4c773143de913b488c892c37d11e80c3126b76bd5fd60932c8ea9a0114fc46ca42b57e13eb9dc7c88febf27c553de71ba0b722cfc5d288315cbf4a6ee753c3dd390b7948d1a16d3489295809a9d3830f640546c0c8db2fcb7ddd0ae7f5a1e5bdea69b38f2cdc77a8387116e1c360285e922739b764c0ee762eab5b19def8ecb6efc010b3093b37ef6d7858315c1978e032b092bb80a99871a7ff15f79f31547b0a84edede2204affad1bcc3994b3aba1279cd6d149d1d870cc312738a0ec81ca433ba4b39920a4fb98f3e849d1485998ccdb088f1cbae0ab8e8bf42f48692413157362f2a5c9731581ce2f91cab893592d11c0b2a7becb17ea222c3aa5d83d2c7a0e54dead59cb1c61640201976af28707138c0338ae19a7732c955be5ae69ce637690211d781dc81659052a0d67cf5521e8c58990489e25904585ce31606c3a8941519e144e6d7963753413d0bf54ffed1a8c223b53546acf8da2abe1ef8c6b43836a6b44a12212070dbea0d4c9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h88cfd33f2d98b1e66edfa12cd7bd6bd282ae4081b3801ed1dcbc6dfcaf7c28c2c0272fe520e46dfb2546ce51a995495186a71287289fedf248c1d30c53a480d28a3ba88c6da047f4f72b514e83234101e750719942e5eb0b2ec27887c33b6cff2216846e62df282d10ebb07ab534505853ba3f49e608dcb863a594c2fc1de5bf19bd98a16b782d952ba3514bb4d6df4159d36eef39c0d943f26c3216f7a7d7572e1c99f585fa3f3a359999687d75444ae8ea165b729cb2d2823adec50af98f12681bb6e83433e7a03d3e91a4f790166f19df234be707bd9e02c5ca2b568f1be9525537bf4063c5b5e995f35decfa9148f1dcb8463656f869d37ec91a80f369b3f63cdad50dd56924114d2c853fc2ac75269f08f3a65c6b7f5d3afeb0104e8a8623c5c2731173bb362caf02433fbb0dfe30835001d2ab2b77a721929cdec63579537c3094862ad6e74e48a12b118aa3bdc10e5988c8341c801664b39e3392fd2fa9d96a7706765b4e4611e91b2b64044930a89fe6bfe5d12028b66205b180d5a1585264241a7fcdf49943c98ba54b1e1874adafdfa83b9fa05d2a86ded9ad4698141cc679c8a6df9030c165666300ade51eaa1ce30ee91b3261ae3e5a4267b8c0eaeb876c57f52a28e8a7ae2d30cc35bccf585c81ddb6a72edc52adfc5e3b53b6ea6b8cc9c40c9ebc18211392a372f732f97aab29fa1e3b04e70de8a320f3d4d3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h1cac8bc28f0da6c668897355307c188ffca9d4e95dbefa1bc74522f0bf2f5e1d42afd86e0587acba1494db795f2716004300c91ca400c9f45c20a9d692cdb025bc1307326f1b311804c704c9a8d3611badd16ae14fafdd362a65d17760cb9c14a3ae02289c502cc848b13b8710dd94c521048cc40fd0a9863391f95d9d69a9b9c9dd814244d9200c96b22b5d01dab99e59d0c99641985117d2201e0347bcee4466dc1b4f0cd0e8c7d59ef4c85baadfc49b783ea2899e72f2888c10d41f12b9e1784062f718b255edf49ae83e4ad79c6963371eaa746b0f2415d6295a799c7f4812c54ebb758cef8ef5ef28df62b0fe314a0fa3a21c7aa9bcb9e6b62a344b057f210b36b5ffa23d77129cb37004e1a2e5be344fd7c80b7cb8b71e350729efa25835cd0762f76b09818c9556be02107fba73a34cc8b892dd3069c2a1970b8237c5cfe14bc10528b5df448aeeaab9edbd6f9e0d63c2a7fce7179486cc5fb640c5670b10edbfb7555d6c08bc68e1fd62519451f37bb9ae632b3d55e6027116e8b34b10c9af33de2188cc55204235a0f75bce0a87494361d0b65b39c59124322986a26e3da977296bbfe36c5ef356275020dda7377169d8e5d2d363e90bc92fcb05883880df9eba90fc97b0377cd5e1c207a94fbf197ce9734618894f0d1f05fa9e6854bc8528f4969fc820a1e9542dfa5f4dfec82fe9ac5ded4c282a8a9f6a4d0f1d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h970381e77d2fb194f511ab6f6db411aea432ed9dbdc0e50fb8c85dbb7a88e9a52258765f9ace1a3b134973e4d720b703d977fbb268a26090d4cbc082ae7f8b755238b6fec4d5f6b63220f158bc244bdc793c7240f16b3d9a587ad855336baff3c7cbfee0292a6916c1151f48aaa2d625be1d8e17eccebd81ab14308fa8f7e3f134bd54801706e18c3e545843a179767c8e46809db4dccd7888fd5e76b374cab15abd8118905d8960e82727ccef271021dd9c8e9a3b0e74bd679d3da01e8ce8b649a76ea8ef66d9e10583187c2a5976e356cbebbc8d8b9d79375444f6dc3422da84cadf7082096df36d31eace0f5cfe56d2efd34adda21b750d57949de98bb37c60e5edd05431a79484a8014dca1b0ade2a66f40f6af2710535836718bba35e5611399f76bd97c1ab25dc67c8a0b5fd77ce2abeae8c2b2e277b453acb8ccbad959bd42b424116f9cf719edf71a1654a624c737b27dbb6b55a56b04e25fda77ab431bce151eb3f038093405ee73e5f9d6ab721f24ab44c0d1219adc920f266dc853aab90f00c57022e03aba1037fa393a6fdd986d372da4db20edaeae466780fb942edf2380f1b61de29906d49f5a5abf6d6a87d8ba6ab15dfbc8b41149c0613ac7e3bc8c33f4405fe855e8b06056332e3a26679bbf708f23738cb1d86d79790c5133113097a61263639f61c24258db33a99276361148fab51b87a30ca7cece23a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6e9e4754e82c0ded4c09734e999bec42a1748dabe0c1e5fa85a86ad1d3f34fcaa0316de78c133bc6c65feee071886f1e901e2c370ad1bbf4ddfd7819a315111b5b2c8080809d8b6d5211615c1b26a86c0b9f5f06171501c356ec63051c1f121c65466341b09d9a4af4a60ffc0a8c1b7e199001291ada2f125ea30be09a809796a6d476ba243ac37de606f4f7923c04d1d9cd0c78a08a2817603df0e3932db4412daab4cf33b95d6c70bd04a0971ebb78f4e083d4807e0e977ee01334f1fe293538f2074f0ace090e28b7c2f8df25d383365e7653b05d8680fbab43f9ef96fa9ef838cf7880c93fbf0fb9d5900379968ae45164573bda200c6147f0c8cf6e8e406a7f5512efd6169b3a4d6177f68559dfbf9ec81d1aa940377fa410b25cb9c359b4026a00886b48bf94ab00597b193c9c65e39e1cc407268b2f4c46caf6656419976d450822d6d68e64cbbc40c7aa5f01c7eef7ba3265e235d978c32dbcbefc6305780a650db0835d0fa5ca4c5bc26066f5abb2a3bcd5b90be2396a3afbfc235acaf4ade327607fe9ca1f625b051270475a0b09ca663277676a35f920815b16814983b7d3dfe426082a1dcb4528057dabc5ff3c86fcc6fc699c7e09420a720deded5f6b021c947efc29175c7fa2fa2ce7b6630db96f49f346d1eef2e151aa3eaea206f5fc6f9cf173e9736164f062d3ed52c3a2d6e2d43a908c8a580ff7847d7d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h2933b9a5f564b810cc8787b6bfbf2da3a7a75cc0729d9a17f7d45727b75f2c1c78814c2dcb4c7ac930cd40595d2d0c0e55fb396033816b4dec6156015d7838cb8b0f3dd5dc9126cd7336ccef2192bf96f8dd6df9a3213bb21348a5a22dccb58cfd8f72b7ba4c451b5090f25825bfed1d18e763fb1bd230480fd4b71a55c50a016384b99ed513a4a2ced1db4d330d85cbab357bdf5ba799b358a5f4bfe99d5c41aec913436027adc3df8dc1b87c1b7fc56a5fed4d595a0d0346c1fec61dff95d67b5f3e4b7d347134bf61ba428e5e39762628144f03a9df86c3c5eab928c0dc9adeb6583dac1599e0e46edc076469b5ea8e38f59d6900d9dfffe36aaaf878d08b2f8de1e14b5582d347c32880b8237a0aff5d7d0accff7dab45c9d0ca11a3f4002713dd38a1e0ec2e85486fe9f68a2eb4385bead177ad3de9d63860ae4a78ee90f77f4a014b4221537e8b0ae65c1765ff919c5d7d8667251c85c244146ee807c4f0eaed37a329a43103119e4a13f615608c6ff69c0d610a0ea7d17d095f505033856ec6896fc22315e40c765b00f5d6895ad8c711c12051f830941bd3f08d3ae3f2692c382daac7b198ba9401ccd8177b9813073fab6416117c52a1d755e953f8b7f761927daf3fbc9b45cacc83b6f16bc2682bdc3758817975f75150675c8d8a00cc3f1e199ece0d36b4e0d44aeb8e3e64d5bcd4fc118d8d56ed9dd2d35d2951;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h48db7a89c0fdde96ec61fb1dec8ad01d21f1d4e380daf44a34b3ce87b0efe1be4a5135dad4bb5e02daef811b285c0ed9ab0e9168a4a6104e4ff51bf02f95e0cc14146a031f490a8d712d9d65118c4e5d1b41a0b8034ca0641406078e6822add5eb51713d50c95a5082c57374361faa675168e71f1190082f0a78c077a160950f3e6f28bd44a6cf52c4b45e38ab798520882fac18118986d30e39afd406a391f5351e072f25ad405f3e8b50b14476807934f9dd8625d53f77c674bb19cb6b16cd444e4a5a24a92441dbc1bf80632a041c08fc956df5571467bd72d0a4a995a71799133e2f55d6f502d5518d0ca217b68243f3e5a6043fe0ca94e16efcb3e60759df578a71062921dd904539b1753a7b69aa6ee41d22fe689a83fb61f2ab16543b364e33e5a3eae65323697ea4bdb8b5b6d4c094bbb84bc2665ead0fd1ad6760c4d3bfac2b8d8b055f3668811dd9add643dcce0233281e67c0ae9a20fd09a588e299bad1a493ff6b2746e59869ab1b2ccbda712084884992bd528c28a3b0d21c14a795ea87836eddee67d5f331e77aaf2d5c28ec641c08ff5ab0c196fc5e5d29db83954ee63d2b35f0163385b02021bf5f3a72d569f7812b2d872d876d6155b7925e2e110124d77dd1eb551268f3aee6b0ae1cccd49fa928a790808b1048dfded89da6f05664ee64e3708bbaf146663da78efa0cedcde7b4ae9d30436a9d02760f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h1ceb43d0f4933e84f0084e70e704cf2f1dc4a3b5fa3606b2a0beceb4f821aadf1caf95d3d8b4701dc229e854500032080b245f73951d8190adb760ee3b472c1f0ede2d3a7e8c47bec15b0d7185615d2ea9883b6f34def8f239f0726ac34cab2b2d09d53b8191f51567d5e55134f90a608cbddf0922f96cc5ac991670cc5402340cb96badf30c81400138c4170a577d8865d232f75629bc3fb1e83b7684b1715ae58cbd4cb29668015172a715a3c35831c2e78b4f720cea57450282bae3fbf6093cb0529e2b9a90bb77e8cb6ad0cc1de9c15ced524864f16e323e3e5b2951699b56f1e8e5ff2e6e2e5d9c37953fa791ff02aca07d106935c5492177f8fd6cd64d6884dabb4cb0cc30bc06e818e7f5b6de2e3177634b5fd684fdf962ebe0b5f1b6f623fa6cd0602a8540b9e0bae04621f974c201133520401f35ee3728ddc8423a8f491a3056cf184d877ab42313cf9537f1bc13a323cc3e7b8d038194a7f3872869641ca751e3e94ab86593c951b55c94d2caea4c935b98cc8e4287f4edfb4180a864dd7c81cb422e1394cf4e5fbfbec44c7c783e44ced03929b81cca2762ce0f603fb37a872d01eb9c5c88ec204baaaa2f05707af6fa9b16f65810739f995c81db1e370933e0a772537bc8db6d84b60375328859d958753798b3985f160d4ea34fb2e4ac55c9538191d6bb73c8ab0483ecb9039ed24bd957910cebee34860dcd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hdd6e87d2bd11b6d5ec9dca20609ef6b779598ed1201a395da3f500faffa886d4be6dd98dbcb65fb5cecabeefe90b523b4fe4c1ab99388e3f6450877f5f617bfb298fcdf921b8132c029bd6d1cd914b9653642684fd5de5c2b4f08e8813d93fc8176f30d4ed1fe598bf7c154c066f0ec7bd8333d0259ccb13280063ac7d0bdf7ec47ba048506030b86119df1269f8b067460ac40a8848f333a99e447221a4ddda13b41327ee08aba4e2d69523eed81bb36ee511e63b320b0110d3b10840f458eb7ba6963ca5b48e7a4d5d910683a970e807e50b4cb6598538db65ec2fa798bce3c930615aee33b457a48a673341b4da4ddd42188bf37b102fc9666792a2a21d14ea7df5f0ba1fd0818ccc97fa60c765a78291878271911f7fb64f157789fd78fd9b9961c6c8a400027831ad98c7777464ade12edaa1a1f4df3666202327adc6753ffa3df73676be905ca4a0de30b58ee5e36008d3269b8de2f63b3e9b73dad96e9128d57d18b126b7a19b1dbfa7589c781f1e55934293cc993b64b65cbe2723622333cc137760cbc9de3a3111236798741ddf81f4732cddeae1a3d48464416f643e83718b980f2a09117370168bdeaf5691a49d1ac439a05b14c90ca674206791fb3dc5b7a4f9396f8b0463a03d7076ec7b5d5e052840fdd1b9277be48a76b4bc598c82dff593a108916201e079ad496ef165b6d0ed57ab972e855189c7d90a0f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h58837756103ac72aeb92ae1a33ff6aafe768779bfb8b8b80c8a1953a319eaf1102ad3d49a600730726e7baf8e9566ba75b08d3282a1df98727987255e8274f37bc0ee0299fef859c789d7b0ba5ff5efa227041ffaea72b22631e35e448f77145637bfc24350f4219f1ca5d74de180533d704c6fc69358636193f9a02b0b241197274acedea5f7b0277d62b476b4cdb64324844a24c56685a70ef2ba655cba1ac4443de37e32f1dc3f0170470bf50fabccfff97af2c234e25f0dde34debe8abc6be405a66915b67c84dfc67eb69123dac12655d21e2a0ba9c5f25836b54b498a9d9c4b1ca6ea998383410e993927d15a1db1c4558d8ea234be5cec02f56ef41eb1b87702ba43d29ad052fba0a12e761f2cb972a5bc88892e5b58bf5b953827eba2250d4883b108666e6468330048262cfe0a418484731cd4667a863e853b604a4111c563664102157ae5e7929a4d2559345a0f3b4bfe8b5b790fe256beb2fb730eda95916055fee3fc6c43c2dda528f104c9216341b45619ef68cd60eede394f622c6a45bf8cc80461e424dffb1a3bbbd53d09553dcf58a2615f1318585e48d8a08175b1b345f0597093e946e78a9b0634abb2e949ae10c274a42b9f4c1870f26653471126bf9f80cd164ffd8c04e1b01fc17c2c4f7755a504b490537baebeed7cc95df3cf98b0142374db45430676f82f3bfb9da746f3759b47bc0212e074d39;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf49f76ff6a8a4d28ab07a43e6441a9eb912d89fdea1d947c1d45ddfb5c4c2845eb7e18779db4646fd675c9daaf9516b88ad61b87b5beeb3bf84786ca270989a06f656cd5aec15b4ab466b25803649f1ea1e266e1b0b69f5008230ff662c12300860d08e71d36648ffb67dfbdfcca02ae13e2e4564efe77deccca8bce413d337f315d1295c2d8f74ea57b97d51d26e04ebc81d26d79d87bb2f26f6086fa52b8fd01d3d4184952a631fcc44e97d5da96a3fb8d79370e5b9ef20b7b1a6056b54af6561aad5330fc9dffa6ef592f6f3782d7eb5860b589570a03338db49050456b67babf4533291382f3b316c4054ec9a2015c268e9032c6e6a9897cf3970be0ee71907900ea9dddce396fdfee814ebb8e6a71892510846c5923cd8c7fea2c2a55c7d230b5e8c2f38323b5b05c88c1429dfdd2280e33ff413827d98388e46c1cf9e381cd75092f554915b74faa86efcbeda730ee36da62ec551344ca806f42fec33958a547051468411e957ec032a1f5d567b1604ed39b556b1eb4a50f50d5aad752eb98754e26a21ac7fe5ddd8d02eda530d14083a130dd351d82e3d7d1c7cc520d4d2886d579678d9b072d936d967399d4c469f10b1737a6b7a7156d4c2fd679e26a0504eae242a3d3f99192f6ec4bbbef926e87ffd9d61fc8e9f239e416bd8cb1fd4fd2b7c87fb03f047feec51f27d53bf9b7e018a5e74ae1ef4224a7e706c29d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h5b9a9067b2cff3d3eeeb81a6d32820df5e06839ce6a0e477cf70d64366d43f0812ed9f4e5c498a1dc13b24175962c97a3621dfa0d764311be7cff329556fe9abfa191c2c4026a80c43fb826831bf5d6d2b57cf8add3d583d65aa1ac4b61389dc9a2e50b5ddf7f119e5599ebebeadc0a9a0df295182019fecf3e837dfc6d35271f751f4ad7a3a3724e84a39dc412d02ae0e11093d2fa913a41bc5530f63be62ee060da6f1ab9da0d7e74f4f61a0afb794537cec0e580effe5eac96b6d3d842ee25506e0b7620065ac4183d17b80beba40017be970c11e32c56d4bac334579f0062985bd4173055a15d257749abcaeedf5c05e9bd5bb48d05adb25022e30bee00513ab914659720a0503916d8fd8b76516fac907ae8cce75d6aa957b0a4a83abe7c5e3080aff77d68fb70a5adf6a24cf9976f23f927bf17d8470e3c2b7e74284df93e37348b3f013d92947d038c93f5868b461e0607dc5752150ce23c96b28aff85891c71c620a1f1457f885e90ad2a70a3c5796722d0b724897d6156db200e233ffcdb4b7b87dd97a20cc8699505c248cb123f200ae4208be5e4cb5350473f4bc5637c747dda9bb54e2774a318486d6cf53a81d25b3e4e82dadecb5de7be30e9239ada95dd4980757ef2bd79835d811b3aefc2368d129ecaacb86fe96d2ecf07f24f6577152c317374d30201453f711ce41e4db4bac1b675734267e83f3ed0b2e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hfd577fdb324cf8409a5c75e2f9f0bf56c06a8e77382b4c5fe273027e3e37717a6540638bc68f1bb652ec44ea24a9a8327d4ad5b14b50580572ada7c45df6732851ebf89893acea5406a3dcb367c86620b3251d5958bafc3206330add3ba53be3096046cb211725d8a89937cc5602c9d0aca7cf67d08b74e6b7d2a42aefcd3439a7779909a908d9819b27d495b0a478bc9abb05bddc31164131d271ea33259a1d9d3a2d84c7abbcc9ee5fcf9ecbc358637ec69ecca0549a477613f50f270d4b5c522b7f5f3756a0d00315b67a130e70cb6d717a14689167d1d3b7c3e1c5728c041784ace3fecfd405cf2146b80888668c266a9701c5e257bfcd45363fcdb07ef466e4641e1597b4d4f02647ded411904b9500669194adfa30c045a1b034cd27911fe0355aa199285d649e5b2e90d206fedf2dcb1f9976628a65deba1b690dc649385900de6ae8339e3334d3f7a3b667008dcc66bef36dcf152658489225e76aead87079d5a92778ed6cc261069e4a1d0841980c4e2c0dd4c49701a9902800b45094c635369957c1c05555917f3d1b08dc15a81600a2b0fd7e059c384093700c16cacb34903395704557636ddaa932cf7e51e042d0b3fc434b43c354b9460e0c80a7ed303056e4c4f3bd86d954ceeb86555d43c97038fa669ae8904cb797c2d293e35fb59fd91e4112b1c61265c8a02be80b465bc45e8629e80dca1dffb7828440;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h729f0b2d03ab0e1223283666ad435b82c1046b6409a9b25aae4108e04f0d665fa761c3702e139a30093db08449647008f1ca564a462b200f4a1308e0f6bb369678204d56e8dd01f4c6ff729d5eb1a8dc404e5ef1bef1995430b65089b32cc592431d2125475319e03987ec2f82510029acb5253cabebc97153ef0f322410ee84a101ed8a183e57fdac856f2d9d6cc56c1f4512a31094390b45e8180896e93ab2c25f47316ec211ca5b25eae7b2580f092b8af55f830ece888cf5c736ebfd8c7d24bbcdd069b6267ce7873134c9a0fd474150cb116a38c4b89c50e9e4c04e59d183883903e8bc5acdd6ce5557ae1a6902422ef1e05579650fb11469ff4349bad9bd3957b75cbdc5022b591b90729781ae107468c549d99ce525abef083763924a274f1ea90fa5281fa4d676320110793ec1be3970e4b48ac9cd7cc212aed7c2913b01378c343c8d44e5b47ec713a69ccbb9a8340c30a1cd4d0f704dfec41023039b8812448891ddc95bbbc140cb7ea901a42324cdbf1cf04f738fe97b6588c5881d1c8fa58dbb5193d712a2aad393068a7b94b642a30de45718a69c1a0f61abca9d6578e1ca4a9be5f4f9ed1e8c319abf2629571ce455efd97b09425b6159b9ad59ee22a890c344547660937380b91b73d9142420a1af628d3ac6f457588662272bcf2da18251f7cf3ae979f55f7b5aacc9d2c88a825d5c70a7d1e84828ae380e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hcca79086d7df12caa63b0546d5a3287acea7f9d9147fb4187850111795d6f233ca35c1549e5a3ec6b2c87a233cf19637892d864d4bb73ca1b7bdb62873d93dc00269ba7a37a38cfbe13ef52f643fbd53b751f1a149cc77c7b24138e49f54dc33f4fb5169fc1698038ff16b03628a178fbf03081b7fc5c99ff24f75d85fb0146ae6b2f79a4b1257a48ddc3df47f21d765a32cfc0ef467b6f1b705a47b687b0c59f0f22636c94d5e8376620ea6a6b06886507c02427e33675a6fc180fa0ed8e6a716e800b68f9470ac4916664e9b3e8c542cd07f9a1200c453ab3cdd0dc079760ccbc98135317884f8e6697d6529122ca9ecc37716b4720855b301be8eaeab03cfa97d0f127db9c950b8eb3a47f09b988fbe329d4683bcb5af384b54fdcb07368734b4bd5936dee11350ef465458ce279ef2a3af2ccefcc1cb56cf23bebf7fcb3f78fe1eb632f5540a86283649697080e41b8c5cf912804880d3e4eb82667d3e5961bcc0d84c569d5a06f874d464b853ed401bdab2116aa741dfcd1e6730b047383a240f9387a0ca3137261a460d8afe21b9f80a47583f74932c107aabdc8d5be31a6d9e9a7ca0958544b23f2516d326b876afdd31c32afd8cee689c92375a0f1ec05dd4996856e7ed6f3c5c9e5d9c96ae5abba89c6eb9ffcc40d7512cb58e98b8380ba11a2c1fd9f2bff06947ca892dda5d8352118023c7f84ac3e2952d4e5147;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb115023c0c51cd172c491bc0a20ca51121dc0498595a651ad9afe559be65e233f1216771f8c96f57a9ee5a78185d90712547ac3a20a5ccde351f35105444ca36893a8448672422c46d8b498bb12516e94f62abd1cafaff8e0b2b93deb774445434577df80cc490a0c90233e38cd310dc1778ed0a1a7a560d8b832614b36d9724c9f303a2fd89cd04daf35fc572a12255a730fe40c83bff8bc54fd6aca313e3549c828d37fc94f6461ba7dddee16b8359c612d065c1f96f05d2cd69ff2d4278766ccdf3ae9ec3d6aca7a847d4d0a4351d38014dec5ede95a4a7526db45aee2023155f684593eaefd0c55e3c5f38d43967da35e6b380ce33353ef91cc6109542595d033ed0c0e4da5b6019cead2803fff95e1c1aed450d72473d9b7571e929efc80f0e3cde309e7b4e469a6c2bc0c2315a0d03c6e4c929e070815ec7395b50791a4643ecaff8ae5f032beabc86c9227c86a92d7cd9219076e938426b09fbdce83171a8b6c904c6cfc7b1d292f9c71709feda71ffccea78f5f046387d174fa0ed3f796fc01203b5d278c8e06bc14c7e67003a2e0f39027ea41a59fb04797792420851fe320a1b981f5c3d6c1da51e7f640b1b749914e1ec96de47924334c7d6de88044fcac7ecf49def7573e156ed0939f25545d95574580253f48147b7bada72ba6804a82ddbc208c65be9668c51e0ad70df323c40c67bc6833b843e8e98ce19f1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hc5e6a6391618d253c54b519f9e013d975c7557f349d8e3f67d79f3e0e83381bc6a945a1e48f25816419d553b179f88245bbdd3ed5b4cdaa7a0f069f5f6d2c6e3fa0067f584de4a06f577fd4e7e21c9cd11429681b9c83fb542d3d5b9b050a1c7780715f11aebc1fc8071bad60eeda62977fba93956a47b0788532e9efceec69a1f1a307748b9d6ff2477a757ba379d429cebc969e80f077031d49064dea4dbf3abafc96a2beaf33bf6ab7ad91e369571d7d2f17ff2022cbd25c30e97bf34f4e712548db1f522fcbd6271688ee683fca1109d6c74ecb4cfaa4130e976917a02520eee5b1d06134f3e57bf19b43b52573e82b76f7812f52397d38c697d12d7b69fe610eae1c773d25a0f340eeae9e282aaa57fa35029eedba18fa309ee497cc6a8c8f09143c956bb5d3466dfb2c600c825deea33fc991a31cc7364ec4c608ebfc973190a05bf64822c3b2e5d62e6d7e81337c2bcdc9f81e35311a56d764007b593a5ef8ea1c0d28702f5ffb155bea4ba70f7e687192560be574b3c2300e8b2858b190d766362c739ac6e7e9352d015d0b2c308a42952b1e0b0439feecd752c583f09e1ef0559676a752b76856bcb8c2e3f0e3f3c30011b2ce17f3853e9cf9b3630cdd5b6ea0a5f412921b14645c6e5118f8318be65eb5b88a83ab5447f77182026af186f9b658d205fa9cbf92da213e98a97fec2eae8ed6d3bf52c21d097c40b7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hca90efe7a8056dcec8c1511423a8f5665424db8fed3518dd09a4f70be193d90706796dc1e29cd3ba97cf00b986f657bb7ff8911112cdd62b134fa8b014be23c065ce2f64f4b4709f2633e6d7b37552a8979b794128177ea63779ad2dafa01486ed7e006decf7f716750f8004ab5d011c19c28258f6e346b8457d757543ddfe864b2773526189931d05798d6a31772941e98535d5608a33d21b1ccc4439ec074d7d18b2602890936e0ae4d33df81a7db5c5f3eac870bd6023bee2e4ed8516808e4ee2edcbee654c677b0bb46da59596d08b3a9a1fb23fa224c98a508625d08eca4ccd9fb15060cbedc506384780d0a2ca378b74278e2bf8df21fe183c39f6fd00e365266650068a2bc00ab4346e18409741c7d4b417f9ec8cb1fcf75c801b98724b850b845d5afa62785fa21ca76b10ea1e99a2b24d366c5808cab9210b94476fcce16532ded48e1e2ee094fba76092cc0c5de9f609e696beb2c50a03ac48723ff2a89d084221b0957b14e1e4e60f32e491405dcb163b42a7c6f69609c9b950b5b99fdee6c4d5a3dc4ea1bfdcab59408c6d68bf28a2bca2f05459cb76948d35e95b7ca0bcdd139228105e4a1ab131747408c2f2fc92a7df6a748642573b9950a520fb243be9fe1f99b237182194a3cb8aa990c4b3d4ef8b7decded9ba4eddac55c0bde7bff98899b56ad6f559e0e3e9f6b2a3290a974acdf3c4bcec75c9d5bee2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb83356b28de15686159dff0737464fafa8822bf710ba5147aa52fb1ea95871bfca710480dfa888d0f56a663ddb07a0c06d706b2cc7ba3fbb52d52a2b3ec05aa4e0ed10134b899886e508495b77eb57023adc5612d29443509c2f688ce8f26335af7962565563dbd673d93525a48c7841f7515286d658566bfd7df6d038f53fe120ae5b17aac1e9b0f217c2a7af0030a1e997f017dae9b8237232170e011b054d5635e2d692a32fd39b61f4371a789514e80e80b7bf79e6f85a487b85a842318447ca5afe3a8104770f87e1a898181cd5f7eeb9cbb11bb11c433c83c0a8913c2bd722823d0f131237fc618663f841c9e17fb6d55ad061a2330575db42ebeee6a146e800a152473a600d805a3297381ac05f0a4d106855451c4b08dac87def61ee626a508a11a418da9eea7942da216a697561de738ca35596c4c13de85655f99d098c408a55073c761fdaac357ea0afc9182281e776dd97560fb05a6a4b4719c45589a2f7c0be22feb5eba448c0d5666887f1e739517a5e244852180c0712bae97ac1b47f18a2ea25dbc948f4728b7d7171604b0396c5d961a0d70837c382bb4c07e13e491f7feae04c67e847f923715571924b28137999b4c81e5cabd276225fc54dd8f0000335d20defbe3b863d33d070b614e564c2f6629f5e0183610f1adb357f682b1870f8bfd80a5503d1531efd2d2f552cdcd76e49291018b7e7545b88;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'ha60de9a5da53fc6f7e6e8e00d778540c13936152cb19f137d13c7f9429af48a8e73c74a7da35ff0e62af81321370bc36d7d5d122d4beb1101c9fa60dd8cbc6eef0fd1b8cf7fa7fcefcc9c6dcea81b4e9eb6434337b6f054972601cdcbda754e4a411f1701a0445bbd702664e4b38f515cd27ff49d8bc3c33edc082f39c733b89e02bc8e8265b084c458f3ac42309c315fe9dde57ea339efd77aa27742cd7e771d71874cd23190539f52d4fb2341fb8a222620f6c160f54e9ad3db9f645749cbc934bf6663a25ffea38eaf3b4190ce7b6f171dbd30a82216c43fe1eb8c8f5d520ff2fac865529bb24f0c0f45d1c9b73cb9e067b84fc25ce548f5f9461f4f8a9f3ea0a25e426cdd55a21c92f3b7d4ffd8cb479c33626ad2adfd35401a5c8cf86aed6431582bcbba461314df2b73507130d5d25c49ab95305c0ad783639aabc777a397e7162581a00576a71b0d3523e0593a9597234e1eca1e05b65779bd17cf5e59f4113cd3ee09ab6875cd0244371de2365b78e693ee8ed6bc1057fe5eadc444f8b12202e52202507ff461f91d19c4daf9ef55b1dfd649eaa4c112730afd15adaf760ac6dccf37728f4940a51c123990fc7ea944f733afddb3de4d696966e5bbc4dd7c4aa69861e1b8ade8d05d9269bf416a75c2f1f258d6bb50dd8bf95b22cd0d8cd0f3584ac57bc432df7fc03046d38e4109cf72193c02ce77ee0436e8fa3ba;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb56329345e432b3df1598d8cee64c1afd4ff4ccad7c4b148e07642aea7983af02667a59ec75379148ea93c930a0b4ea344f29347398eb39714b76dac5b1ec68d81b11028aca96e0a90460bbb1b7f97206676f80e40da0b55a243936413db0613417b9f709bd7ae7a109860534ff278dec979100dfe9f3d14781abd42be139e2c99cf09b5ca9756fa24740873b209a6e40f6fb4ea5f685419d2457aceb27ec8ccdbe097b49579ac5494e3ab2f18c7a384ff3d7f2b54bb492c43a85889321a5064338f25b99bd23e89e6e0b54d767ae5f4cd74226ca4b8b458acedc3848deaca0c38796bc650c4bd701dc2189f581d88da93f62bd29fdf2b07b56dfcd7f34a7590376647d478b25a03ab12935ed40be1b16a10b43ecbc978ec0867cf69c1f8d8802fdafed77ff266574fde9057ce1e6f03e89b3111a912b2b656398f149c2a18c5cb8c9482b7c556a80d9569fbd1453810529e881eb796157d3a35c326fdde417e7387b41775c671407e485391b95fb701ccd8340fd28a0b8f29374ff3310d9b681d45115175902d7223cff06fbbbb04b265946a1f6f0b4fd329bc9d1691af65315b6dfcba86bf9ea38a95851845369fdceaff7ba629003f1f07e37983d77c62dab12d7eedaa22f04ed945201ed65758d80eafe2c0adc8dd7a7ff86bb2448832feb727f12b01e751cf0aebf43cae7276d7a1eb55d980c48abd8b2b7db16abfbf86;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'he745709a227275885cf95836d2db28bf66376ad68d045f791375f62d2f1a34e97e5834844e37d4f70260f1607f0ec2f5d7a6e854884f7d970968e54fd57b3ba0aeb5d65a5fb1fcb775ce3817295d252c8acb134364045621cb5fd0d215e2e8630aa9f1f25db39f327a061fdf8d383e0ac5a26fad0352c8807deea7faee34a0da002a15caaa7299671fc00ff1362e271070a82f7ef50a84161cfecb00365839d21634f79f73496883d1b08d30caad3d562b01b438ab9e847cf5db12c25b1d5484c227d71e20fcc2acd16f3461389c9d284dff1d6f0550cc3d77a47e46742632a207aaa38951b3f5c50a017484818da25a876fb54564a87f8c61c29475bc76c6ecec068e0b6fddba28a27d5290413727d59a2be542e48b24331c4259e0b1ac5e2982476d33d9c4bf4ff8c54457faaf28bdf73fdc237365f70a00f3b55d1edbdb2503dce529d56c093c797adbfff9220a5235248e5a9b4ffe90f2b977ccee7fd7e1e949ffb9fce709c98b1f01ed2b5cf407a6e31929138b308ad312abc97b22971b8495e6b6188a89f98d2dbfe369434d4cc15df14e1212201b07b289f73ad00fc766f1b37b33a847dab0efbca30463c7eeb58e6a97561edd685c46344556eb552f58ddc2b6d8bef9bcf1b23fe0c2ff2d97ab14e8cf3d5fb60e7920b7a682b5ecc9a40bfa7047aaada59919d5f72aff979571dce84d8387659c2aed09826fb52eea;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h804c72d4eb2991334c028d6ba411ec383c2e79f107a2459e01fc3a357f0f63c8d94f8e692b5ee92a612d75a0f09af7bcfa15e52bfafa919aa23c666c02ccd5977c096fcc8ec3a3e73b7e3ddd3c21b541932f677e56788ae5c54a9cdb389de32efa14dc7ed6ce27e546a8616f1c194d4b71d7b06bc1e2f21a2f39304985b15a24dc82bf7f78f3a01e4358e0ee3fde6c1d74ff4b374667f2e6e962ac9017ac744425db0811e9f41a1dd2500dfa5899c52eb6b4a4f97a4136ad26d5bcf6f794f24919446a0ac36fa0a3bf828d5ba31de5a519ae3b7e03ad565c21c5f1a39e47961d29f16a8b2fc8c7e601371fa99fbe09026226076da969643d2f566e0fb94a311646fe1b63e24fbb967d8f7f848e40b5708fde6e93426bcb3e23c5d59baa9e7c51aa4be3b938d0620deb5fd8b82df1526da03cc800c98965e32b79864f891529bd911e48ccf2a2a5ec3936438ca3d0307a1e3ba480499b6ea58d043b8c345fdf7354ce8421e8bf2079454a78556b9554494fc9b131730dc59130680a229b10c00a2ad8dd69b05d5a8f2db22d4042cee21734ea4e73862f6a9077c0ab5b800bbceae7cac5a5c47d05a2c19b7932b36ea27231d4f898120ccc513b9c369d8cd03fb385e389768bd577d4e3e8c37ba655fb15d626d5ecf3befdf86787b43962977a0d20c584ed7e6f10343c772b740f00f281d6a544b116cf222a033b1a14fa23b241;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h9b38bffe9a69431d8d69f456f4a4178cca36389d94fb9039b7fbad43fef471265451e161221a34649125680e856438108ea740078fdad7df1e8d83a350ec6ab2988ba32deed9deba69623e2098320b9cea5dd4d6fee8b57900ba8dde46c96597b411eee9486898566fed72c735cccdbfd985e9c3877ddb41124d7e617833e987d0d40e334f6a9fa49932af373a5e3c06b00dc794043deaca3f5087076e2e35b7437ee32dad062ee711273ae3f913bc77b1bdcf982beb219f6937d598cb15f366f805e37650c9a195e459acbc25cacad2e929aebfe292c592eabd0954346d82fca8ad1414d2761c67bfe297033dd8570eb0a2692a144ca25ec77efd597e04f465498d864dc737032432172766b24df21c674ea6d656f6ced447a19060d66b16785d3268cad5cfd435012c4dfc64cb6311892d6adf39d989a9e92ec86bb5c2d725e8fcc829ab514d068a6c7b22c6437e88bfe60658c1eb3d130b19440bae3e2a55488119ad8ab3b13d215f5ca3fe4cd567d6fead392cf5c1abf3727ce7ca73a6274e1f495e4620813d111573203d93b8e0bcb389bbe4faa269badec0f884742fc99c058fc0628be7569ffb2b06416efd5526d1f1559d2c25c38de29cafc200d641d74c2d43c0e8e3706bc70078b7bf9961aaa9ae2221e02e3049dd5961a8fe9dea873e9aa07ff4df6080ba0aadcf2b89e4c04136b779dd601409530bd1ebbd8d59;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h39c419078ec78b1a0b0b01cfd7e74e01e68d21073c08d9cb4d3d9e1adb760314e408efd7f6832f4fb6aabbdced153286894b076169b3db4a7416bbeb1b0bd66a6e30316a34db43ae6d99b613648432d67e1b4cca62c787803db865e24d0c2af353d93f8f6b7b8f47f10cf6e9de01e90514db0b0606a0b8961b36a0598aa0cc052c0e85e15d041a19008d3180a038ec0750158dd58bc1f042b9d8d7b6842aa7174bce2ad26407632d94feb37d107a1131a08bf21fed3d80919745f8ae66bafc9327d7b71b7f1f809e36947a589884306405ff52c7410d7f5ec730832f791311ba9b347e67db09922c226bf6e08226fc46ec6ce1d2139c84a29dc0d37dd71d3ea8140baef1a9e661d3e6705e542ff19f72c83e92d26f546b51d56c0157fb9dbac3176c4d6b00f3b0066cd4344a4174c1399469b77784a6e58a6411737deae1ffc0f7f30eaad97cd20a5102a05155df234ad1a3fd899d7fdea903b528c8f49f44fe75bdad94121d66a9bfa706e9f2f7e0ce01b53e143a47b7159d966067fe6a22948e89376b085df7763cfde1a5aae7e987dfb435115698eb414e2b46dc7fd6f6ad50f795c5b1b51127b7aa10c3124d33a624c8a32a34ef21ebc9e83061d1c8133f82a0eb1851534bdb4a2e1a9b3b1c17bb72529e3d169cbb89a3ba59562ebaadee9e76b2caa2f1c513ac7b54c33cb6185e432368df153704a649f59a894d4d95b8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hc38383461a775c04ab161746736b9ade26bdf4b713dabc2c7bfc8259daaf644ce6be80ce8c2610efe147a98a5c1a15807bf50d0ffdfb944852ec47c48d51ab59f85a96208e550f96a941513cf44559755da64cec2e89156db8fe1e18446f89b5119aaa4b0adb82675f784bc12ffc34bdca2f8312a466588714d4544f8008104f993cf643b5994ab4f664e2a48db41b8766efcf9fb7aeb0b5467872d04d30a40ddc05d05eb4cfe314cc4f16e72e5aee6aafc30ecc273b01fbaf24b91c5484b3637f9334d6a14c807c6047f1831b6dd43b94c28a34149c6844683953cb57291d0818389d29c481fb723856f04d2c836c41f310d5b002179ff0a697c247036582de1c562e2dda90a40d28995a8ff4b53e725e966fbde8f8ffdae4fa8b2363c3db5c0d77b0636ab2caa95be1e2d4fccdf9a070f4dee0f02c67bfe958144144b66d352225d28912bc79a1f83fa27ef94a4f13adb4d8e0ca846667c1a46223031de03ff37f09017b99fce628be73704b612398d8cec40486d04dfbe50da3c15b87c5caf0bf400caf401a3a18411aadb4decce34d7b09d18ef18ab42c24f1e9b15c0f928ee0f1320fc6e461b0eb91b2fb3f62ebdcc60bab27e7c651e00195043b25a872092e78fda29a51fcf639e2ffae1cd7f9a78c20503b6951a6c7fcc76f48083a7d46c3f09a79be6f4998c8f90ac6d4383f42249ff369cb1fea4becce089552cc2e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h847472b446ba46058833686aecee47c76d27ee2aab46dc93ae0a3bd8c728ebda30c178f8bd1aef59ee63d700a7ba44aa657df8469ec7a72d53faa05fae31f8a2b90e2c9b395a0ea4bed824c0240aef93d8f0c3c12f6e3fd0ffd9024e942fa2992406b76695942f7007445ea656aa1bdc78ecbc31f4a1a34248da0214bd05eef3611e9ceca6f61c94075b5edb31f5c043fb8cf3130016002c7216efe7e94b3cabe468e55331d1606b74ab6d2cdefa6bb79be17030f6209486df65d9312d270bb4033fe081d7778389b16d14685fcecc7558ebfc1840de96b5bb6091e79719ba9bc6d07f22b70cd3af8839b527fed809040beaf12daafe8263aa4d5dcbebb666ef8d35b031ce74e8a1338ef5a581b2a13dc4ebf0c052b4ee2195db124b522f8da0597dc719f490edddf552c8ba644c667b87a109d79c8531733a017b2a142e3a24be26fc13102acf9b4dc2882be9f34b5f1955f5132a68fd28cae8cfdf8b4ec885df0044f8695f8540412b9bda528cf599fed1729e54405d8d597aafcff7cc798ce2ad7ffdcab3171841750a496f95027d2d56b7c30d78d7c74e5dae66aef4c28fef4d80d53d252c9b5679f3277ed09c37b302d1f700046cfe79bb7ac70868731172a951d2756dcfad17b2ad414f5324c938d0a7069972216a0aabd249e3c8289125f5f5040312fc2868658d29cd5c32813b40ed0169e3586c63616353e565fd1b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h346e7c109420e79c5c1467c8e8e65415c5dc73f18544535c7e5e827c6debc299922ff6e86b6a3fb2a9a83a6fc0b7bad4b25fcaef94e48db04e6e5188ae54d31c2961cdc1688d1d050b505472e588d0b543ca1590dba50204b4e400fedb8239a72386178ab0f1d61dd7e50b2b091ed5f2f7f568230c371ef42488db51068b74fa166bc5d20b0ce108bbc35f12a5628e6fa7201d8a1b4e298d9203889e160b178562b003c69dccb9232a2175e5954391e8a5049325be9708565b287d524311463a65bbe0023e3f559fa8824be07a9ee6dc48b97295e818bcbb660e82925d54f28d31f33e14ef50ace21c6c6c2f267eda7e204fc6d0ced5ecc0ad7eef943efb350fb797af1941b177f18e764398a575dd16608d7fe9f0cc6740af26be4b5cd28d27a0a5e663d6c64c67f263b7ab2bc0ba6a771271f7ad185b9d742eaf29956538a38e48d57ba79f21e8774fa45460f4d0f98f3537c5e6618a55b5be71a5f1e3f3da2272ee88404c69bd0b53dfedf3a40f8386a9fcfbe580a7492acc08f23eb4e8bb520a71ec34beb4f14503115b4fd59169bd93a4f83002a61e17b335057ab108834098a04370ed0a59511d37bf25510ad65238b0faaf75ff533ad22054cbfb6cec99287aa1da7c30f7fcc8f69b63fffe3b5615eeea9682cb115960906bee1d0da5ae43a33c1bece2e09210133509cca27bf05be725abe87448575340c2b667e835;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6c8faa9c8ef119811c876766b80952695037506fb2a2f72e52d9bfcb9eddcbb933ed52d15762a181f0e26eb4b21967de6054ce0033a3f28a4daff28492944cd074b5440fa9241d66da9b6351a4a69232fc73311c8e679a7586de6fdaa01493c374afcb3c20bc97cd4a749efc07102886b6459fefa050e6f3358655566167fa9f81ff4a623dac6c818d2c5f529f932dde2b2b8b67bbfd83e9487b77a1fbaa971d5a45d078fd0a1e80327575ac57e6282394b031f75f7a4826a4d66a320c925bcbc26e9f19d941e40177ab052eff92931645d84ea0b22a7e44370a7fd9217878b436bfa29d8cabb6d42b3435a325fe129ecf1848b60ce07de66c102d8d566ff80e5d94e715855fdab13fb5e34b065a6a552e6b53d021311757c8da4da3537110cb0aa0d1106392b5bce8130e4e5f4c3528a631437dd49ba14322652dad9c63b17577d4aba9968b5bd7e2a0b66d9e9d675efe44bfb8695c3e779532d6d2d14a6a95b124724b320128663cc020baf600e2e8586160ea51211b55db5b5a06efc1fdea1bae6498b3bd688f7e675c0bba609d7aa3c5eb33364104f343bfcca9570efb036f74f6cefc42df5bfd192d506b20899bc8b1ff58bfc72a5b7fe651fad04a47a7361db14ab52e9b0f1bbb5b558b75505fe53f34f186f61b8e8d596ce5d5144958cb981024bf9fbfe3d32f89f1d26461fe51f394e8d852de6986359ebfc1cbc9dd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h4cbfb1fc1159f88e663e118a160df6d9a19c5fa82b7f07e3e4d51a5bb634e152df6fe7af75410a74b4f14e19430b7ab103a8dd78bb676573378fe7e3c602d05cffeae70cec211d9a1f32dce2331d0cb6a4e3ed5d191ddf5aa7daf97d0871d185c3622d6fef12f8333a4f752fb27f623b1e151ecbf8b5702037f5a3c8cfba836da329a7123b14efade27c86be6d49cbe182909d97008560815ce1ca3fbda24b1242c141828b8963abe9aaac3667758e4ef70200b6a14c7d04a290b8f53ea3fa257bcb192d3873fc2ea8e212013feb7019099fdb3138d3f1eac9d8934d8f0e56b41c5e6a46e76810216d88fce0f1efdc4e02509338ba21374105302663f119042985c7037149aa5715ceed0e363de307179b42c0a580bf65bd5fd319868e88d579fe73079ebd62cfddc22d82d6f2e9110558cc35179a0171813940b96ae581e7bcf3fcb17627074ea0d7d6016c4c282fe5739c3159e08970d0c9f2e24c8ecb3918d257a5bfbb89ea9c404228bed1bf4e34aab07a0dd0c3e9db6ec1e53f402f1a7ce61ed04998f75687a5302ed77c441d2c8ee88f5daa291cc1427799471bc5dd973002a1ddc80e1aaf5922365accee1319b8e6def28d11c012987d12238dbb1cc63bcde9230bf2168ac253f33ca2d1f61901b5f2f27394aebe518f5fb04ac64b0723450022c29923ce99a289af3308d249c206f4ac179fc3e3c644bad9fa7004c6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hec12d5cc6357e1880e35ab80ec4b4a5b339a6699dd6a69e714311180abd9513b2ef69e6424b90abf726550eab7631b67709e699a34534b23be986cbdbbf2e66663823a95e180f1b0b2d6ee31978aae91782c6c88512ead03d1ba64d8f41bbf6d31998a8788e0c2a57389d80cdb3ce88d16a998d7375f83bce31135ba562d3bc9e0abfe1c1fcd6bc1dd05715f574705b7d059ea599ee9f0c3c7eeaf3022ea9c8386ab972099e68097d1abf04a99af73484db2aa2d09bd95e36e8504a1db786fe53c3f46807b816d8d67397dba3f5106217ad827ea7607bd401e06992ad371c3ee0dbd5cfce0308a3616c826518a2dd2da1d29cf6b44cd348e42ea7200553f247ad8bf9333c811b841f7ada6aac18c7ef73e47f34b580130090553d85ced5381fcf37c88b45ad42f797cc69e76b3b176290ac374803c784af53f74034fbd34539d7968b491e19bc45bb16f7708360a15e700d2f51661d1fb7718b15ff1395257e84219943affeeca7009470f9c61a7e729523c95596910904d21d8c70f3c87637373079b37a701b9aba01d591d3b9b7a01d0c67abbd7816d41f9d28c1edeb441d2f4f60d66fefd8bde1edeaf484c97243b87a6ab69d3c14bdc39703b72560e23c1cb131b247b32d13ca2e7f2a808b6e550e3222d883115c9d0cd960695dcac404629cb5f10593fdd8bde564833f418ce324f509cfd9dc53c3fb32b5eeb4607350a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hd64742126ae94c1b41fcb831e72fbd3efe393654d9fd7bd0bc60f4d3571bf5d1862fdd3329e3851880a4705efa368f2bb9de6122765781d08de9f43430ea1a2bbd04bf4c198f93c8541565bb24f9e286e7ec660875972c25d7ea0ba00dad46a8231ae52f4a299a21d4e520f9120830b7369924255214d9ed34a2337550293bdd20db9322643641f26ed729c6054f6e53e19d9d3a42fa004b6c27f1d0d72bf5e80e57ebd62e3731cd4d8b1bc08f2db85340acd98e643fbe10faab3f783dd5e2f199151e4a477cd492104e1ecc7f14008fc100c78e47005a679ef6496765572cd7507019226279b47e705c98a5808047e69f6b758d8726f9cb0080bb0dda6d0f5b2632e5ee2aba2ab20400094b72ea7af39435a4dbfaf2aa427087d98152beef26afbc9625342ecc7d6b2d41643681a41583b8e14b350be427612d6f6270d12421eeef8121639188054874ca63c071abad2f60f0ef44e743b272acc1c16897ffb80de21fb2736ce0fdba4fef31d5799229365b92c06e8e5de363c9c5262b475d83143952d6d89f27652a9783bd7891244be81cf95154d9c3f8310fe3751783273ef6a0f3690af38fd24346bef279507444fc27f5406e30f3a048663dd88240abd208bac841694d929173676ca800d2f658e0ac6a52c2ae7bcd494d9b8e69d2f3a3953d3352da196cc3bfe647c83171a129d155aeb82b5276af10fc1173c76f564d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6fbf5f2f4ca594aa5ce97047ba7dba0609681ab83b69abec170309f35c5a13ac863d69bab1d7baeabb065c2c5096d8692575b28e1b8c151886f63a662ec8501ad02efeb689e74a0abcda9f4d58ae48e9a033a87c9b8eef1edbbfb5ed39e1312a1af33a27fb3f154fa69e09fbd5c8454af13854b5437a80cf8a1c013e374347aa5bc2c627e425e32d2c08e1e3079cdac1212d2fb3ab758d0203bd3b50d914263ee6f982d4ccfdb119279474f99f3dcc672445f07daad302d78065f2dd29a516a30cc75699aac18dcd1f5a45558cbef8bfa027035630e1b0994c296f45cee958e03c57520e73cd65b48e880f009e6aa0709ee38f283e9ef14e8868001421050f1db88597d6b51d523f62806cacf856df600746d84f7a898791dca53d0d5405995c5d33524605fb023a90a6321edcd59417751f574d655274e2dbcaf74ad52b769e027f3f84303817b13a0a363f6751d8b303a97cb7c4973536f0f5e8c29d1a3d3e680c750db06fc651dc9d8e3704de996c1b0044afc0ac75d907be58ff23a490cd46b6c04d5b2627da5eda49c7028b84f5e57e3a50bfd9baba83adcfd7e725372ca51cce636fb77fadbb6842d708015ab39c8d85e47c478a1a9873103f740902e9c809f945e590f924a36abf63a8903290f426b287672e8eeb07bf10c53c48ad7a6713a220fd710db4af35aba6cf8224c2e6a77384b98f7c2c50279c5287096d9c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h2a0dab8775acc187932452fceca9aa2924cbd90925f3f160a96aacc26f14fbe243eab7692e1df196a2ce5e734bd88c78983900c3438cf765a880acaaa315862f1f8a933a5f7c5d971f90f712cf7896f741122b8a70fff6cfe413c54b3eebbee119671bdb4b2d3bd511fe2fe4bc5264edd8e0c9820c5a853e3ba2c0c649cf933bc34ef8e0f62219232e8fe8a4d784a3d82ffe3ecde2a3a11f1791f86d9dfb7fa3393dd892db3d7d5b61f0edb152df7689c923f121cb940582ee0cbb1bf5dc578dc3f5563073a90679bfcdc2cf98f98cf2b8d6e9be087cd3f5db49e71b1f4381d283e0adf7ae6b4f3c0f1878509760dadfad47e4e50ad5475057517122d5e08f5898401624a988d79b82ffd779ab7572aa00a2bd3e30d8a29d5e6737ac14afabfe697c3743151ba1e0945687134ece2affce85891e7d3eafdb37922f6e77bb1ddbff5204d137f7565fd708220212fb25360e78a2e2f5bc61b30a1bfe52d16c9d22a029ecadae690572ae10b3cac164fec49e8575cc88c420224acb771b4c4b124af68773ba8efc3ed8c934b1691e9571479dda49c5421110c82ef3c244f151aa000d150c214038334b4ed357ce2997d12e3ba24fb90b5b57f999ad5fa87fcfcfa4dd38fb57c2fc72eb8d850224371314dd84caeb9406f7a2a267db68bc4c6359aada3d20c8c3a12a4b83c86a250f6d30edd332e5c244369bab890396892ef0382c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'habc0432a0e0b1f5528a64ce76a8ec1cabd872166f424325a594315fde23f05800d88804ff57230873b55e01efba30495920605ab2fa09a4949b4b9105957cc702cd52d8ae3757191a9b71af02b210dcae8b1d15f1006b1e294e63525c90230450f6582e469c9c5c4445b41bf8800b3b65d5fa7a65fd14065f3fcf30b415e2ee350240857ad71b973e6562f35fbc4c4e1b0e9bb48e78390304d304f643de52aff34edb7bc7423275d0458eca14572ff31fab7d286452665e2ac9d7e3014438814da368625241e1be2d5c19111edb5eb5eaa31ea1247f7fad05d212e999e14def12f92870379c3c26b12363dd3cfa70c200348b29f44c7378eb491bdc428489a48011d883d9e076d4aa95e44b54f8345d41995bef28bef9df95a2af390f4aaf811dcf564068baf5d4aeb8987f2734766e2e996dba6f75f470ea9a30b8d4d4c4ea788db567c657b63481981304753286a89a407cc3dacdac356613f25b51f309fcda439794df1ed4489d8b8a90b9be39eb3ab81309ca903a67bf364a89cbda2226705facdd95e2fac9e8ab053492b843a0504d9a90041875c579691a7f5c0bccd03fe56ea8c93680744c886ce7fc499f755c1856389ed4cae57852fcad20c974fb31f10d4378fc19a4b7231a72fe6a7abf5c5c0230f08fbd48a8acb816e61ae04ed621b63ab160339390c1ff9b1ada8a3e0d02b594b68680e15c4969214cd1de26b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3c36e6260fa467d0cfd4d5b9abf090e551a9bbff6666964c98b8881b2321d1aaec95cd9f8fc0173fc565a977996eac7e303c791e5dd65586f6862759b5383554b8820fa57ce5bedb2dd51279ff225b8412d7217361ed2f30e89fb9b4f4fe1ef79cc33b752f2d8e64a9790cc0d599e2d943db3dc05c924ee824edd7a99d1223e1cb89db0e7c6e4d3047a09ea11270ac0479c5fb8ced7301930bfc44dd0111b7f38420fd7f690f75976db2828321bcfac2d4bbd76b7358ce47aac0c3315e063a9a352767e1700033026e3c1cbfc74965bf8051e35042b78e358c73419e59717b81e3cd14ab21312686182c56d72c0410a7f898bdeca69b5118eb0746869af5911b877b4716d59bc4506bdc4f6bd760be98b222d9c3c07c9df4062c9c260ee3b788cdd6f632ab7233b1070464fbd9215402aa2fc178b5721d512ac5c934eac40795cb6b321522e0f85123b905498fc54fc5372f61f98d47c2531910dd2fce29917d0719f446ea4ece68dca81c44011b0ad44fc178ff73068c524ba56519d3b7fcd8f0800853bcffadecf65afa27772a442f4d213485fab619f4124fe2c630178eec0cf0bb90410047128db47aac1d6b7fd92e9badd9810b1fd0237125d6a4b124df2731b47cf9152eed9570891a077d9e7e744fc1c09fe603b9100de599588740d7dc3c02967ac1fdede00fe177c1351a4c6f6ffada157ab742f8b5ddb5050f55b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hc9d2a4bf810f9d604dc2e3c70a35103d81804dce86d574a22d69a0cd7add5b9ad725a47b7c63ac6f061959bb3ce83c2da61b1495a5cdf57ad94b56dc8551908599d97c77bbe819e08221ce827c9695f005b75ae281d07724cf2bbc8578fcfd00e3baab0f0ce1c2271f23e6bd01766eed7210b992b971a484baccc314792b2efddddfa91c6336ee17185289ab080ee108c9d5ce134a2069e5ed151d5dc75c6e0e28b04f717773fd343eabc92d4e760dca9f4f07478ee7399d436128ffb8eb10ef2d64c299e5d30f6fbbe43d3239fca5eb349d55b435e597f4588fed332979bebf3f648a2e18f37898476353dcb2e7e14c48a86f6490c981ee1b5baf048a7f6718245526b3b9bbbfa63f67442a1caa5262c670150c68d3a18735798a9a032a33154332a1fb216cdd3af5ee429ea31b62bfe582666401fa2fa6b68aed436e7947f7ebb3d3816d712c40770bb30651dd9a9fc6f0f86049756f422ff986c5389760bf99f3b93f5a0166952b00f408dfb19863a92477212eac4b6f0e3257959620da19029d11977a95b1ee4af32b0848f797fcaf5ab0677d7595ccc26de8e649bb24db91ad82503dc27a4d27510b18ce3d302c06a4d2273c6b9b42d4a66a910f9ad62ee4467b46398cd08a7f455f65237e688de2e8216cdd25160ea252c42562924689203f1a0645122114ea92a303592e4d43f9ac74fff35862b79772b360709707b7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h223104728c33196b5a839b20ac979ed36f3a4649b3a7b13ef2969a1378ae40f082c0e2aeb02e519e223ce3d272c953ba52b9a68e5b96516e16e7db8d56ebd75bc013ab14a88e78ef33a5fa1089a5a0b5a319b0a19f0f9b263d2e8866a767576b8cbf7d2653cb5a0e27bce5b8271424cd26ed82d86c5bffc35eb4a3aa539c28582802b3e6f7b3d3f6f97c49ebb6caa3db378371e31f14ac3d12aa7eeab268ae57f48a9f60c98694e278a063f39ec8dad241bc9407f5efb1dfecdc3368f4bc58255cc42c72ba17a307ca4621a4e46e61864f70031b1806192bd08d08f9fa05f392a469c610bf4bd4b313d6dbfe906a122109d4d4b4b5c523db4fe4cb30233e3a3bdebdd1961af79576f79eedbb2dff77b5154b1cfccf357c2d5b0d9ca575ec0c8e4a48321fa9f20e72dad1e5181b84f95a161cb94ff906d82aa37dc4f425ca485c054b9bc44c0dc19de8e1fb18e81c51e5bce473e9a910818854e83613a65a9fbf08c9e66650d66f2218d2574cc2943b985a88a724399e82b761919e43ed8d83d6c92cda99cb4fb31a68651e8ca3338eb45a7719f1e07c67769bcc7a5cf1b7c8b294b96b2228ae4799532c9171fd7da5d08e36c2f09a0e12fbbe6f31e18eb9d2125d492a8ef7af909d39a439dd470d19dd3e5f2ee5cb9b54176fc4d24d15d916e44fc5850c73a64a649d125e760a777affccd3461cc5488cf202b456e2ebc96dfa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hda15b7fa6158d4ba6e58c6f6010d368e89ed81fa850038c924ef6cddc34900685c201fd5960838282ac87cd83ec15ff746401064ff9076404b9077ed79bbbc6fc7b03e179b77849b2bae0a85a587282e7b16624ab041fba9c6aef64c5bfe35eea3ee931f3c28439fc6e89202eef25f835832e1ec5ac8c05ec09d5a0a0a3593746c56207a8317298b546040884dfc411e7e126014040437affc2fcb56cfad912d45233042a680c375ee7034694648c4486f3862b49287c9da53ad610dc022f678c7cd640bd6d95968f64cf5aae636c4a1b93b11209216eeccdb98dc218661a875926b1b580d1c1f332e6518d50c659c972c1a6d35fae001271f7ffc879c8e412390f85175b13015cf24fe19750e5c48707d49573f10ad00fa0753aaf430af4dd7af8a24a44e68113b832ccfe5ec9673b1355cc00d28a8a5e68113f2f3ee6171f7fade8d1714e844a5ecd6006003346e7eb7e753ab5a5e2557d18b9bf70573e564d0cbb0b46a396d372a37881cf218f0176bf4d552c45b7038655bb690454437931a839104a691f216fedf97a783689eac9793f06358e2670e5b59c2c3ad4f2ec1d706b0ce506b89ec9ad50df4036e5f98a25bb637499739d13d31775ed00fdb3750f2703ac3ce8ec2410280a531749f54bc2d377b742ad0f7a1c89aad9619eba3115e3027b6b441a65c39477f2b481cf8707cde63c58b1690f36c6a50aa5fb22c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hbb1124da795686eb5d614ffbee09eecf9a5e6af1492be9000c3ca5ba720aaafb75b5f2025f79af4bb4363bb2083193bdb35175acb6f216096ef300990607b08611562713ed74757c748018a7acfd36f40bfd0ba01871d70733f662371d22882d82427b032dca933f0f7bb417861fa747492ea7bb22bb9bd26a35849c92d901b2365340268e7982b5b9dee2f3e4be81a3b24ca4ddbcd41332343865bdc40fb39a71f5231bb093df2de17e51561423ae1db2f6d37ed9834f3676e6ae0822a5821ddad4cc40892cec3432ea1afed32f6c61117cecf5e2de6acb947424b0ac2e0a4b90ce62b9869046108e63a0144929a15ce2467971980537809bff35a1046ff2009a9bcd6bd51b8f74cbe6d5d2ede2c0fac67867aa63f5668a5f8a748d6e168542af854d58e406d377e4ef9121f2c189ccbee1ae027f8e7d7c8c422f12ac803dc3cf662a4cd7a0466b4cae54699042bc9004fabe5717c9d97f00afa2dc89b170032a51efd959a07f806561b09ef3b5cbc78a4dafeee90f8d34ad7dad4d6f6e7c607d7c406e2bf583cb3199fc4aa795d72d43706c3dc0fad823f7d5f1ff5aa012296676fd5e9c4fe2004f769fee8236e3d1f3bdec3796b664d763f538ba7144e7f2476a1f21c1da486d102bc9441507bf38365ce552491a5312e53119ecc8f311df5a6045b2995be32e843bec0757481b7516dd40ae99231f943971020aafe7eb83;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3020f0c6b2aaa6ebf90273adef87e199cc619cd28f286cc6cb0f4de1f28a31248dd29e605d3f6d4c0cdafb8ac4a063ef89f6b9e431ea94c8da9f4b72107ad0578a1251f6d0f4e4bd0a284dad3ad404b6bbbdfbe57d0f209cd307dc14de91562f58e87df30c417f85be24d0da02a87714e3709f1822d926280482db32609ed7e57cdd7ca133eb359cf263df6282b058119d65d43a733717c601dc4c1ad2582318f8342a50b75fa67b9bdf82a8fb6852e5faa6520f813d0ef1ee06daaeab454dce0e34d325f40b64866d9dd8fc355a64a3247ffc357ff0abda504697c109e4cafe25b94347c3a0d6dc9a997de204606e97177ccd0f2812a9ad6166c001191fd58149e603349270ccc717e1415b20ed17459cb6bfa1c0f2dbe1d447ef1ffd1986e4b70fdc584e8643d7120d0a9de9bf24876951ae174634eeb215b6ae116140b7d9ac19ed7fe5fb8af4b856fe4456bd0d81351c0e73d5f64f7343345fad9ba4da74e0d91335e507f042420a5c69d33655aed6c12513335cab7f48e0433eaa0cc640b66248efd22981438ab2f6a96e7c733040e79862639829853b6a51f13ea4a8186c052fa159f6ce7068c8a7e5cf368824476e51d40b0cc99374a7e41a7d6469f9e5a8ace31b7fd1287a98b0eb605fc6ee27d5d0fc1c84f624a6c0692d87647b16bd94048bfb413871e4c5ae055c8c3a4e678290a0497d0e9d44c3e5f2d7c09a30;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb4da82303e38947a2edd88227e8b80523e286213f770a4811426533c82c8cb0462def6048ef263b0e9cfc141e490f27ab449d293c0f2d773ac2faf0baa166558536949039e67f6000fe6467f0f326174a0adf6941c85bda67f2c96c1b6ca2c60c49d759a2053993948b4710479465d38e094d395acf9a15a20337e444d5689ce5a096a3fe82bee04a0928fa6948ac73a6977d2dc87f57ad617ab8618eb1f9239842942bec85fee854c47ab189c5dce5b7b64bc588efc2ba2198123926fae9eda1894eb7934945dddccd2ef8e09d8850ac44292996819666f63f6c8484a3f7928965517c897dacbd5940f0975039c40bd74fc2986ce9adc1eebc72536d215e270adfc48a3ae0bd615bfe5e23021c8716c031f1df67d792c0bcd9af214bda06d93b5c83bcb6fe05d78bba151a9ee07024315359a19873d5d56bd1d7270be22395327af5d80f263840d870482a4b568827f57f908740599b1b6a4d8abd4bcd4ec54b3800738e5cc1e04485035a4c2066e7910193a3fa903faaf9b8e764f106dc90f94022605630d5d2a973d089cbaf990d486ae2eed17ab965aafeea389f6917c79b6e5c06ca576c993369ab8e765c6c4d22de1b384a02ca8228bf46eb7b0311de9e3644e5b3edb68a6d01c023ec87f0d75fe1f36a3e0ee54ba58eb9d3c54d7bf6f86ce38b892d92ae6be26e5e96ef2ab4dd8dd5ed53fb3b8a31be11c35cd173000;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h689b03dbb3bc9ba0f5294e3173002e93ef1e86a41bc25c90a25108c5ad0fa9e3bfaf7bd62cf3b3bd71f9d1283613e0b4f3fa6cccc2ceb50a3ae213cf0e64e24d3edb371ce315c163c231d046a319d7ecb9738caeabf8c04e56050903602caeae442a0c9b6e12dfc9abaaa3d4e26cae61ed1c3bfad25c1684105bb12f88057ddc1205abf241b1f4727327ee48b0616c75f23fc063e97ff252002f4069b56bd5616691ba5871257ae9187449a95cdc30cf539fb44e6632c151262b0de4178bba83ab268e4ac0a7f09299eb364af49ba93adec0a4cc13de7483f628a24b2b806f51c505a1d81b65561fe25ffb1ee5a0be0e70a7fc6f05843c83b55ce0c9254d0b98ccc1b004814a5a26a6c1cdb11c23cc60694a383bc97c3430de8f36dbe8d9a9708a0913a9cc9028f2eda909013557395ffc9e54ecfd08ec4436b6f432bebdaca116a59099274480b8045260b7a16e24f756ae749dd426445eb8617bec7914e28b63758d30f62d9d8c156cb8a0173e57c305ded3283be6f2a5976d02b1df057cbb582485c9bc8bd21003e64e90dbe4d88db77625b6463bddace3aca4a7cc724e9fa5e433365d54d32f3acffe65a229c202625fccbd52fdb5efd788f2ccbbfa7ee5a4eea44ec07280e58173e76448125dc192b7615cf703c1ac254fc824fe16cc5c6d50a6571453ac26d284faab9dee2fa3b0cc822785a94f561e9845f0c0dd4c71;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h279ad26d00086c1cb5537dafb42ffa67e0808692c99e46dbff9009b613ff010c25b10d5cc51a5eb8355d7093379e7a3f7e60626b5b91e6ac87edf5f24df14e034655680bb1c2a9386875a916e661118fbc5a3cb3f032bb517c6a869c4a778f299e29f5bd50be8a64eb667e9fedeeda1869d342d0f177de529191c5979ecea38f13c137a859005d98d67d0e408caa2bd9eead5f28e3cc42c6dedad02f80dd3c4ad8acc0f942562d4b1bbd41da80056f55d34d8509b8dac3441422817861c49bd1cc69c1d5909f47fb76b0c0649affe3cbc6d867c6088009c3a3274a27aa14f22722ef418b5a5a7bff89b635e6b555c8ad652ef1679c0ef87d429da55d56a6c3455ca314d97e4b2385c3d96f48edde7d44de023393fbc8a8dfc8e65f1f793f707167bfda42316e2a55de8c77070e9925d5e585d454f6825c4d555d276216cbdf2b4a6ffbcbe7a85fdd9dbc3652754197b8eed333ec2df1d99775e2012fb4cc280efc7a1000cf6e226dfc60d5382649c97a2c54da70f08245ef5416abc3305fba98f79c1055c9a4611cfaf31f35f53f0d79189fddbf022d16779f66beaa55249d27591f51f93b2b6c7fc8dc4aa7d9b66121581f6ff80cec54e30f14a0c390cc354234246f9ce09ec4bcb0f9754a27105326ec90f63911aae27642e0a30d7f6100915f4229dc3b218ea4562462212cdd6c503e0661c1f53305be8aa80ec9c9eb39b5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf9063e8b2bf3a1feafbf5713696d401ef8c042d460862fd6e6c018a19ab53ac0c99882e1213e343f519cc4bf9e0d41d596a5ae3e37731580e4d5a8a6dd62291a56442d24b27f1721297b77fdef4e856ee2808a57d36f6e676cb857093079441fb75888dd8a4cea70523cdbdbea6e85fec55b3d043ba9402da381eea11fe5283d9811fb0383fb956353197c2a2518b593982190b43fbb9e5b0475fe42e48144d5b308007fc5f784acd800760e14fe71063dfa2e7af0749c7d698ae80363cdc0bb15070c94fe5ed568fa250f46330dc354f3b31095df0fe7c855dbee953fc53641c6b849ed389f3f6d0dcf061071fc54c73ee9858577c915fec868bfb59fb70b351e0665543f6091a1c687bd1b06539110e5e7787cf42621014537fbd732553b72c86698539ee3ab7ab53ba6d7714b2bfce42b642b2351a5fe3af32172b4f95569e6c8049ceb22d3ad963223ad4b135f685780c0204538859a0cc79f7de4aa1e5838b2d5e17705734554441231ed873fa74437f24a11398c0933f908477b731e6d5499e6d18228935535fc04af6c3d7059d50960340e13710f4eb73a2f97013f67eb42e1650794aadabb80339f4bc2c6e4e8be2233201f23c2b93d953a0bdc85dc2fbc120037110f85f55b04e2b38bd50d580010f41de3b8a560cba884e5c4ecdbe4aecaf4b37e014af14a7fd0e98a9b96b9930f12446b5a72dd3a226bb1e6402c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'ha8dada06e98281a734310137d2243495f97a9e5385c20701a199e7ebeea394de4aa4148ad01760509d47069610c2f90d67736308fe7bbe8cc0ff68baef7935fbab1a43ed59826c3ab9d228d6dbc809511e91f1fd0b96c37a56dbe29ef44eefa8400543b7eac963e668e61d3e40106e5c5a06a7cccc6663553903f08b2131d3d4cec4849baa0e23d78d3bf2c74a23919ca7c71c6c64467984ceaed297c6e81b4ce26a62a1a7bb044d8f171de7c6fcdf05659e1fdb4f59b079b484e602abac64c1a82ef5071345c11ff2da4b920717a212c52857265cd0d5c0c6ff80b5ef7c03f840cc28c522a55be3fcb5c99dced11f89adb3640432b991ea2e7437f29903b9df39b0ace7c317b5fbc686b5483242c756b068b473529fa94314a18e04c5e8f33e678587b5c8eb6c232f41364510e1dd0adf539e2ddf72e4b893033139626c9c9f44b739a0c28d82c08744ad9d327bc79113947eb1fa35dcbde38c55c2f6a7dc2a008b7f050adc48a82fb6cafcf3ec6c5257e1631cd1fc92077d217bf21611d1aa9fe208fc9c3d928123238e4cb0a05023171c804e3cddf5d27e09f9064941ff132cbb933672267f7abd2f1ff384fa3fbe269cb199707010a23cfc978c731d4499bbef5ab2721f231eb4ab5c8aff0e2988f424148284eed649e06d5d620ea9d99ce426c924c62927029effa1a743b446348c1f8eea4127f4826036762d279994fb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf569c17847c7598ceb4ee0b6523efe694f7381a0d86eef52adb51cb18345b29823c52db880953d6bb7f4e3cdc592fc0983c192ee023f46d7a95e8728cbb28be8c3848b328e00c7a25d4b9e2080e8f9b9ea738bc2f8ce6e008c126c2aa82dd2d3820aa5169939626af53c4765c7a65a2849b1ad92bd21665b61464ab4b088142a101bfe5d34f269c2f2dbdb77a366d30b2dd4495d84ed393f08757b974848ec830ac9c8e72be4c0275dfec80f31e5bbdf08f3aa0bff36c98c723b33412ba72ca71aaa3c07984011d25a9fe275d08888653b62ccb9f3061fa90e73a8a1882965c70556fa59110e601fbdb775ebe63250483e14cb2c188172b42c59c495cda919269d8d6c0b032d7588a5d902dbeef56cf894ee12e44b773fb01bc4e1be65919887ab8762bd0cb7132aed57b64bea1b0c2238cf91b2da73d7c08bd4b2ae067febf426b98cff92f8596c01314448b8c20aeb34c98e24b57b97ec9975f5ec2e22286ff5a486ff05f3b3e71e68fe5fb0ab2e88bee4a79ea94d1ed0380977663fa44652bfc860aa8a71a714a633c3e9e2301fa04e3024b72fea168e05364335cbcf34a1535ac39bfa1e3593e14381f0ee9bbc7b776cadd5e2068d49667b13bba4e8fbab5710102c061d56e38ee1239eb6664e46f17f443f3964a1cb323aacb8a459a58d379b7903b721d3b750e8aa5f2f3a9128c071c1a36f7c91f3157702352fe30b2b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hd3037b1ad471196a634d1cbcb08f1e8247c7b53bdafca7b7d8436e6aff97a0220825f2025e8fe7a1f47f8bcb5b2ca2dbc5295e99cfab8851b63e887106d1dfade96c9a98114020259d68062c74a7af1ab33a9f61bbc981b5638fe57a18d035818bf152249bff78234f0ec57df84477ba4b2724d9957b1b56520b673ce8759a61700a25f0254ed791e972a5a504b919d7d6654d23ed80cadc65a674077e0fda07fed772522e33ebf5233b9d178522d019ac3d2c2b96fb0993fad53ade6fc4c0154a1f7fc5c6cbbeb08e430b4b05c9a0e4fe684dc5add58aa7654229c66d9874e28895ee57de8b4c40a4371ad0be98cfa2caf821278e76e57bdebb285a56f12ca6566a654360a5c5cef2c5e9edf8394ace1eb6fa98d13c9998a7ff2254f70a937bb9f5f60b009452a5528b9d9bc69aec84764d4c591c3d040c5da8c570346cad4bbb7899973f67aad44e1672c3ad991c9fcf8c0dd63db974fac81269d0f728e659cb24a1e9845da5254098afc3cc86d5ca694c34fff3cf22bc2ee4ad0a4e795167e7f0364f1d7c3874871d4b92ddaae16bfe12f4414aef781b116ce52842ee7bbce5f3de1da62a441d3d2a18b7733b71f9f9a8698ca6f2136f25a59fad40fadb8b529dfc86a81416f9779fc991e80eb2172700a03a9470e624d1e58d6229c0ed830d8318d0838d28af3379fa9dbb7c6ec17cfeb7f097a263734f045a05ea03970c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h84ecd007fb59da380c9833ab1e8af7326b9ed3cc4458cff5d1c6f03ce7af5e29bb7343a836bb7bdf2697dccd0127cc189c5453da17669ffcfddd7ca4644ed09818fe6a6fb871c417033a0be4f904eecc85d81672c53fd4be40d4d155217e454a03bc8c244945fe63a54741c67f66d012ba01fa61873be34c753d980c2c4edb7727921c90f944da22a4dbb54e7306596e380078e26856c34264d047cf944aa69fdd9a62ed5085fca8c6daefa1eef5ba95febf9f499fe2021a484d32cbf637482f018929edf7ee9450087c240ccc6b4da465a41216d5a8a414a131124f724282873a43481e784dc4f967610b295a3a5dca9afc404661777a84ad6539adb4cf126aa1d6ae0dafb75124ab399ff2f6c4578006b7e743c09332e46bb1e879a3d3f6bae11703e03bab2dfcbd408152233544964e0d1a48d240a55629633088942130f16fd533925b39c4f368c9e2a04492474ce797f4abe61d19de4ac7b0df7f3d300892e261ef54b5956b874657c381cabbd4287f83758517fe7f3fd8de8f7fe484412d5d955c79473d6ff7411258189d15225042461e4fc03643ca7bcb825a521347dcfc007b38dbd64b3a207b4aef92893d4faca7e7cae5569929a11d162e15b8386da6c9b354662f40bd6b090191e9ffd3268b89f28cbfbb19a2c7e3b9678a41ae889b0b1ab789bf2809638dec3be6cc0c60de8e0e42d3b82dade1bf46357a6039;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf3c035e13525d66f497e74547286ba3de2b24db44fbec5fc78bd02337af2a0d9aa2e80d1927e78f600765bf6e94bc3dc638cc22d6e48e302ec5f09622a16fc9e60eeb24028ef2b2731ef2b820d62b908812d5237bebdadb964d1a5ae124fb1dc1b733002fed328ac8f975d40ea10c1889ae12b5c485e8b2d88e1b8acb9ae5d67b1d143eb6316fd2d3dbc84ec95f2fbd88791d6ef4dd924f7609f8529944e38b37eebe15759299e21b263d59a63e37cef2f3f029cbc2c060add85121c317809fa3c338441fba9283fe432b5025aa0403646b483731a1c5616f88526b234b7965c83f2ac21ac3ba5531eeda48b7f8a0cb3285540f1b3600ba72135afd13594b049c0a84a5ee6d00c8c8e52667b85e7c1c7822d5848f19961fb09b1b6fd2847113bbcd51d160e4789ec78b46d3e64d0dca9a59c03ad3f0644b957502dfe150b6ebccb711402dd9ce0925a7dcc4e843a06affd623ef7e443473ebdcbb4a88294a8fcf1d095a1e41c2e93ad9b3f58256340936070891ce4294dc75ade27943ff985aab722e7359d5f79bff8cdafd32713b9d3d1bf82aebe298e32fedab2b8c10728e3b54211b3a241bc1d9cd6f3e8a2380cbb92c8b58fa5c6d6e82fbf014b9af4b710c6ce08c789a621e1ef730a976b09f16ab9c2fbb52e954947be8e2dfed87b36fef3e66c99ddde61ddf0bc34f1c371c04df4f49bbd835185c43196a8f27cec3478;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hbe9f651c8f3914e3c7208ea04d759dcea9308fd8306bc8e8b67732008073432a16e1452601ee0c33075b683e0ed591287194ecb16b836a95369474be9072ec750807c38c56bdbba031e7fe3121341f4db71c985c537454cda47110dfa6b79d3246a2f0101bec6692795b28c5e6a37b706da6139103d76446a83a0ae8b5bd974c46e659e46ead626cde3a513f05aed5e35c979a2108a186ecbd6999271c8157005f2095245f441c4a3dec2c497af1afcff32fdb7b6557f9d341abbe8c8ea03fc75d2e7f3674549f487eb08eeca0a53fb95fdcac512d402008749d8ab6cdaff667e4d3599ed0848f0156b3320c8965ce406ee8e0dbd1508aa10f0c9351fa303e7572b3b65e1a922e073431afa643b39c697b346ed5291fa798da22edb289d6676a34d5afbcd6cb1d9e4802d687b377133ae8e6fdef705976ac89c3ccc162b84b2a59e7960d0453956a7808cbbe34c670860772aeae3f1a49c3a3a35c7a5b9c035c3528dc185fb0ecbb74e24d74e12271528fbacae1407689fe08cf63db7faa7f40c676665adced954d2fdd18dcd812c4791c9ca13036eb056cf1eab0e57aa4a053a486c7b3bea388b3a0461837b0731d4eb44e33ed46eae14decdd63120bfa7c94db360e7799e19b08aa483422486431bf91002a0dd12df752afeadcaad648029b33eb3d0622515793c73ff2419dcae745d57e31a98c166066f04717840cfbccb2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h29065638621b524029bad53eefa5659984bdca0346f6d449ea1c03ddff51e91bf628737c31a1011ecb69fdff8f3749cbeabf9a7d8eeda42c715e46a15392ed35464f02a61f80cc7992fcc8df90bab2b3f772883a0f04321ab08cceb21d26d3f52ec073c91e2d56ac7645fb82afdfb55916b89e86f36cb83dde1d40c3c177c1cd8c87166d6bcc22f00bf39200073e308398e30a1dc5643340b39b076bf29bb9869410e11f4b4e69a80f1fea5e3384a5054e8e84f6f4858e87faca44c5c821d754b1329ec63eb74441a5750c05d712d8bcc0cab3323a51aa79dfb4e2dbeb898694a0e42c9d2b72310ca4d397acbdbbe21d73c13fb42ef8c7a1f836b23249fb64d4c90f4907751e4f65e6ed2d8d2ee096ac6aeb97ce91e178cdbd0c018bea6443755ce61fff18da4a7f1f9a6f1e1a89ab98c6702556c46a42a517d32fa0309442199d17fd3ee147c55d226fc6c01a46cebc08f6a0566bb3da72f6a15fbc656cf7fc87f3c5461c4efb0a0a7602168e13bf02c175da377aa93763a3116453395da82aa923b7aca0729eab42a9287111f448b6cc39031eb8340bfd00cb30fcdbdfb7129895cd7b9b54927acf09c405506fe61b76a00e3a7105d82b91b14e02e0ac05257044181f3ae6bfdd4738dd7027c963f304e2f5c6ff5ccc789002e740faab3563b395bb1b6d7991690966aa79a73af0d78bf35a486ff5abd42ba80b4e7757716a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h64ec6cccbe0b384f58c4497887a9d22529ccae239f572e9499a73112d035274fb1ef7e280b8e24cbca8f35e345dc7099c078b21f74f92ce7084f2ab1215fc6a039c96bbf03120d996f053f330456e06c91e37d02944d922c03096ed35342403241115dc23e7ff0d957246a95627098438b56f12276a862c84d87ab4e2c4dfbe7237cfbb79c35e1730c1890b6f31cb574a93af387789541f6dda37e55342ddd4d868e3e8729483ee88025b7fac280b04e01143ba995e3429e94045f9d01e70b8b380acd98bc43020a8bca3403d86bc4bc98036e922e7592037b2239eec9e59d954f879613739428f3234d5f5830b25c1e4e4c1ba94efb23c9a46ced32af5cf979d862b3261df761c13bdf4ff3e97c4cc3b99113a8391c2dc50553a94e7453fe1815bae9b0fb60a2ed5f69382190b6fea72e3bf5eb647c5fe2a960b075503698162db81e63c4546799d0b0c6ae78a753150eeea88a7521ae47efa042ff2bf7de6fadb5f1331306ac5e876bf045dd7fbd4eaee03b9424f741e01fa2774c57b2cbe7acd692bcdf2cbbbeab687a7aec1ae7cb4b2773f1358ad4f8b657fbf609af65da695721010ad5531593b4b7cbfd834bf54a43bb76a31d9af190be1322bc8e8630f38e5b8a5f442cb9c123568d92d6d5931f99b61602ae0079ce9c556ed38fec0d039a609e02c2ea478913b6c2e576af93ccb50d00a830478ca7f63e842f28b4b8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h1a71838400dd5396b74ebdb542cab8ddb26d0a78eca5122572b9dfdf8ace8f6e2165bf5ecb6661506f5225102b67c906051463d6c66cdfbdd9533a92c00f5a4cbf933627225ee353da2f6ed1825e669c524693356acb2f73812a4b5f0dc04f2a75036fcde927f8743deee1b0d4ef604c5d7b708f95230fa08ffb9e851cc6b1fb47ca730aaa3d3dc8bb2481e13f79268ff8ed9300ead7a74acd239cbe278a5b76cf4a0f0f1d90490c955fe087da4b70183058124b31918fa169137a5c09b37d64f2fd52b9dea1fa955882dde20422586febb5b0d167470f4635ddab9a2885981aa87c051132c1e0f7a04fe6c0fb05e3ff5d9b324a9f852c5745a307aa07920e79eaf640c2332c08b0cc554acf993e8b46ccdd5653e12e1aa4068f6503217f8951612dbe3fd28778d40718288e8f2e342f43582af064e1d25c4e914b78e2a8095ef686586a200cb653e8fd81a234ee2bd6ba65d480f65cd86ec2396a11fd74397af5dba71e797b940a0f492a08ea200c75d627dbf6058d005fe8665966b8698613a676c721843592cea8c8794b2513987dcefe04a829396a2b969e60441661dffc4840770d65d46d1e33794a0a90c16cc22ed8216f631cf2868bd1af4592148a0b575cc4c43efb0919c020a0fd3dc30f67639edbb9ed7392610266797c062799ea40700873e680c0bda0206939f47744a42d714486afdbff8308f9da84c06097de;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf7d042c454a83c136c04d6a30d251ad2351cc2eac49d3d8d1e0db66584071eb51108029f057d0e5295b0eaebd7a5ee0876b990f28f14ee7d4800fe81e0ea628da11bb07f1d0a4346885c111d32011926203aca74c5df38bfa2564c2eb092f2a6190d958f508bae12f96b9303ad2221c432651ead561b9b12eb58990b958389f719dbe6d899a2659bb5bec08438685c95384b70541fa7010d2e2e13c8aa1fd2b281b8867ddf649907eb9a77fa6002663c03208083c41f8a340a2fc1994fee540bed6af3fc5ce8a52e2ec564941ea7ba9811800c0207e27486f84cdb34bbc49b1bbf890f353058a163253141b6a5624b6c4a095da658d49082d65696e2452ca834eca2be408665257ec9ae22cd94991171daefc5177cbbdc3e21fd4f7b0a76e3d9a08296a314b4da615496fa551f862c23f2b37f5127f7d046031271bda92b90817be3eb24f4a95e822671784b4bd2063d39c0f11ac45eae2dff81e099f8da74f592e0852007ed5ba611656f5f04a5e014ac5e7dc82864d6c3bbb53ea1423f2a1890ee8a992a77c158fe5c6fa83da3e5898688f62f59490eb709e4d204f5777319a8cc56ab0c95a1a57f68968918d4df594b219cbddd4b16d408298c15670b1a34421b785a4a1fb0ce616cfe796f2f1f6db8150d6291f3dfe3e847e9b2904791ad089e91fbc38d7319c803d6ef7b204a7f5f1626d2d54821de6092e4a2b8ee499c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h4820fd3d41ce82a8de63348e0718b6acbf5dcfe386aff152326435b5a8b52a8f21656550599bbebba91d4592bc352dafea2561613552229e96a525ce22d09477dd0eab864066a2e9012f75ec3c9c8344242a0cd99fb1919e039b81467d6bc8431df70d73ec7309da5ee44f718fbe2899484573f3e28070e9af377337d171bf363ad5068fd291c508dcd6aefaaac95f13367ae12084791f8e5c7c5e18362c4e49c22a0d33f48a4de8700ffcafb6f20302933ebfe1abdab427aff694873953038d52102889308c67e791b7b2bbe2a9c4fdb4dcf254581de1daad02acbc2220938d67432e939af081d1bd9a100a69d558e8ccda18111216336e3b3d2b81f934c8813eb37d2ed0f5b6e7c914f0b7c161f879e8e272759e062fd95a5ce88f7bbafec543b14d61b4ff171ab211bec750e6141bad368f93672f6f215af842e43c65ddbe7ac1fd8839b95fd5f7547159c2392c34daa34be04ec8268ac6069a5145231fd76a65a40c4618d4dfb5df6bf3465497a31631295ebb2da8b69b8dc9d41686bcf37e47139611e832f4b57ebab3698ade503d40ad95b14db7a4b0127cf7fa35277ff0c976e3730fad941dad797a4bd3385441a46f0764743f527895f10c4d98f9a8df485c4ebc277b571726ce918f84c815da34a5b6cca287c9107eb5cad1b02dd634d6da859ac939cdc2389a7bc19665ab0411a9dfd2971b21fdc3e21f99024e22;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb7dbbbdbfc9932abddc1ec2f08a11f2d7f3f4311bd72686f4225f447d9c80a1b828a86d87149b4bfa1fd5d5b5cbccc40a7d98b28c12803d1c34211796c4db397e1c06b52c74f2c9c5df34efae67c6bebbaa310356b9f729f30af9dc23cb1d7f32984bde736802dbfe71361231c05b05169f1ce72eab63caba914416b35f6182279a9735a0a3dc57a9878f10bdd7768d18d0d77b4f4e349a723ee1ec84fea2ed65b5376685239f66c8ea238a9abc5d5c72337adcaad34f9b5da226f3dc7f74ae64a56b26e2f74f5a6da1549cea5282dc2ab12400cc5f93f598c2cebaebd1f20352b3c3dfb6b7114c722ae69927bff729b4916097dff2c62c15f9d78edf4222dec89a8305785e4da676a7f23f0121ef1177b68e18bd59916f08933e1fc0263fffbb2bcfab54a586c398a8004f45b4f13e11939e7414da0be08b1aa4c771f8ceeaa44475154028a822051e7bfedd15a2012e7cbf69b367ab0260741b9157551bc4121e765548c97f680a1262ae6283345f11847137696114e86b7b835a753305b7c2e21db300f60921afebc9f0941c9b26a53d3b9e956bf8d2d3eec1980840dd3cd421f15c68ba40363e151c81c64e203ed6aaddfc0028506b2bdaa2d73e2bb64dcf90540d908f2b1ae9cdc40517537eff9ad55c2da241e47b6ddfc06e145eb01e576ca1efac433cd4b8fcab695be9125a5ddee8bf2893d2cedb79f49523d15c26a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hfb726098dbd4b47903de98c60a3edd7c3952cf4e2698e1969900eb95f160189bc421666c86522496239e615760a12863a32e982d38ea408f3c47c52d8e04c7083fe13a1662b6330a42fd70f911bc042ed0a2a1e11bab79d60aae2e6dc83c71c2bf2edb098c19438f936173ef09ac18650a28b54bb5e966a5f4fad625ff01c76d0c3f6b1e431fdeb32623585e070072aae6d656daeebcb797e1a9b34e912389b4fa1b9474d848ce1e742ba9ce5ac1dddada5208396ed821af8973e2f1be1503be46fd6d4e97884c93a17257298efbc40058e53f31e60e90850878f6337763d997caad6bba6d4ec1b736099237b8da27f7320440f7dc84bc96e1d0ca11acb1eab39ab8486991a6c75ac40d437bd8226c329026f943465131caadb617c0e7271a2519a9eec4189d6efa35b9f3706ebe6aa6383713b8f18bce4c69f837320195dcce20116ae73a329722d81bf5824f9fbe480dc0b97e5410f13ada6ba3ab2a02f2e17667914857e85c3a6c64c7f19015cc214d75f1bebd0319a7e4560c2eabfe045136be57c2e4caece0774d26484d9730bee4ab19b662499c1bacb5017089b01be1a90e0afdbacaed4f8190a1a61a7d040e5e322854889bea557c156bca4beb65f083dda1485a73ce5852315e1f9ae4d030c4bee8a6f0ac831e473e84f46ed7b4348f2a4ee7725496e5e852a10e5300e8eaf07a9d7ec81b4e43d30db754374f1f7d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h1335bdd385488390bbc2da965aca9f9c4995d9d806b610521f68f4c4741dcd8d15685298050e1db02338c5ef2d355e8a5e62bcbaa844af0767e6a0eda95d7d69b95de6b98ef3231938f81d4c5c3a3dbd383ad536b5381c64ddb8f78370f3e435b8790a2cd69e96606a91d6db385f30d16f56eafc479a722de11fb4f18afa4c930d9ab6872300c3894eadec7a150d544519af2b0cbb9dec02856ea13c94f980bbb71bd6222fa73097795586e4a3128931744b8a8623a8d112dab107773e8d40afb902a685c7176931d16d68d45fc695cb2047f07e2f19b0c41ca669b3c0658a90625b6144cda981b584e867962f457e5b393b32f885ee8e2ddb01746cf29b84c9c96b37783629946d78c3992bc4a6f5bf779ab12a0713240df8605d464e5e9d623068f7a26a3929b47c6474982435e48beca8932550f4ce95f2f8f2c9e06c7d93e72b8562cfa4ace4a69fc26cbc263eb20d29e449be5381bd0a809ea3273b6037c4baea55bfef3d1ccb59cb8d53cd6500ca2cf2e5f0005f6210aa7f493cda459da11d784a16472fd80f08046bbcd86c6aa7c315e779227b9a58d31cf4d67abe226bf80bdc3ee753b72ac8bb04aef268a6222151982b9f3f92b887f1c779dddf52771cfa291f899fdf2aa16c412b2be4a3d50510670176df7334835320c7db51714ac6ade15ed48dbdaa94b9330a310db5c72c487feccd08a15f0fd8984a32e1b0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hcbff195d440441ed9ad2a868c0d37cbf1d3ea9eacecd6f20c1a7e37fc77c594f8c4eb5fdde3603d5e9a79d5dcf567b2686532a47be4a7e751fd65b4d3cf60bfe483762b9d558436e794e577c380b806f2242de5c25e423159a3bb39b99b90df3a652391558538af805f3fd94670564acb8cac6a0d4cc079f97fc2c112f2c26b85343cac01db93deefa41164537ac6af1c14038a78c6fcb408398b9121af5059573036809a36f2701215e035c7c3441d3f88ef0c45794e928cb99e74ab15e0a1e2bb4dc8d7275e7433a4eaba4f2ce7344dfe158ff3315d21ba2afe1ea721dc898cb820c79d0a61016dc335194e3354903d9fcd9246430123e3597c83155a311e82956ae61d5a5f356507e193b2b175faacf82c4d385e65f5dc3a1a807cae7167368b9508cc7ecd978ba063060ae9636c0f185df652906d9361fe2c75f8811f270eb1661e2d2e0508b91af00ec6167c118cb52262de27ce9fb3363f7410dbc957fb3a8bb31e70e1a094bc931c19739366fe55edf34b2357926036ff5bfa28c830ce7b436080abe05024c6f992337672dcf64b261b5b08fca456f4ce4e44fbe138279d32c3e9580f8006317895dcf692fc6e7bb402ef66f849885805f3578ba47f9a504b23ddc5719a9ddefcdd67d2cf74769056b716ebb83ffb5592ceaab3a5919411c6bb3b8243d7f4016862674d92d6c50e50e176aab3a247257b663c781e139;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf5d0f1c38b7eb4cb61842f060ee290e210a40a652cb3957439168812fe0c17d9650b1e417bf9126c3769500a3a81559c2c647186796cb3145c034ce08002545cac85f0c7b09839c0d880ece8817f52d7b82a43fde715d5b12e423ec33d473eeaad42c715c7d3cbfe0f057058a94422c7d4addba4b398e1b2fac396585ef692ff8e96433c978f809e6796be2aeb3018f501a64457ad23c72e2cd138338650a5f18ed6af096bef4fd991f7de54fd8a9a36662c32a41a6fdec2255aa7eb949854b5734f17a57de241e666e67868679d20951d49f6ec0e4714a47aa068c84ecf155a6009b4924a4d9bdc4e27938f988f5b2ae28f27eff5e1cdeea4ad0d6f65afb9da9f9c5dcd54363b2f1be24960f64ac9c350e9baf1854287d9aab473d6707146f35f7b29b69a32dc8c591013d02cde2ab7bf635df6218016c71e63856c3fea95b0bffe20d9c4ceddfa9a0ae857b5ae6e46bd5eece48cf29bc616103e7905a1961a577320b04bb324cc919b190947b980c8268102a0ea5e33bc99f06470e4cf5ea7e7f7b9bde3e05657daec83776c492605d12de77d8333197f2df5b7481976fb6fc97f0ebf1b7e7d1acdd5b2b0e1ee08e7ae146b5f8f6a3e1e99fbc5dbd5830d9fe62cafbb85d4a5e4a0d8b0d9090d01b3b16c83ab8774d6bf75bda0e11f2680ee010d7983de8a055362accc0d3c0ede2ddb14ce8fccd92fafea5b27df9ab85cd5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'he0e4fbffb3c5506abb45c95d47bc02cfde9aa2a8ab5a8d7d4c5d0fc4b4324bb887029e8b5aafdf68df14bf6609a86b6d4147c2e363f96da4d1e94ea8fc71eb9b65491ddb57fbbfa648cbcaeb9de6c717f77c3eee9e66d38e0799a893070a9741cacb5a8586046b46e20f1f944f04c7fd1691f60f2190cd1aa2041e679de2f5f6ed0fdde8768e2d54e5f140d593086b2b8e43b90d1c0b298f36a8eee0a829233a43d1805777acb0721a61dc1dc5e1fecebe91724ac2a8f074f33a7f8d3cf970eda24cfed5086c6a7594c72821a832f1b908f2f3b847de3d84ffe5cb45a1b61bacb382fdf7e75037ad782fa4c94e97eec0d13242cb8e5eb160716f05b05f635190dddc143660b31a70bd5b03405ecc588117f7d4531fa68e1f6d13ec97181a60981ea3b53e1b3ca39e2e53dde4bbae0246b203b883c299800447c50f687fca1abb8f10dc27502bf15035152c1094c512ba2ef4a9750c77e0df3119c9cf11eb5f752abce1d1656c4262b0e91835ab47ad3ef3316ebff5bce42993d9c250fc66312d10ebf4634e48662382673d5836e8f0fbfe4f99512ac0d50cabeac30ab1db6d1e606c88a7960528a24ca26a1e895d947f0fc8b8cec04606d88f2733eafc70d73f4cb7ddae69f890c9334e8e44ad4c318ef326c2ab86e4262ac02504baddb872a7eab8509c12f353f5f2d2feb886baa415e97b02c8ca859c081b1b7fd36a335ba1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hcbf36a788839f9cdfcc6ed2cbbeef194d22139ee5bb8770369dfa5e5265e2d317a21f3fb8ad715114091d41ddc2bc77e0b1daa7e0dd3f638fe8cd1082156a4e909949129f87d1a82c48b25787c4a8400ca5d10461b37f2653768753fc51846288c838055c66b638fcd544758dfdfab43d83bf28844c54cdb98219f80582c6eb02c6321f483967603950f266d347c82367f4f59b881fb2de48b420bd558e5ea3f18207b6021ca10311f86f61fd1db1da09283af676dc526911cd3a31c65f589a18878f2de1da48f7dd8b23ad57d5404c21ae25a5fb3a05b83b46b586e1dd5f38ed5137cea70e156a7aa34761cb6ec0f4fbe0984aedf4ea2eb93d2bb63fa018745c1d77b140c2fc0dc4707f458a097d58cf2a0bef9adf8eaa3da1aa2f78ddcb4fa3208251ded9d7f5fd9b5b686633853539688be47e18b15185567ffa94c746ef682c29511050b5a2f1d993c644e91f3b2bbee7ec58634395e42628b15b5dcbcdf20fe995a82ae4ef96cbed284c39da8025e91fd21604907f1603a6e798899919fd807a2ee136c1e4a7d0db66fbf963ba343eda9f3bb1d2dd3a89f51c53606df7e2d7f7e2ede94e30101f65027d5a885b25e7f9c4d55c964a7fdafe9c69cc9719c4c12fb930368417e5d338b71383df44a8360a030a30bd7b522ba8b6ff700cb407fcffcfa4c74825cd8a1af801797df2584875f66e4f416dcd2856f24de113da7;
        #1
        $finish();
    end
endmodule
