module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17);
    reg [63:0] src0;
    reg [63:0] src1;
    reg [63:0] src2;
    reg [63:0] src3;
    reg [63:0] src4;
    reg [63:0] src5;
    reg [63:0] src6;
    reg [63:0] src7;
    reg [63:0] src8;
    reg [63:0] src9;
    reg [63:0] src10;
    reg [63:0] src11;
    compressor_CLA64_12 compressor_CLA64_12(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17));
    initial begin
        src0 <= 64'h0;
        src1 <= 64'h0;
        src2 <= 64'h0;
        src3 <= 64'h0;
        src4 <= 64'h0;
        src5 <= 64'h0;
        src6 <= 64'h0;
        src7 <= 64'h0;
        src8 <= 64'h0;
        src9 <= 64'h0;
        src10 <= 64'h0;
        src11 <= 64'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
    end
endmodule
module compressor_CLA64_12(
    input [63:0]src0,
    input [63:0]src1,
    input [63:0]src2,
    input [63:0]src3,
    input [63:0]src4,
    input [63:0]src5,
    input [63:0]src6,
    input [63:0]src7,
    input [63:0]src8,
    input [63:0]src9,
    input [63:0]src10,
    input [63:0]src11,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [0:0] comp_out17;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [63:0] src0,
      input wire [63:0] src1,
      input wire [63:0] src2,
      input wire [63:0] src3,
      input wire [63:0] src4,
      input wire [63:0] src5,
      input wire [63:0] src6,
      input wire [63:0] src7,
      input wire [63:0] src8,
      input wire [63:0] src9,
      input wire [63:0] src10,
      input wire [63:0] src11,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [0:0] dst17);

   wire [63:0] stage0_0;
   wire [63:0] stage0_1;
   wire [63:0] stage0_2;
   wire [63:0] stage0_3;
   wire [63:0] stage0_4;
   wire [63:0] stage0_5;
   wire [63:0] stage0_6;
   wire [63:0] stage0_7;
   wire [63:0] stage0_8;
   wire [63:0] stage0_9;
   wire [63:0] stage0_10;
   wire [63:0] stage0_11;
   wire [11:0] stage1_0;
   wire [19:0] stage1_1;
   wire [23:0] stage1_2;
   wire [24:0] stage1_3;
   wire [27:0] stage1_4;
   wire [30:0] stage1_5;
   wire [23:0] stage1_6;
   wire [21:0] stage1_7;
   wire [28:0] stage1_8;
   wire [30:0] stage1_9;
   wire [25:0] stage1_10;
   wire [21:0] stage1_11;
   wire [18:0] stage1_12;
   wire [11:0] stage1_13;
   wire [3:0] stage2_0;
   wire [4:0] stage2_1;
   wire [7:0] stage2_2;
   wire [9:0] stage2_3;
   wire [11:0] stage2_4;
   wire [11:0] stage2_5;
   wire [12:0] stage2_6;
   wire [9:0] stage2_7;
   wire [7:0] stage2_8;
   wire [11:0] stage2_9;
   wire [12:0] stage2_10;
   wire [10:0] stage2_11;
   wire [9:0] stage2_12;
   wire [5:0] stage2_13;
   wire [5:0] stage2_14;
   wire [1:0] stage2_15;
   wire [3:0] stage3_0;
   wire [4:0] stage3_1;
   wire [7:0] stage3_2;
   wire [1:0] stage3_3;
   wire [3:0] stage3_4;
   wire [3:0] stage3_5;
   wire [3:0] stage3_6;
   wire [5:0] stage3_7;
   wire [4:0] stage3_8;
   wire [2:0] stage3_9;
   wire [3:0] stage3_10;
   wire [5:0] stage3_11;
   wire [5:0] stage3_12;
   wire [2:0] stage3_13;
   wire [2:0] stage3_14;
   wire [3:0] stage3_15;
   wire [0:0] stage3_16;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [1:0] stage4_5;
   wire [1:0] stage4_6;
   wire [1:0] stage4_7;
   wire [1:0] stage4_8;
   wire [1:0] stage4_9;
   wire [1:0] stage4_10;
   wire [1:0] stage4_11;
   wire [1:0] stage4_12;
   wire [1:0] stage4_13;
   wire [1:0] stage4_14;
   wire [1:0] stage4_15;
   wire [1:0] stage4_16;
   wire [0:0] stage4_17;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage4_0;
   assign dst1 = stage4_1;
   assign dst2 = stage4_2;
   assign dst3 = stage4_3;
   assign dst4 = stage4_4;
   assign dst5 = stage4_5;
   assign dst6 = stage4_6;
   assign dst7 = stage4_7;
   assign dst8 = stage4_8;
   assign dst9 = stage4_9;
   assign dst10 = stage4_10;
   assign dst11 = stage4_11;
   assign dst12 = stage4_12;
   assign dst13 = stage4_13;
   assign dst14 = stage4_14;
   assign dst15 = stage4_15;
   assign dst16 = stage4_16;
   assign dst17 = stage4_17;

   gpc135_4 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc117_4 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11]},
      {stage0_1[3]},
      {stage0_2[1]},
      {stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc117_4 gpc2 (
      {stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18]},
      {stage0_1[4]},
      {stage0_2[2]},
      {stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc117_4 gpc3 (
      {stage0_0[19], stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25]},
      {stage0_1[5]},
      {stage0_2[3]},
      {stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc117_4 gpc4 (
      {stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32]},
      {stage0_1[6]},
      {stage0_2[4]},
      {stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc615_5 gpc5 (
      {stage0_0[33], stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37]},
      {stage0_1[7]},
      {stage0_2[5], stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10]},
      {stage1_4[0],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc615_5 gpc6 (
      {stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42]},
      {stage0_1[8]},
      {stage0_2[11], stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16]},
      {stage1_4[1],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc615_5 gpc7 (
      {stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47]},
      {stage0_1[9]},
      {stage0_2[17], stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22]},
      {stage1_4[2],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc615_5 gpc8 (
      {stage0_0[48], stage0_0[49], stage0_0[50], stage0_0[51], stage0_0[52]},
      {stage0_1[10]},
      {stage0_2[23], stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28]},
      {stage1_4[3],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc615_5 gpc9 (
      {stage0_0[53], stage0_0[54], stage0_0[55], stage0_0[56], stage0_0[57]},
      {stage0_1[11]},
      {stage0_2[29], stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34]},
      {stage1_4[4],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc615_5 gpc10 (
      {stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_1[12]},
      {stage0_2[35], stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40]},
      {stage1_4[5],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc606_5 gpc11 (
      {stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5]},
      {stage1_5[0],stage1_4[6],stage1_3[11],stage1_2[11],stage1_1[11]}
   );
   gpc606_5 gpc12 (
      {stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24]},
      {stage0_3[6], stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11]},
      {stage1_5[1],stage1_4[7],stage1_3[12],stage1_2[12],stage1_1[12]}
   );
   gpc606_5 gpc13 (
      {stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30]},
      {stage0_3[12], stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17]},
      {stage1_5[2],stage1_4[8],stage1_3[13],stage1_2[13],stage1_1[13]}
   );
   gpc606_5 gpc14 (
      {stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36]},
      {stage0_3[18], stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23]},
      {stage1_5[3],stage1_4[9],stage1_3[14],stage1_2[14],stage1_1[14]}
   );
   gpc606_5 gpc15 (
      {stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42]},
      {stage0_3[24], stage0_3[25], stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29]},
      {stage1_5[4],stage1_4[10],stage1_3[15],stage1_2[15],stage1_1[15]}
   );
   gpc606_5 gpc16 (
      {stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48]},
      {stage0_3[30], stage0_3[31], stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35]},
      {stage1_5[5],stage1_4[11],stage1_3[16],stage1_2[16],stage1_1[16]}
   );
   gpc615_5 gpc17 (
      {stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_2[41]},
      {stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41]},
      {stage1_5[6],stage1_4[12],stage1_3[17],stage1_2[17],stage1_1[17]}
   );
   gpc615_5 gpc18 (
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58]},
      {stage0_2[42]},
      {stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47]},
      {stage1_5[7],stage1_4[13],stage1_3[18],stage1_2[18],stage1_1[18]}
   );
   gpc615_5 gpc19 (
      {stage0_1[59], stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63]},
      {stage0_2[43]},
      {stage0_3[48], stage0_3[49], stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53]},
      {stage1_5[8],stage1_4[14],stage1_3[19],stage1_2[19],stage1_1[19]}
   );
   gpc615_5 gpc20 (
      {stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48]},
      {stage0_3[54]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[9],stage1_4[15],stage1_3[20],stage1_2[20]}
   );
   gpc615_5 gpc21 (
      {stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53]},
      {stage0_3[55]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[10],stage1_4[16],stage1_3[21],stage1_2[21]}
   );
   gpc615_5 gpc22 (
      {stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58]},
      {stage0_3[56]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[11],stage1_4[17],stage1_3[22],stage1_2[22]}
   );
   gpc615_5 gpc23 (
      {stage0_2[59], stage0_2[60], stage0_2[61], stage0_2[62], stage0_2[63]},
      {stage0_3[57]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[12],stage1_4[18],stage1_3[23],stage1_2[23]}
   );
   gpc606_5 gpc24 (
      {stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62], stage0_3[63]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[4],stage1_5[13],stage1_4[19],stage1_3[24]}
   );
   gpc615_5 gpc25 (
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28]},
      {stage0_5[6]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[1],stage1_6[5],stage1_5[14],stage1_4[20]}
   );
   gpc615_5 gpc26 (
      {stage0_4[29], stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33]},
      {stage0_5[7]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[2],stage1_6[6],stage1_5[15],stage1_4[21]}
   );
   gpc615_5 gpc27 (
      {stage0_4[34], stage0_4[35], stage0_4[36], stage0_4[37], stage0_4[38]},
      {stage0_5[8]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[3],stage1_6[7],stage1_5[16],stage1_4[22]}
   );
   gpc615_5 gpc28 (
      {stage0_4[39], stage0_4[40], stage0_4[41], stage0_4[42], stage0_4[43]},
      {stage0_5[9]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[4],stage1_6[8],stage1_5[17],stage1_4[23]}
   );
   gpc615_5 gpc29 (
      {stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47], stage0_4[48]},
      {stage0_5[10]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[5],stage1_6[9],stage1_5[18],stage1_4[24]}
   );
   gpc615_5 gpc30 (
      {stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage0_5[11]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[6],stage1_6[10],stage1_5[19],stage1_4[25]}
   );
   gpc615_5 gpc31 (
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58]},
      {stage0_5[12]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[7],stage1_6[11],stage1_5[20],stage1_4[26]}
   );
   gpc615_5 gpc32 (
      {stage0_4[59], stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63]},
      {stage0_5[13]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[8],stage1_6[12],stage1_5[21],stage1_4[27]}
   );
   gpc606_5 gpc33 (
      {stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17], stage0_5[18], stage0_5[19]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[8],stage1_7[9],stage1_6[13],stage1_5[22]}
   );
   gpc606_5 gpc34 (
      {stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23], stage0_5[24], stage0_5[25]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[9],stage1_7[10],stage1_6[14],stage1_5[23]}
   );
   gpc606_5 gpc35 (
      {stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29], stage0_5[30], stage0_5[31]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[10],stage1_7[11],stage1_6[15],stage1_5[24]}
   );
   gpc606_5 gpc36 (
      {stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35], stage0_5[36], stage0_5[37]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[11],stage1_7[12],stage1_6[16],stage1_5[25]}
   );
   gpc606_5 gpc37 (
      {stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41], stage0_5[42], stage0_5[43]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[12],stage1_7[13],stage1_6[17],stage1_5[26]}
   );
   gpc615_5 gpc38 (
      {stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47], stage0_5[48]},
      {stage0_6[48]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[13],stage1_7[14],stage1_6[18],stage1_5[27]}
   );
   gpc615_5 gpc39 (
      {stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_6[49]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[14],stage1_7[15],stage1_6[19],stage1_5[28]}
   );
   gpc615_5 gpc40 (
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58]},
      {stage0_6[50]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[15],stage1_7[16],stage1_6[20],stage1_5[29]}
   );
   gpc615_5 gpc41 (
      {stage0_5[59], stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63]},
      {stage0_6[51]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[16],stage1_7[17],stage1_6[21],stage1_5[30]}
   );
   gpc606_5 gpc42 (
      {stage0_6[52], stage0_6[53], stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[9],stage1_8[17],stage1_7[18],stage1_6[22]}
   );
   gpc606_5 gpc43 (
      {stage0_6[58], stage0_6[59], stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[10],stage1_8[18],stage1_7[19],stage1_6[23]}
   );
   gpc2135_5 gpc44 (
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58]},
      {stage0_8[12], stage0_8[13], stage0_8[14]},
      {stage0_9[0]},
      {stage0_10[0], stage0_10[1]},
      {stage1_11[0],stage1_10[2],stage1_9[11],stage1_8[19],stage1_7[20]}
   );
   gpc615_5 gpc45 (
      {stage0_7[59], stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63]},
      {stage0_8[15]},
      {stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5], stage0_9[6]},
      {stage1_11[1],stage1_10[3],stage1_9[12],stage1_8[20],stage1_7[21]}
   );
   gpc207_4 gpc46 (
      {stage0_8[16], stage0_8[17], stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22]},
      {stage0_10[2], stage0_10[3]},
      {stage1_11[2],stage1_10[4],stage1_9[13],stage1_8[21]}
   );
   gpc606_5 gpc47 (
      {stage0_8[23], stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28]},
      {stage0_10[4], stage0_10[5], stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9]},
      {stage1_12[0],stage1_11[3],stage1_10[5],stage1_9[14],stage1_8[22]}
   );
   gpc606_5 gpc48 (
      {stage0_8[29], stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34]},
      {stage0_10[10], stage0_10[11], stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15]},
      {stage1_12[1],stage1_11[4],stage1_10[6],stage1_9[15],stage1_8[23]}
   );
   gpc606_5 gpc49 (
      {stage0_8[35], stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40]},
      {stage0_10[16], stage0_10[17], stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21]},
      {stage1_12[2],stage1_11[5],stage1_10[7],stage1_9[16],stage1_8[24]}
   );
   gpc606_5 gpc50 (
      {stage0_8[41], stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46]},
      {stage0_10[22], stage0_10[23], stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27]},
      {stage1_12[3],stage1_11[6],stage1_10[8],stage1_9[17],stage1_8[25]}
   );
   gpc606_5 gpc51 (
      {stage0_8[47], stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52]},
      {stage0_10[28], stage0_10[29], stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33]},
      {stage1_12[4],stage1_11[7],stage1_10[9],stage1_9[18],stage1_8[26]}
   );
   gpc606_5 gpc52 (
      {stage0_8[53], stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58]},
      {stage0_10[34], stage0_10[35], stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39]},
      {stage1_12[5],stage1_11[8],stage1_10[10],stage1_9[19],stage1_8[27]}
   );
   gpc615_5 gpc53 (
      {stage0_8[59], stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63]},
      {stage0_9[7]},
      {stage0_10[40], stage0_10[41], stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45]},
      {stage1_12[6],stage1_11[9],stage1_10[11],stage1_9[20],stage1_8[28]}
   );
   gpc606_5 gpc54 (
      {stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11], stage0_9[12], stage0_9[13]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[7],stage1_11[10],stage1_10[12],stage1_9[21]}
   );
   gpc606_5 gpc55 (
      {stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17], stage0_9[18], stage0_9[19]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[8],stage1_11[11],stage1_10[13],stage1_9[22]}
   );
   gpc606_5 gpc56 (
      {stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[9],stage1_11[12],stage1_10[14],stage1_9[23]}
   );
   gpc606_5 gpc57 (
      {stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[10],stage1_11[13],stage1_10[15],stage1_9[24]}
   );
   gpc606_5 gpc58 (
      {stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35], stage0_9[36], stage0_9[37]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[11],stage1_11[14],stage1_10[16],stage1_9[25]}
   );
   gpc606_5 gpc59 (
      {stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[12],stage1_11[15],stage1_10[17],stage1_9[26]}
   );
   gpc615_5 gpc60 (
      {stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47], stage0_9[48]},
      {stage0_10[46]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[13],stage1_11[16],stage1_10[18],stage1_9[27]}
   );
   gpc615_5 gpc61 (
      {stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage0_10[47]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[14],stage1_11[17],stage1_10[19],stage1_9[28]}
   );
   gpc615_5 gpc62 (
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58]},
      {stage0_10[48]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[15],stage1_11[18],stage1_10[20],stage1_9[29]}
   );
   gpc615_5 gpc63 (
      {stage0_9[59], stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63]},
      {stage0_10[49]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[16],stage1_11[19],stage1_10[21],stage1_9[30]}
   );
   gpc135_4 gpc64 (
      {stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53], stage0_10[54]},
      {stage0_11[60], stage0_11[61], stage0_11[62]},
      {1'b0},
      {stage1_13[10],stage1_12[17],stage1_11[20],stage1_10[22]}
   );
   gpc117_4 gpc65 (
      {stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59], stage0_10[60], stage0_10[61]},
      {stage0_11[63]},
      {1'b0},
      {stage1_13[11],stage1_12[18],stage1_11[21],stage1_10[23]}
   );
   gpc1_1 gpc66 (
      {stage0_0[63]},
      {stage1_0[11]}
   );
   gpc1_1 gpc67 (
      {stage0_10[62]},
      {stage1_10[24]}
   );
   gpc1_1 gpc68 (
      {stage0_10[63]},
      {stage1_10[25]}
   );
   gpc2135_5 gpc69 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4]},
      {stage1_1[0], stage1_1[1], stage1_1[2]},
      {stage1_2[0]},
      {stage1_3[0], stage1_3[1]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc615_5 gpc70 (
      {stage1_0[5], stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9]},
      {stage1_1[3]},
      {stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc2135_5 gpc71 (
      {stage1_1[4], stage1_1[5], stage1_1[6], stage1_1[7], stage1_1[8]},
      {stage1_2[7], stage1_2[8], stage1_2[9]},
      {stage1_3[2]},
      {stage1_4[0], stage1_4[1]},
      {stage2_5[0],stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2]}
   );
   gpc2135_5 gpc72 (
      {stage1_1[9], stage1_1[10], stage1_1[11], stage1_1[12], stage1_1[13]},
      {stage1_2[10], stage1_2[11], stage1_2[12]},
      {stage1_3[3]},
      {stage1_4[2], stage1_4[3]},
      {stage2_5[1],stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3]}
   );
   gpc1406_5 gpc73 (
      {stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17], stage1_1[18], stage1_1[19]},
      {stage1_3[4], stage1_3[5], stage1_3[6], stage1_3[7]},
      {stage1_4[4]},
      {stage2_5[2],stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4]}
   );
   gpc615_5 gpc74 (
      {stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17]},
      {stage1_3[8]},
      {stage1_4[5], stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10]},
      {stage2_6[0],stage2_5[3],stage2_4[5],stage2_3[5],stage2_2[5]}
   );
   gpc615_5 gpc75 (
      {stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22]},
      {stage1_3[9]},
      {stage1_4[11], stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16]},
      {stage2_6[1],stage2_5[4],stage2_4[6],stage2_3[6],stage2_2[6]}
   );
   gpc615_5 gpc76 (
      {stage1_3[10], stage1_3[11], stage1_3[12], stage1_3[13], stage1_3[14]},
      {stage1_4[17]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[2],stage2_5[5],stage2_4[7],stage2_3[7]}
   );
   gpc615_5 gpc77 (
      {stage1_3[15], stage1_3[16], stage1_3[17], stage1_3[18], stage1_3[19]},
      {stage1_4[18]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[3],stage2_5[6],stage2_4[8],stage2_3[8]}
   );
   gpc615_5 gpc78 (
      {stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23], stage1_3[24]},
      {stage1_4[19]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[4],stage2_5[7],stage2_4[9],stage2_3[9]}
   );
   gpc7_3 gpc79 (
      {stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23], stage1_4[24], stage1_4[25], stage1_4[26]},
      {stage2_6[5],stage2_5[8],stage2_4[10]}
   );
   gpc615_5 gpc80 (
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22]},
      {stage1_6[0]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[0],stage2_7[3],stage2_6[6],stage2_5[9]}
   );
   gpc615_5 gpc81 (
      {stage1_5[23], stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27]},
      {stage1_6[1]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[1],stage2_7[4],stage2_6[7],stage2_5[10]}
   );
   gpc623_5 gpc82 (
      {stage1_5[28], stage1_5[29], stage1_5[30]},
      {stage1_6[2], stage1_6[3]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[2],stage2_7[5],stage2_6[8],stage2_5[11]}
   );
   gpc615_5 gpc83 (
      {stage1_6[4], stage1_6[5], stage1_6[6], stage1_6[7], stage1_6[8]},
      {stage1_7[18]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[3],stage2_8[3],stage2_7[6],stage2_6[9]}
   );
   gpc615_5 gpc84 (
      {stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12], stage1_6[13]},
      {stage1_7[19]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[4],stage2_8[4],stage2_7[7],stage2_6[10]}
   );
   gpc615_5 gpc85 (
      {stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17], stage1_6[18]},
      {stage1_7[20]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[5],stage2_8[5],stage2_7[8],stage2_6[11]}
   );
   gpc615_5 gpc86 (
      {stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage1_7[21]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[6],stage2_8[6],stage2_7[9],stage2_6[12]}
   );
   gpc135_4 gpc87 (
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28]},
      {stage1_9[0], stage1_9[1], stage1_9[2]},
      {stage1_10[0]},
      {stage2_11[0],stage2_10[4],stage2_9[7],stage2_8[7]}
   );
   gpc117_4 gpc88 (
      {stage1_9[3], stage1_9[4], stage1_9[5], stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9]},
      {stage1_10[1]},
      {stage1_11[0]},
      {stage2_12[0],stage2_11[1],stage2_10[5],stage2_9[8]}
   );
   gpc117_4 gpc89 (
      {stage1_9[10], stage1_9[11], stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16]},
      {stage1_10[2]},
      {stage1_11[1]},
      {stage2_12[1],stage2_11[2],stage2_10[6],stage2_9[9]}
   );
   gpc117_4 gpc90 (
      {stage1_9[17], stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage1_10[3]},
      {stage1_11[2]},
      {stage2_12[2],stage2_11[3],stage2_10[7],stage2_9[10]}
   );
   gpc117_4 gpc91 (
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29], stage1_9[30]},
      {stage1_10[4]},
      {stage1_11[3]},
      {stage2_12[3],stage2_11[4],stage2_10[8],stage2_9[11]}
   );
   gpc1163_5 gpc92 (
      {stage1_10[5], stage1_10[6], stage1_10[7]},
      {stage1_11[4], stage1_11[5], stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9]},
      {stage1_12[0]},
      {stage1_13[0]},
      {stage2_14[0],stage2_13[0],stage2_12[4],stage2_11[5],stage2_10[9]}
   );
   gpc606_5 gpc93 (
      {stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11], stage1_10[12], stage1_10[13]},
      {stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5], stage1_12[6]},
      {stage2_14[1],stage2_13[1],stage2_12[5],stage2_11[6],stage2_10[10]}
   );
   gpc606_5 gpc94 (
      {stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17], stage1_10[18], stage1_10[19]},
      {stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11], stage1_12[12]},
      {stage2_14[2],stage2_13[2],stage2_12[6],stage2_11[7],stage2_10[11]}
   );
   gpc606_5 gpc95 (
      {stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23], stage1_10[24], stage1_10[25]},
      {stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17], stage1_12[18]},
      {stage2_14[3],stage2_13[3],stage2_12[7],stage2_11[8],stage2_10[12]}
   );
   gpc606_5 gpc96 (
      {stage1_11[10], stage1_11[11], stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15]},
      {stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5], stage1_13[6]},
      {stage2_15[0],stage2_14[4],stage2_13[4],stage2_12[8],stage2_11[9]}
   );
   gpc606_5 gpc97 (
      {stage1_11[16], stage1_11[17], stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21]},
      {stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11], 1'b0},
      {stage2_15[1],stage2_14[5],stage2_13[5],stage2_12[9],stage2_11[10]}
   );
   gpc1_1 gpc98 (
      {stage1_0[10]},
      {stage2_0[2]}
   );
   gpc1_1 gpc99 (
      {stage1_0[11]},
      {stage2_0[3]}
   );
   gpc1_1 gpc100 (
      {stage1_2[23]},
      {stage2_2[7]}
   );
   gpc1_1 gpc101 (
      {stage1_4[27]},
      {stage2_4[11]}
   );
   gpc1415_5 gpc102 (
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4]},
      {stage2_4[0]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3]},
      {stage2_6[0]},
      {stage3_7[0],stage3_6[0],stage3_5[0],stage3_4[0],stage3_3[0]}
   );
   gpc615_5 gpc103 (
      {stage2_3[5], stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9]},
      {stage2_4[1]},
      {stage2_5[4], stage2_5[5], stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9]},
      {stage3_7[1],stage3_6[1],stage3_5[1],stage3_4[1],stage3_3[1]}
   );
   gpc615_5 gpc104 (
      {stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5], stage2_4[6]},
      {stage2_5[10]},
      {stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5], stage2_6[6]},
      {stage3_8[0],stage3_7[2],stage3_6[2],stage3_5[2],stage3_4[2]}
   );
   gpc615_5 gpc105 (
      {stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage2_5[11]},
      {stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11], stage2_6[12]},
      {stage3_8[1],stage3_7[3],stage3_6[3],stage3_5[3],stage3_4[3]}
   );
   gpc615_5 gpc106 (
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4]},
      {stage2_8[0]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[0],stage3_9[0],stage3_8[2],stage3_7[4]}
   );
   gpc615_5 gpc107 (
      {stage2_7[5], stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9]},
      {stage2_8[1]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[1],stage3_9[1],stage3_8[3],stage3_7[5]}
   );
   gpc606_5 gpc108 (
      {stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5], stage2_8[6], stage2_8[7]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[2],stage3_10[2],stage3_9[2],stage3_8[4]}
   );
   gpc7_3 gpc109 (
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11], stage2_10[12]},
      {stage3_12[1],stage3_11[3],stage3_10[3]}
   );
   gpc135_4 gpc110 (
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4]},
      {stage2_12[0], stage2_12[1], stage2_12[2]},
      {stage2_13[0]},
      {stage3_14[0],stage3_13[0],stage3_12[2],stage3_11[4]}
   );
   gpc606_5 gpc111 (
      {stage2_11[5], stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10]},
      {stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5], 1'b0},
      {stage3_15[0],stage3_14[1],stage3_13[1],stage3_12[3],stage3_11[5]}
   );
   gpc606_5 gpc112 (
      {stage2_12[3], stage2_12[4], stage2_12[5], stage2_12[6], stage2_12[7], stage2_12[8]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[1],stage3_14[2],stage3_13[2],stage3_12[4]}
   );
   gpc1_1 gpc113 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc114 (
      {stage2_0[1]},
      {stage3_0[1]}
   );
   gpc1_1 gpc115 (
      {stage2_0[2]},
      {stage3_0[2]}
   );
   gpc1_1 gpc116 (
      {stage2_0[3]},
      {stage3_0[3]}
   );
   gpc1_1 gpc117 (
      {stage2_1[0]},
      {stage3_1[0]}
   );
   gpc1_1 gpc118 (
      {stage2_1[1]},
      {stage3_1[1]}
   );
   gpc1_1 gpc119 (
      {stage2_1[2]},
      {stage3_1[2]}
   );
   gpc1_1 gpc120 (
      {stage2_1[3]},
      {stage3_1[3]}
   );
   gpc1_1 gpc121 (
      {stage2_1[4]},
      {stage3_1[4]}
   );
   gpc1_1 gpc122 (
      {stage2_2[0]},
      {stage3_2[0]}
   );
   gpc1_1 gpc123 (
      {stage2_2[1]},
      {stage3_2[1]}
   );
   gpc1_1 gpc124 (
      {stage2_2[2]},
      {stage3_2[2]}
   );
   gpc1_1 gpc125 (
      {stage2_2[3]},
      {stage3_2[3]}
   );
   gpc1_1 gpc126 (
      {stage2_2[4]},
      {stage3_2[4]}
   );
   gpc1_1 gpc127 (
      {stage2_2[5]},
      {stage3_2[5]}
   );
   gpc1_1 gpc128 (
      {stage2_2[6]},
      {stage3_2[6]}
   );
   gpc1_1 gpc129 (
      {stage2_2[7]},
      {stage3_2[7]}
   );
   gpc1_1 gpc130 (
      {stage2_12[9]},
      {stage3_12[5]}
   );
   gpc1_1 gpc131 (
      {stage2_15[0]},
      {stage3_15[2]}
   );
   gpc1_1 gpc132 (
      {stage2_15[1]},
      {stage3_15[3]}
   );
   gpc1343_5 gpc133 (
      {stage3_0[0], stage3_0[1], stage3_0[2]},
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3]},
      {stage3_2[0], stage3_2[1], stage3_2[2]},
      {stage3_3[0]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc1415_5 gpc134 (
      {stage3_2[3], stage3_2[4], stage3_2[5], stage3_2[6], stage3_2[7]},
      {stage3_3[1]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3]},
      {stage3_5[0]},
      {stage4_6[0],stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1]}
   );
   gpc1343_5 gpc135 (
      {stage3_5[1], stage3_5[2], stage3_5[3]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3]},
      {stage3_7[0], stage3_7[1], stage3_7[2]},
      {stage3_8[0]},
      {stage4_9[0],stage4_8[0],stage4_7[0],stage4_6[1],stage4_5[1]}
   );
   gpc1343_5 gpc136 (
      {stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4]},
      {stage3_9[0], stage3_9[1], stage3_9[2]},
      {stage3_10[0]},
      {stage4_11[0],stage4_10[0],stage4_9[1],stage4_8[1],stage4_7[1]}
   );
   gpc1163_5 gpc137 (
      {stage3_10[1], stage3_10[2], stage3_10[3]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage3_12[0]},
      {stage3_13[0]},
      {stage4_14[0],stage4_13[0],stage4_12[0],stage4_11[1],stage4_10[1]}
   );
   gpc1325_5 gpc138 (
      {stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage3_13[1], stage3_13[2]},
      {stage3_14[0], stage3_14[1], stage3_14[2]},
      {stage3_15[0]},
      {stage4_16[0],stage4_15[0],stage4_14[1],stage4_13[1],stage4_12[1]}
   );
   gpc117_4 gpc139 (
      {stage3_15[1], stage3_15[2], stage3_15[3], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage3_16[0]},
      {1'b0},
      {stage4_17[0],stage4_16[1],stage4_15[1]}
   );
   gpc1_1 gpc140 (
      {stage3_0[3]},
      {stage4_0[1]}
   );
   gpc1_1 gpc141 (
      {stage3_1[4]},
      {stage4_1[1]}
   );
endmodule

module testbench();
    reg [63:0] src0;
    reg [63:0] src1;
    reg [63:0] src2;
    reg [63:0] src3;
    reg [63:0] src4;
    reg [63:0] src5;
    reg [63:0] src6;
    reg [63:0] src7;
    reg [63:0] src8;
    reg [63:0] src9;
    reg [63:0] src10;
    reg [63:0] src11;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [17:0] srcsum;
    wire [17:0] dstsum;
    wire test;
    compressor_CLA64_12 compressor_CLA64_12(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63])<<11);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h5014a82c90c8d9233649ef073e03613fd9bd2e1995f5c81465ac309cd315007e4a6033a161644906097ca3205b4572444ae95ceb0e3a8778d58fd1378fbf0419b9e781492d7a9f31feb55d83b2624a21b6e45ab399ed720117d5205795207e37;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hbf6ec63f306599e341d553c08176f43852181b7189c29b19b454422cfc778bbc63f495c4ee0788ce7b55ef193915e7817e3f604f922f8588fe3a07948fbc94b36ea1ad43cd8b9866fa7047ae1f861b8934724c4f661f8181125790ddec6b826c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h14b1d074ad61361cd7399f3c664f483fca8cde1773339707b8adf2f8ca2566363ed8abce38c883ebc129f0d0b6525e990d1c44224575b7b7aa76a57fae05712348c05555486fc4d124c3a0748017bfe368b576b72da954c7afc791bcca586446;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h218b23c5ffede9708b6ed1083d6c7f3499b67ba5e05e676eff27277eae0b117816688b2e46f8d4b64de661b3bd2240fe4e03a76308e557743d6f3cdd2a0bf2334c85b121b4b45554a69701240e3b51d97bf4c22132f42593c41779b3727e8c6d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h89f57c875ab898b15060c3da2e5eb4c0880ea6ae6da0156880ff3f16e873a105203b6cbadd002137df1c3bac817e55788690aebcde4a4a651574c8b0391c632e72c75aabf62f0fc93614d3b2d68cb442afb6cdddc50591c619e4bed9465c7b33;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hc7c00eb2beb2e7adc0dc7e8c13eb86166ffe6bdf940eec974244ccca960db4549f086f17b5cdf6e616fd59d697aadfa45271202bdf0be1cf5ed4c198940f9a6c0333785dabbd11888c34f25bf24a420063e3c033ef2df829415ef44c61d1325a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'ha2ef307f6f03e35555c35af37f6cbdc1b2fcb8774ad730976b96b22e901b8892f7ecb1fd112b21331035acc37d8fdc3352e51dc921f6055cc06488c5bf29ce3b8e3108e4b3f3a5394945374f30b95d409b67c6d9b811e2f7de41ab8e9fffe998;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h5af28ce74db60657ed75485bbca0c5d4fa09201e38bbb207091daa05f8a7f0813a892c59c63a1e0b96cf91a64fa0173ebbe6ba789c2d243b8f137182c966093e000edeb9cc121826dc27df676044b88c11eb1509486545bb25f8eec419a251bf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'ha55e85da95af70d6961200ecfad4d76f70404637cb032fc3b9465d59fc4e38e1801bd875953a12ce464be70b37cc952761741a4e74bbee47c2b21d929f74d90bfd19902c08a293023b0a5d3f6e4928eeed1c6082e20b22ddf97499eeba4cd35c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h2442efbc24882e5fddbb31c520be597b8cfed5d8817b4989520cc5e565f14c39282473764158b471dcb2cb368f2fb1867966f77e896b3f98cbd7b767f3d381d3859527174869d261d1a04cc81a75c69008f4fe4d98f33c6e1683c57d328030ab;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'he7c5fe910507ce93b7574177df3afa33a9a98dad2a2a497c1c422e457a6af118835f574fbfd59c3ea3cec0aada7935fcbdf6ef2e03ca3110aaded184e669ac9cbcac979443eb83e83bcc9978953cef6332f17bd84f47dd40174c97ac978fd6d6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hf514445f3bd969438d59ff59e121962abb71a790deef4feabc366a9109444dc3291cd4b6e72fa261be760454ee7d1fdce9f329e459b5870e0ae6e5233cbb4f75bf0ba6594f5c760f45e3809a571a3cd5edbf094c8188c01e73864f0a7d14e544;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'he6213b67ee5edfe2f1f2a4a86346b7a074b9c06384d9b17ee821f40bc9747d854e1d452ec7d763b826e19eb3ab3f4262683f9660cdb416c7541db9dbe90853c999d6bcfc8145a13fade0d8a5a41a95ca4aba3dfe58a973b2e31adf0bfeed408c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'ha0359f207da67625ebaafccdcad538e12255990475bd80b5167da8168cfefd079b741c5d8284232e01bd6b7bf74043ce80b0fb8c75e7a3fc9fbb36b454625b3217632072c5b79f5e73f3ce3abf94398cb396bb46217c9cf524cf2519552e48d6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'ha87471f14787e06d5da13d71bd8d74ccdcb24d77547bcbd348985218b26a4b6848470a778da3b66566ebe811218835d0c803ef1ce99d3b64d873923504730de676291fb5bdc8bfb303bf6199f327300133aa11b81f16ae773394edebce65fa33;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'ha40e5e552a52d3e7d4479f3bf8c678352529a6ee561a412d8912db5582bca461169e6f08d2b1ddb2badb92d2dc1bed97d314e8b50c651cd4fa3e874d8220e824dca32e8c43c56a900da2bf548ed5caa74c8adbefdfc209dfff09f9828e52f542;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'ha6bb306df35c4669c02d4ec0e7cb3eb011ebba44dc70072969b49bfd98cc6e26359bf072ebf685d5137c56fbc5d6ddcc88f076dfd73af657283fc785cfa65efc18e50c91da957a720665c5d3d3e9659864926b75ca8dc9a5d65898659b387c3f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h8b527c137c2f8cba2f82536a32a09cb22ebd22dfb41078c077f348b69e312deb7ffe5f059554fa6d48cec30df1644df7d4c6c045af43d7a6e11a31c76a0dd91e9e1b73f85fa4e242f6418844930a06011a7b8c189bfbabdf95a7de1faa32ffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h2474f425efbea6c29e7ae86637cc176d6e46456c92039430bd92ba83ae6a6279370c1497906d7cddcddc6afc87f7532c283ad36193cd37fb24fa5660518e12803442a344be9e4840ec977bc2fb575708bae33f88ef5ad967fee89202580600e2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hc49454f5dab0d7f636f7d30d7b46c74be56dbf4f4c92356a198cd9baac0c29469366c069c703d2f5389431e6dd16214a65504b3335d3fab00ea164d04504a07d9cb0b7bc1268b4844526ebab56f16565dfa826eb49728141550ed444c2607e4f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h39ae7b1a637cbe56c951ecde4033a0c8b43df8738b04320068c48297ec9fcd78367d68b05df565d455a93e9a554af45dbc5ebaa14d7eb961b902baa3aa5168056057b6801823e3b3edf6066c54ad9cf78108e73b053107ad35138587ce744ce6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h9a3cf63902c8716993d522abfc6859c8be4ab20435c9180c53e6c5a8c7ebf71bfb08e751dcf9fa3a59af0b19743f107150726cd13ea73236004968392d5c949e6e5afaacd8cc56215517938912cdf9a7241abf55bb88b885f4701240b8742358;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hed64bd750b6664d0a55edb0ed614c328dee68f14303d0d92d83f8515c28a9e3075af5508fc26828ce2126c5675ec8db87420bd1c56b4f1ec14a63434d3849e9e75c7e53511a0dc8ffb2a6c279c064de83d9f9a215cbe818b0f599964a7974f0d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hf2276d0c294800cc2ef9f4e655b89a15152be641cd5cb3e354cce085286b1c2a72f476d42ca1dd90e610cc31936951e96b7f646ef5b71951d234b7b52dd5059fd839fc18efd13e2bea8a15bcb6a740633d5d24bd8b416a36368e0a47f46c2ee;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hea5b594696895fa19ade83e743d8453bc0c87cb73019a09a246954d10d9ae448a2b98bbf259f09de9a5dcc49e6cc84691cdbfee43518742d739c001a6d696f925fa53e235d61d0250b7ce27bb06cf33d3983daebb0fc8cb410b07127b489e17e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'ha9f9a9b4476bb5071678be1be341bb785312c7fa570a0d6a10e0e3341c9afcbd9680baf3692a394d43555aaf0a43f4c217dc0431c5ba7f87f140c62c7b369b076ae0e3b96d67cccffc867c8ea8b7748cf6226b07eb46fcf5d987e3d038e1e478;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h60485e5bd70bea64d1a32b679e3286fc96c805a21c058e19b3cbf986b790f2217b723eac72864d621a5c4c80ed33e82c75fed41da734c51e3cb6eb1295bfce2cfa41bba6128f5d84e40b95761abd64076ef290d68b2164b24f83c649ee5723da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'ha46291819908b6c1963320ad01435a54d8174b77b869164ab97768283d2acf23fcdde584113c8f94314cd78ad7cd900a2441ca7e4befe56d93be3a22bef9e0b02e066e23f2a460f1ab73d18bbbdcf4eee902ecfb3eea6d99f1622fadce451334;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h93d989b345707f9185ad92481e2910a03942c65f9ef00c37f1e0e6579a61981c226f2df3625fe564d375b50639fbca112f01062607b88ee1495f8b1e5d03f919f33a90cf4ed784799d64966729b71dbac6169494ed29361b1e401b608dab055;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h87d106b5e824c453e864ea9d957ac6fa4d3b9c299af1746ba3fdc64248d4fdf23477ed6b18a68ad1f2f3d549cf427b92408a1fb10a6848f7fdc83e93a411838946c8af80cde60ab5050d7c1bdb7c1e4c57ebf08cadea7f60d2fe3c485e5c6b5f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h8bbc448fd43dfb6b50e851d7ae47429b7b9239c37a28ffcc72ab6d24d1b2018f670c029c943a4cd7033e97def94150afc3a4d94f121c0a533d32c17e5768f72b7ca179c9ad30a7a0c85c9e81e956fc3ce5656bbe89b2cb483cf3c919e8802672;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h9b6d353a1e37630dd1b2af01730a6dfc303f6de52a150a22854bb637c0d7a854df8bcdaa5834960a758ea79fb0a4c70c0b4e78733c6cb6645051597b75d1ebd1489cd42f223d207dd78db56d110cc87886afafb9dc7050ce0cb169c2ec832369;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h28cf1e8e5e3405542bcc187f4861bcd6bce734f81196262613e616b7df844733b8547731c7f49eacfee07a398dfe87066f2293f23d679c7bd0bfa46e51f651971ca1d1736f9a62ffe374f19db197002c723170966043e1f1e32dfea63a57250e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h6c742c9704ce7b22cbe7fd6a4f7e513f2825bb3a57f37e0936ae9f5af3ec2362298c11a4a22ca4f54731c42c8812cc4e98643e1f90c212004f321dbad95e96ad0f905e135f1e2cb8b154813d84f6fb783f2cf324c93d0fd73f96adee06502de7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h26d4e96e70794d5742f7090026e1814b88fede425840818b28cbc019c2522cd3021720e1f6ff8fde108610524fc5a59e1b4ed22185d725d7bd86dd56ffcd8a160a927a69d534b28bc26e9747fd210e2160ca00a0ca471e01410142cc1d7bfbe7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'he28f1b4a7b1265f8a84f94c442466fd97b1223a1f5d4d990513bca3bd3c806fe72ae879fdac90ea2349b8ea4421d78a8eed8ae8fe9db5cdfdfd9411d0d5d2c9617320356e535aafcba00ed0cf99cbd8d776ac765dedb600dde67ceb7970adc51;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'he6b51b5ca5e0f40bb6164b275ebba98e615f33333b636f40e1750c3e71ebf2c96de6f8ea4051bcfa3f85fc53c149c98a9e1f34d4d1834157b4c44b173cd3d45a8802f83028649aeadd1be14ff0fa36809a98750b4ab1b0072be2708862343a4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hb0c3b0575386bfa866219e2e9f9e2816d70d8548d7793769a83b50ddbc4fb677ab99c9dd008eed7da0658c84382d1edf2aa6037ab74ba10d14a1de99d0319e8467ab3ba9577c2ff5db0414701cf1c5cb6b232bf90be65aee66f86726eaafee8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h35b88cedefd8d98626eb8d2498a5172ec7ed6ed938970ce11ea40b9b2fcf612c7c1bc78a7565cae9c937268643604931d3cd6f12dcd7ff37a894a974ab7fc4ef3f2d6e0c9d2a63fc0a6983a25f5f4ecc1109f2194971c1ba1fb8d78564ca061d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h5060e27d9e11b6269a9d319c7fd16b1f92f8f1576515f3fea7fe9a99c6a89fdc61e082c00cedd59fe95e792d662ea5c29cd2d728f067e3390d095b8f0b409309972918f7c086151fe7ef3a43333d6c3bdf934a1c28fa470fa7aea1fdeee34d11;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hbe13105eaf2df87372fb9e4fa502eecf6b3b5a5f06a51d1cf71044b8c3689137664c188d3be147af003a4a2fe2ff97217a7fca8ca03d75ca2911c3bc17ccc29d9d310a49082ea895c48bf1a09b2ca735fbcce20e2563e38fb9b9e6147be494f0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h221aece1f33137367a9be62b23d271d0136f094fb582b18341f9ac48ded2fceadad54b12bd217d70a92fdff329b8e0db39276d04e7fae91b500e4fb9cdfbe4bae07e3de41e000e0ea9c214aa9d4eee1682d880cae94fe5d32798caeece7d5688;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hbe31f3b4f0afddfe4172ca3b810a3bed2718b9a59820fe2593e4276dda4b679faf05feff844da7de02ee1c18b2f77a016fafe3ecef2ad559a882a564042d5d5ea15ec884d7ab85ffeccc9b1ebcb70cda97733deece1491682c74f049c6e6dccd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hd2d9263281cc98bc06a64305adfb0a23b2519df95686f0a8a0e03119c7e9b28c400c7e6b8a99ec1c479e21d584f9979895dc9f53a0e1ceb41f225f5e36f75ee5b4a2b6aab46ac296dbdc2284f28a9b9c366248ed6101dda215d49e45cb93739;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hcce6f7d44fa0844e1964a11193984f1d737733f62745b27e25ebe7b6feb38e097bd7bf26bb9cd9b32d232402a3904cc9dd88357d9d510ac7bb2870e26183a8ae682c00f9d909a022870220fbe78dc0f2830276ab6b08ce13a8d22fc1c66c772e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h1e06cb97976c6224804a5b6d6cab18ac38cb5a4ea69ccd908bd2fbc6afddcb699e0cf9fde2c65ea8544d018f80a093bcfd5a03c19e405fffed9da17ad827e3085c6a690531c8d8d3cbb73d6f27511e687bac04b00f097e90aaaeffd48e43cb7e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h7c7c59aac0bedb536baafc4a48f6a1d38d7e88b8ac8ecdc91a9690cc839cb4ab1a5969950e2259395eae8fdebff8eed5eb316933ac38ed6a00369cf3ddd6e7431f451405d18525e3aa5a45324cf608f939eec6f0dc606b2f83214084fbd63354;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h716a514b50787f90de6ee681776545b184abcbd2887c6baf1d7db8a608173f0fde53088f841364e53cab41794ecb09c9344cf4b1d7b9918bf8666395b4bd3226f8785c3db988c4216f6e326e9bb2fc3772b2c529186becc14968ed00ba483cbe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h82406479405512c907a1274c7930a9d4ea2b2843a4231653735ace6bf24c4f88c704c8777589b5e625fe125df7c658f14cb2b217e5244432ebef2253cb31092858329606de7146a83eb804e2e5cc9985f57e58d5b07e127c6caaa0957be6c9f8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h7eb530710c4523413ed420084347ccd302916b909d4f9bede510e85e7e42c1de0ca54b2bedf60a319a8dbf08fc7146a561a031b46e6f25a5a8796b77e836f71bda105eec7d29c1edc4f19a025c08e691520adf776b1c712ae5e5f4b23f827768;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h27242208a804fb59a36f4488a71eaf961d2b85d1e6619cdf01f9978862e740e886a2a793029fc441df6755115ae88a24b4f55f0d0d03fc998133107747345564fd7c29eae153eeda954e97765c405f318edd6cb0aaf68381ffe97a438b56ac38;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h4f4f46873fd2f2f976ac0403d45146237d7c930a6ef1221302123b0739ae78002c80fce99d7ae7cf32a861c97f483efed43f3aadf2924d5271079d0455ed076e1c8eb0888c80587e6706063d0af32795a7aed0ff37346bb19e426e2746c9f1d0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h5a8e809c74531e5d0362e540b7a0113b0d0e1bef31eb345da14b601bd13588103a5d029704cd580d3fd0ba51b68fb4bc10957d882bbc3d19cc091be430db7246300682110129410d02c9e286e255a2edef0cc8526b5cc78475846c68d9e49595;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hfadeaaf7747f795e00576a3a8bb42076ce9f31eb563a83f5ed16cc85905e58bac071866ca58c68adc23a1539ad5df29cc0de3ae61ab2152bf5380bfec1cf681098923a208d2904cad49aa6b2ece394a4593faeecac9a2ad6da264bf66de9ce5a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hb4749bb821b478e147ec213040e592619ba21305430d80aee9bfc52fff5d728d0bc343fb731c29cafb8e45a70b6a47311b2b7965dd58a219bbbb656319eb546b97215ed699dbd5803499a538c63b603566dd1b6297edf46bcd85df2529af2e02;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h2a8a43429e088ce86a0d71b69208204df7b00b3963d6eab14901bd53569b41c12b064cba7a69c78c5f2ef351a7d19012920aff4e71bca5cd49cc8fab97b81fc841105bdbc7093b492aed206d59f3a703a962be46cd7c56d382f8d4f0eb46a1c8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hd1121b941fce3b143781348312aa07139bfa40bb66b237a7dc38fe83edd2f874f9e47300828e24518b9cfb2ef1c8ff933c5779c1a6160ffcb911f43484d2d1070e7a6380a6a0bc9d0f191eb62f558e4aad5db9f4c2bed86e1c727cd663a47aaa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h457062d784d5b6b7f1c5a4db0ac807ec4f046a3f03b6e8fe13f0689b40885d2365cfeec62009207636b28700df4fa0db8508aef6e3e6ccc0541eaf1e62cfc031dbf4ee768074adcc850a84a56bd0ac481a3a4bd426a60a78debdcfed60586910;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hae73a5e5fb500ec7711f0f67f9bcbab4d424c1f93de7d241ee89ee6732f085421e9be19a53d7fcb18d311cf50a7e3f1e2c2c1ab7bb08b65f502cd5cabb8f7f9998a772be875c887df0c75bd21f196641371f61cb434c4640d762b8a7e4cf4fb3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h185e06468fe96de5e2d71c706509dc4fe778c7e70d83f0ca86706d97dc242eccdfed8ee9e6b904291e0c7e490b367e4091c7e66a4379cbbe3238fe666bf9788edb1494f17883710384edf2302e494fde61478ef29500db1623b7ca4e0838b310;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h78a2e62970fd55b18f81f4594ea50cfdb8287f469d879c380c03cb2e802af87b42d97ae136c2352870f6178fbe5dcc518d46f06102b70fb5e4b482fdea2771b4fd80a1bcc9d0702c5fea6aaa1b1e08fc6b7ffad2b5b93475a7b201defc18770e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h485815206664ec83a98de5a0cb2b17fc5f7d0448f70d58da9970eacfad03ae6e95828bd27b7dab6fd2545353c6c4167f1ae94f5c9765fa0fa7c7bbb7865620a56d2954e02a0f6aab959273c35b2108f232b2e7dc118fa52ed0f044b4796bde31;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hc7a8579e1d8273ecffa368f54ded5286dc57c8a91d0970fbf583af223686b7c63f69c5f3960f6ab08bebd1d6855dce1a31241b29ee0b25ab79a87d940756117f91daff0eb905be551abc96192aa9adf69d58b2af24fb5a84b50e6a61d2952fe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h7b2eae97fa8283a3b9a97d77cc6b11869f942f5684edb861bdd17ee27b1ae3a5b6ce2f576bc75b457050b804875064ac7800ea689ef573e0c111079ee54f24b02aafcbe792333e7a6ebd45e06a26a43ed289be1e9ab9ad7c38860e741e95064b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'he3e04a4b0362d7e2e270e6b9e4300035f97cbfef5794c819ab1fd0b66ebc8183df6ae2c169c9cea2c5c5f03004878a17bb44ca1ac5dbc66e15498aa6366807c103d59fb44fa45c6a1e2a3dccb782127205f5d0cc9e61081712cebdbf0a38ab6e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hf4836d978f55c61b4d4b924280665fb78aa70494be04099ae52f1b575cccb80a2dd46cc699e6b6028a12902eb23e502beda94e1dc6adba143223fc18cd0c3de771d7b40905257480efeaa7862be0169e0ff9cfed3c6413ce7b79f92c14e5d098;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h375cd88cd62c7dbf231bc42d5c099e20f5b4cdad7466322e8b53671783f5f0ab7120116bfb9f6ebd8b254e84d5d6f63f56738ac8ff748a088f4c77997887e0c53a9cacae8c79a95ef2294ab75fb51d55b6623d62cafa28b866ff926ade0910e6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h69f4ce5f2b93090da062bd39fc95668a3149a38a04a8825ea53374aa3695b9a5dc91a3240cddfae11e16dff1d2448a79d10ee5cef3cfcf492324d1adf72f5653ac8101d6d1f50e103311c59ab41dba74dd2dda721e19e099118b1e2e4fab7ad3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h315400e8a6a48553665c573719faf79c7454a296f4647857cd8fe1eb2b8f07a1999ce5df463996fa9fe1a18214daf2baa3abf0970100a37b0815620771d78ff1b6ecb693ae60a5f792bed8ae06ab885c42bf27db40729f79a6fb01b17f18fef7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hbed2f6579fb19f27e0c7bb9da31dc4791e5ab51905902f097799421d94dbad2ac9ef7ff65528a4147aeb36c1a2d42a39d86a8423e61ad141cb84248657468aff9ea6da6e61cafb9f9e8caebf94b5d05359b9986d7969ac9ffc1895bcbb0a840;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'ha4fc5280edad24805fc6d0357e28ab52b2032dae01d1b17197d31942299f2046b2c54bb94ab1644673a23fb286e70fecc5ecc21727903a9b3ad0d482c3bbf635131a224c00596cbe35202de9e3dd7e9a79cc9d8cfc845f44d483040309f4f46e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hf488b8849d3b4d8c2e7017d1a85f40c9faa70a087c7dcceb918295bcaf5353cc02087b78f6b5f8dbb31743335d8291a3f5aa8b80e90f3658142039aa76e4d45f2c723a4f58015aa1b834ccd9e78f32976cdb88e7f49efbf37b02ba721fefa420;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h628c02f3af74609429f8800f1f3e8a9526081a021a722bc32d392d8282d3e006fa36569d65702338d84c20b7ab39fd02ffe9a33ce8946a4c004c82b5be720c094e5bf6a6b4d228daf5599dc092502aeb893dce8eee10987bd01e32c55987ba3d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hbfd7a5f0790e43544c10fce6f6a6ede8e0838d43ebcc1094b8c1eb7e1e3d0a0f75769b2521924464110497754b7bbd7177520a2bf79f7e4189289e2091d9d42a20b76c061367a9827843c955e0432410fb36102d675ae6c8f2128ffafbab6e60;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'he5d409060961ea313c423d3c9bb11d8b4ee57033db7c4e5490c7ecd45b8a8b44dc5ea19be87efe1daa5e47242dc4700ada28fc08709e8429267f850f8605473a5fb3919619950cf9ba86ef4b5a2f475a3706758bc85e54069ad9cd9a24052eda;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h992aa2602f93515fcaae47558ee014b0f9705a7d42d91457f4953e4724cc5d8939a8d6151453f145d08afcf765bd9ef51e2ee6827e13d5c234d9d9ef879e0e38a7efe9e76e8414be998e278fb7c74240efc3975d7ff59096fdf36f926e78bf10;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h10fcb37f638fc7e8dd35504e3f72fbb1a7df7d13d6e1947c606c95769dfc85d59e302e9c10871d288c50ef25da38306d91aa9d3f17e833234b6661e8190f87abe2fd2dbb2ccba591b04b7a1cb43fcda80396c5883745af938629e61d584178f9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h219eaa17ea6d8276f848abd60697f150721d3582f14a62162e2699f50da4b763383642aa62a2c7c9e256eacab758e059e2aec3b22e11ce7c63977ae071f93793ff4c1d7aa8e4a19defdf13f94c766bb9e42515adf3417bf6006abff2d5b08707;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h49ed8a4055dafc64d5ab54badf078e32cfd04e050f06a861f36a4c3069234cf7e689a3b7bf840233d6f0161cc7c000f8145791a5c996c26f0bed26317d72f87e1663c9d778b14add1aee947637576aab36e0a99e24709ce3a8c2ce8c4e47c00b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'haa4c1d0ae4697ea554c084b52a205ac44a8b329b8876a5c99c64dcae14233e07c35c4c2e2e134bc7499fe1b59f45bb9ec76e8a42ed1d36e3fad73ed6fd9b4d96d5f881726445825552af9b1a0123377f634a48e86544f57aeee33105e982abce;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'he605aebefc6beb49376a8549833a8d86ff84a8f179ce8c6434e4a073c927ff4ed64546567cb8589db0b7e7ca64efcd79cc401067a50a01ff962496bdcb3e7fdcb1e591e52ecfc97bf9340e93cbb2685db30f2eba4d6745a6e5c2294dad22583d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'he2cb1485e45410a54f5cff8fcc51346d69394dc808c5fe5a9af7e6cdef62cdbdb6a5a954cee0632e5a7448450aae0b3d91c00641fb9903b999c0b8d6b69073ddd7d8d2944a20a47c10443ffad4d4a269581ae970c26a4e820aede3bc0ba896ee;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h3699778b121562911dffee10b923b57d1f9c5e3ca03e66b8425127d554baa21a81fb129a94078a6f2d9804a487af329794ccd3c56294000727759e813546dab213912f678880ea3f070455c93e246e77eb6ccffe1fb7ac76d4d5e8be844dcc81;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hac81a1820d3e5ade09b598bf6b2dde8952a9049381509dff7fc57af46769c13d50caf146fe4bc9c980bab7526c5b6ffc745b34f7cb95266352aadb55dbe08be51e031f395622d8dba21111669dc084789b71850d29d9821fd4eb7a08d82fdd9f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'he8f6b27135ce7e02e56087646a7100b8fb4df389143c5854ce2139ca683baf8fe3c5100e15af6d099c3fa3f8862322c36e281b60c2db52be67daf82b4bca2578b933d1023aa35f932f77a1fff66543be22e413d2c84be9607bea663dbccff8ae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hf8f16161290cfaa1b3fda253b21cb1474152fba10453dc07560aed3283cbcc9f803ca5798228b15f778ef72947fee7a65a4f52114b8440c6c55ab8ca0756b55faedf7919a1672969e88ed1462e8dc6ff40566808a7668493dbee2b4d80168b07;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h3d4a6057f073fafd77dd471e75de43c9e247f36d74d1df179869921a60e2567fc11b9295a183dc3cfae5837bc40081d74e7bd838a94dd6d6eeb70cc1303dae4113a2164a930b013eccbede979042679535a0ce8866934fe298a5ff71214b98ab;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'ha765dd82ba6708330adbc1000173e46c0bec12365c70339bdd5a3ecc423a028470ae2ca04e1fdd0f7605267ff1cee15909e9dc457319405dcfd46adcff244646f413b0df6948cdcaafe22c9ce63a9ffe2642cd5240dc9d5f750fb20e266b9dfe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h7beb317539c00557aac72e933686580a2dd6334d0ddec09a58717e66395bb9cbfa82a38c4aac3521ce01d78ea79af32bbb705ce11f60aac3d22066f45fa2927897db35bcaa4954035bd49b1da663a4b280ed5256c857d050e7ebc8212bff45b2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hc23803b344f10d07ca607dca06cbde48fc55904038879f1685770499c8a093707e0d59ff875a5becc7539c1b25868e443c20c3c3486de83417cfb3bcf8a0f24eed294b39d4f9161ca6d83cc1ac2bffc823a8dd730ee5c29806b8973ed7e7f9dc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h9934cfb9840b0c9200f2459f665396b657099785f2b11835b348bb69e392d8bd691a0f51132fa4257b484bd781966a7e25297802b5b66ba725fe104a42a8d1ef3582150157fe616fe592dc66727d099f4e0715ae6c741aeccc472aa8f1ce1fb8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h7ca0f426470998ae80e6cec42a91cece60d1f5a8ac2d0aa6601abf17b002455712abccdebf43ed004cf6f6c3c6afb5ae0ec4c88119e62823883cff21dce7751b7276bfc8dc78a0da7611101d652b5e82de3e3fbc642387b360f1b3edaa78533;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'he2b2bf01b1d7c752c827fde133682f4d76e8b1f493c7f1e3088c0314c2a9751c945ffedb2474be4286bbcade11352c172808bb3ce8c031d17b75b9d392bd4093aa422dfc6e56f8dd9031d1d8bfeaf5500d7a8f8c80bfd37b9efb6e0986bcfe7f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h7fcab00acdc9bae61ceb6d34a65b9b9915107383459ab58507c43cb69d3b92573da16d579fef0218a49a0b36724902c0f2044bbb60fb7acb5fcddb3d14e9355452a6d2f42cc235e37a4d0c95d9095565ba4334fd6fc7687dca257774f1695791;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h8af0fd24a3a344c3f5545bf6e35cf5c15e5d5f7f0d922d592c25cb9a4aa536b126d2aaffb49a1bdff31aabe9827d1f8c183f59bf8b057b967c86d09993320424a215a6adc80dfd61753c29d4f31708ad9ff5644d157f4b8a99e7e9736ada14cb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h5f51c6c85eae9f309f4cf861d5a8d2c5440f6c30f3dd2d0ef0227873c16d3d9fb3c01fee28db484cf2489fb920572ab64da839be1aa50e7df33ea42e205a7ac835493c3debeb88f448cfbb7b30f95786ef0fceded6ceb3f8fe2053057e4826bc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h7f840f6d16ce117fdaebee18e6d397ae7181db036d117cdefbf94cf25b2bb796eff758dda75898e83b8366660ff52acde9b2658b05c29be29a85c031b9959d7ef1cbf6a78ba4d6714420e34720ac696096eff37e29fa4b83acf92f5b82590ed2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hfdc4b53d65062969944082b947943d646803272641c6edd8f4f61da8c9663eb2b1b592312294ab0b4d0741e54706827ff877db684aa24644430e77da01743575466c4070c01d3a379210ece48045fd6f8cd4db46c7b9901b7554e0601cec8808;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'he3229e23ce8ff19cdaa65fc0e89990ecb12a80aa4935c76c99376ef3d5825911a871b9ff82ab185dadc1baa045d52458f6475146bc34fbd705c823b2630d3e42d478c828f588c190699e4eb2b7d0ff43815bbb9c33d70f2a85f892985315b0f0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h11ffc492aa1767a5052c60be64259e491dbf5872ded1bfaff89590583029eca233edd718f6aeaeb3a77d396f5c7449079208b5b6be816ad6e648b127d7311bd15192b39935f06421a9bb57712739f71917e7542b649765c2de610cbd2ca1d295;
        #1
        $finish();
    end
endmodule
