module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [27:0] src27;
    reg [28:0] src28;
    reg [29:0] src29;
    reg [30:0] src30;
    reg [29:0] src31;
    reg [28:0] src32;
    reg [27:0] src33;
    reg [26:0] src34;
    reg [25:0] src35;
    reg [24:0] src36;
    reg [23:0] src37;
    reg [22:0] src38;
    reg [21:0] src39;
    reg [20:0] src40;
    reg [19:0] src41;
    reg [18:0] src42;
    reg [17:0] src43;
    reg [16:0] src44;
    reg [15:0] src45;
    reg [14:0] src46;
    reg [13:0] src47;
    reg [12:0] src48;
    reg [11:0] src49;
    reg [10:0] src50;
    reg [9:0] src51;
    reg [8:0] src52;
    reg [7:0] src53;
    reg [6:0] src54;
    reg [5:0] src55;
    reg [4:0] src56;
    reg [3:0] src57;
    reg [2:0] src58;
    reg [1:0] src59;
    reg [0:0] src60;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [61:0] srcsum;
    wire [61:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3])<<57) + ((src58[0] + src58[1] + src58[2])<<58) + ((src59[0] + src59[1])<<59) + ((src60[0])<<60);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf485388b3908d6656690ea88de2c1032940f8fb9240c018654b950f155813a4db7f05856797699b285b4088bac89fddb73b487289cee411ba43aba3caad9c9881e9ae17c62c73a435e8e50ceee8a676ba6572af861cf260a6447a7797623ec3ed7633676d98d00368c044473d7fecce89fa1efebc2e5afc1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h145eb80526cf883517f195bc79ad6327c3559bba99352c208efb7a631a1a87f2cc5c5f5fd4c5a41787836f96522b1962dac8645263a5bdf617e1528200446326dfce44c1abb129acc537c09e0b279e7ac73f64934fe6988b8c6101a9c80f9af221972036dabff884cda599557950804c96906e4a60123e155;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a5f74185a97416ae0b507b2395d413fb66774bd9813ef31a728697c3782cf4eeaf43ccec6967ee2852d4d88ec85ecf1699f352ae76b33bec65f376f3694b531c5221cd8187761349033672b0b7fee9307fd78f3cb60e1870dafd1e7bbd565b7d6eaadd9e2eb7085de4be5e2e973a414deca0ed956ff671ed;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h36e922cd1aa898a09507f6fa19089f800020c4da4b520ab9f71ee164720e87192b20e8ec87955fea7681285964df36a81847beaaf1ec4ff3f8f1995c24ffbf0c7e1b9bc7e84819427116181811fd5d9ec91e0c0a54d5dce9da4858ab6b40c5b2097a56f840ecc39785d652351acdd63a4b9655ffa64afc24;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf0868da41a20a4315c921eed326c49f93d35be6a62bc79837a79a1be2149f93f7450cf645778533078a3f6c9f6dd5323cd8c6adacd01300695c7e90d17c01780dbdbe5a55d316083764efea6063ba76303904d3f3cc29effd2d9d15ae5a949c2558308210f6b4d37172cc86c39e6ed1412a6f4680b3f48e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13c089581e9b375dd51ee5ae35f7426b788d723de8677d14494ad11c557154e1b7e5eac84ec3cb3362d9420e2a0e725695af0d936b5d019b732cf189e761b1986ca3156c5380885189a390d96f7de6de0ef5a05f3c4026dbda506eab93cebe05ff66a2c788aaaf23066603f7b7bc136f5e0928129d8821f5a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7ae5cfa38b96885eecfaeac92f294d4e0033ed463d66f0e5685d3dc5c03628b6465f7368234048f6d2d0c549b86d064842a1f326e7679290583f056699105ef5043412fa7b6580f4bcd21f2699160da8dbfddaf7751e03a05fbe84b7244cc6c595250e8b148dc1168db7ca3808efd659a60f4c6794e888c1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1947951c7206598127a4190ea8353f3206f9d7b99c0cecf45b1bed8652580c011be1f2c8726ef74b6290178b4f5a66262363988549fd1f4ebf7afb4a5789ce04b08a57417a6652dd342e016fcff47e4a1fa50ec51c51aee6359fb33a97a26f83a98fd38fdb5df312892da64b03197bfd032f541c3e805b77e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e516d0c7925e76a022aec2dc1efd443989065ebf87d694334e3a28a33e5c76c164cee927af341202b5b430d77a89826ab6d08f9506ff5cdf3686c412fdb6725688c804437cdd26f315a7a760917cd40efc403e848245d2a407aa5acc177668a66d1b94ac33f7e8b8b5c5b4baf504a6ff9c76e5990d66fdf5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e0132ccca0bf02ea35459fd2c4df86897aba4fe20e8ea7af989a17a9eb633590d0fee779a2a5f1de40f69670b57160662cd7bc886ca7240720e0dead11e8ab774ab824f36e7feb0220d6f4f2b0be8a401cd1c0d630f68b3cba1ed925199e0a7bcc001211392e6a8fc3620f01aa070d4bdcf34ef94cf55b5b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h383b23666477bfcb4c8346b1dcf8130eb3745b455e0cbbba2040b15052c47d88d9b0c7144209021947282d5677ebc7c6dd7d7bde4e386799ac6298235c8684c197b28e87d8257d4aed13000fcf8c79a8249ff810f2ad05e61ed2d62c5fa4a92714a68faf9e810e2b233264cc7396f56d06b17e1f683ae0a0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd320388eb27bca9c7776fd6b58cc6a28b3e798f73632d38504ff79616c0c51285f2d17ffcb89b2080e4a9362f2bfc07a113c4e5581950d9eddddf606ead2e67e487cb967057b7b6f76f05113057bbd0a5294cdfb2d6d21e8776804af11ad3f087c3eacf78b3e8615e9c7709454e4789711248eaf53e581e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16e5f6944c40533e2e1660ce80044287fde9919fd35ed6e0ad29ad2a3cf7148c707b659cdf418c443b90560b7708f8d313cedbceb00a2ac2f15b013b92f7433289d110d596f6ad5a51d1363552473e53d6980db1cf2368e0dc5a41b247daed4b25fb8cac99a6c0c267e9f7108777a1dc7e0b2e17cbab1d4b1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he923d7a14c0eafeb39e9d491db968626a80eb1c2a41d85a42b782a078378d201b0c450dfc422b3a6ba7fbec0590c69abba061509883ed559ee3117aa176dd42b5cad5da3eef690aaba05712cd4ad271732b33c5c6011aebc642baf17b68641c680b03191916604ed467426926cc7ef8897a564a5ba87c43b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbdc2eae391c9738c12dbc97f9fd99d4746559c5a2012cc2d9d64a68f9eacd4209e1d4b3cb32ad84e13fafe92c17f4204f10173cd6b09493f1d85f0ca3385cf40e3b34537ef321d18440153d1fe4f771c0bf1b65da271fdfbf6f109963fc8bbdfd8174ec950512ca46bd3d00b8632d4754baa415103099aa7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc2686086da604a8fde3c276441b893eed74870df94285cb982c3f2560752c89edb5b971f51fd7f139b56e095e11373ac6b3ee68f24fe4a20a072010aad9a2fdf4de6681ef0d2ad47d9aaa37cf01667c5062a47712400c4a6d85ff79694ce8da78d912b55c1235e515042f47eb2a40dca695e22df7dea0e82;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf2e96f2ff1d8a0188eae8c21eeb5d0123c10b97384546c50c3ffd2b607ebecda3e2dadb0ad0f1cf8e65311ececa14a8736999e706d707cfa3f32bdc4d5e76ff3f87b85c49a486229c927c29920f91f54ffdfac2db0ed56fa68e6dfe802cf9b95c8bd8f0e1b8061d7974fed5beb747c841d31e1d27826663c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dd8f0806983dcca361323ea97156b53b99e312d9ff396a3daf4d269ad86158ffdada12ee42f150259e30e50049142710b004853b7be5a42e0f50c3730f2902f9c47c02a19c9a04a0726b3a99823e8ca3888ff6c409779c64d2c11cdc8688e5c60f52d7ad9f9e0926dee1b2854adf02ff10e4ab1f638b1a9f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a8cda5075749ea3539eee1eb6f4c92fc712e9cec881f48146ef199081c3a3e2320c3c9b4532c5016ec4267a0cd206daec48b4edeabd50e3317a1e196c5bf1b37b960aa3bbc82c2d97d905fbee8a61854f5555f83f4aa8eac9c15b58434317b540dcbf623f58c0f082fd79db88be66587d05edb358859819f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h186e8f45bdbb2dff1e22237b5f56ddc33f7055106acaffd5a5c11b0182bce432e22d6698cbf03fcb3c85b75ad5710359303ce0f54dfff62a99e03c041cf313a1413cac39f598ce187ddede25d5d65183241d1de42f72d7cad5642977002b364f0e7a4ddfcac5eb08a67f65aedfcd54504e0a68b8ad9a09a7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hebe7270a97a0efdab07183f40ffab73ede834aca3d7b65577b982ae2a9a465afaddaab74a13d83301ee130e1df7964d6e1d9a12e88409099e691bb902e6837ba24bb48b92925bd4df86ac9dde4c7cc818b3e4fe9eb78345da4b7aa6c131e67d396f6d1ef3fef6f1275d8c39252137aa9b025ccf0fb9c6c54;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h106eb209d77e8dde178643aaa83f350fed739a89f0944847afbec06bbccf4713494e91f462aedee8e85a761a7b3a2287a8fae5e19e867db8d28eed13dd64a4a2e46d774f3805f30758bacb4fa72fb36a9f185bb24dba3797360993b67f307b32a9881582699166a3655ee7c96853fa013752fba3b15d7e748;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc6b497f09ab6c8cad8ce3e9d1e16ef6cab03f261068e48a95420a17fd37189d13e8cd750c8da4e7ba388f2679c1de69362774088950ce2f7f28361e452ec9fe679352bd0d895e28afaa9e5d21375b0e456842be35bc64077cbf86ab7c68349b483c854ca582f75224366711c5bf7e76110d764f57141e107;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb372573ffbe7589addc67a99ded521de2a7ad945ed3d2761325108f5fc4c0734f4ba465337d5d1645cce52687feb2d25a108c89564bf3068e96b02f227511f4cacfa624082392ecb12d2fc4b6574c5bfeed7ea7fdd427e91d829730e531946e7f180a5e478fec207210089ab645eefd50d1a01526a65bd3d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h53886a0cb2cc401f9f4603bff33c5c905d4bc12df541affed0f5090ce9c6e685a02a183e4b10d58c576d9a73571fc0f1aa3cfa96f8653fedb8ec4fd55a445dfb4f831777b3218109a8b34ac616715a1feedc79e9259f5d37fca1792b88aaf2532acf0d74d35faff2a13579efb839df964848145e72b96289;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h616a13c7127c522cdb49f1da34e3ffe7558d7122ec0bdf8b96be9e3913dbb46f58da40a3b159aba04a3dd873f95cdbc43122fd91ad3b6c3e5c739007301bda07afb2efaea898dce3e986c9d2e9e680f2e33367f92d43a711ae698e909552f958637e4e61d310cc8847f363a5699bc561845c9c9defdfa80b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h160db639b1170556b98a648bd22bb136846a63c00d16dc8993bb3408dddb4d6a7d30c2354337616e3caed630bc19615cde48e27f2b4f5f39158f65e4cde85b332ac4540218a0dd04fbd96454ca70967757f249614dc80ecec5eb1c7377700bc55df0594aabea4670dfa956ed521f2a31f490864e9044117f0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h196bb35bc0334d5c14a37759a5fb0687e2145650732e4cf5692001645b0494d06322083a621605e5ab0e4eba0a0e31bef64fd839f3f0f78c2fc35eb8651c3d31b0396e4e17e445c2b85c041d83a36e5575b10265c83bedb43dcfab48455a782794d9766e1fff2ba2c45bbbea7c4c03f5b5868bddec9362446;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h25e6b93fc41593400d09ecf5f16c0ad7ad7af0a6039f6f6eb30849552a776ac819ac121324cd43e4f69aa7680fff3e8914b93b62980acb40fcbf51c43877ea7fce33b50738bd73ee1d5603cf22bbad203c4bc454f775f894affc15c6776e6d8cf59bc330d3610c31441b405e175f87ae2be611cd841fb42d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4f52f8c67677c477ca2b24717399979bd40c305d40265ed95a9b2f236859b14471ff0909004d0eabd594ac0f284698960921a99a575160053e619a8c0aefa845d363faa0b92a36899b74f87495d069d547e8a76c12f3bd38870cd068b7801c650eb23432a3eaa1071100f9a2f9e904b82f3f51051d945394;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c6efbec7e3150b21c4a3a983de65e529568a79b894a0b3cf7ae6bc46e0961bf261024c03608c06663d03096d53af108979b6f891c8b15db8545a4d7104132c55d4a60cef9bbdce2a3f4409b497496db13f42908ec844a1fc6cd1e724eecedaf4306a7a6f1b2a6ccef0162790fc9f45bcd446a24707828d00;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f47ac16e24f0227f3c22a6ee4e3731f0044e86103e731194a34ba1366db2af4ada640c86a3557734ed98f8e698a086294c1d065da90777d3ec7c46c934551fda467bb375ce9e6be681312332a811c6fa355e9ce4534ba5ec80d05f170075344e8ff6c84b73184ae18850342f70561dd9e485df75b8873f8a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16c3d0fc68ba76f16d6971525d9367b518e82815b6b79129dbf660da8a7eb6db8d78a4708409f744b600254f2c2c2649c769ccad762e406b5dc498f5e8e23838535f151cd14560baa868dc532f7d8527e466d33cb31077a5206b6d55e5938b7d1d35a526024a1b85deb23b32983e8b24e4b3137ec1bd898aa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he636bc5188d5aff1e38eb75063232105b0600de3222c7e5301859e2509528b0a64fdcabacf533a3785687fdbf78ffb6435eb8d811c68e770ab65ff6cc5734b7840538bbc1efc4b0f458fe3d73be8d7321e513195038de1014f7ff9d213519d7e2a332cc9d3757c5831bb104aef0d13b7972f68072a98881f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcad34e5fe981ca6c3b5a38def9f8669819e1f889ccb8f2e428daca9fd116785c117a3cb2c17d792c9eae1e8b8590a52e5e331020a3219f1683b05245cc1fb28a58f67bb09e96121c4a2027f1411ca7b662046c331e68214cece90335b156d3078c74166f2539a5d6d7e4aac57096363b95c432533d20725d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8fea0da7d608595090014acad012dac6eeb35599bcb5a1c5f82248897326891760a171f86606debcb58a9960b1d081b29c9a4859547bc9a71edddafbc8e63d6ff7045aef2edc6297843f28e5579443b125d27382a92b7115334426329cd672ef2dada3c3e7382e508279232d9c6bc20c93d17223acab7aa3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c7d6343d817a05f2a85747904741f998a1c3dd068497805f2c246e690e05bdf4cf8cd835b113c59506c9393affc734964c7662654b23f860a57d4247cebd637e4b660f90e52ef83a797b4744a739862a120164861bc01cb21ac27da778576c789b938144ff3a6c9ef7adcb24c0742c82f18dc9ebff879442;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h56b8985e19ac67a215184811b1e383e2a1ed1252c22cd1d372ca39596a3849276e07c2aa4af243aef0cc57926535dad0b025da7d77376b752fb1cd8add395a9ad56dd8ee119e0d5cc71c82acee6cdf4fb162ee57c6c5422fe90982563411056e44705719fdf10249209bd9b11c22686344c314e7d756cdd6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h23c85f7b106193c5db7a999c8ef093bdc893adbe4d1f8ab37d70187cb4a343dc5279bc0bc9f1427a22e14644929f4627c0b398c2dd3d5f4a8003bd71f8dd208bef835b34f3ef6531971833743c827819cbee212895b2ade64c89c4c1be538920fabd49bf4bdf3f02e2713c02ac219b3d624ec50a6bd656ff;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1675c4faa24ff29d90b144cee371a1f324bde1ea805953185b4445a38a95b70a5c98638c440a909f9e0b1340dba5f2fca7afd21c3af409b5f25d979491b03a0d7719820009fd4e7f98cbda13a5a44e4f2b0f26a6b091ff75e3147df250ad9003f0658a6268b86e9b1def78a053f721da3758ec12e16315e72;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4ea2e76df1a6e8e8a70d122d14b46df7d7e4a883641e78e29fe8a5de48a42744ae62cdc512cd3313388ca94e283cb5552eab86b9d1f1afa8b09e81b30057b9fd906da1d9a14cb3ffeb9245d51a145f2e3f19b2a6f1eff8eba5d0afbb20fce67aeb2469937fb3f43697903ae827f499fbba94e7e4a6f2026e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf881e84d2a57e10cacd9f5f4c1ca6b74d156ffe6927f311896288a3144be2a726d700984105fb34756f6faa3b9f07875056fa9cda7b2b15f5efe351cc37705c8ea77147b6b9fcf3d2bae1f07d34feb218d5aa0ff402e5f05be37a560172cc1e0580990494b6a037b432e62947d7fabaa2ae61deca68a8ad1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h111e788c49df1bffe2828c6ae6666f3ca7c0e47e8b178130b0c1bf62459381e62c4d9d9e3751b6790671f4fa8e8466af547547209552dce8955e2276d28bd1e91142e5b43dbd9cdae4c9e0cb94f36110212514c4dd3475048a060e1db1814fa0ea21c4fdce2be3d485b7db61c23705e7724aab147a881f48e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17b6c742e3ee068e0c795c230db57e5199b5b9f5ae27647cd178535e15ec25ba650faf3450a0d14a7cac1570402a1d2f3d7d40f3b96bd1b3e716fd5e3375f367d8194692076465b7f03af0941bbf01b466f2d56cc6821def1dae3532903a7ad3503e3753f8dae2aa96a80d89e6cbcd62703ba8cbdc49ffb19;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h129e15bcf8efef3b7da2ddc13cdddebdb13d1149d868c0e183b91554a560416a536cbd7f4c9c1a977bd0e3d6e78417c8f9cd1d9323398ff43509d87dcb086bbedc61932b3660d43efdca43a42387237e3860b4b06cfa6ae343f838d44a95e5e97a92f6832c76adbf58b268930340b9062baee9df668751f08;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14271132cf7d28fb206fe1fddb4a78cc4e74b91fe31b6b3927ea6efac721a27f8d32099ecf4dfeeb7648d1631a18816289550832f570e0385e8f227a6f2c7c14f88b3a77871e491b658b5463181abe6171eb2e006797d4a0eea2ce7ec5f86c8215190387f885eac2b5efbfd41757c69c3eb323ee206028e67;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h400f5d0e0df05df3bf714c039b2f4017e629423df9fdfd967acb688020b1642bf54e71f39055888e23246e3d1a9514bec62d9a2ea636aa9569784c9257bf94fbbb5d737101deed4f5a4c7479e5ddd62e8c3626e23eda1dc220442cebbd10b7d73ef91faff376ceca1d6842a421d6cd0f375ea80f3c4e3a88;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf5b2efe96185681364cc3321afe8333f8696b0143d6027c0b994dc46ef29f7e4f68819a941cb2e9a93e5d482d8f2aefdd3e71371beedb90a671729ad5b3b440ffac04126e937ffc980ee2c47bc7fe285e99168d6c79de92a50f6a43a0d8b191cfbc02ac6c357bdd08f6c18b2f412997e57daf0c991f0d852;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'had078d4bb2e602c705cc0ee834292d6757a5ce19fb41c794c32de07074524e015ead01fb64584ca20f2e463e7007068c30ef822f39d07aefd33b377c1e233f817e8ae5fb472aabdc96885acedbbcd177221fe1b6b72cef9e4a926c9cbb3f5d1012367b7042497a08cb748511d1615e5913bf1bfb1418a355;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h420ba1066e938d92c3b32617b75bfc76f4417b6d6612c25ab38fb42e94c56e42593e3aa2c143211072c4d78de219d7f41df2f66cf4be5dfd65f356678813db49f72284cbd441893667f3a95a9f2227f9d504e325cbbf4c72aac5199a51a291c50ea33e8f0223bc44bfa624367876793d8db10e6c80ae24fc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1554abf9a725b4fdd0da018a9e2e368bf3ae650b94be5eb93b9424db0a647cf987bf5e21239b92e8d28b7761bc4d31f880d85c4bfae11b50304c03bc1c5cd1fe8605fb8ff69e159527c1b86f4606965d172ada53dba9060d8fea09c6e8f01e1e02d0edcf5f553a7c1d26ad41299e4b3c5e7a9b44a4afba48d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9c0cfa102ba678eba542ccecf91ad2ddff8d1fda55ba221afc8d47689a6f4357b02b5bc249b20c5acdf8940e8282bf6084587f3243f636c077f478f732648a56bdf8eeef54b4b86faabbcb86394a8bc05fa7fb963c25e3e6d9a8327944f957b3d413de0c4ab5f1f5f64f28dd77402d5887c7e216f6bacc16;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbf89b8d03cb5f64ae29a29309c66d2b1b0a398340d186fce6193d976da6c7a6dd6524942f7d918c551ba8e66f27d4140b5db5b4e9812e7f10f5b64c2a05d74d7b50168267e580740f75dad40868d521765a42e52da53bc6ae4b0b11fe925adde8b5a03a8e5d4423312ef20bcda86e4f19eb43460445709aa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4429cb405354becf03c2dfee7c44306981bf1960e0c57104f677d26f527aa3ea1e761dfa238a57d75c97e0c54452465bfbd541a3dd6cbd2d940e4c6b1848bb6a0cc9d673549551c9379e9a1355f520ed99e8232979aca7fd8bcfe7d9c7797f179a5b949aa6cc83d2354a7ee40c26a905846f89431db37a9a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dbc9376c8027ef8b16c88b3c9bb7fdad6aef206373913555d85d8dbf51a28794ef79189b1be795479e525ccea316db522af68f85f13eeaa698857b9a558cca3878aa396064def488d42a593023a2300207a048263be0f8e020832a289264a583627dd62b8333d74b94f904656ca330041b6b8ecee3b4d2cf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e2346c0b1373377181e42bba95c70378c5a5de8b58e5126dfe03c3ab71a474b1d75f1aa0174d4451a4c00d1380cfcf887c2fffd52139a4c51a696dfd20fce7ac8c04d49fa81b368a478cf3549bb2b9ad0bec41a0a7b4fadeffd8bde94ab8d713dad574f60470b1e006b7803ff6b73d2f41048d20e5b2fcde;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd67301bc97cbc5ab27cf480bc8860148583e956977aaefa56de332109e158f221fd46cd28f41d0cd5c2d034a8b0be041506b4d166127a7845c79e4048014418417145316c1ae4f315db2fba89fa094343cd78bbabc98316580b127e3b57a5197e997d4ce54b9323f3f4a64690e5276000be08bac46920a50;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4a6fc764c32ef0f02f63375a4a3a5904f018754de9ce28c1e75666f5237328c26c7d542582b0c70896dcfff9c4b380e6d09d14462b5805ae56b674fb422f4203cac24d085328ec2ec154e7cb5d35eacde6d6f928511b1cdebcdbf7a749f17ddf07a9602fc5bf173fe04e06b1c4ce5a35c1fe40cd4afd265f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f2e67030c68810862c6af838fd2a53f13bf869a0e21b4fc00b11d5bf025954a5acd72d71b53c7531a4d947b311139ea7da017e591704026dfe035e64152f722b6ef0945082df2a32493c50ad1381d9f27b2c3f0730ccb6e26d9cb104f6d06bdc6165bd81b88d59b8387f3f3d3ea5b120fb7e67a9372a6fb1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb8a6d6326cc3fb490319a8b01102163c40da6c653cc9f16a2dff3677efed724ec81b94fbb71799b1bbb33de1b33b326c9d8f9d509d11f422b22cdd1b32b554268509553cc64578e54050fe9da0f1cfb08e80f12a0bd6bcf06749cc70af133b5c0648176df9a563485bb934dfb26ead7ceaec369fdaa74b5a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf00bce4d4e1b3eca75477491b83eaa024450cc62fa7b8a9ef58b5a4bc1e32ca682753ae18028ef7040b37162ed2421fe8bdaf2000733d757d3c4ff37050b651de9ae021a9269259ed4a8b851342cc58c85cea1026713b6479da26477e46bff033180614b75cf5414dce47685c40fc22295a403d5e5a6a363;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12e1dc2c61a56f56354511b777808954b819d826592054d4c777145e2ac98fb52b3ef51f912b6ffad02421f02d9f12be102782d1326afae0251ca62c2d460fa17040e1668449964505ca074a0213599b6b839a9cf664baca014486085d61a076afeaa4c64f2bd189e0188d345bb0cde4cbed508695360729c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h703f96b500bc3f3dde8f8e09043a185c18f0d1a9bc4af7e460d33e274df8d22d45d51d09a36851f86bc3255b5a0fecd54c95f5bcaba9dded3a6be6d78398cb9143064aed7fa22ec75675dc790f98858d8623fccd7c73e2b6bb22efd19a0cdc7736453dcd0b63f25e60f6acc4189921f9b926fd1274b3d0d0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1befdd3a4ef314757409b2b232a229c2362a46fdfd50ba6a4d27c569783c899ce2c47efa62e21e4c93a5eb5f9479a075512c35caea8c83b2869b8a78b846551e391868b5677a0d0adfde407deddf882deb353fb8df8fc2536dfedb76f59309a4e45602f880db4b30a895aca26c76c471c472353f0c6fea686;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haefddf4dacc7f89feb6dd4f9b90c9bb405b8895202030848fd82e84d7af3f69090cc88f448aa9a7b293a27dc87ad62ae977988019c256e8049e00f39db91cefd1af5e14d59592239e185d9df9c3aae40e9ae4424796bbef566e5613bdee727093a1f6ab3527b6c912563c207f332909e27c025f0475cf61d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4c7c2aff63de045c000a249c06675cabca92cd27e2f7243a4af3f35092a61076d71fd5d2c4eda3b57cd9d2d4631512c5baf9801694e7a3304a1baa2971e2cf131e31160a3152cd953005324da5f6cc7940f8a5df402e97838bf2f043b6c55b337d087150304641e29e6de0e9330e0ffa6f5d9d712e6843d4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1badbeddbbcfb80c7d8890cf904fcf1460f17c01d3faf0503bc5d241dbb1c314052aceb6392f4a2de5f2d68b62e7371c27a7f4d9452a45f20d59af35aae15a211fa01e7607689f3f8506ae0253f1da1065bd9801233bbdabc711655b02f71e1d2de45b50719876569c73af0db950a6d364df6e5eaf6d78115;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4120ed7426c1e1b0260c52828b3d782866e94a41b53ff34bf0b1c3b2e31a9e0fab1e78ad55e6d718ad4ae0307237285f2d7cca15bcea558ecf6bb89a6eedebe0d081295e35958dfd03d49d6fbcf7bed48505519f1b19c0a7863038bfbdcfe403bbe4877622fdeb460b4b021b59cf1f0451c0e9e1f520e77;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h654bbc5afce25ea1f7989b49df5159f2136a56fd13b38204bb9b92bad90042c94112894b415fc400b7de3c58d674f57a69228349a5261af928157a6c50bd307505dd036d8b9d366148962e5f5018a703c592ea3599dc83157649b0a64b5917e65979d64d96d6d6efa4d3985cd3e297aa8ee6dddc2206285a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15bd3b73a8e16a7e49d22ef81fe9aa561018d2b0979d23aee015c43000773ab236aa55d447793ebbc6a8fa57c6026cc73e6433fb0df661b1b301ad9393c89a9ba06971bd707e07c0d2f7be219810ad4840f890deac7c9caaf54517cb76dcff002fc6915a5fb1287f4181d18237c517de55cbd3b6bf6d768c6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hccac8cd89ef948a01844e78f3faa85faaf97abc3d202e5ab352786f65f6d2aab6870a2d145e9cc80504258899f4ea82e1dfb8a8ec3ca1533ba48382663c94a976c10e1d60bfb996447dd6529616e1c6f7410c684e5d20d136f88d4edbf17708416b6f14e92ae7c29f1dee6d5d6dc5e5ed529d669a5371382;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hde0ea9cde3de0aa4c1e5ce3e9997eb9b2a7fc82d4d5a627dae1e6f0b19abd7fe00ed72b5cc24674bd8f20188d9eba96a5f91f6e4db1c943ae6c06ab037b959de6660a6cf2861bc3fb605c287aa770be2967a0b5e6b168013d5a49388d1f6c4dcd607493a35e939c36de2f9dcf6e7ed914bf6958479e3c440;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h377369c9cfe626a6b41cacc91615d0df6dbfafa2370f0a4611007199bf8a53e8ab89e1ccca71c228ca53beae091e513e373210bbcd830db7798de98ca2892ce6653f72ed08aa8ad5ca4cce0a77004a2cf7b1b5cc7e93a503d662381e25ea335e342bfd4ffed54b498371d43d49044efe9891a65376ef38f1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcb626f1e142a3b38d1d3bdd74d96b65169a4c0f93434ab96a0b8da9b7a59285b6064a1972af3d4671142e91c8298db25c5484984ee31ecf7e6cff6e55a84f4fe5dc8ef9d04b2b424f4a5e7e0da6cd23eb9217d2ce997d9346b9d7f992fa513b40bd757549b2b55eafa52e157444f428741dca5417a0cbbef;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha4f5626d8221650088d9e85fae8215589939bdfafcbfdfb0524c4d74a08b2e3670ae75891bed779f4567b8e19ebb89ec72e818c2e8aa1c9c288f70cdb845fe47b3598f6a3d1d51b67dae30b74e663f6fbe23c8ead4339fdf35d942fcce107f6ef387438e2783f9ca6f7faa1d5ad5da24aba98f6c548b2653;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2ea83903866a72305be425b3687e3aaf9a3deb64a4fb003d8e7597d44b330e6d00b0504fe0234324e00110b18006cf9b7e7094b78ddf49975a0b984d27cfaafbfdd3261ed26b71cddf8068efb2e49269949f074ef6de673076ded780dcbb9c947c1d0299933875474abd6729fe95fafe9adb7142d976b6da;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h62e7508076544053d0bc39f8600a96ae33307fc2f7902516b710e4c13cd70bdfd6bd8370782c4e643b30142170e6a4d92496ee020ccee3eb26428bad9ebc3bfb38bfdcf4567ed96f8a6c54e488e08e08af35ce875935baebd2a7238d17b7a836aee13f640530f4cfcaf022900aac97990c1838c1d0d35edf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h91be5334f6e64481c0af82fdc2a1942239b52a1a20c88d7efc573f8a5a1fbb30605b63869d433ab2d58ec5d97ccf8d6acc6d33493fed473fcd828dc384fed45864c64ca4bb2125962c179d338143a53dd902f7794b00188dd4a50d970185408a4a5e58729e3c67d4309e74fa9d7d847ce10fd47f61835e7c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b2480aa5c9ae0538eb9685d2cb7fb6e17d9b168406dc48a5d095f8ae9a4deb57cc15791d4422918ba4544a38bd8a8b359e57d06703f6853877f29e8f52c922a51ba5f4364f2eb9c2b99841cf94237d6eb9bde2bf47a7a432832ad45020ce24de5f69d9c45aa22d88661e60a89a0e8868990d4bb53b42038;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h72e6364a7b9d0e1b6afc757a2f2301de11b19604c06b8e39cd66ba3885c7cb88f7bfa2e8f6800a8d6124d1135fc484302a24704e9f43e723933459c5515956085d2d0c419fc4023ddf1a9a303dd63084dd751983584ea606c3a41281ec7600dbbaf9574a36908aba98e485ddec7168c7ebaef36141b79b4b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ec9ba80dfaaec108a5429b007b010bf9f9a3112ae6f91fa361714011c80c9a654252e12a0117e8e923927a0a36da03a5455a59877b041865b74f0f6b19f9a4c030940866cbc02bbe3809c3edda891344969634e6b5b8e0675f1b4bdf2184aed9e6faf1e5875aa388f458dea8814697c23d5665852c583bbb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h27219acfeff59b61578bc408e5258dfaa13462cf41d7f697d2ca0945aa69b90ca08328e2d7dec79efae3285a0a4a7c22af601ef9a0a5c1021a2e71ede15668f5f023b28ef1fdfb00f3445ab18189b6980622f71a9afb8c882ada9ccdeb765accfcfd67fe4cf78cbd3054f36f0de88f68e961b53844d8ea7f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1118817407f60dfddcf2989f4d8844a583bd504541014262b52afd4624fa03dff3a63b14b5c8c4f01b371ee8a8796bd24a1470068e5d8cd01e53325cd2cc4003070e190667d4e4f250df90c1bfa45151dc987cd551c3d81d677943b3dc7822e9a004203cf0e9d8879857d514c436a5a97f0e799b4e49920c0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha00bc57e3ee8f9c4b73ae411e6635c10803358ab5850ed318d7fc12c98f60e20170b4276030120defbc2d93f6ea5dac50d075747d65abc11b71a0ac0336711426a737b572797ad32ec3eb2aa4a26fd3a901c87b91b351327ff534a2d9015064b5cf5de0391de4c189f2ffb695d8ba398c483329396ead7f3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b49f79fcd2b74d694881e089f0e859053b044586d332ceae8f04bb0a23eacf570c219422eb2b2aad0189cf59b9ddd7367fa18af3adc135ba9b77c5f584446e9238f220efbb8062960c49605ae6e547e9b1d86e3281eb3761614193b20c980198e327cfaa0e84b93cb003ff4b729df2262a19f8322ab3901;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1758d141b7a96295d6f3679617ce4820858bc3e26c4a889847d8c6a485deff7a2e1cdb65b8ed569edf0c98894c5632945eb623d0517c10056950c6706c72886273ae45f98ad6957fa9091fbe5c74b25a44b57c0c1a2578c67c9a33c5b27b1849d2a83d3535ebffabf7bde335c409559e18d32a0496bdf3cbb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12e8e0a34997341d7a2a2ad7d9a25d75aa802189edbbd14c916f324036737b88afd1af78db41adbd72cbf575bc4aba55592a97fcfdee8987f67ee1d6f54fc5dd4267cb7d9be719687f2cc3609fef0b873be5466db58e512305225a7c7b334c8a9cbf2dc14628f0e0210979e7bd4c9372a4aac0b1759cfd061;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h97835604c6efcba8e06457d6353879d1f6306f3806d8ce55ad15d07619f8b30638e596e031c490a9b91ff12836ce0dd345e4c3276e2dcd60c8b4a657eca07d8238c8948e77f833abc26baac166f7fbef2a44fff2f422074b4d49246a764e680da299aec1ea664f070dba87ac12f1c7e1c799f768187c89de;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6cc994d27efaa0586c206177f561a80ecb9b260cdbbc676c34f4c08f18371fff473fd1ea22050e9ba204aeb92b7aa147e6b53a93c54668107b31be215e2e6befa62ac50fe7f118ee369d4d8ef74e4e7c03e755aea80b010930d10adfa15d49e99d17a0c5d5212be5281ec193a3231afd5642f5f67ede6baf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e71d879d938a5f6da53ca2ab07c1607e21f9d7568b9d030bce8885988a419f5031bd989db8bef252b4483b73440396874fb85ffe1a2e5e51790431c019362748009dfc029f59aa2f0ddf19e39111bc0cf3153478f1d54e5f40a26b6a42a3ec0b3ac39a69a13eeeb65b8d60e5f21e809fb556e39e807d06f3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6b4757b59c0a5e5c0fd193b6230904311050a24fee2f032106c704353da508bad87eed028637e0bd48910523665e803162052c47e3ad9054f42decf5b0f8fe55d4b648f14baf56c2de4374215dedefa1d8cf88cc56300f8e65873679a6281caa60bff95826708fd2fad69dd9f01244452add1b3563a9f87f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1593a6034355641f2d8f1d6c7695cfd481d9d90089fe61195e80f32b9626fc6b3828100e75f04df0c6d835ae81afaf216df0b4091eb08fdcf3db0098a65598c6ad83fc7e94b515b9be632bbece44b1be8aac2aed78817ea1c515276b2ccec5f2156cdbdf5e34c377d34e29b8dd08b52eae677c7d8e95b5640;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h325e9fbd22736a333ab8cf9cd1906104785b1201f63486e1e3284ad3b5f5d049704a3ebf02a6553ff41daf3823c32eda683d174f1ef8300ca7cbf567cb59195dc4cea76e67278998e0a18f4b9afab12da2898c2616f4ee24442c2605232bc8ee4b503c11206a46a8936756af9824484cd1d2b942c856ff4e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdd28acdaabcb7ea4ef0803bde5e8f45ff3790e143374dca9da81d4213285942ad6d5d4b7846c4f82a965d020c3f46764aa750386bd03022877eecb2b9ab3c3fc8fd3586ad17fe54cc5fa87f6b5e8afcf92347d361c67eb84e65163979518cdc0bfab0782f3a500f2fa27fe40de7c335294d5f65f9db24880;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1de89740105f357cf8ae84c323cb8be4daa71ec2106128ec2285351ae6e22731577aacb9778ef7f995ef736f03dc2d6971bc41c55b3e0c8179110d37bfd64d2db23c83d4c6544d2efc6c4823023af2733b46c8129fe05a4d282df995e874b735f04babc1c9d8e37cc671b111f29eef616a04a9f5863480b44;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15b6ea4be2cae97378474a809f23f36713e30716280e016464157f1931f3bc32b856cbf4a67cade103ce00df4bbd3cdc7260b75043f8ab4a74bd7f924dfcc52c3d13deb4b800ac2d91616584487aaecabcf83c0bdf9530461d1c08e61b7e52a1a501672d1eaf6fbb3f8e1cc3084aeb0729b719af90bd3611b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h159895cbb5696922f9a8a28a33252783aac1da36a6489770289fe91ab50aa58c9a63307cefa89c8ff9efedcbb5b605ddc905f6a68efe38a016983eae2d7e043f9dbab9091dad3eb6b6464ea8b41cf5c404aa2b6d9ada09be921453f8608e1b0a15592613a2f7f281bf9c9ffa138008ceaf9d5f8784f48cfaa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hffa6858e1267dfbce18b1d998f4074d75c3f3ec777eb7b7b07e3d0c5095c0761eac34aefffe668e80390f68c3f6c466872790a56dc814799bdd0ab98d56e7e24b0721f84ddda02870baf1220e6915df9988829adc79eb626a92a65d8d4982698428cd9bcfbfe0a5b67667eab781b4cfd47ce3f15b8031887;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16909270138793c3e1c3d44b813662ec54c902b00cab88fb2ba565eb4276e7d77ae66bb21d7b2514bf2cd3c5b576579519e674314950997b6006a91ed2baae74072f9de56f0ecaf1362ba896a2ae46b83d6003a8f68f3a5c5f5d5c90048eca0441b6a55a2155efc87919a9364e3ad6b1868d7ee8d48a1086e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha477035ea9a6c6f91f3f750fc5cbd716f12eb760a8f57f8c5e5be2935ee7f916f2ac4d3ac9928916485bae8a939716adfed8acea128c61687438f3ecd5b06bab41fcd8c1aa3af43373f0be2d22546c85b74b71940a57dba59be5ac2c1f2590d614c9f4fd40c6a91db7b098dff22466ecce5dbda2cff6bf9b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b5be6f1e54c17ded794f4527f70c7b80b55612d6ee8246f2c7c98e8b42c0d77d95a74c9c1474e2ca4b2f12c79a07613143c184a25d14ef0b1f0e54dc24f5d07d6b7ff22338b25ea946bcbb0c24b0ee651752a10f7e5eeb12150c586c3996491f63f292cf8bc51d348072a6986e616780290947f4f3248f3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2bc357bd757e5fb2524fc40d5cf82c94f757832c0d149d184d282bbd382abf2fb6c6fe5bb4e8bc4fe743ad2068e0b0d0276a30d0a0b38adfab58368558d7dc82e6c373abfdf31ba52b075c862b8c3600ae39f1c65f2dab8eeb233f7d957a7157975174b1c131129f86b1800947cfd714701d3e8c62934768;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8ee86a1ee92533566aa54a9f0adc7368370107650d57dea5c46b21f535d8322d10c293d29512b04fc37dd267c3252aefe38a713fe7b4d9ad69b336b5363b786b13d1522b367c0d6359292116ad1b2394dfce40b8145e3f9cb001c91c2c1fce298eb2294d7ec5666e41aed57b062b9ccf647ef30734c3cfcf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b8c01748a5484435dcf2db135244ab7bef993ddf8ac5656b150ff2ce8ca3b1b56cb154a6b462e17bdfa097b06797946f35ada25ebb02e615cae18dcb13d7befaaa3445c25772830bd9ae8413dd85a0501af59e465e3499a9681ec61a26e4c5606bb9ae029af0cbebd3175f1fe36d057191db23c85836154c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d79aa27d36cfb9dee60af98d51392f0348485eb5234bae770e09bcd1e4b410bc75652e664202b22f00fbba168d5ac742ba269b39d75b9be144e1e3bfe0b7f13ef008515f74f5b46254a82853a9faf023a59b270cedcd40ced0c363f36919a9f90502e353dddeb08ac6436172b09a0519b1bce697fb3290df;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha68aee50ca35faca99fab2ec8037a535bdbd726c82a6749bf3bbff7fba01d36f49bb28413db364c59ec3b4fdcc1c45997eb59d950e257775175660b2048b0a7c5072a2cfd20abb85878b68ae4c2157e995912c5160b6b25b28b02471df99721e8f836f1915b9ff8793ff11eebca6732f27368679576082fa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h170a59bd55e1cb974f477de848abfd206ddf6d33af4984b36794ceb009bf73802a65f413b2dccb7c5b7b1d1495fee1c99fdd947d964951db952e198503860c6a2f4171a907ee180cdf059915074a9ad4e06c82763ef281d25e63a13bdf98cb350a8cd0ac9d4bbbb04193b34794c2f0aee5f270b8deb6a813;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b48ccdcb2cda7b37c9094a4f4483ab9b8fb518b290d5cc63c5dab2c15c81260eac757b1dd2766faf549e12303c3b92cc4758e85a813e028da4f43dc30fddb331febaa858effda78df8b22cc3dd08c6e18641d9f8718f68baae99e04f83a7a238d1e01401d3d20832ca72ee9a837b1a55758855d5daadb320;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1597abe23a5a44f9b42a6131bd2079cb3c7c73dad2e56e02df91c6108db22c8dbd7cb732025e08cd70da6a69ac8575ba3690d89ee7d0096671d505008df6376c9be7483e79f2dae24ccb91df2a7007a564f6ff99c18ca74cd603e1bc0248f75ad7208f06fd5030d64eaf3990d980671e7d8f8c2b5bdf50b24;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ef5c8314448ea3991181eb388519b1ee4a75ab17c5afc154228fa8f8874c977bf8e775fe6c9e398a67a272dc67da1c3ac6188f4476906221663a624d0f898704a9ef96d7f7bc780df18e7ba3d40fccd7510f6bf005efab7374372fed7d700f9eb0bbf364ad431b050c85ce89a2c912123383fa8e7fb601fc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1576c8b711b9cdd7ecf561f96fdb741b98ab6fc316ec850f3425a67ca240064362667bd7e1bad9f742f8dca973ea8180f6d84eea65b3eed4faa0121b7fb5ac84540311743ec6884bddf72a2b723161a9bc32db1c5c9c07312c6f19ca87459fc7a97d3aba788fc30b4c865dede460258400ae14171ea570a54;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18d4f3897c42235e5ee3946c3c2e254a19c38089612216c5f0a614372f2b89d2d530af91bea5fc7dec46aba44ec957539e77c91293be42b5efa4d3841ea104acd42221aff5f91a43db30de6bba3717018e2a647417c34780a8c8336c6b9dfa1e45c9567249352af8b972a3812d75d1c996cf194f833e21ab5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfe6f49b1a8bec639b2ceb3e5aade1dd505ac81c6be1b7f9d6e251c05f6df93190fd2113e327cbbda6b1fc8cce7bc6aff48838ab556fd080f0b018ec538a2cada869e2d3501eb0b4c54f0ee93f2038a0cb90d097e1d62f78bf234e369786018bfc5b6e25ecde4b7e6b536c4738adec426a35ca66ccd9e27fd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5d88f1e68049e407da0a0571d80bdb0ca7f6f2a1759b425a4cd5f527c81ddfe0721634ab912fb932b554f666c34aea8bc749193feda9e05d748f26bdc9a79082987523979a88b4f61671b15ab2dd249bf8e9dd6d937a9d25aeb292276b3f12d2498736e1d9ef6e9bf1ece34eed82647106b9bda96476bfa5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ee0124b6db031d6d8e46f7a8bbb74a732d7cce10480437d337d7af023a6e2439321cf6d9fb8b69d8973aefa15e6afa353afe736c160add7015fc1fee6cfe406910c79906e68a6654e78e09fd0beeeb8d932c0c60562844084169ce6460b8776750bc056f5166465210f8013d824d07cb4f8da78daa9191b1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h64a143350739d2344cb387fe322e29f9d637532e571c9b88415fbc86789a69e2923b54bef4b450d92934fcd16827af266402bddd811b51d48e4a7d09b78689da38ade8ea61cd1ba6dc7ee295dbf708a90a832f3754d9927ebad5163ac98571ea638e178a92d8bbd63b5bc094957223e29c1d15b3ea02fee;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1edd50b7155a8713f3db0a0f8fee29b5ecb30d752f0d9a70299bc999375c2286960231dc199ed76efb47b94f669c6d19248be940a2c30fbf774998e91cfa2f90a22be0fa341545c85cb2b344cf78f28e87b3ecb46578ef62b392de5bf94658f395a73e5207e876fbbfdec024c9a25a909cf07c63e26d316e9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9df807492dfb227b77855219f4e39a0e58dd563cee9838116dda9c5ce91f755d92e1795286ea2dec9584a63ff1fbba9d9eb3d1c6d83976ce185d5ec6659fd8c4c65faa384cea2516f4f228dc6a364559d92c9de10d37affa41ba82af3ab96fbf9adf174ec6e8762e761584b50db16f5003c83f81103f42b8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e7b3dfa128dfb0dedbcf056636307d6d8416616bc6053e5d41dd8da9100dd9fed8810129a1104438521e137768fbd71a43c96fc8c46bf7652f0b6430c52b6c3621bf371e5f74f50ac72acf19902b82c1893ea4e1d895c08f964302718d0f2ce4dc4c792e167cdc4e087c21cd08ba42bc9cb1c93e86aaa95a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d522fbf378ef1bfbb0ebb042e8bd3b8fd6f5fe3b834b06cd5f2aebe4978fc9178041ae6feede1a4efedce3b40e2f65f603d63728d9afba103f2ccc3270de5e8b1024311b015fc33b75f6073fef58e83e6a56ddde6064d2e110c43a8ebcc07340955455dee4d21eba6e85c698f4dc0f74db57c8cd04b5dfb4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h149e974c36aeef6c7b272d244dddcea09b893c0046c71c2b668ac32199503d344cb94cbaf9f38c0bd4d5328dea86f0588e29097e4a2c41e342a7a8a16df4e344beacf0755129c25668ece096e745e6d76e0d42dcced899e2b46967a53292496a1a0cacb9626cf633080eaa384137646cd9ab79132a8f1c822;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e57a290c25b2a0160bb61777706e1811bd4055b02d994afcd58c0da67ede73612af7643da082b7a18aa134c85a1d4cfeb5b579d5db749672b1b926acc2677882de34dbf0b8fe4b3ed0dab7f0758e22fb5c8ccc6acf33f9794793bdb75938b3eaaa79c61b554645dc38de202598e7cde459cdfadc9320ba87;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2e3149567f66ad38d1902fc67c366d0ecec0fbe413978f06017d5e1ea29d957a117a91a5b054e9239bb8252afe8b8b491b30979ec40dd30a81b2d0dd6ba5504180c6c5dc454c763f5cae32738b676aa6b474fd3e9053cac89c641fa50cdc90fda58ccae2a67e2b136f32829a51f468eeb99348f111fe15a2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h172cccce4935824f195942237f953d78e50e6bd3817a6f82fa3d7512c75792219a2128c0f09352f791757e605509c64e25c6424003a0b01cf0c2c094bc5e60b0a4d4413abdcd4f174c8183c2c530896f5438b61b465a6714a9dde7d5f721669554fce5de300a960d2181c4d2728ca63d08977e26861b21672;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h70156970b2f1cae965318c88519ef4c00727e70dfe66c5cb1920fa7771eb8af1a51b10bb930cc5eaf7026a00c8830a82604db78347e4278a3bf276d74fa09c884674ce3e74e84ca98e92b2c50f815d315579ae893ef15a5814cee022252aa1752808b611a892c941bb04f8c2409518730f19341f2d0d590e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a0d4b46b3a0efcab51699f1f717c95e2b1c6ed7d930daaa308b31ad6272c73d5e3b5f95aabac4ce68fbb3b063620751f4e7705796f24ebd5e9464cc3684b9a6796f8fdcbeaa968e3c030b5b37e5ed3474e4cbb483cfc87d8db2d05dac40e3a4ab2de4fbbe16e110cb62017f33a7c655727285414a1911c7e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h550ecbadd79a699dbdab8d4e9a73ec9d260b0709975e311b58fcaf8df24550c5494ca6000fb2931859164a797051129523d9de5dab65bc40bcdb9756bcbaf863bb61561c7a1cd3ea44f3d1e753a88e31b023528dde680dd74b847f9da312dd90cc28575d0854ca1094c5a7ce450cbaa80ca6b2124e966115;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbf0d983d9aec9d164b05d905f69cfda5b1865bf4b7475e670ddd0806a2273fd7a5a2eec6a2ff1618a6523c4515d536c6bba4db6dce1ba24dacd47a1b638bd07b6ae806de6c10eb5bdfb2c48960ced3cdd1a2b1c4f46ce69e9ced5caf373d73127694eb68ffaad3ee59eaa713b6d02a0e7a72b46ec697616a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13bdbf47cfb52362b730d0be9d04f021343e1f8a61a35c46a9f71588b3b5b52554a3ccde0dfcc6dc1fc7f7795c74e922a72be5132d406b925f4e02af57d10f43087acbfd812498405ac2e4b4829b2fa857b2b30a517575ed7f4d46e2ba1c9d08f2c1ce25adbc74ba5e5f7017ddb4dee86719c98eb2c8c6755;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcd76b8ad8144fee9eeeefc14eb17743729c464b3cffca6bb2635ab803744538cf0f36d9b31c1c5be694fe808d9ceb9dfd3ee0c031927b863fbdf08604ee0ebded5bccc5c5660a39754379965aaa9baf33ba9ff887ab763a932a256f5e8e072f6108806e2488ae0f6d06f7c12a25d4ca241d5b9a769ed5b4c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h97c405ddbc2c0481259ce4b2325993acebfa13fa4777f4ecdf0f81b2d076a31fc82de79a5348aae5f3dfb4e1515af945225b1e0d5ad40a80e834e94d4be68558996004fe09d0aac317725618c0317a91a8af8145e8d27ec927dae362c238f728be533547c87aecbf4c2df9a04a5c8001a5c3649b4d4ec38d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15de4f590d7f71a87dfcdc099ef66411c74d60e59b48152175976059765a28b8e7cb9bfbcc1552cc28f29bd15513982917261f1b048c7f8ab0252475293572e3899f8296ae774defba55d2552ebf071c065beef6a39af54d2deae730e6f388d83df50815317c2748728a810180b38431e47000f3c8cb52fe3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h320b3251f599c3e01e78771e6f0cefc0e30150b0950e1e51167406fcdb122560fcba71f34f559fa5fd10ca2bb4f224208052f71de08d8e12a8a097170651b5eca68c2d1cfd071ba561eca68e527fb1bfe5d47243d37c031e588a16b8f720db7af9edab16e53ce27307683376658575a5e90574515cb497e7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17cbcc0734d04288a5df1f9c71f3b4c41c659b663b88ba193c879aef3d3bfc164094d0319639a76569ed2c62c21920fc17c05734cb4e3b68209f872e8c631e02be846e314c232c9318d888fdc28c8e5c49627992f1a54566cb45923e1a952afd8551038ef655b84fb6836f51f39f626603c63da058998b256;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ba4de1da4e831353263f16b2ece848901cb2e37cba2f6468d7a3e31a0ea3c75953d6f1d7296afa3f372b233ab90e110bff708493b1281ee3d6d766db089289fe834152edfca7760f1c27abda63097f2431f5fc02ec2bb02ee42ba18aa48e8a0e4fc1131dbae93c5fc06042ea03536992317eca6f3662f5b8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h105665e2e8f8058c3b9829eb506e6c054ecc7b1de86112b4420ba8fbe1a7f0ff736f243fef60819fb627503efa10ce2b25cf7e35635f4b6872d63f725910288998c627e64eeff7ed77ed0cafeece408638305d0f18f1747e97e6d591b3cf70c825bedb89e37c274b219ed66fb1affcaf405c3b883033b07a7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11bdaf06e8dd73133978224ed6be6fda0cb9920aca3fea247c063727afce30076456ec6e12cf962a4fa73602c07a5d4b558c9f7707fc6958d8b7f4e89469a938600ceff168936e48a6bb69ce474c49a3a7a3731511b1877d252a3de51035e08a24f06fc2c81042a0ae4e62a8664c1923f2e23c6e83301910;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a635060475b3a310cfef518f9e14ccb0ccfe43cea9e8e844dcd123947306c9ce2d1fe77f4e9a543563f1c0e806b993af4a62b9b0c29d480609b2e76ea06e908d3025911f1572a0fe1aa740d13841fc876bc76ec5efe7a24918adc3bf9e02b9a6f5c3c7b08bbe52749a6af19aabf54486be2d1e58f2c7f0c1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8710a3d3a6cfc4167b8775bfca8d24a7dd26e0bf525c5d92a3bebd87b086fcfc46a74393e72504a29a5b17a53a5b653d5c70fc0c52e9881f68e8c1084a5807a1a3094a64a0eea54bbea25234805dbdfc98254fa0a4f6aa7f182bd2b66a251f9e9d2e13506ffddf55e2a091807f4ec4c7da5eaeb320cb2b25;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf20ca879bf0d9843462169a3c1def27d4ec45a57d97f7de1b3e6abbd5b8985b4162e914f8f6d1b4584e0f319f1306b3fd0f661c8fddc33570c40d34e07333ab433ed23a2c84a9642b3c20bea001df6ea8c58c901f88a429d73b5e9c96ab235c79a09d24a04b1933d36bae2e1ef61b57284ca7857649a14da;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5e19fd675bd6db88792bbb302c46e59a74d9fd081928d2239b1ae469382de97eeb9a6067527a91b4cd126ba574c4cad3d7af0e22f3c9ff18bd33e60bc165bac4eed1ec0fc98f341f5587faf5d4339ae22b4cde78a9363b1612754a7269582b429dc199a4212dc4d104fb9c91be4c7b8c6e034c08417d80de;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d11e72b01ddd15460f74b469a99f759345720a13c0c02155b15b258379dccb53eab2c7cdae047db6824857bc131a9250bbe560331900cd684feda1cb0582b7b63a64b491b6b96cb49b08e4ef9c67254bb1254f5360c620b2e0573a2b075e31accb8ca20bcee08e87b7d9e9208c90decaf4458c8e6efbbbdc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h142326af76e245abbbc4690c77dd6e75bcbc3c96b24b4b9266c92e7f222fc9af8c336dd865870e58ac859c60d60a8bc64bdf5f90110774da01f4c2e834f24b6ed6b2dbbfa90e8b3264de1cb6083d33819e8a2e13865627cc2b0744481007afc04b37129790593b1f8ceb62c496c0101b4fb228ae31cb2b399;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13ed9125a7d104b55d545b705dac986b9dcf01804474ec504422b465b66a1e0f58ac23c51c461ffb44de02fca72d673d25c04be78c02a7603d5ca3f788ede24cedbea69b16a554eb49a9bf4d6d3a0d7cc5f97425c18dfcacbee2b050e9322e0c9025871b1d586a52ad4a2f328995b45ed5ea779c2c9285382;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h117e62e004fbfa2eb234b2ead328c5f8cf71b896bec9d3083f1efea25a6f51d3be549891dcf3f25cbef295eb676013306d2bf5d984512619c6de7630b5cb7a307333dfccd34ac6c66b1e45f3863666bd06f3475dcf3311e6c4eaca57167fc20f6d9db4727d154d3d6892def76a846d929510177485ba5ef9e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b291181e16ae6bd4cd620af3412a1617ce19ad57a164120a94e071bc92592f4032202fd09c801dc4e71e8d57e9be93d1eceb984be6a7dfa8a40bcf7e1c1d53537271f56328f9a67737681a18b2694fd63fa04351452765cd38928b0d72303e4e8dccf7053847c0615513cca176d25d24c6fb69ba28fe2eab;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h578c0eea61b7f343f8c46e9d9db1b5d10e94922d2ed07156528e756bd9f866a5dd2a8d82e7c329446753f2bc01908063c8aef74310bd39216dff964aaf381e7e9d2b0f03168017ec74e8bd09d7c61aad3f81fe41e932fa31680961d346aefe09eb944140489fe398c02dcfe4d8684f22d1c5105c00d7e1a1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6a963947e9d99cf8a508a10f35358963ad5d0869c87ece67b9261e7d50765cbb9114acfc6fbc9a3eea4e956792fdf30ea356a51b1d3c48977dd21b4dbe5b2db459a365f317f37088e6bcf65de06ffa110b0a0aa7b6af33c1f79633cec4b0c314cc4de837a8a68fd16784d4d717373486b7cbd0854844c646;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h167b4d2aec3090142695311d010c2927cce177a6626a745ded5bca76a9d3522c41aba1bbb3cc5e9f0c2af8ba9e9ad202728d2767c35ec3eaa36b066884c94341dc67f4039120dd08b6defe0498671371b9676b6433055a8e7bf62a73485615de51e3531eb116e745208009e3e21777b3ce2000b17a3062814;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb299ed8faa28b407a0015297e1dff730bd72f0db98a8502eded751c62442654af7ca36d56b77d62cc6cf33e0fd9d2f6a8cdcc63c542f8dab9c8be72793d5805e9d109f5b11ad406e0faf087256d2b2a641eaffcfdbc19031e5cb9170e789f2c2e330bb224c35f7192a745b5396e139ef28a4181385ad127;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1995efc34cbca5c4e45e3313aaaba2e9d31d570af2a220ecfcdd65ca5bcbb84979581a9350e37e2f03686ec5a0d0f5d817f2d0a72a485b2880d8303838a686f6eeace62b3684fd799be96849f71ce0c239b338f4c307c6fa1976fdf62a5cbf3d68eca72cd49ab823da16a4e36f4b3a17804403eed97eccd33;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd912eb6003237e29ab8ebac8bdcf4d5838e6f33efc458dca190ea169969953ce0411548065b6361165936c396778f81df7eff7c9c706ae15dfc3eceee1a0ce5cc6bcb382dac4e191ab8e85f3bafee09a77877fcbf9343ac3670ad07e70bf29419c5d5f6f968310b6538444347cb1bc0567a150b31352e074;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3ee4bd3decf2c5b0aba1259e3928fd31c78a106acc94cb7b39f9b3b914f2cdf5c6e7cf4c0d71a2c7a8bbdb08b206b9cf231c0c0bee75f258bc8fefedf2db4905fd386ff7cbeaf94da46305558bed98f77a5e75fb08d19824ddadab4713b26c685d04a9593286cab7df8cee391d2871c4b7dcca7f6389c6be;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf9cc13d80746d9e09c783a428260cbd317aef1a2fa6d35ecdc016f0239da69252514e44c227b1edcacf6a6d020c6b44b1c8e03f3c8c1cab57deae73c8023742fb498200bcce72b984a16f8cc72c3618cd9291d180807e5e0a7ea064d43f60d2642b816a90bd78ddaa7dae59111b182403cba510fd1e0781a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d7069bb1d98ab5c67fb72e10f1a3c0890d327cc49e374ed44ac9a824384445afdc0c4ffec8c1960045ac09ea178d6008289014123bc68f1ac557a53c16039645955ec7bc75792f4c4a25fe79d6ea364e7e4998c430572d36ee8ba94db27cfbc3a58330054a8091791334e63129422d19290c15667bcd4813;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dc6f3eabc7e602983dee824ff0f0afa791b0033c49466291f0f0f6c49cbb139caf12c0d62792dccf526c7d7dcc23641830aafdac06157a8966830a1de99c7659730083cbdc09a698caec6f6e4fa92b596e6a02da6f81b4bd03fcb024ffa527fe2423d926f7b5ebadee7bcb4b69c2cace7203833a13fa79f5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h159bfc9d30ee536092d7859f2197b9e05431bbde4f725dc483896fb09e2a5cf892e85acf993f87eb24e3d04eb5721eb5ee73ec1a0cf296ecbb21d66c9d0fb6f12885d6724abf0cf1aea4f7e7080b40746bbe94ceca8be544f4302fca3783ddfb85e97e3fe211c1324f04ac6054179c3b39fffb8302dfd9d32;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15e2aa0c057a06ba4a3af3131779a58825f3ce1541fdaec7094aba6cbade0c2bf078f4f9063353f0bd153f790fa0989e0704dbf0de94f80ff12fa171bdfc5d5d302a2b017e7d6169ddb46c245dd1f601d294556fd96111cdc05a18039190a8b16a1ca5f71facaab25427370a44722696a6a320f7058894959;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9879fa8118489e741405cb8fcab626eb0c487e9fec04c5a064025eb1206a97bc340b5578ce0d0ac3e1cbb56a0e885c123bbc3f917e736ca4a5c228332a80f5a00f50a386da9aa17ffea7a8bbd2605e99815c16b15aa29ad84bdc7fd961aa76488642ba47255d4648c18baedf7210afe21a4a0cf2896613eb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8da8db35316754b8be5ddd7ac2367540c81d062c5272d5037fa16002ac7db9069ae1a0a65a52d022c8abfc1bbf01576bfa52db5ee0fecf0d87a7e35c3713339e73230ae1d5abb1f75d9acf75b200cd3b77269abc1c7aaa3c19becebb00c473572724a77e512d6529600937291f25c5f7db1690cc4c9669a1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1636a80d1a04ffffdaca248bcde59d79c48af9ae1fe310f6ab9b05d3658d2bb9aa90d27cf924f2ddc7ca4e5de3662da23cd4c80ace0e328dc03a91eb5fb1594bfcf84963ca69fc6254681609642482ee0be274500b4dc5a213eac0a744b59833a8522e7a73598ccb549e8aea20a7a415791d05510f95306c4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3dedfa2465bfa197ad8110967b556db1fef5565d627190c689d2016f5bfb688ca3a7656722cb13e6a2b5485ed2a1cab5fde23e2811bd603bb3e486cc1e0c9a38e2bf0e1281ac42ad4ba199b5002150588a7bd8f53bb063eb716a2cdb93f1a05a414c597142bf39bb539fa0b3bc3c08b6487aceb2158dff5a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1816fc9e312c78c14a72b1501e0b1b240b6c53e5e391c4c9b7bc4a85b205761dc2dc9292f6c6e513cd85057a923016bf653f64083f66f0c71502083963fbe8adfb4f44f50647c07d590466d14f9e9b3cde671398e03ecb60181b45bf9d6da813b00424a07673c9b224994fafcb1b6f2cb0761348dcb2f61d9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4bb4deb134e618802b3d056c1089117c03280382931f9a8f8b4e8f19145ce9ce6935319ffe69f7c01573bd92c3b418928a648a72f02f1586c869d53ddbcb123312f761c6be42cf7127d9fd9673b5129b86453694a2e31b0bcaa662e13cab63e0329561623040928625cbab5caa28a447980fa665065dae50;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a5b51ccc8812050b190505210a2c631899e3a81832ecc18b3e02411eee3c932f13ff430dbdba0849aef1fc14c05305875d3a51293531522ada5ecb2c99179b733dfde9356b266c37394df4051eb78c351e0ed551c4139c4fc7cd502d46075a43be346a26d9d03654ab5ab50dc93cd7e0b971ea3b80f1e0fe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haa8349823a6513280db5a876808c2bd25bf5ab9665abad9ba64713bbdf44c2f479f29a227f49c839a13b782d7bcac1eb544966d796a9095973e72ccf76661a8baea30c6b2b69f08603ac87012c513a5ae20b39dfc69869c552eb93509eaae86d6dc13220018be424c553aa9b9eb0fbff94af378a1f3c4ec6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfd788f81b7494ce240143c67d6702800cfc5deadf5acb61495d55d20785463650c2ccaeba945992035000a2900b600895b2d70d0e9a6d119a795e4d7321660f5006947d04b7921076be16de42d9fab455db4c4dfa1f2297566d63f8e6b24056bfbb5060b369e8f241ce8c48dc075f81fd94ad24516039f57;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4a032d2e422546181e11d16f1b14e81b5dd4565b155ec6149c9fc3feb31140253210e35afece6802fab05bb0461623a85b18fe6eb729bd60581b0966cb02834585ae31a34328890dc017200006b250a06d31cc26c287388e722d6f0ef8143aad8395ef567d1aaff422b4c17d00a216c035e5fac1cf02ec06;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c62dcb87b2a352638bb8d409d1cb5882923c6aa4ec790184781ac46aa7318d80db921679fecbf1dd4c900f363cd1c3918d2ba602e165bdc25d8559b9cb985d3eb7c70c1622028ced412b2654369a8395ccb262fd4a84c5590a3a6246e660bbb931b37ccd6514842addd0735a03d6517d04865e6a5c012396;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18f459c795c69ef5459148d050ab7c8b10256f3ba1047acad350dce2eb6504d1953e0ca4a43a36a24f942902c68d512bc3610c5dc6bedab212f3211a2f08d8fcdab5ad1c7e8d2978a593c3ce6770eff0824e46332f8deb76b349c638d19e87ddc87901d8a6b6f6e4eb903dc97132ef66d676433a73bb1bfc6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a2aae9a5ccc8c62b7f0388af81bc86f322e2638e84ed6872e473755f674a82916337b0b5a010f1cc3dac50f12b1a8953b0fcb182f2b612cbe35258e41d67c31dff0edf6f127d778a2aee482b05c21f2460526224d6a60dcadf5af0259f87e5afaef7349dafce342fb5a94ae6cc20199fec2e99936bddd4b1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cd0c8c00f0bf6f344ae2f5273c5177dbf184d6ad71b94e9b955ceeed5b19ca675bb5c9076669a1198f7b227ddc55c26e7f7f6d77e6d410c4cddc4b5cf929a61633135bdd2942ad6077c14ca2daec9258701f4eec22fc9a05bdb766ab609e23f1fd883660d1eb0513603fc0d86e60d0ed2e093e415bacc97e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h455fc79a47e02af034bb4c41a08f4fca935cd51a3a6c23fab1c7a1fb88233d4082f0ae601e30c116c8385982e88e4aef2b164d5835d23e558cad2c0752d7948e5a12cda7a002f0f3901f8b11948882aac1609a7a579ebd133a3778bb4ac12985cb112f6b9b6ad6b65aebe99ceec51bcc9543f9ff14b84fc1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h56532c4a875c199758dde7c5c8e9da8c21a0acaeac2da315bba42f20649828b91359c09c4ae64dfcb072ccbf81074d5648416e2c77a79866c836d5ed7c017774edb27cfbefe00a3d8b22d6c1bb324d75cc4885a31dfdf600f8d34dc72bb7e013e6088713a3ce48818748edb0cb75b49585e0619212a8a1e1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf668d69ee3a67300024ef7c8e774b252049de0231a0ec98155e3b09b1a378beab46040e9df3ed1549c9e9ecf93f5d60763fa7d46e43c02f20bb72439b2dec7c5bc1c7efbad09eee21a94320f797d2de66949fcbb38d693f7919d5a6ad924ead98ded19c06b0940c0eebf8554b053125b3ce912fa317cbeb5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19b884c8358d58c195faa5afa4d83484b4f79d057695f195415ec3d7dc65bee3a9f99bf383f20907d3d99d27c2dfc9e0f5f850746f67d69cfd3dffe7da421863ae9a5e1cd7160267348bde7f425570a5ad3c5e249cbb1e1556f26e744337658b7aa85bf210a7763ad43a76909110993698aa7ecec3f5cc3fe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18f972b3911c9f477114bb7ddd76e6f7f2c4d979c7ad82284fb78b05d46c01e575e14bacc435556c029d8b8e8c52e58f741c4572fbced1c9bf853ddba03d4a1173b8c5d2f718b86d72ba358d6b751aa8bc7ab4cb11fdb137ba35785faee4009ba5da4f726914fa08f92ae80ebd3f2d0295bd102d8c4767919;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6f3903775f7830de9cc9715003ca39fc1ab2f99795ce2065ce44608301f7f14cfb0b58b531bbf364ab8c99bd956f856d307dd61179d71dd61a88a586d4b90762a52bd7eef4b0b5e133762081137cca78438f0aa442f9f419e408bd88c5207df9d507d1c796b20dd29b098d80d512ad406970a741c450ae8a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h70857073631806ed2a10b0807d460f4b0abdf69d658af3f057d9341d9b2252b5aaf600319bb078be6ee5f2f80554b0f88eb3c21fcc0e1adcb1837adf60df96799cbef723a97a8cb179ee4a60d2052abf6479481c2ce8929a3da9c2feb8f259b9ea4c2ee46fb0916be4059b329b5a604083b8f90c0ff9a6b8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14801719de9210c96ca241a51c20f38f049ebba488e35904f8a3b5cd23a679a0fe5c830b2aa126b0fe9371004129aa84f182c05f78c2aa405968aa8c76c0551f69c888653a2086fb92fc6a57090ebd7ce21b19b7d9fc96905eb2930a244f81f37873c4ec1a0d59efa365fcf773b8f7b829843bbfdff53d3b2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a5b0bd5d54ba3d5bade8ea25b42f38b0ea1e67b59d2a40e2318fc089a6f699aec178ab3ebcfc2f3bfa3ca325327c4e5eb9ea7d7d7b4bfaecffacc174fbae3cd0b734caca8547bb87bc2713ea8072ca660b241ebb149c73ab4d0f42d6aa1789e27010a09d88b3297f369a2ff7e765619fb8bcece3aa7ba52e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hec994d0f68a7d01b0669f3e5a8cbcb2fbf21bc67a8223970b5b6f5825999a27cfda67f208e21cc949825207bf31cea847a3ed99489c8b3df6ba316fbf0fec08b0968999ba6fc7f7e0808aef659dfcb279337302a256e576864c081ca6506e3eabf8fe178d593b5890f4a4f11d6d75a9290ffd4a7b351c816;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12d19e7fb3eca14f83cdbc853c77b1305fab053b2ac510378862576b0da6d43deae43b7cad88eac99399a26c7e2d8343ed891335d90963461e6c357d0e4f673554d2a40abc87bfdde4ea4c44d081c8bbcfb019ccbf50877d048911554fefbb4730817dea2333a8921d2468dd5067b56856b3517907cab0e8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10296dca3e8969bdf3190c1c0d43e516f4d05a1b1e4f621e33fc4539b4174fc8c08aed234adac9030b3d3d19b49254a170d21bbe23c6eb41f8865d878e49b7bfc9d5ae4c03ef589a7c670f9d0d8dd8ca4965b1dde357b95f2511b64ee55c4c2bb78765ba9ebfee1e2725b95ac3dc0cfa87195cc85af22a76f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h125648eb7ab53c25ba8cd9df54b5d49cc468baf9e6c9dc6a562fe654f3fc25593e780111cb5f44fdd5c5a39b648fa9d55e30d3ecc166a111655aeb0b4c9feadd0a0f675258d70e7884d69eb6ac96b0b5fe4b0d47fbfdc7be5fac031433adae42aa2dfba49e24127df4c80296cfd23abc2ec5a7aa6f6c6779d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hedb451e90d6b25f62489dea6e5665a9b363112c545b623ee4b4b11415d895eb6b9fc00ce091bbab24f55b77f95ae78ac8de4e85a8a599dee17d54d2a24d645a27a2d7d8cd5baf0a097b6c353545b25d53ad0604e7d730198319afa0dcf6f658421e952830dbd54c623149a7718ea721c8fb32901184b8a6f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha12ad122b052c5c8084b48f0cec0d7ccab8d6ff14f9d3b853a19ba9d8720832619c60bc01284e0eeaffd8640dd8adced6a8243315d704021706d063640532c959c5eaef862ebe61ff9bb05a6faef2c5a920d19831d410c06ada5de15dbc3bc724812d78752722de43423767bfc1914833cefe4493d4802b7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h790e452f1e06ef8bd755c30d0719bf25605772ef94f6181153777598b07a7fd71cd33fd390863733ecd7a7d13cebfbda036d7d131a33531e0db0d72d8abcc30fc65c36f4fc0467b89c9910e822e4def0873735b9a53851b3aae868034e9046e855d332b50f570af40ed93f8534377d35573cd0fe85842f4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11bd1f94f1f9f470b8727355f2c9c582ad9adcd87c7ce88b80651dac616c9bda90459a0f87d4b8531d5fe29fcbc3ce34a1c72209eb1aa4b59710a9bef6045a3c1a855a6362c3855e9188919dd620938b0fda268086e821c76fd727ae8f17b44868132c8e32344c18df72b6f1206b91e6f9d0634783c5a9da4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f273c5312619471cc8516b75b6b02a94fc8ae325b1093b67e49d306ca619e0677c7bf172891efe031f4c75715c1e1151dacf48fe12718491392dd4dd47894565fef9c39ff5f6f5b8c809163543802b11b20c64a89e0e8f9e9985865eda218435210da3dfaa08c40c07362ffb7d98c9f55ea0a31cc23db4a9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4bb2c3e5de6196cac7673adff33e8020c2aecadab73cf882e17e2a8816aaf2f9259645b3696b9c7802b2996273090ca88788f502359b6ddfd58c99c19dda9036179d2c71585f480d09577745727ec85a8b4913497813aeace646ca69dfee14ccdde837922b6c9eb76c1cd0dfe60b47a940a40ca816d7adcd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d45245f75e7e9716ea0a074fabd0f93f7f4420c761cad62e8718dd2e6d1769ccac142e705c452a62305a04e1a13876b92b87ef845651f05c402d68859c82a2b72843b9926bce6b29efeec7b579e06720e374655b621bfe89f0d0bbb6d5ca344259e46fae08d2436f7b2fa5311f2b9cd399456ad4c6133ee8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1355843d7046db1243ac434e70d1705ef7c3760471be10b5be4468d4ec74ad249bd3789864f366e48ece1536ad836cd567897686fd551029852907b65181f6e59e8483b517383fbde5f4e33d1667705a962624a4c454061aef0108d816261fc2f1175eaf3b56d5398cbf2f526ca5a88aa77bdca689bae879d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14bd530326e31754aae9c226404e1d245f681270630af113a5deb8d95a85b09f2e8b4aa856722944585e8607ed89cc011b1e6eb5fefaa3e91ea6d518867d12d895d0f75304084071c7ff46367dba97c9b827002ac8624bf5ab2a6507ccca4b032f2d2d43749f3ed3449f95de98f2adab991880e9460e8aa7f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19d2adc39b8063e3ee8fda4e143453e2e0033d6a10b9c7c023ebbfb73fc3db32dc57dac8b71c9ebc2c3cd443d939ecb2b9d2dc59eeb40a4fcd834289c819c32cbc5b93a8010b1f696646fe3c6440f04f8664e7c827b7c860f1dc7ca8fc3d15ce768de3d3c966b1eab4c997f3fac27a9aa8afb5e6d3613de08;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16caf540b6bff450375804dfd5577562ed20b263c7d0ba3fcfbefc0dc71287ab5dbd7a4723b0bb66324c19746f7443a45e2a18bd3c3c422712f994186731ef102f1b40f19e2af683bb9f4323b23240539ca87431344ed11937864b0d29c5c4d25d98a07fb8490fe2f3e097d5d2c85ca44642617a0444e3cb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1293494b9fe73b10eb08e89b687bd34372a7f4be6b26237fbf9030e19a90d5f1adbea9cfdf86752fcd115347c45d6d33399de8bb2097d4e0dd08cd45383cf23bb6bf1af5654c8cb1270e37e023ff98a69f9d08e8da979b576fc77a7736a34aab8d417ca16588d1235daf726ecf46edeac3261556f5c3d1afa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6d56efb9abf3dfef09a3181af8e2fae373f382e19f2d3b492b6b2ef7ec918722441dc874b0da9c190aeb6f028531a1168beae7d4b5da58ecdd1dd9109efa4a6009702293f0a020eb9dee627398b9619de7b1b518d4296f122849e3f75bb70374c095a625f03d3c27aed22677852cfb2de0f7995f13209da9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h44b40f95e0bba44d39c791b791e62aaed2a7307b6c61a7806ce3472afec06b8baf2255bb7b1c7db674639f211315ee08df0267cf7bbc69d17e6e70e6ba9d30d50f2c87a473ba5e47840cd789e791df3ba25cc0ebd03be7df808b25069011d83b12852394053a82ef756a078f88d66790c5e73f1a4a76da5c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12987c64220b49c0f3e700b5471210b847c05e7d1bcbdebc5dba7f61c5166f0bf2e7f9289c5df427af4f3f59bfe9df0542422d5a9be01cfa4a020bcb5c0903e446c81ac14becdfc3864a20b7a93f9cc1eae540df931913a830e2047a74cbd1c6e85d9dd083aecd919fe6c5f50fc521c50d71bbefc4089978b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd726d50b40f795a1bc51c4896ebdb7e9a362a6af5cdf87f79e69112a42823957d1f6d886cd2eb787cf78ab22c067814cab4be404f394aee3db69ce7651b28fb2863c2d26d4a7d95d824b67ebd808eb6b191a1107bfacd4877c736942a965343d6cd50b1c37af2ec329e28c881dbc460c02fa2749cd240d41;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1191ddadf4578cd73424009900152d6dd5c9a3bcc6b4626ae194a475f57f454cfdd0ed24fb1a740eedac395c20353dd6c6f4c360a85675ef38e14ef232a4e5e4795eaf0678b4ee15f8c4123320df623ae485dbad9fb36207b0e2185009e7dae83f68b88017a37d46eedc7918e675cab5216c3f410af79486;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haf3b74107122cea119a6d17b223668943acc38e80577bfa08a8445db5d66a1f120eba613759618d16890cd814cc387d8dc42f71459d79f5c30102eadf6aa7dc2a5ff93a974699ba105b60e59060d71b55cdd9fb70a3d399b25d00e7977e36f1d849781ca029aae68f24be3af994296944a7a4d717b3d47a8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbba0f395e609a78c24efeffbc542131b8741fbe002eca0b9fa5d5141f570c2eec484f8d0dceae6225eb102f232c9406add2512556ea5d0cb2c28e1325a00274e0ed30ec31594170f7b770abc8123317d7eb41d147076984958b49a93822931ebf2f197b9a8f9e97a9c0b2f7556a26a6a24ead1396fa32235;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h25eaa4053646b19ff5d6809504a3a32f78b62062de00968f9ce0245b53088d122b7823ba3bd08ddc83712ad36e39788fa88df90613e89ee8c19fa8d65694a740e63de5f56788bfc2d677acdb46372b53bc7a01d6a18c04f8bd16d93de3ec7da5a7ed8073e847a6e30368e3a8d54f6c3a1dcc39fff6fef5a1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b242e9e0fbd16e9e99b5805b7655ba2fef87be71a98233d5613b9140bc82e7666e7df2f3e6a22153ce8d6b99a56986598f3e76aea27f2619fe67327acc868b522fd361150b1ea6bf99551261a31aaa917112165f2673fcc4b07017dfb2066d730e8ac3d1345cc6fe90b3aa61306df1c111a1ad190c94c020;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3252057539ca2a617dd1666236c1cdd3ab3a5fb2f8744e8dc00ae337dea8e64e151a2bee2c0ea09b98c8aa61542f2b9913f6627a5c5c2e1278796f198c1e1daadb22bd34fbde35eae0d83c17aa202dc3117e2f6ecab3a35853e869cd619d26025d638ee19a941c0a31c7ef57433f9c034545b818d5aea941;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h61f6bb812e2bfd707b7777e6fc1afb3987031b346dceacd59144776bd27cd2110f5769840334b4df544fc730cda6e583463da6c179f0b68348caf7c764093e0453a6eef638835d934dec3881bf606d6c888574f5b0d90af991e77742ce646043c26a02cb5873cfd838ce9c123b66cc4e49eef96151d20be9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c4ffd7a9afc5ba6d008d28a252a88c5217ca4c94c64f080589f1c2393bc0d818ca1624e04f425c4be93d8956df0ecd4cc9f58da169dc4b377a07a989fd2018d21b09f21cef6276a2c4dae400f82053d5251eda0e34ffd18d93fb21a22f4c8fad8e54b1ab117d860b66cff3d31ff87c756c1cd8dc0df8ba03;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b10c3a15a1e373d187a2f6a3c2255bdc3e3e053faebf2d420bcb021694ef3bf42e9ed11eac9fd82166c6405fabade0e0d1ecf5b70ba51883902f55f7e739b4b3734af778bd25de7575bb6b5ec40cb6d4f03ecb1088a86ae770dfbc49404d9e0892f2be4f4a4bfd6d7ee03f3f982ad60a1b848f4c083f793c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f7662b9c03571f82fe327e9ee865f2ebffa4a7e5dc92250233de2bda8a8af8dbd664e1aae6387e89d2695b039980716d914b4d2a07d857e095bf77fc271038f430043c4615394cc8ce8775a6fc6bf1f0c85fc5d4017b3b3b2dd80e87174944f22b5f5fe770f9d417ec03c17cc44c5981b7247c719585185e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dd11348d2922e1fb1239a6d13b134efdfa127ddbbdc2e9a1e4d35ccc179f1c2368f21765e6986a859cb42bb8fbd6d09975de07cfcd6f11230821d67e537c36374b3cd3d479197f892ccc25ff67bc1ff169ff479d314fc15c993f78ea29a327c5c4a926000ffdf34bc6c93b42059ea884a0cd8d7abb438ad0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h73b8bfff13036a558434f3f398db0934b61a6199dd967bea25893b6ae40cbcfd8ed3fe576e8af3dcb642018cdca63b2a8e088c968bba172d07ef873016b016c8f269f355e92c6f4b41b48702df9b30d0ebfe1965cb5cb5dede1a7d7f3eb847624f929d994206c936d5fbf0ed583cdf5ff2e294781667f554;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16c14c224fdf2b408cf677fdb97eae5bd1cbbc73f4756446a4d77257c929271bf83fbfb592ce61181ab3b38e6b059f7a1223555e18e4880912ac572280d576dacdcc6a01e166efe61daab03273bbdd19c48137e64f7774a062189747bdefd1884bd9f458f8774c0625437726faff7d6c9331001f56766d8ae;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10361b7b0fd880fd1b0555925edefbcfe2e759db5352f032fdb95376e3ebce189ba66d35756f63c9da4f57675d50ed7650ee3c516c64f484d19b0e6dbd08dd65a6adc46e788f2e63f927f1594efa980c7da488eca6a1f901c330ec3954a172508d63a98407ff262d375e1dead013b21ac811f93338f9ac070;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c30ff523309ab448af12b34fa505e17f89c7b6e0163c94bd9f31f6402f938c566daa3e437762bf9e48f832e1c65e30aaca19c516a2347817a41e58c2794ed72472ec594f43fbe244feabb1896812f3502ae5789f8d87516bd46177af511f6df9d4436c532f266a9e286c6cd3936779880025fa6f9f413745;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haf3f64c01eb54bfa903a622450257efa53578f8d2b1781dc7c9714e4eed9a4964c5efa132fd6ae703fe7b657017d42a40e48365ac4521923c85e9704031e5c564a2950b6257b39beac5adad0cdf5434c747247faf9e2828c6e0036075383640cb270e449165376d6d23256cafb8e03b649b6acb198b54902;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15106125e5fb5daa7960efd85ff30e867b1cad62f4b3d2597da6910ded57cc26ab2f633e21bcb1cf19ee80ba3576d2291340fdd06288cec056e56e06fa69b655bdf33dbc40f922eb5c71d3c19a3bff06224c554695b67a2edb26c75ab2cf5dcd3031d4d523def02bc568967bb5b39365539b602ea5d934a5e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2f5b599893aeee14f0090ff0590114731bd1bb4c56e8cb7bbccbce93e1a6e042dd9362abd093b5d36c3809a1581a76f3fa04b328720bbea3e7397b61dfd35f8e735b1fcaf1e2dcccd5897f78c1dfb8c7691cbefc8c5c135bc5722221236bb5c4972f2f30012a74b8ad393f7679012e356ed2d96cd628daf0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16cfa627a4cdc789441bebf91490e83060fc23844ab58c2122197f25a556ca5852ee63fba1f026617467d0b856bcfb6b0f7a3ab91ac7393ec52df69fc341ac95ccd79473387ebd7a97d4e41e00ca874f30b8ecfa5c1b8a43727681b8b629444e431a8bc5409994e28eae57ad2208a77ead02965735e559f72;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfffb75e2b5c0d426c844870f80fcd1f293e1e0754efb17d6ad6511035606c5171ca53701a159aa3fb216241ce44d930279713b299d1c23d4ee4e1e534eb26a0780ebfcdf456bafa2cc4250c752f2d16010c2a152da8ba8292ca91f59509d3ded02f93b66e9223d3dd22dd275e1680051b912afcfac152795;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9592b1ba6fa6d7c60a240696feff04cd1f0b7cd0c29944295ecd59f0c7d27999d6edabf72d3b1a388f24f32ba10445c275b93ed2f59c40ecd2efe2cc0fe9092086d95597311d2a9f5bfcf1dc9b9f2c4944bfb17b7c2e61cf4ffb79502ab86b3ae6dd28ae1ca82c83c71da9149bb9cca1053c52aa59de320;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17ce00e90421c1f6b1137d223a33f4e308f0b7d14eedff0b17efcfc45e1d1f35957d87d297afb2a5b422576fbae93e25dbc2101157f62fb3d7a231fb4fda3271d3cfd55682389f05b5b0737534c4e50b5662e5953a7a7cd4b1562696d2f5604893318c9b37f51d64275817df8e289ce66729dc8d1052b5aad;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1330255ba802b9b1a96b0b28fe63f8e4ca85494d1b89cf39fabb1021c137e3b332139cb82406cf738e996ae4612df22307fbca0a0ca0f391ec297df49f9d6e286b79d58602864496b88ca99dd22d79e6987c7644cf79fc9d7cdacb09e5c7d53d0704a3ecd735c4dbb750ee8fc79f530b8a679058570a5d963;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h181303f326965968bfb809dcc4f27357ad500c7770e7fee501d1d5ead472272534deb4e34b0d0d8d30d7c0ccedb277e9c1989ca00775fca8e7f764f37c30ca34e73476c006afc260b396dc969b1fff30614c82855509f1a0d4f57d5091ad83f146115cecaf0da3b3d1dbe512540adc2e7af09f934ded296a3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha9d544e8e9ea0e813aa3c59887992b3e990588961ef723a3dd233f1788dddaf10c60cd5b7f59d99be6e3226219f61804d34bf53e66b6f50127bb4e4cff413a225c2b61fc2a9db91097617370e0fa685a69f28e273ac76e33d17207d8a8f7dcf0bc67220c3a4f3a2b9dce3222d3018f12d341b044f3e1c4d9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f3d861352de58e36e39e8161f2dc1a0c93a1d4a2df1efc4f92376140f43e3d294ccc01b502f30110910f6ade2d81eca4f632f277b2425c94377232a0376dc4be7195827b79075c96bc744311880a45d82a4d77a93038b7c18228dd5cc1e6d3977d328a008ba6fc331948a59601e1458da22d6c3e0f9f5b3b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b35e9be1b60296203c267feacba56e1fc504c87727ed7a2e51351942819984116da3beeb93eeae2c8ef81c9009ed227f6ec1f63255c972f0d41d7530edad99681bd5cb058689f5cb6ef835f68d8586b3900da1e85deced06ece562af6d24d4736c43d2d330be90670c3c8dcb3d199afc70b6a13acc56cd7e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h24e0cee0531c2359817921f3e66b8afa743c280fcc03700cd89648c267fe88a5b9dea62b5bc547b1ad5340209afc095bb844a06fe35cc3876116579cc598026a7417290d9dd84d676dec7d102d0917b25bfe291f2fde587dd7836a8268183f364f254549f9ed9920ed8228db0c1a45f6edb99ad3d26e5dfb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h107d086c1ff8ec736c5fd4759cc3e15ff995ad5a2ef0e4b7be7d492072e23a8e6f1de135370418d560538c2008390c5ea3a8cdb6a6ee59aebcfe0244d9f9d5e16d337a79548089cb32f4b7f7a8964e4ae67572ca0f0572c576f493a093428ca434392d80d40ea982613bb1b8538156b204f5cb3fff35b077b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cd0ce0bb46fe98a578d93a04a18c4710f9dfa3ebe8f72a2d0a0273d9a32346b390aeb3a01f8af475310bab360815c91ed8d29328a22042bc9791b513b3e04621b531694c4d1d2452c7044385ccddcc7c35b2d87df87d28fc4742badd2584ef08ddfa75c4c4cb8936deb77cb55c8becd48db1b7b4a0369f6f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3378fc4c480970068a5c7cc1daee8a1f351d1d8120ef222c82e28fc30e532e811d2c1ef8b5ad386029d405f3f6c8e17cad44c6a09dd00cf1d6117ea012eaae5fc73d49f75a6859863d406c2c8baf8d036281927cd21d1210a6173690f9295892514bae033aa54360f7c0b0e62666a1c311d0a0d8c7949eff;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h189c3cf99b3687a864b9d462286ba5f7e8802e993728018d30221ff9a646fd614f0267ffdcf4a9ea854f2f7e948e0791c0e9da374bc5ef04b464adb8ed4c666bba12e5ca56836ec85f946c6860c52ee520aca294e3897b09e3ceb747ab3edd9bea9c6739cf0c1e06dcda70f98f4baa57910f536db7dd71bb9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcb740a3006674b10a83e283487c49fb09bf4c3077dc68a8f4797e31faf8d5f7e3418ee28e3fcec4ce4b973d3db2630df12cda738f30ca3cbda2c9222819ee233157908f3dd2376845eabd9aed910574824bc3e80310361f2b433b69c93f2697f9afe0d607c0ced457e925a5718a86867366f5baea5d72295;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8669bde790aa1cb67710c9d6d011f8c62a3f7b191cf33fd8060d2910a35f31dc5c28303d7b12f224f20d651ed5c94b77252e32d6765234fdb7b090805fd35d19f8c1c006962817e5049e30bcfb1e8ddf957b0704e128076fa7fd5efd07ca0a71d109290082f124526c53889b0f9c16fe459828f6e7b3acce;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h110e312bfa05c322dd5036b64ba2a0a0c56baf1a9a1a8c2d927180806dc3e188421d3c314e719288ba5500d20458cd98fd56cf805242977be2a91ac962ccc9a0824b682c2166a982c61e1553a170acd80e18c084aee8d2a85ce4f278c3d4dfb048c5b1999959bec52bba3f1a8b10fcf2ae12d5893953ae213;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h151b59b9e6e6c3767e1f2731dd2cb4646eb5b50dddcad2626d1904873b3e2a8b19bf663e41bd819a761c224be8389538b205994b99d887949d4338c8e1d947abe44eb84dfffa4abda03b02a9835af6f6618732ac920aaea253244747472b5dcbc47c3a8a5c58f0cba0d7706da3871d090110e0efca22198c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h63017092872a797c3919a705800cd86cf3dfeceae1dd277e5a6824dacdd970f6938f2c0959ee5694003b3a65f9b30c03cb8974ef6466f91496ce7611e81463662a8c52fa4625caace7eb3fd7ce5d6a497b6623fba91e4ad8e53806c9706f2cb4728d48d5c480e760d283d52e1a685bdd62a72b0df9b41fc1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1beb9a64c29350a698c47fc3d04d3025a52c351d7a641029f86c94f40b35e17a7b71983f2478b9842f6004cca4e6ed82fb21ebd33fbd511b4623c50998d1d4abff89974754769adc561edf5f3f4680f861421e833d1a9d7e9469e03fb372789780526d27619fab57f9d711b9a1dd48f541dbeab939019cdfd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd2d0376ea919b26347af36797ae0ef9a14d40b8c79ad827d2c3d102819499e18183ef8825a0debbda3d6e0bb643b960f8ff6e2fa965789585ebda50344464a430485766364bb546146ea0deb14ed9c611284d268b4df94a5f34aaa71d6bc11a8528172947d8e960c3caa5168335f9dd3d915ca6d8c9eac33;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcce1f9c34463ab821e4de280d35ebe354094944b60cb99f287163f07410c7e75f065b2e9bb47615c62bbf5a9c8b4162458fadaf56f158f4cf7b6609a8993e2b8a0de013b0feca082c98e2fabcffc8dc57f25d8ffa35af0d4a0572b69196ca3e9816868e2f38dde295b40692f7c462c3a39e973c8c03821ac;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e3a0dfdcedb7dc12eaccd7d3716ae60149badbb60c6317bd991e96bf9d956db1f500432ee505a4ea7c87dc1a61ebff45cfdb2fec0dd5e4838f9569e2fc60a3fd2940aec2add8c33c3497f495e3da0f3b53f8a484ea4ac80e11c20e80487c21e2152e649261c24409a1475594b62ca5aca8835824d63a05a0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha108c795ad07e168ced631d3ff9ba7c512f11003f0146d84f3440eb3c2f6c3b089f51b40f4c6ebe1a7dfba74b361b5a4424961f4279d57ec02f9e3c336ce1ca4912b7364858a53306c1afff55b2b1cdd5c715a80d7037f5b28b44946932500d8a2574dce8268570d708b2c78376580bb19b5ac7327a9f318;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12bfb1265c900574147bf8a854418cb0e0a9eff95180609c0a7486282b7af5b69d2ca6c4bd3f94524baa48d7955fba75fd9435344818fe9456b232cf491e7ad827cda21ee9617d06ea473ff08682293e6dceb057eedb92d61a73ceb9cbe33fe181f92a5daa3822028ccf239db0696ee9a353ba8677ee79d45;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb73951cc5457c6f130339a4ecfeb1d78d56e90f7246c8d9189b60dabb5348b88a209276b7a92c594f126ca5888d1e3920843e20e02075c7d5531079c0587536739181ca99954b5949b17f83a1e36e4c3b74f3a86dc7efa444c7355461eddbd1d2b4907f3df28e44a87af6b05e2564271fdc9f3ab5861056;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8f73c184ca30b477715e21e7cecf224d1837d459fa4ea2df0930d0c63e59e55d57b03bc761755643f4497da3acac2ab1311e49afc29cc91ca1b193ed6ab20099cc5ecad69d3c33c1ab3ecf1635eb5f7b656c0354af098cde1cd710ec3b86dd18cba9e714b4cee2856ce15b83fc29fc22d76c23bf7909fe6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h198341b312507d50d04de0695832d25c33a567cc425def18ba37aea9110ad5994320a64241f9bb3b10fe8d369581cf008c612940a3d3d7fa51893c5abb377d760eef6b7b060ea66275eb4f6bd437310cd5f5970c4f8b6f6ed8a03c0cdcda352338e4bac786e3e46456b2c0cf55c171b4e904db5ca16354c60;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11f5340956f2e5146505c7ef0c0e64595b513e2c9f27690527acf8c827247c9007f448b41d8258de5c89aa4177f3db79cc53ea4cb41f48537c40485dab667f0172224156cd4b34e1c363ff0a1665ce31099424a4c7f11e116fad7837ad37d4972a9aeec7b8eace155ad3853d24f47a281b6ad5c4f62cc4ede;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h198cd7e255771348c6bbcd60366195591f6095129c6f84bf2388402e42b8388e3dd9bbd2a9f79a352a176c51139d146b8b4722649d6d0c993b238ecce52dd49378379073da10881dbdf953b78d197f7cd72e20b47ff2ff32985c9617717fc3f9e2bed07fd89a2df6a623aee22183c26181a0c73304ca4bbca;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7a55f45aee7be284edb433e765b136b2efbc47b13eeb14fafeeb36bcb26c2b3861062f3b4308c0a9687b95543643af2a20723b116a62884b7eabd10fecd8ec22f2eb6dfaf19fd984714d60d7cc4d5082df019e67564baaf6674016c4ec77d525d86168408f240b0fc9e790a7cbe449336f5d3f414dcef043;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dc8da247a75e0296bd71b05f7a9eb2244c5f1158a34a6f9a606778eaa225f3619d2bb3e44f2944d421cb3e268431a89d864397ac07eb78cddd723c644c52e488cdfa2966dd6e6d018c3f8759a75deb707b3b9fe6c76713264128458f7512b9589a296ba23933d315e0a8f1bc3cf5cd8612cb832d50573b7a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c184bb87084826f99ecd1cadad31ed183141af561e890850f7466f2829c665315db4ecf47575cd6957d36815a1cdbb7f1f6c8bbf598d8103dd55b4df051cf0507e5fb4b21f560a8cc8319810b98bca0a872dc34d16dde99d954ac0def38241e82562b549a71e30e8b51ba8ce944f8eda0ce42b66b4784463;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19380258f52723055d9fbb85a278542d095372ffe9227300b8548a07fe0a7d02afb8d8c2d095b631f0b36728d40e2a7204c9686e9c9348b41b6b9595533b725c2fdd0305520a0f4e5e5208fd94361595121219ca0c3b80280d43470cfdfe56bb22a9fa5731f37780b6d2df74b0ad5e35d939bda75844429e6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h195d4ce15f036d212a77aba32ebfdeda48b7c6e24e874d2003b508b76acdde4ec0ad000cab593c040477675ae849566259c63faee7981bf9d5c2dbe4b96702ba67bb54a9b1e31a58d00e03698fdb60b85bf0db5afe1af013e97e85dff2c2ea6ae6311bdcd484a0ce8e48f14de0e9f48bde17fb7710319b035;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1076325b933d2bb376a3de7909840fde00ed34b57562ce45ccccdbd393b0f97eb7f59a57907f15e0fa34eccb2f14b2d57d9e9a042feea47928159fd89ae5c19241a1370202781694dc15c6cfb6c071662ab4ac882772237c8228a4ed6e44497f0941fffe6ed7f0cdf61875d62ba5ba30dcea4bbe1457f4239;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he5907843e1178a8b22cde23c4f48f6a50306b699016d24e16a8016b8c341711f0eeebb52169d6fc8ad126245bfa5a27b4f414ba535717ed651abd5421bc29443da74d40dc6ee4edd85f4bf2c543042f670595d552848c7c45e965b685d74e243e03868b2e1fb2d83d0a89d7dd9088866efe5fa2d0f6d1734;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9d9578efc6e8706c2bea5c096d2de534c10beaccef6e121bd01ca53c2baf810a936ab73dd6956cbafb4562f994e5096327b92d683bc1f84a23c7ab388a66cdab8119b737c7cb32dc6d1d0f11e1195943cf1193949adb2929df0841653313bf5a0f2b6f6cc990f95c00cc5b496abbed5aaaf286cbd85a11cf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cb785248311cfc18c8df98335c7eae9e741ecd0720949ca311633c89f37fca56709338df6d59abff148e5ddca5ce9c9ec6316f512ad60ee6e2001f0b00ac69e9547b19abe17022aecb551a1a6886c45de3b6764c014ed840da5fe8774b4e140fc32f986f0cd54863e9eceb2b6899a7795b47fb205ce078bc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hda7c02b343a7d243704598a77c2d465ef0ca0dbe92fe6329b225ba7eff897192cf48952c61ec0d78a47422b75cebf56953ee2bacbd96f1d1df60873cb00761019629ac7d7e5f4446610cb56cb24034f35c016a9f406cebc49549b39b2d9444f70b8179b7b179de243ff9a974a046095ca7c9c1c25c523815;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h131131a8048d2f60ffa2061bb2b505d57babfd74a4a925165db66802c871b98a37d9311d476082a5a00a68d5c883ffa34c0096aa0c2187bab6820c2c4c2b52609690e03c4f725ca0b65f97e9051faf8aad849be31d143e8dea5b69faf83e9d57dbdec70b55b1c3d604f6047885243f8491e0a810709679757;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbdf9ec534cde03b70d88ddd495106353a92d3ef18417be3b6e9c1d4e5bacf776932fa58786418f118862fbf33ddb8b3029c142b5da81ffda8335bf1dc25f6bd5e86904c36612e29b4ae2f2a0090e2fe8ad93980647392a123860609bf41b4e3a6095b4a7c58bfe92f8d924094cf671d0a30cea131cdc8beb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h59a2106938f2b98b9f3aea3291e9e4a7db5fd59f822e9e8a750f15c56b9529f9931bbf38a7ebd0a49cbe31831676144f5736e429f1a22356903a036d6531a3cf9eca20dd1c6693f88473dae45bc9f3ce4085797018367631d65c760a2ef33632e123dad82aa1dc478142f8f88165b0d0f6fec8257c6b3915;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf1bb8458a5c8ace1b9e13c32e36d0cf0914b816d65098d9614aa8b196eea55c4a841ebc273e2aa61f8a1e8fd56563e21e34d554b28b0a912201bb68bba318d47fdc20603f8dc65e725a260af99821f2f0776f8c9c9804b0b7a684571387bfceb440db4c6907e113c62dda3e6a6654f6bda61328fcf5ca861;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h110113bac1649c6f6e0b3c873b37ba187313a8fd58cb4ad3d2f915c609e0bee92bb659c84d6739034137043cf9abce1e3606918af1e9eedc83d608ae10eb25515edaa2283f70eb267991bae7210e4fd36ab0165250335beb5960bed08236a526cf10c8431db4f16f58d0dff9f931bf2bbe88e23f32130c53c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19a20ab1b711d4b74bcac8a3c1231fac3890026b328421df7528b95206316f00545a6c4663b162a3dcb96406d1d924e2de103973404aa8ebd799065dca40d286075225705a28b8c594a21914adb6b686af1be4e605604c3971f35b28d1611e9134cd150b2d3a0424ab166d4a6175aa759a6c8201320c53904;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19029335e30b23b32ae7a0c099e6181677f4d186d55be57eefa3875cf8c1c2edca1c1f5916fabb9ea38ec397a8ac911c9b6b7e60c406c1ce89e0ce1e49eaec17a2b47e0a46340eef808c8037cefcd9f8a2f16c196a5d9f03b29d17e53924325f60acdb4152befa49163400e0bf36aeb909a9be3d44b4b3b96;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb8f5c0969f1d6d7a8e2dae61863bfbc60049a8047a5f96b9aee9ab8eec977511e259fc314e7a08c5f75ab5dfce708ba3ffd7781b58875b354b5c5dd9721a8dbb1dadf0084b82ebec09f2ef2176783ab772b2737882a90d9a07c704eee99debbbde5b7d52211fb64f5ceb0cb7985becb26acd8b5c4ad67fd3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h173d4c004812fb31052285725f9caeb026302552bc69eed2ec1341ab63e17614a3a9df61c6fa8fec6b948d2d07ae142dad04b7dbf3329a73b9c0551e84548da52878254fe78bfef401f7446d1a81856044cc3e960d239f329fc099b47b41d22621d64ca666c15c0c5d7b0b915a76398dc1bcfbeb3845cf6c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb6b8de3e95702dbc70333b55cc46133f23cad907d310ce7e9c8d4dbaabfe10854722e6b2224d1e50aec0fa5cc01e81d73052bb8380daa4ff15021b088fcab64b7d06040049ae9db548016674f2da3ead10f806a789fa85d414899345decebe618ab8c74b0e9c6a4ddc07f7cecde9f7d869648e5284db3def;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h570b6631714c9c2c5ddbd23a012ca5aaa04f4c73e6fcf0871e0d2655808d031f9fde1d09a6aa2d4a41cd28732b3b1e56bceee18eed75887bbedd64c16ff99a2031e0080245162e16a31439306ca743c622d467c9c2daa2782b50fa6b7528a94a86c939dd39cf410514166bf934b516b6f491ed8263f7d043;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12bdd26f4fc9490b0ecc347b853c65b2c6b370f49e32c9c7ce4b98d62d84c39a5afde95e7726490939208472f2b8c3cb19233acf3035dc051d7b339382572bb1e43b3ee31dadb03fbf62b022ce5720db9d8dd1d33b00a7d51e563b3d52ee554cc24552c5111dabe7f040c444480994e9b0a4036b1754db72e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h117bdec7736bc22f7bcf924d335d404aedb4be80a677902731c808cdcf7849656f2aacaead6a61367b499e757f7140b6357383054edcd85e48500c6e2a55b3620a133a216d4ca736850d6a82926de302e969f48397e7a266ab7edc9aa223d7f2ecd6c26badf861d53e37d2a63840b00dc76a21087c4d1f302;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h593aaa090cc2bc3a4eaf6e5038f587c6f81f95514dab4f617de14a5b41291a9aa208d382b66a2ced8603f5a1cecc0c05c15c8d4e29aee130d1f358534fa94858ac85dc6d892a79caa475d49db1a4f4a88689784be48488561fb53f2ead0359d9d762c9e443a96276124c18a5c75c9c4fd4330a1db5ec15fd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5895ee7fc1164ec021dc4d95e459b6865f868e22234e81d7be69e8ff67462264a40205894d54fd00623a4e7d49e4f3b81421cf1d8499b1d46f4ac13e6721d4ca5c026f20a48561ed6234c73a5659bf56a4c6fc50c5917ee94668afb9108558cf26228eacd88593f9f51c2e440853a369f11bb91adb5b6b19;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h175273ebfb6e0d77f1189ebd72f63ed1ebf22e3da860316ee0895d75fa8787ead5724e141eff91bc8c88c47e6ee2a26fee59baef15ebbbe9d00cebe01387dc50735cc8df33dd04506b4c1b5393f5e54ba5d37e06f788f1f60556dd20eb660c025e69cf7e5d47b5ad241362f555cb2bbf2989ecf79c40e844c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h800d31364f85a275d8271ad09d047fef0fba4564ce5faacd095885b81d8df362fa611ed9162b9fe8a1a13cbfd61175bfa4fbba307b0ae4894c0891d27f160c35613d03b7e850ff540b2e3bcd47589791b195500ede238eb4b12f140863f2e67a56230a7f6ec914c198d657258bc2cfc1c00e3a7734a1bf81;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1793c58db3e791039973c213afd00698263a93098837c8d78c5d547e64488075b5cd675b4a34c63976185e217812a425f0d89f117258e39820b0f800327b093c852524a800e0d6628e9dbbc2965acadcab3e9f99dbaca48817caecbf977a3195d4ac349ea055efab1c2bbc2c0a6de1cf3314518e6f7c2aca7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8befc6d4898907cd485ab5e8a77f25a8f5258007aee22215f9ee9b37434fdb0d67d01d0de00a7b8c9ce27312e2d139f546b90495398b6747bf1465775e5c0f8899e9caa27656ad518ffcf013e845844678157938eb4f57d854cdffc205dab6156f0e5c230497d910061fac289f16d8a9a5f251709b134be5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cfeae232dc071d604d23ecedca2755c58be98f2ca429413e852cefb181af3945ce6dfa33b29e891318472b4b2adb601eeea0a622eb3fa34ff14f4d5f9138e1eb3f6f90b23bf715b98f40ab4a7531a213f732c2f2ff4787eb748eb149dc7478750b09c5138659e7c94f303dd0087eb6490fc44e6c02d55167;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16b4a011602358141cdc3ba400855a960cd71cc0b48225814c79cbf5b1c1a4090cd51ef9d5656c675c3cf4979a1226ff9bc5596f7710b4016e13a8820a9db1ceec32962e7c464650dddafb570ff90a6a2c7db3eb66a0880482a7693fdafbe3d3ba200f827ee06dfd0f791045a1cd1f1bb5fcb75dd6c633266;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h22994b2592fde20e4db7d37d18d16437097e2670a0bb2f253146c4f57741957fa060fd2c22de2f62191cfcaa3b880dcfd59d3d2596290ecc80f671929ec9a66584f633b3cad6f887adce75cd74ff1fe45d5ec91ec59404f23d5e87975e18aff62930745a2e2ec88bc43eaa59af0a1435b72362d356c17566;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c95995d0952da6c26bdf0399066b4b2e602dc58d392b39f13fc44ed1c79b4275740326bb6497b7777ca17410e64d27c0a973fee1b23011c721448d24b52fa5413e3c1373bf095c36fb51eedfbeca5845c0628a857145e4ad87e4224b16e13a15e9667ebaceb25b09701eecd9850a66c0d31f14d98d8ff17f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19e3ac60a393c84140966ce0e56d8e873b5765dec015de2cf99bef7ee11960ed7a64c58a83f4a7bcf464069c341d36223687865a14c6d21939609d03cb04c4d7627890233fbb95afd62e96e72bc7f5977d03f83682aaac5372bad63316a804cf915cbc3d413e7d372a629ba0b4617c6e7eb9530c6a423b22d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h36517eae4a0a2a4a2c159a7bf1e7500f4b797e2ed954f57bb25b9182f880f634e119c1583378ff82f69777bf5f39753f34df2138949df807e05583db80a991c176ae44eba8a4b618f7772715dc09beaaa4b1a5c02c4aba646e37cbd7c68fc4781b847de98f7f9a93fa8a4a00ab3ecd99ce68e23571783ccf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1282068d8d9ff6030a782af670891eb33fd5cdf908c684a04611677b0a3e0f5d3dc48cebe55f0f822b867f13d9d315845fbe477603a631c4e8c0710d7388986ab28693825bceb3130dc8b880b31ee3545401cbff012a55ab3650492f574590ec643bbab4a4c074a72e9ba96eafb5f80fc6eaba478289fd0e7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h41d0c6a318d07aa6ffc501dbbb3a255586fb67c49332f658ef8db4622457102a338ca11f49b813711b9ccd01e14647352d94428f18e1c906fe5fb1ee711e65858234778f6ad322a3178877a1ddc23c6ea7508f480133e44984702ae489d65ed0457b91d66c2b0ceef12477ecf4d415332b3b301fe8584f6d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h316f75d078c011d10c051fa8d63db086ab84eb3acfc3f59abaf204d8c524a616d8236dc44a544c54211d4795fd885abcdeb9a928b264323cca3521d2e3373ec8ef026983ff84e2fffa6a094b59d947bb9fc848e741b8c51657be954ff08a7de261d46b800d818029706ea96c1744278eeef63d41e1ed1ac0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14f5f3ce1991cfec7c29b90895459ac3af23813410f804e31bd42aa96b916b72c99b6f4136d541afaa9c21a437ceb9d172e07088b9efe5c229528d1eaab7b930e9d8ff561f02eec33426ed46c2f4ac70fa5a151aad4040c2e4aad86623b90a86821c095e363b1cb1983481e48bf24037a9363dce6d371a371;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fb6a5eaac618b509c61b7a4c5f2b21ef16083f041c5d554fff2272c5e77539639e469cab519a37b4b5cefb225d6e8035ae99e2f4a4ff6c1efedb0fc36ddd135a9256e79f66354ce821abf951515df68104d30830d5bc4e2a3feb54d1ed2ab6c5d451421c5d60cc798f70c4f29583bfbd03205b5d296dc416;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h104aa765a14cc0c04ef5ca1d1cf5fdd5bd34896dbcb0b4a5b404761c2c82e0c3640ce8e993216aa4b7d0773986db31e6820ffcc10b292a52d78e7f41694f2002919fb28d2f3f54f6b80caace9d75a41e9d3fb4eb53d28de0c8adca0f00537da7cf6579eb7017e35da05cc0658089fd2c29a2f755f89c30851;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h198516a6c0fd2bf263f471f0715ebf1a81488919d8bdf97db9d57244e1819abb937268cd2e6c2b58e9549b71cd9c32f1d9f50f8f89f82def3f48caa6b840ccfe53727468c7d130b30dc9322f5afbbfe36b3fc332c9d723b68683cace08526a70a567f2eea7576f5244d52b950d594132b7b565ca243e72525;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cebf1512dc46d3a0b7a5177ca7f7c26cefe301f53f040f2cf1a7140791c620c8c0068a1f0c36b7d31eadf083b4ecad973824e646b80828b06c804d56a1290470392ee901cc838b0b3ac2990cbdf9f975b1942ed8517686e9bc77d889663318de55e4ebb58837dc543558f6e717476566595c451eedff0087;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b133a9e04dd0b14ca5a5972bccdf18fa229b15a909eaa2c901db3d6415bd83d4a9ea492577b27a173673218265ca742da729975709e0b1a2a520fed7c1dd69f406e1285880019ec005d69d78aa7a0dd9cd2258195ef56ecf7f2961a72763c9115751c35def630eec8a49ee72d931b412de2d39379eb3728f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd4d189236cb6eaef9f5ac50a0abd3226ce4db3fcf52eafcaa593ccd95b59725a31e5bd5ca7b345f165983869bf81d3bea62e0ee5d895a793c338080f14049e4ecd4dd3851692d78f25faa21cde42ac4b928df9097dab388fe9e2bc158afe4aaeafa228fc8f117084c05a1e33b98c7485be411087000f6184;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h79761621d10490c1a2d880b849e0457d3e1b5a43a0812fd2005618ed2bb4c03e8cc389e0f94558b51e27de8085d1e8cbae89d4d38495677d8d480715ff1c446ee582828f01de964c2a926551f124d46b68a397f4f7ffaab1492992567e670277ba00e1fed42d3178bf0967fbb210d87314cce9888cfc7252;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h147c4c4843b86a2814fdfef2c261e7173e10c826b3d3ca39c9e58e00283ea45851a0a14657a3501b324fec732cd2d682c214e5e5adace744a8e3b4c313d90c96eb3e53101bb5ea158cec81f4b047f302ff8e3bedff3d6237452f4fe0a2d9bd961179fb82d64de7e5317e794d0f7ec2d9ce07ace31fd1f86e4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16e59ec881458ba29acadf06dd1dbf64dd594fe261e98f4d0916c83e2ff239cfafc35b2d5d4e038551b0f8e5ed97b4275ff408b3665ac7bd62c414d048c239e53e474b47628ae140eb21dd026b4981a850ca66d7899fcc3f27e609abc36ba2ead97254129ec9ed9f810b0278aa359f2d22cfd104dcabfe447;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e09a243e0996d56110133820547554d3dc2e9113215772f3284ee632bd8c14b1f567853c19b61c17d6aac498a11ee58065b38732e84926771e2d66b49bf4363440cafad1eeefc9c2232c2a318fc1bc638ea05714a31bf59c5ad55dcc6ce1cfe8ae3a7b9aa847adede11a3bbeee27b5363bc27c64b5d272a1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7662248dca862f85baeb836aa423134bda99abe75b58264b8c2514c459c0bbc168728feb3de97d3e78418ad1f5e1ee4e1e2dcd7b58d516133d9e9f52d262f099cf2cdba82fb6ddf747db6ede290142625f21923c84a26f726e337c80686dd7580ed71393a1aacba614e29d5e941ea63f43d4cfb662aab5ed;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1eacec92022c982b0aec70c7c1b4ddbdff9d0fe320da0d1e79f09b3bf4bee3c93dfae05f7341ee6412c6af7e575f8d6cce80980e28685eee6cffde2e1a0b30e5f503e3e524dca74379317dc1d57b8c5e0f81fdde80fd96ce10ae99d21457a14d1d02547a7583854e0a62a9ca1d488fea882d91d9a75153bcc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3dc0d33b8d766037a7f87a0420bfe21d6f0187e86251b96226f35c19ee8f767fbabb6118b544464d51a9a7a1d1ee794ae599ccc1b23ccbcfa9e3d6f4093367aa8f7ff25ad58b3e87274143f912aaf60e198544105b53967ee187a9529e8ea02e6e41bbed5261cf7a3650328547650d73d8efa202ca099401;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2069e4905e3542ce9978f1dfbdf1a4f8eb0f35f03e39a27a36348fdecc1cd3afe5eaf50fc1b8c2f40f0f63dda548feb32dfef9726f53cfa1dddc4b6acb1fb913b12b0933a089822fc25086c85bc2a659f1987a366e91e01bd6e5f99354f0a9a44a2bf5b4df656d82e07a519facba4c9fe2450b6b52a910cc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha1f8e26e1d3bc05228ce1dc53f422f59c47b49576b35772685cf47fdc61dfdd7753dbd21d1bc30c63a3eb436062efa91e09677dfea3f49aa331a7b43ecb1b918a0a29503e181f8a52bf19b4ac883a44657aac5c1217abcba057dbb416749a7bacfe88ddfd8f074f26d525a9e74bc0e5db51e2ca3317c28dc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16a9bac9b42442081baaabe7af3871693aee65e47dfd325a63fbdafc0317be7df21a059af75d24e8260414cd35b245a3d24ca3674fde7eb88843e357c9251d9893a5d12641e467ff57b586c94d0a4d7aec5dd53672d8add01955b53c2776138543b7653254fa1f434b72f4ca070954b89d5b3d6ca61246e1d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h814fc6bf957c6b838d20853290bf39c4b465e0ab0731f13e599c41496987fdd5877dc26684119d2a4b803f6139584d3dfa74294097b6610aaa425f72ce89c507e59c108c9345e17786ec6f430650a1ee669b378b70775a426754dd5abfb9863a6819e0142ce60d2e66c7e90ddbdfc8906eda2ce090a3b13d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h591e86d4917ec2b9f3e608c4e21300349b55d72536d60a1ffc1d6548113f70adb2da7efc4ac98ae776dbfbbe893bb41114a534be2e2b540db98c4e9c98761dcb70c2ab537896899a7c5299d56ab7eed3f22e74b6bf3f013cb92f72a53c200b866a1d73eb19aa0121e3682f0e758b1df33438b3e173c35849;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c9ead23356183d5d13037b0946174f06eb3704ecb1b508d2234f819af99d41d2fc45923e681a8c14b957e9b26dac85aabd91acaf174d2d7b76f188661338f60c675de40a4f2fe0d3804b0c8f60bac4ec9a6ccd587d553dba417d59498bbd5000010dbc5d0d5faca188be68cbdb38f424f8c36af1251e54e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h29e06ebd75f5f145849253717f8d4a7cf01eb81d3cba26b67f6840414962ddf318d6e06deff8d1f13c86f1609844109976c8651c075983fa2f1233c6330eda3a198d3bf064a7030aa92bd49452e46d42753d4d248fe99d0157201d9697ea52143db0b400efdb3747f4a91a4298ca7d9e6efbb7a65eddade1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e0880f4def80fab3e67249918831f692d5343cdb48e919d7094071c76f3fb8697c917b8f2e1ef01f638632e730f32ad9c062a19b899f4b5819c6aa6160d7e7ca85cebdae0361c25e21d4d9fe09304a408c4a063d44c7dad769c2ea52b88620ee08f400007521ccb0a067a241701c0054f8c67f8f0cb8f8d7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5e4b107ff99ae277b33393be138c789aefcea297e5f5ecbb54f298b27a54793ad05e74c5fa766c73f246581f81a6fb3f4b994391362032e08f758c3bc35ae9f31c10df20d2111a75c1f8abbb39c5621d38154f9892091fdac43f6e83ae6605009e2841bea6eb4fe0313508b657b6ba80fa002511e9476fff;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18aee8def7dc73ed54c11ab2ea57cd60da3d3a8425e9e32e802f617b54758298ccb99b2ceb7480dc6d6cc143aa750193d09bcecfdbc74311a07fe2ccb0256f1c9f4138e54a79af1d7e4915b127608284502feedca2102842762caf64e80912052afb8b45a732214cfb1b46f89a66875025aaeb55da7fc41b8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b1d0df96b819dbae20ffc5776986a22b7e79477453e6fa30c9eac1459769c5b792815fad0bd4d05a15dc699a75bc2116afbfef57c47310072e6b064418cbbcaede4ed4af55848b378e7653e7fa3f769258a8457b65c5e3337c9e54fc09e98471a301417b20b2895ef99534e3aabbe522012228426e65d34e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f7b6f44aedd62545b41e1a3d74975fc976c04ef16defdff8c77a2b5b3fad4408e970936f415daa3d54f31a57419794390edf948fbe014f9a801b8d50a8012e9171158bde6eb16fc72c672ee2a23590ac54222bff5c1bb3f0488bded47872f10b009e2967726f29448cbc3121dd7d5d600ebd678c3a93415e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15bee340eb7b3421576f7e29fe6eb45aa242f6fac456b88d304e7b0b741ef4b8391751f1e1988b84206d4d77380cbee248b973e0b79a28762515b00b191e5e24bd967ec49d9bed4a1a8501f0dfa90e02db7cf956828814a7a7aab2b6144bc8cbed76a6496e6378116742b9505a60e919cf13c18c7bed59dc1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1291c6ba2ec24b3cb28c2bbad111c38ef60c3c6d9292b0fc84dec0db189e8a6d88a4ae0708751b9c8665de066ecccd4f61a45a04614440167e1da17b775abe0b6767e231eb8648ec07c0372472604ea578397050470648bb2a05daf9f9398e2264b15699f151b160e0c5c5d0da70a32a99376d6f1629f5fa8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15458790ab7db2a2bc99e9ba881110a46e5c6616a2bcc7479f9425cb1b861d36dc39bc1215c27d317c6f8b77cf3c005294ac9af114f801f132e5c6f7046dea6f395762d052651b73be5e03520c9b0dcc09a85e5bfa945ea69201bdfde4243b9d1a27aaf6967906de62f5635077992684868009467289ee376;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h126c4b5a8650fe84b676d89cf26fba0a6a36e5371964d82e6bba1a86d5f8ef743209a61aa08410a5a47cfc02e4cef0697adaee2269dc403d4d7dc5b9455250e56819e464e41e78dabf00671d58a67c50ff322223a863dcfb08cf3ec3b2e043be741f0960fc2e90ce2e00989cb6ddf04b4b56b597252e676c9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc561990cff05741821a8b2e82d610e9074b1f821a7b4df56c1d5d0681de702d5b9a17daf9b43cb9cc6627a06298a29b2a6ccb28455cc43a3e056ab45a9f2a5714f342d07fca283481afff912974871905a93ba3f4b2f36a3fdd8e515082fc8af8707bb177ec9d47772d226d378087f5ad3157cd3182f3a77;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha88aebe2535d19371179352b0c37cb93a6a3386ac2e548a6eab2211d8347a9a18a878d9411e2ecfed8d47c5726ee90696b1c0840b1eb900603612f9471d44074ed0ece24349dc7e3a6a8e0af684fdc1c21b13fa5b7da35ae5995824d6f4ae75cb0c6ff42dd1bb60b50ee181390cf211bb40940aae720b68f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19d97c4123421838692125ee5160ea8b7950b67998093676d4aff35f2fffb5eed5c44252d1e6a3904fc9fc3996629dc2967e93c4d1af89b505eecac22cd3edd4b2248a6c718fe66033141b7462411ebd30f83afa7cb813c4b1cb02960bd62015610bb42d76ca930d29db64a114453efd397df26835e23b83b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15f0fc462c5ab3174e4156b2be9f9ecd5aa18ebbbe4ee36cd644c6fcd202d861e76b5bd1b6d79fcfa72af90a49d43b255b06233840ba882d7c749e9d00f1e233dbff83101d7e8cfb7e0f650f0d15a98e0b452fddec15962509be553c00d60342a8d7127a8d37ff005ef86863c40ca1900ecd7c25c81c2bca3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1374f72d64251974885e2f71d9dbcad21a7e07f7009e21ab8b5fd1b65173ab23ce6c0ba125b2ed2590e0117c54374ea15932ec27c5ba64f86eeda1ab70400868d6daffe6a1bf597b03d012acede8075b65041a879565e1f9fa180d511bfbacfc9f26316214bb18db68efa808e06dc9786f7f151585e3b9b92;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf8ab24a8f805474a812254aa415f5c4613fc303352a9eeb129458860d516590ca8007b2907c1a25635e1f130a1495f2705417d53dbf974830a0d5e099ac195bee145b0f91cb2fdc010fada03905783b3e8655886defef99cc89ca0903eabd10865d83284e3c7bbe6edf68d9f46a8ad9cf2c5be0068135ee4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6846fcb38e466e6067f4e86a5018c122dd0f7f7e2a68d9fe65f1951689210ab662a8ff08d1ade3a7ae306d99a2057a777d652cf7fa58a0b7b4ea81e540572f25ac4cf2da549e144db5f57f8ee29693794cdf9820fc31b74bfec60996d096ddd650b7739991d628bffd4596d65c4f0672e91262c4a4be79f8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h152788bca7fb3540d1dc209420cf60a2d0055807edfc6f840b3cb194483ec2c5bb4b378e24c0bdcb420a99f87691320a319b2518cb8f9a905fdedc91d6a7ba8157c36fad8f7b45c4c2fc4318912453672c9f31d732b95ce09198ff37ec1868030f6a65abd8250b59c435205bbc903c5cb1af4414a14f1f031;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6fac6da01544fc0084a3c1639d45ef309163b3c6f3713922a2f2edeed1a3b510eae9ca6a226daf1c95fda2223b79c2aa345659df80c9fe0302654ffaf9905c978d53bf08d5647d310fb475688b9a7284bdda285ca5cc52f9c6605230960b033450d0f79058b87135318c178e53b6c3be54c1bb282e6a7f01;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h355f2488a86cd922ae1f16bc183c53e2208f5344f3580c7ad26f0a1364fadf01028e5275141007974dbadcf3534595b4f44a4a05381acde3b8dfdd2f58fe8311e349680bb20600ee06c50ac210bde260317f03b197074063aef1f98fd0912e8b6c4cc7621da44ab65c4ad34cb2acd71665d5da39223fe122;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h201dc90bd0fab3d52637acfd7b91f368fc96a794f3d92a5221d05c9fbf0cbd6a833ed7584ee5ecc865f49430c227742a16640b7f67e121ff3da5b0fa28d91083fc7458ad79f56667d2bcf8093b83ff02f12c081b2c4dc264552e05e6c1706ee06cb73defdf96a988db317d628f9e184cff3b9eb73cec78f2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6e18c571d9c620986745dbae3f21d4705efc4e601f9151b7242f15b5ab0c80ca4e7947d4cb790c045c2e1875ebc01b0c40d185e629d6da3d915e696efec55fb666cd8263dbab71f0edc32ffc7f77bef50ef49d83829f96d8867ac4fef66c7fdb30405401be22b2ac1e9182949908e309ed66cbcccf83faf9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4a028898d77bf9d2614ecd99fc30215cc7439748a9f3d21399bd9c14da6b5e9292a4d705770fb5aecd66161f6d1df73adecfc3f7577559a352f1d8fc29921e97827f6ebc7bb2e0706f6be2ec0de955e3fcd6b9b9b7d1c603fbb5cf4cdde6c5a59c83ca2f4604378e883b56099d5a693fd2c469f20980b2c4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha5f23154b1af265a1a220dc8151d1497aca1ffc308317ffdc78f8758ff5694fc8b55b9f01b8d53c7f0ee3993e4985aa0986f9806b9fb7329dbe64c673c57734db7137c4c70213516b4b5a757faf7f8137c08f0b2f9fa96db4f5b7d18baea64724da261a8e271e72f6b83754bb8713e270f59caea1e9fcabb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c69869d96207121bf7e371e728403700ea5f71ca255afccc0b74215e4769b8e49d62f52e0c02e9a02c0d0943c2f308064aecba953f4b748f7a9202c38c6f2928fd6b0039cdd897fbf86c54163e888220fc40062acb184ffa12ec271b511cd2c66b3d7191fa6fbe7b33ef556661386f1d72b7858f09034339;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hee3eebdc6c16a5bf2e4f3be65318770fa54acedf8657eaebd2675c1ce9c494093dbd0db6b5d9ba3f11f934fb218f3aba712c10f5b49bc318b4b522d6e7387c77539ee91d9c8ea928d522ee6adf736556de3959689c8b0ce9ff024fac4631f59f4c07b544fa70c8da81f8b28e6cf7a6148e28c2a11aaa00f8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd2f79e4be65a786c80ec9e38e647ed8a51c5e1d3ad88b22d4156e61631574fba077530141195ddd20d036aac5e417c45ab5f290081bcfefaf099c15f6ef57ba3ab07d560b082619bfae31ae42e20b009fa70acbf78d814ab58e0c13c40e98bed9351b96b8379474afdc028bfd54ca354da7bdee017e2c69c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14a7055bf47e76dd2d78d268ce8c09e45eb9cc102c928bd17168b54c24d88dfce733c0d9dffdae3ca51b67dc21935bbec0241238be5ab0773b04e28acec7c42b0e69345f21d0d2349185f0ec7902d79fd732ba476820fffcdb93582b1eaacd452e696e1628a1b0c3467498497e7919ed569dbb42a2e9c8f6c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fdbf77a44315d6bb97645952543d8a746a8d77698e10f521b2dd1494f5d100195b498c301c80d20a662345ed5088bbc6235cba1097e2aa8f1a12bf7f2bf4b136a3f0e986dd162ade429f1c1a994f272e4acafbcb7c5cf44e1f54e149261ebe71058915068f056f5a4b8d540714f9bc3c7f70f36cb38981ba;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hef78bfbd91619e10794bc72feb654a9b7ed88d1b1cfa6e0c448649dd7f2ba3fe179693703b15759546b1bc366a346801e3e33954dfac9dccc6a11ac524f852d653e57500ba0748a13a7bc8d12a1587c37fb9d58547122c1ab38de3ac617577119fea69493c26ea32fd08c7f444a003531be8f6fd3199fcd5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc032974f33ddab7fcef19d50879428277d3351a3c97249eeec55905e2dd867d237c97c41e0ad811b0805046dc48054ab2a41fae6c5278a8239a310a01365bd4c026ec753d76d86daccf69e2422940fe1659b1e2af953e400aeffd94fdde6825820502f9a4a4cc8ec0abb6ff0760d6cd6a58bcc9a4ebbb5c0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h82a7adf67ca10601d2131d8c141c6dd7367cb0b13189cd553b07999d67fc889f4ac8f0fa61bb725c9d3ebb1c9afb9b52cdd50e7b83dfafa607ee701d3bd1c1d29f592d2fbeffaef4cc7d768720523cba7b5754586bf771db393fae599d741101f973b1a6a6e5f37e0ffdea6aa68470644c1eb21756f465;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e90cc0c7c947b9cb928c34278c43eec38a0e9b13bddc3c673823a775a4291611dbfa5fb5c9c041a819c060e666c6c5778066635130ffe7cc71229a0dd7a555a14329fe052c0bf3560f5b185db6befddda046a9537c79ee712a485ad7ff40c1d2a8028ea68d1c0949d2a2181e2b032beab9509674cddf0cba;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11dd09c3589f26c0c4bc74d31ebba430e278e430d2db8f2e7ba9fda47cf783002e295968bd47a7af6736a998d7d1d25e6824d3062b6d3a161891900ec39518095ff26523ad1b4eb4068f7b31462d9adc3acf851cf3e6c9dbe47724e2424b14e4efbd3ad169a153932cae840bd60790514c65153a128458591;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb73d08bf536c97792704e88089bad7ae20e7498ea36d03165240ceb46eafa5a952d794dc06239a692bac081d3d0df835afca9c2d38c50b3af09a7fd56ce72b335ff85c25d7253397be524ecea057d247899a48db7ec2f39dbef7c16d2edae7681f1b29077a4fee354b17050622323620773552e93d68cf12;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h177a368650c20c420dfca78c39811934bce282e10975b2a97d485b713fe1b9d1000a01069f2c4a8b713a469863ef38124beae745403cae8616ad40aa9f838438b4f379c82251f3564ad0c7b8ecf2b692a836b3d863edeeb8bd285668a166b66f6547e05c901e51c579fa8941d0352d56bb548b08df829538d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dead240d33162f3abe8506196d2041acd981018500cd2add5a7470658ca035bb3aee8facc5f063060dd9d5bf86dfa5f6ab5bc86f6dae25d17a3ccef64c75d6a7ca3a9d7888b91c56900ab3ca5be4d093b5b22b585c8bb467c51ff0e951a0bc0a697eb7141cd76c8a13986c9f2fbbb38930a4897d71142cdd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9aceabf158aea7a1eeaf385c29f3d94f2997d0ce4256104c67f5020fe34d9c1fc305fb5d1502ff2335cd4e912b9e243ba6699c0744ecd53d93f25c20847e890f749f0966050aa860bf9dbde0b8eb9af442a3a93234118217419eaa3986628c3478f65be71c306aa697dbbef96011469233d139c7c6f8f69a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fd11773bc0134c71b0525272e2ef266e6792fd1a67e1a101c34b4a37811906a28a097ea1d63b46ea0c649be3f9d072d0444d387353257d596e58e7f5739db07d85ec78aa0ec2071e63ecf3f1e84fc41f0f9ff60a5ba31aa0ba46e215454f98c9501d6a614e3ac544a0b7efd5233947b21533a765e755d0a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17e6c4fbfa636b340680d51f93152b14dcf4e0d4e2c8a3f1a358a46a0b0cdf7a6f9975986ca06956d085447bc4022d3bc1af782a7f03cacb588d8fb03a053caf65f76cb5b63dd85a1c236b2b95287aa49cd3127084b8ba974663f0d36ae1ebf822908c619a77707220c3445b5187bdf23559ea6a7db03a53d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b2ad597b51b42a2640bbad7741b7983725164dbea6be97318acc04657dc2161a6fff25b4fec5ad1e0df385b33355f8d6d85ba5c27378d6a524932e321bba47ce485a3870abddd9bb5c6eff191793f5fa42271c31c9c29ab6adcba77e93049aa689dd813e16de5f801585a9751d289a9d2431c421bfae039b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9b77950f1491455fdbf618db50c8e2179229617ff35c22fc01fc45cb5d519833f7c2276c22476c492d33b47beb07cf7678a6028fc50229e0f0ad56954d1f89e10e125b35e360ad3f95002db18890496c29d69065d0775cf50b2239a5605e8301be2c5085273f359e1b23bc687fcf86411259a0d54af48127;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16bb7b7294b8ecbe8fabe32025511115e7f5638702c011e0f425c9c98d825eb9521215c452ae9d0d2af8b968f444db1f2613cfaf5098748d891a8b5e522b98384f3448d9e90bb5d2a488a4b32071fc5c06c83b4106f96a5f88b5bf8df6fab03d7506f35e3e7fb7ba1613ae567bc35f876243c3cf5ea9d1e70;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h196a9ee12365f6a8cd074030d72c1876ca560064e37881e7fd2510e8daf749c522e17eb201eaa0101aa6c5b8430e43321300cd17fc377ba59eb56583767a05c6e43fee90f3f4ccda3b9f9c0bac7ef3e2baace52f18d4047840d05b2af26eac4038f88571b8582b508799b0b3f110cc387b802ddcf0f860e5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc72ad83e70a66c800a0d14c5b0cb969e96def297ff2b1ca94e8d5863ec3118193a32c1324421565fcd2aa59bcadf8c4247f2c223ac2c9b4779b8490b5428eedc9d32ccbcffaa47686bc22892bec717120e85377b5f59ad9afd29e796d1f20a2db403976935a697ee5d01f33c658bdf137e95f7238c473b23;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd372c1d08a0ffe6070504b12015e9494bacdeed4dda76bf9cdf106ac2b9f9b31e6342cdcb6fb3c298cfbf9ede715f4aadc22225c3555d3d25426853f2ea8d90047a858a459c96a83c29c07c7d06cda5460ef570be757cd748b615cb27fcdbbfb816cba907ab335c050afb0fe12ad2d6903a96b9abcc40524;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6ea5340167ecf211097471cdbdf055447e16cedf8de9bf3e246e50e00d80ba253e1de9d628f80821df18f4ad5e8a2a9825aff56feb60e229113286bd84748d3efbdbd667daf6deeb7fed87f2a6174e8400d1ef1d1e012526326a31b5997bdb701fb709235c65fbcf24a5792239f595a9b5fdb410936ef195;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11ef94bf65a8896dcc00fd8ee86fe38b0f458123bc29ff351d1efe790210fc6d71a245df2e60df250e387e9806d938a7df14ac74970f746682684e3355f1c8b9a40eb02712c22dfc11f609d2c4f42ffc064bba59122c8a57a77ef4b47b0ff31b09caf7aab4c4af400bd76d1c521b106294243ce31e1f9a51;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b82b2053674a7d6135d6778a19463a807b38bf28e129ede378a581deca222d0394905c97d3c302780c720f98196a59031462d96b83eb284e6cbe5aa31f140c5337b8151419c485aa45f05e9eb232873a6466e02f078a17b45218ba02b900a7dfa6846b95b21ba2394cbaef218c7e41fc3368afe8a65a0b89;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16187febc3622fcf2996e7e63208ab6eade2d27362a30f972c3f65c7323125979df88d46d669defc19d53c4d5b57119a7437a1655a901ba8bb9545a27852d857a9444bf1e3fe230f510be6dd390e7b07be150bc7180927e8932023ccff5e13d29e7151d0e7f268fdf2cf776b0541cbdafde554eac51d8d93d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6c7d345ba1f8eed50b776bf0a0d4364a692c1fd8143825cc238917aaaba4b1fe4fa0a95c285c3305b570b2c7a11d3e4497221c70c52729c06ea4280b5df5587d851afe4296566879912a649dfb1dc7e741762e44767f9979b2e56d3b1d77819d5856193d65422aeb48c7a3384f80ab7d391da253ee71970d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha1d7284d3380a1fbb99307acc8acb299f138e786486006c661f4e32bbb49952b35ea429bd06e77c9be7b18ce1c6ea03f1b49f056798aee7fbac36f9a0e0f901364cf429cce04fcf9d517c82eaf35fd83c6bedfe1c0b2eeabe5858a932f2bf6520d578f9243730ce57a5e50e0353c442b06595e807d9b70e4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7d0a298f0498956b1433e20f0acb03634cb168e03de49ec4085a7207de8831c865d4f433c71a46f62078cf5b0e79c368076bf3274e7d191662807f1b25a1890668735cd83b8cfed651ed2d400ba5c6d44fcde42b677c3fdaed18f5c4c633569b958eb884d103462fd37e9046bb5894ec782779073aff2df5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he4b1b7ebb5efc30d93c40fd2c6b89d19bb0f25995c4f3e5e35bc7e6985c05c72ff11a39ec677ebb0bf2391e59f6181fb1f32bd5cd28f62db5fb796febc05d86a60850fd35bb44e64cb33781a2c14c1570980bef2d438ba212527c67c952e03d806b84a5c5bcfef60e80df5b18f76ea64006b63e86f41b17;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12130759d50988d4bb685104deb7bfa547d1aaa323274922140727bde08afe08b4e8dc2b49e8339f71e525f8381bfcd9bf411556b160fbd906fc4e0c95737a25718f0b77b533bb924d970f11cc079c7c41eef1c1af9c2bbedbfd68db52b1c693d6e2ded0c3ca7e89b4314b78e3ee0eb01e52c7769a7e200db;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17748b2ea11b4641f9605029e5194e6da024a9262a62c1dfac0df3c2fe80e850de9b377b0cb5822841e96c5d870447ca34d284c0e25eedf54856632eba23781a10db39cfbe76d8f4b3c466879e5df769d33753e26761a86c895382790cd062376b6d3155f3eaa8b8b4c229883666760f2533b4d97c810682;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16e451a594318e5c2ca482afa41393383f2a760134319db2d1bf1090ab46b6bb756428fbe28dc5d6a645014e798d7a554c1576c42c02eb7b2ee51170051f7117b5a10f6dde7b606bb0af42c320ae124d54af2d7a71a971e769551683b6d4abfe9475db8bd693d70d87795e5e16b3cd2ddd93aecfc27cba4bd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h663af32dfc9562918babbfda6371a7d03954ca16f1fc70f92e2cf1b4af24f591e852d0542253a02fa3e2da5aafcfa1e27ce22e57adb539b32f6945fd46df78c1024ce65ffbefde764ef76dd505c1f35ba52fd8131d0337500beb62ed92eaaf94a48a449053cb72b87516438e346a3676d1689af3a8ab1772;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h188a4e53dcd97a532e9217fe972d704c0bd82341d0cc051e2c71a2226e91ce2230273405b24cdf7d1d688115c84276f31ba08b69b57f76a7da3e5593863b543036c8b297c8c276b03f02927ad150f84ae03ae98dc64af07d72e4c2710e27f226c97bbdb382becd01bcb142106acf9b1555c2c46c71d433d97;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13d6d043a60036b50eedf80c91bfaaf1260e22713fe1086833f75e737644664abc3430b526a103fc552ce529ca98db62a6df2c73bef34e6baa3ed9918e3ddc0e58c17d8d797800ab6f996d6cb8dac611928522495fc007db1503a5bbfd422b9b4ec8acf5a6eed3417bca281845065b3a6335a2dbe7565aaa9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11589cb0628bcb0af7c91ae3fe5a384704c38709eb3cd442754a629a679b7b44e2c27faf2e5df3eb658e035558e86440af4f60f9b669c9ef9a3437ba632688a068ab1bef6654cc6e79442da176608c0916dd7043cafbb50d3530408f42b81f5e3238d51895f1f974e2c4c2feba26160e7c87009ccc20b82a0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a2c17774e4b5206e2e222fae624e489786966a6bef89dfc575df05c48afd8cc84ef5595d2f2b72b6db766e7fef6c5988f8929ab89263f3bcb6a398f4f003cba8bda18b1d9e34a05d2dabeb034aa8d913763b280b425b5f795a8b9fd3e710c3c39d72a770a5a5aae60b6485ceac63931983c7475eefd94a96;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11318298773f4357ff6d70d039108eba2dc223bb79ddf87f859fbf3f64838ff1a7823b95ba4b079014f87ead095a683ee6cf6ce20fee9ddc16616cdb53fd89a1d4d7036d30b52b6fc31d1957fa0b99ba3f587f8e2c23735e30a40c179f685fb45f71d742f3d40e62a99e860c4470211a597eca4ca35c57ffb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ac5332bf7aa33d2ed812970c9d5a20130828c6f8a98a3e238caddfaff690ba24e1ae97be93dd6fe7d90e1e829dcde20b8e28f24833c7ef46e438493b677c3e66616fab40a7e318fceca5ef558c592fd88a9cf1db4274a4b198cba12caf7469c5cb12f2d96b4ffc21973a33b81c7c08bfd022c0598c6bdf80;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1be4a726a8c466f38ea4d5f208dffb17d5aca4327c3124e7d9b259c9196726eb244b80216ea25641ec93567fd33aa8615acf10a93ba85f3c50325a0d06ec5f50609a730f9d1a1609f8762c0e75d8c09f8ab3c29dde43d3f11c952aea66e2b8bdeffb3672ea3b6e667f4a72d1c72602902c0431d4b3bc6d81f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7a95fd0d10ae643a944ca0a24dd0040290037b6fdcd4e9abc82f14ba513d1779321278798e4377742c2eec8b376747783adc7886d580e300becad8ad65007f20bf3c845acfbcbe00a983c37732df2afc50e62c328322d12ae903030011ba493ca3092a7b78b1dbdf28a41a368f797fa2c4cc9f3488b731c7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b77ac4b50402e3a2129a7c152780fa5e08e0bd058740878510284b3e35730284bcf1b3a0f519ad8f71def7bb7512a24501b2beb4330b4a67c98e8a18ad08b73b238a5bf6efc4165a104d9ec4e5f25a6a9cac1e0f2e4f517c5677663a77976b4b4c8a6d8f959e9186dccc60ac4abb7727dcf53e6f36664f26;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15ca12e5ff1fa419fcfd9ded3319b2433830d6c1dd1c7664b8f62d59b7afabd2ef860d0184a371fe09f5cf4da194f28fbf5e322ee265de9a330c02115aabf29e10dcb9bbc06d2040984023d48f2d99f90b93c4b5f3b15b9b80e32e19226be19f21299cdc35382dc491d73b4a7d387f8159c4c5022c7a5295e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4eb3fbcb23784f7bb96997e469d7d6f0952b2a20dcb654035f04fa3438ad65165b767b51d2a266e4dc0febe344fcc310bf66be8dabcff9ce229957d9a356d8a00553bd549ee92e577b18a7771617f32163df062b443fb37d1b25413e06d6f71cefb4e07fd96a54f59915aa88eff2a94edc8ad427503ad4d5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5d05d7bc4bba00e6b4122081053518931cbe5cdd4ad200b8ffa0aa05be33dde336fbca21aaa1799b8e177feb099652175376c883baff813eba9d02178276079deabe822c058d43e5996681e5f714ef4972776d13328725e221c5e8594aa6ce39bb491918a8a3f9e8d19e665a105685d09cd7a0dc05198cdc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcc9ee32a8fd7a49d1fc4a8926d4a202f93f64f31b24411110a041e5931fd6908b354281ca445aa53aa1dd88f19a00f0165bdc6855af5cebf9bf34537011c7c5533852a21839dd0adb2eee30b37e1bf8177928d41ab5bc485ad71cf762b79f64a3c8c18af15d1e28eb9212d0918f7640233265ca29c52a579;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1713e7269fb4ec250a53d0681957df080ced5587d09e764587baf84c5c4f7bec904c8f4e9a725ae9b7f7391a1b4b36454437bfd36bfacee48f72ba7ed38f1965cfe1165e0cd6470dc0c71fef2bf02dccf0d95430eacb6129f3f67cd284559d0cc51ec7928d5758bb57b33f5982e9903bcfa269722ba114ec;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18ff607a2b6c05d83ab1586d2d9a0fce991c3fc1b1392dc99aadc211ef34f3fe9e6ec7e6e159a7968aa22272f0c16f40fe4bd8651e01347c4b9ac629bae6214e0849f9053f271b92ee6bef7b2e50e4749c5a44ec33b50519fd12862340b1b91b58f7b40dd15b7d44e4c69e6d8e49a0bd09455d7335ffb8980;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a2c5c283c410a4083c5501adaa1adb5c1c619a1d87df71c9308f05fe643e0ad84b8d99c69ffb0aba8c96419077c4c12ac32faea0a96e5b7921876a298fd7d1ff394064d6ae35f15adac2c3de9254dbeb60a912de4c766969332346e595781dc64be49b7ef2cc7c515bb292468f84c9a0dc023b54be96f6da;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb5aa7ccb85f5e42ffe3a529c0647731ec9e418c8633bbafe378c4052787010086ee3c5cede82a16f1bef5e1a6ebcdee145e2c6cd25bb4ae26f6a5dccc6ef01157b399e20f39a54b37d3111f1b1c13f911e69da6d5b038c9ae8288ec9f0620044e46836e2c04abda6cbf72aa776e2fb81ea450d29bab0bbc4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h107c367f52b84b1c6e6f5784a21af03333eb56086a948d0376211dcaa0c6c964a9e82638b3a33e494ee783acaba4db51b10f3cec60a1603d192f1dea2a530a59ca57b6145fb92badbcc26efcc68b6576f718baff88425610329b442fc589cafff3dd98e9211d4f4981420370cbf3cb993d5cc23ae8364984a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h125d71397034e36da788a747ae44f778e53ef6df5a09e051952f366415835408b5197bda5d84691ac7c79f4f66e986752efde73be48db7de60e3aa87e6615b604eceb11b11f6dcb274e9517032140e332abe7902fb4ac24469957f169dad9834864ff1a610c554e39b68e844bdc084cd9f1362d8cd467e92a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4e08f5d4268598550071b2f13b14f16231a82eaa4bbf1cb053b364d19f1f75886839861c303789acc4c106746d26893cfbba3305419f77bf1e8e5bf16bc92fcee83d0f107bf3e7873437d66963835e4824bb7bc0623640654e263b0555247a34376a1a8c6797f6df82f2f621ee33940ef577d23265aca1ad;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18dd4e1b038a58a0ed6eab50bef8b2473d824f7325e1e620876db844f31d2925bb99ef532fe62f0978828c0f490397a94bfc79f89ee13cfc6e54ae3ed84f3c086de81bcf830d86104d14dc998af12b97c06508a97b73f4bca1495c85466e18353226d5a6c4101e995be1c859248460984a46f426ae8741079;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc4dc6f68685ff74c2659ea5610e75185758179ebcd005bac393e60ac925b116e2c577347bcdc532004ef576c763a208fbd1017b82cb4c8faf549d6a91d3394f13a424204334036199be22199b330df23baf98f6d504436e450c98a5d9d5835890005af82d7ea1708dd985e96d20737eecc1ff0928e22a7dc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12776b0ded0bc82b0e62164dd24dc199485eb1fea31d0bf0ac444b2227fe5c9b292b22861d39837ee82e2649e279c3e7119d1a373f8d32da030e82cea9dcdfe333fb866ddc86f3170173fa6497324fc5738d9854880cd54fbca91159374633a13d3a4773d74d86df5ccd24541b45b2bc4d04cfe9a5243f3ad;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3249d847c5b1308e8d7b500d6d5577c7c95bc9f4cbdb8ba49e993b9adda37d89a42e9891b232007cdf38a5cd5a085f8ee35026f6c4c991e8b1fb3b3092d916727cca207ab8fad5f045ec4994f3b099c52e2a3ee5d47cead9201090d56e8ea8983e3ebf109ad991fd487400191bd1f679ce31462cf91db68c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h102f74836c62e712ab65b5974fb9c8d0c2cccd4463c43e38442518581698af3ef49251db62e73de20acfdad105e3f52d25df25d0295aa684d8115d86fcbfcacce021c7efa980773f3f0c3e78b790ce36e8a9c1c6d1dbb2f45f2aa742b6892dd6c8a5a083eb16c247a98b63330023f602a987b9b3199d9c519;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18524618a478cf92074c9290e1eaaffa98dea3d42bfd3292882806dd67dc99cfa559cce6c5d04fb6b9657fb41c1cabc35431f4598588f64ac5107ed0366cfc31b3ac4dbac89d54ca3c6065b8dbe303df04411646d3229eb270a3b5baaa640d252855c2ac5abd5851900f43058d09669166e3e4ee73f4614e3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd37d8f50e146e1a0820bf1c9e99ad733060268a5c9dc782f6a0940a09e04a5ecaec94df7464d66b25118a869b86565b9e7754505b62b17d55600ffe10668d08fdec4b813555d6edac0fbb4b6a909c50c0a38daec68f5b966cb2844b372a10e5dc343c22f45014388a5f5148fe251cc23b701eadf865e3752;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h137388657af3429c99df94fe64ba506cda5f5eaf48a189ab46a460338bec074fadae5d9cdd46ab14572c628137d3abc964fbcfd918b39577289f8bbcbc9e1b8b8f5b739212adbc7985ab9a5247f3f5e1d9bfd3ea47c11dbd771c414e8dac19272c06dbc0c105931dc4eb612b0a6ca7590c1b7325a047a96de;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4b6536f8da1b8edc18edc213d1f1082c50f9b39e17a53f387c25aaa368ae176402a0d869fbf602fd25c0211b2d380a9d473d1b87d00566cca0740c82bfc0594baf6c13f7298457662f3ecb16c958a2ee13f4775b77e0498cbf4fd659f4a1356b7bf6a6cf19027e1a5ddebc9f671cbb0ec7d15c4621b332bd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdd190ac871b964002b1fed77504c268b3cd6bbd96b2adfa2555f4ada272b78f745bfda50c590a864beed4877192f0e067c4544e24694c06124d4579333eac2ed08026c783fbd0762568f54bfc5e61f0ddf1da66eb84d9ee86a4c50de685244b72518c201f9b18ca383302c293614609c5696f210c848700d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1df1ed8729a8895f4a7962edb76f7b58848edd0586935c45f45dae7d8a43eeae3fdb9817745e7a0bfaefb6c337f12e28dc25b4d8204b0df6ce07c8d09aa632932611f939864bbea87d04180d1ad3b322115324eb731e7c5a8823d0f72d013146432e035a2a26f4f9883a4cff12cb60a1ee338f7d5f25ecff1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f154ffef91b408f7fe53d830a36e0ee4dd911f3958cd380c94ee268347eed484f4d761017e244db25ed1e299017b957676668f2bf260995239cb2798f7ae775820a660df9d074496dd423401a798364f7fd6cd69b70588430e984614b809ec508328ab736bcdd8571721a1c7c2b26a84bb18ec2fa9f6a598;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1af2bb39ad0dd065aba2a92f281da5b1f18b3133e32f268e63e6c31597952f917e4489299e461bd16d9cb641678f91e89aab415e3e97c57cba8c507d93a1c7b3f5f29db70a920e7a8a21f9de298f78509fb91730bec6328ce1112415ca5e5f5973c26684aeb9947d55d27227cec34efe8a1282277fecad97a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd6c5cdbf22bfdd5e0dd08f63b501d4d9d3ef8f98cad76ff586e8f232bf9b936114eae1e940b527d7952549c226460f74de676ff6aee908574960b321fda516dbac04be23e141b8a7cd16675cd4b2f498c3e0a4f8a2bbe6a2acaf5354f3b5f6c9ad2d9b266a5e4c1971307a23a8724df1459285b10b5dc6d6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha3c507584e0a1398f8c030ee71b8dc58f49b3cb8c3c35cac332331d0bff82b7251a190ba4f1261c4092e23463af283adfddc6b6ca05517c028f6589595f060bc8d3c6699845a6b354f824eebf66bbb4926a6df62b509b8f2dac28a587b51d357b1b7fe178b405d80b3bfbb1fffb3a0200804f7dfafd4c629;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d8008cc7f6bba1347f7775b741e49f973220c047d284928a5793ce5f931908ed6399fa2a22263a560d7eed0e5259146e171a19510ebed8c5348e20d1db68633b8d2c4d60e5104430ed01cbcaa07b43abc832b9b69e7db0115db93cb31b2edcd1f21594bdb325d5b0f391b03842fd89fa27a9a24b126d4fd6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3d10de32a08c5c599c419d8efdf5167d1df757b0b759f2d4ace9906f5dbbe85f93896122d2c92870a9bf651749900028c66f54aa17bf4a2749b0da388502307fb5cb1967840b98431574f9c9c106d685c49ed4fb29fa2f2af22b535269f8bfd327718ad5bdf14d240f123f41c3872ee08a55d10264bb1136;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hde3ffa56934f624ff395859df31417bd9c81a3531ddee3c90629f80629fccc7095c981afc7625f85ae2436f387a1af713edec0a94d39f574b9624aa78b4d170fa45ee3c46d8c7cf48faf3f9e925526543714167f33da35337053ea3bcbced3e22d88a1faf202221d749406b8a25d638790e9b0b6c44cb80a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17972490b4919adda18c7692a9a5a058c7bb5c2613afaa50ab84147e8467a9eed4811df1da5bb6769b6fb84ddbbcfa6dc306b53719cfdff06de188da51ab053f5f62ca8ba417f7e0eb52f7396c8e07b4279bed6833f2ae3a78d2e3e1d69f45c11d10d9f169539a0b72fb652627d277d6e2f7df4e05c02b39b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h69e6e666854328572e7839296afb5d0b3c8de5e606cba661f58c8c1d301f586664107f70a7070034de93ebd5d598cfc0588a43bea2e505e6e0862a49429fd4943c1b2d54d2fa557adac3b80a1b25b1654f6fb9db1581f4af6d9f418a70958202050718624913ae9f2c3681842a76cddbb9f7c30dd02b5190;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1950843d64a811458685a5dc96f2fbb04c88dee97a226e510b34125346d49bd1bd135602266dd538d70f769c4188feff11f7d5a8f0c1543a5af811354086ab307aa9f083c60a71d71bbaa49d989359c1912e94a11333081c5c37abce3dd814b2f80665b146f01acc6c9d9f3acdbfc33e7b64f0f7c74199a85;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h155c68faf70f0dafc865b8a510d717f1194fc2dc910e386d42b9bb13eb12fb679be19585c9ff8064e78fc2de879fa1cf5c0d416e93c1f0ea4bd99a4bfec1d3e6c355cc01b0197f69dca32b1a2fa758ae3e6ad70909c2eae701e7ba0a5183a5a55f0edac2b18055581d7181fbecd309b5b38824e8d3a19937c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hebdab00e6c3702b4bcd1dfe5784a25cdb6b5b366c79886dc7c5202371459d1425362e1db340cac0b253f3e4f677f472002a103848584172c16755cb027f1f600e453fd7e11a5c645107205cc7cfe3489115501828b2a97b20b2895a8c50f3ad01e8ed9496f3d8e3278c84c4ea0c12867211ac31442658689;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2807ef45301a2bdd3b4fa067adce917bb7c81627540cb11b33513881fc445f32fb2c012a81b30556e4e7f1113effb90b0ccf0c9bb4539b863bf46b00a328e977429098adb2d803d0ec83e5a44f04f2ce924c99fefca2551fc9c9e92c11e1145c51f020fbee06f91aea26de3e9f512d3dc66bccd9b5b111cf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17b465c6874540caff8510bf79f6061535c32a1e7781af4cd7d7de70c02c64dd9195b102f9ca4d079e8a5614d1827241fc5cacd6f7b435f98a3463cc4f937ece1d79c9b28db5a1dbff2b241c9422a6a8a6649f7ce39582d4745b770538ba7c785e380da31f605089a429fd9256393f26fcfed98d32f42ffc9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb4f5732f986054ab0b25dab5ca633aff450890510c2bb58159e5e9017ce88a0e2c2f475ee612cd442e6f5f5fcda296ef1cd75857af50759eb697b547909daca2235bfa3d447f264181f3539e3d8913674467f703eb25961234fb656738bf90de7c529a843bfd15a9024c54ed00ba3c4a9ec626639c5821d2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc9a1b722bc3d3728b39aad2b9371b06a1ec34279310d3e42b631ba821252c74e4504e1797ce8bb6d880dbb172d8ba2ddba8e81e150965a3cb5be3cc60d7bb4b72a8986c9e468b62f619d5703d1d38cbe3732c9e1414ce6bbca136ca6ce9e626c141e9f68c108a229b5e20bb7fc15db6ad53e52fa42d2d1d6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d810dc422eb58e704a2852df2a312c63c159193480e23a4b23ab6d5b8519a631d9df0a35202d2f6bda2b45d1baf7a629a149a2a50d39d92bcb32bd2ae4941b1612c7be16670463ed46f67bb574095f4d2e3e92105cf69bb7acb41e489601e59eceecd06d8dadb1cbabcf969d39aa9a6f2e99006635a3fce6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b127d3ec0193bf1b08613f21219bd2b375d96a6f50e0eed4935bcf4f84655f60bd56b9b4d5350f226989e0449aac8e00bac5cd2c06eb9250532ec4b898ad5ef4571c384410320a4d6a246977e03bd2497fb832f38945726eea84d965565e8ac1d68468c93fd316613c9bf3171026141862ebc3a5f9f5d11;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcfa8decf901da057ccd1778acba2a773a551541599e812116a440183cf2a27091e31a441e1397b4fa09fa37d5149607d5452e0a371a3f3e19b12093506c83a0c6e4933a9aeaefea686744d2261b4fbc40c1c144d0d3f6086b754320b1388d0da8d54967fe4084d9e0ca69a5bd1d05aec8692285550321844;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1695b0161a41b586c1919fed83e61b8c1ec388312d50a17bd7b925734c252f5f909040be0be1351ba6b47732961e917acede74f653a8c18f25d32b98b86e249e4794bb64dee2eb4ac37991b04aaf83426ef93438123374e4911dea998b34db46011ba593b8739012a5c93f904c8937eb408135d1e70cbade8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b5a6ff9e85947c225d7d5ac76ac4d3ac75dfe0c82f2780a02900de873bc4dc47f975e0d4ef969b5fad50d861abf4727371dbcc59c68d986cb295dd970eeec83a34232e623fa426edfd585233cbff94feef8029b133da091f419fd6356504659d0660bb627377c3ee5f0163a94bb36eadbb9fda061f2a80ee;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h132d9fb26dcce6cc2b13e2184888445c778f6608e0b4e220e737572bab5bf10f986a952cc6b0aa478ced8cacec29d215a2111956c246cc9edbd62e8d77f0c5763f89b76681b1553f81b3b8f2ce78ff26f770a08b4499479e994672f0ad3c8f6d2402ae975ebbfdd11a10af563dd41d96cf194665d28346822;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12fd2ddaa698226e5b2708f27f8167ee6ea780dbef7eb94bd4754e7f35f672ec0909ebec2f8fee70b5ee9ff391e67dea785dd1337f6fa8dc26173e34515c2bfaeedda660a915ab871e104296bdea183cfe3858a08bb72a89eadeaf708c0b19720121846e80e62906fffac703a687d31bb5a0ac6c8da358193;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ed2da0c41793ac6a6e06102b4d41192306532275c47669f63f3db38c753aaf28274877b4e9466b61b27a016a3443fc08614dce4adde67f596c0dba9fc7662f9b40d6cb1e9deb79ff27dceaf27f46cdd0a640c15171ee218487aa88ab6ef501d5472074ea8ca7ef5cd51f25da28044fbe11da394e155a68aa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d2fccf197bf8f56c0fd2c362ee87525a42a386d26fe9333603872388172bb2a5c681c392d265eff2252034a59c557221220310d505f638b07ba6fcbe05bb26c37268b2a6a0337e80e93e3dfbb14714222bd8dcad866a8ba7d6e1070610133469c5dc01d00b32d581a13527ec64bc0ca2712f9a78d35b1400;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13b806fbb291ed46260de193492e62d55251cb65784afd02460795a00dae7cad372567f957fa51b6375bdf4f8823586758fdafdc82b5ea45ce276d21de802f6277d4a5ee44616c57e2a2556765645aa388d462e7c760a359b0417f89a8fa756fe0e67ae1c8413620c124099cb91e064139b4c8a80f6b7f7bd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a4b00ba18a89baa06294caf2a4bddf0f0962b39e025daa329f14b66022d3d666a7ab06822b4d302892c71423478b14989401b3b2efd45f8cc0ba00daa7f6a8032b1496888d0b73a53d160ed120bff7863f2414af479157f992dfc930cb386cbbcd7fa2195734cc61df64127983ddaac6dbdaa9bbacce1d32;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h289ed963f032511e3df42c97185c5f3bc9793616077ada64a5578c7b54ae56e1edaecc6352d600b36d74a6fc91e22096c088a31666e1457e7e3da5a9f40c6fceb8a27af0f6ce36429457ca1fb3a6903e95b59d396d43ff61d099dfeae59b96065f0559260f2f984bcf82aac644381097efb914993abb9a13;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he8b8471cc55a00d398ea9b7106fd362735768339270ac35862207ee73bb8ae7a49215839e59f02487c08c0467d18a2383bbd06d76fa7f6e84f73574061394e15fa321c36555212b81b2fccb93912188cc3ecce4b92ca8b3ad8121240475af6f99f01cf839ce394a89f015b0101e4b4711ec79c5424dfdc1f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a51106241883f73950b850e9586c93cb4a7acb94f4806477bb763f7f79dde2d823eb42113a1005633fa7d3a32ab1cbcacd1a80d9a18b9cf734fdb6fd8989791ce9de104513aaad35a75a8d27e28801659ce10c81f505c45f4745d3a304392f7d8c042141ec2f0e1c9b6eb121e61e64b33844f803a375d79d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17e1dfb9280bb964bec20104eb50d3299ce1547aa0c566deffa9c0b7e7186585cc110e95e1bbb389095b66e65a1a7da6de332f0cb32e99bfa40390183f2047f966123cea8c69653b5910034f0d5f5f4d52b5b00984471c4f308d48a00a0c97e0c60bd9fa3ff4b62f2af9bd07b06f818f8250ac03ad783b6d5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a5bc69111b9588024428c9552ac9bc09ab5b9501503ca267136955bd960002d0424c0f5f772758dc0e9fa0ec833d780967be31fb9b5ba117da19cc52e8a435c80b4dfad456a4f69a972eeae846a5b0014cf9fbbe3c64dd2219bf304b5ad3338e3ac3ad821c3af71373be0acbed2d4f275e4afd1326e4ba52;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h150d7338d3eb9e1535cfbeb8c6d0d62e238455f2f26fb6c1a4c837411028bdc01d8024f75677717398732079274fda857b1a5bbfddbd7b0d7fbf31772878c6c01d398863bc4c24c56f812b443f3e49b2c131e4cb602713cf61a65f75c8e907c2b4d46822ddc9594cf22a8c3e30e3640cea0b836b3f9675b75;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13cc9ff87b12ffadace950db89f5bc921d9a5db38f08a3573e622a5d450cb56833ca7627c4b1917a6df3e0d9fcaef31d985d042ad45f879c31d8ca1ec67ecf03c7547443f2fa3c88828f8264887166881b08d163e7c6c8836d45d33090a0fe37925f85ff746ebe4fe4c91cc3ec1c5c304f8ff3aac817f90ef;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bb686700c33578bcbc491516def47fd03a96c86874ef3743fc02d24d68eca7eaa0f3a3639ec04665aa678dbccda9df7112692712ed24a6e52b09874785d046898d441758ac8c492917ea82fd2e4f2c89b332d6988878a0fc69ceec570c699f4ddcdd67d9ced5575cd54bc15e168eba81112dcb3cafe57e9a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf8641e54684b2cc56045fe72c3878e715e14bbc1119ac1f659ae5231b860d749530734080197f9d4c59c0ed862628f46ec0244b8b18f831e9729ff3c5e75d0c433d75c39b4e0cb650a94b8d95b9c66002fda573c55ef483cd8b4d214faec2d8c13419eeb97e868e3012bc17a1314d8fe1bb34256cb5f9bbb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6aa86e3bfa441cf2b80b598960d54f896f85d20ee91ad7ed3961d20e0d498779d28fa7187a60bd3f13408dc7f2b724b29e1ed838eea516d8e23717fe764dcc02be212d58e585fe86aca9833df7204b5a001ef922983c06c1b0099acb9a2fe3c178f2ff4dc5605757afad18481c576140ea517a2c3c9c85b2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h22d24a89c359c8335844c76dedd72c64d9bdf80f586e8ad98ad2e000ed100f9dc31d89d4a23a4f1d52a79a805daf5f9ac646459f3b31718dc75de1385eeb6811078771c90b344109d93296e2d4638dc78b637e489919e594d9a6e7c9a872ca77e80d8144142052b18ff6f4175ffd7e3a396f15803ab3295b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11e140b3dcb281dad42df2a053db307807a314f942aeb5ec8edb3eb78111deccb07d994b3da5663de7ecdfaa4bcd7c030d65116fce426c16a22758a7229556460f6217af8a793030d819d48b29536bd0d649e7a1e70070b2fa44fbea8b05995f749bfd4eb3808157771551e9a18b8b96427e44f7c1972fc98;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16e6ae3d4ab7f4d734eea6e347402394daa8710392641f32e285f9ce57b944a3e11b13f29087a92e12d44ee5abf6813bf47875e499373d3c403ab4954c92ed6fec09caf0ddedae657f03b1faaf9cc92fb65c786ef2fe778eb1f653c7ea8237528c083afdf88910f24f0cacf8dd3408b13a9711f0a2ef26b96;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb6b85fd4f36b625b37442cdaa1c74bacb4eed85fdc2c1bde0dac564da05b5f3ce7c369e5575a26879fdd903b0d09ea0a40d137ff5ca1d45b442dc572614b8f4cb35797a2d731c73e0fa7252f565e2311e2d43ca540b447efb07cfc5827888246fdb0dcdf0cb0429d2079b41d55259bb81263b77d35bb6071;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha0ad3a9c94edcb1d5a611cd896b03d4169570f6711416f0c3cff05d7f0feeab9930c325c1eec469e23ee204293be531517cee652159b54ba836bc3b8d57bc52d4480b69135c1af8fc6ef9e8c907f809dd5ce03bffd254681e427efbe486988efa47764fd3dc2fea207d821d1288b9d4b51f59255aafc8e3f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fde42a89b385e7b1df599246cc448769fc1e082462259cd61aad38c687d6182a5300f2deaf202b6a6787df7f984af8ac2eed89dc64de008d043c1f4ac7825a67b0275cd602800ab6d6e603b377f7b0c60ad4d069cf57081b32b8302b23f00e10a53f38a56534022825e780ce98365c94c1384bfe12a547e3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4d9c7929e5e4566dc2d5a07fad129f741998ca3f07f0d79688f0409db02a2b2222b8bbc3e04a505f94a64d69a7cf1dcf156ec59ea81a565abc054146c13d5a0c40f5939077784c213f264789c8fdd63cf7b31c74f9fdd4f1ef5bf5986c850191d33c7fca0e93225258df7166678adcc1bcd7dd2716bb5585;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fd6131f9cd909ffc83142b9eee7c25c3d64c217e57931b4537e5cdc5280abac62c54efd2d1f368834955e75fd34f5dd6fbfab98cbf4a137aa9210a2718383f28749b96d5ea8ffd59c9543014576cf1ca7d6c73d4b2f7f03549bedf942568a1e501295b878b220ec535ae1fe9eba9f9c5fbda06d696a0341e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1129c366916c79aa20b19029c5226feadb21de70275f50b7ca679f002a5f5dab4aa62c7ddf9d2698d1dcdb6946edd745849b433f16941db6119340367c67de9a18191d3b5742a9dd6e8022c84ee83ea6e1685ee78d8ad174f22e8546f6978135692a8d20f8ab44e1af2213561a407644e989b9addaa9454c3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h57f7919e411c2299b134d371873964de4788a603d7be514f8290a64ec4afab9759f8e43bc5b7d5375f2dfc9d34ed6ad47cb2fb6f9353f22e7cbf9f4a2c4dd012d2d2e392476675c36099f338e853cce1357cc2a3cbf3533fd1a614dcbb5bfa5bd9e0b7721fb6fad8e5dd18df5dbd0b740781f9e34fd987ff;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha5be1f382944ab47b1b38b497ce95546bfb4cc8d3c3bfa7ddc214c4d52d67b8209fff55d2a615b37559bf62a63460a9d183b17199b1d72d106b3fe090665b1e421452a1cfd19d80cbd88569d5bfb7bcc90f0a0ed90606f0ee01229275b484e9468a2dde2a1f52a87a1640ec34d4afd1953adb416a56c89d3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h58c251f86628cf29ba4c0a9970ba2ae6288231a72dbe3fb332f67f9a8ae0b0219a32c2336eea05a00c1f821b3f9fe7dc89e201b710c3df6439ca1d2e348f4c0fff4295348dac1122182392b3c94d9826b31382bdd9787f89de4598c03c33e501e09e295a08260c86f1a5df14782626b87a28929484b6b3ed;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h738aa36d11d905c8b4ed409522152a768b7bed82ee7f593d00e822b0f6d9ed29030c877ba80bdfe91e8a34ff19825444bf4b8e1bdec5478c0722da004c1eb83129db13a8c13edae5755cefed8758494d7d476e4cc00fdc1db512ecf22cbcc4514502480a4c5eb917269613f21aa56561920f86f764082b10;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc96be9a11009bbb657f35c8226b1526fedfcf97fa677941e1ebb68903a8cdbb5f6d91869c6a7c18eb6568ceb555c3779165d92dd3a2d131fbf4aa23df563d2efc5925bb7d6e2b477183a4787907af5125c9448b8fae6e0eb33c7929e10fceb875803b97b87d48f648a9e45a89a8d39f37b970ab8d089ea7c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a103633b785c5f658ca20a770ed9f690c505a0596b7be853e6f8e5ef592789869c63edc4186891200750db1ba322f6b1437bb03e8953944f648a2588eac4d06800daf4115c82f09cabe325a65806decb8c311566088d48e6774f390470dfd0e9fc8c673cf6c7149e1e4d43f6e7dfcd8afdd35ec6ff6090f9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbb451d8045e4e8b1502eb1499cd21ec6380097d58da4f754c4fed6ce6019bc4403658e86d87a4ba048ba8ef39046c45649c09f1ceb97a388ef23281a2b477412a2b000b5a544a2ffc108a12b7e407b4596eb16a2662c0dec79711c3493576d5967065204156b4da4d8d223c6e48e0ebe1229b9d81c4dccb1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbad7190b4e52c71c19f64cdbab30dadaee6a7d65945024dbf18dea83a9887d5fb0fe9daece894fb27744c86505904cb97183ec457ee816a716f87cb6feae7975dcd3f82d6629d397aa3783ac581e713f41712ff5ddb12c219e839f04285e62051330c3f53e7403c5061c0813f304dfae9246c03700686857;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c1d67783049820b84ab54afe9eaa9482888a4f935dbeb0bab5b5a1133394f848c8a24cdf005c46b3caf9bade7397ee8cbb54e833e3f3201e4bf35e43f170f78bd6bd61d345abc18dd0011535a1ffeb3b3c276669493ce3a143426a6e5186776fd924de9180a94d456548765388dbb1abd16148e633e2955a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b7334f3d0fc8f43bd71dc61710407ee99bb195547f549354da04f6f801fe4765ba5eeca6cc51c3dc52ea8d5b98d80f282240c939b06440a17570e666f2eba1e39c6e9967db3441d152bc1516952e3f721b91435e2a6d174c088f006a8d3d5dfcbc69e675962f2ab5bed9e271e9131f138e870c46beb5f3d4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1450b565a3abc5992903595831e5d89d21d6c303d261297c892f1789ccd763be4131d0885e0db496dce9104ff483ea5f6fc451dd4b9a5d225e2e1f23dedfda5ecf85645475a62aaf788ce80920074fc947eadf02e2c97c6be5656da82732cf3b769a2f6e0c7a7c0d8b61efbc2bc9b897d32ba68c3cd3b39d0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12921bdeb65cd653ae81c95c13a8a71484271cc5c88b9ed41da45b334a898c702b1889e4f44d36cab2f5896dbe05cfe59ca343577ef395b67f5fd4fea78ca07a154da240bb90d61ca45126edb95e2d292ae8ea72c48e2872c55b7d05bea1f0533eb9c074af5a433c6902cd18d516fce8474e0f4a91c5da2eb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdbc05400017b695373356b865b2ddff5d1c8bfe52f8b0abe430b335683ee2edbc12979fea1c7d9caf73db67dfbd3a37457a7fe1795fad5c99b57913d0ab68cce94dc0df679b9c28fc7e2fd81bbce93f0ed9b515faaf858efb0440a0504a4bc6312fe6c4950f565c103a24a3ed1bd9441db7e3d7c925627ac;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdd1272987b90f0eafaf528102b5b7114048f288f897c3702cc47784bf6fee7fbb947e8cda04660527581583952a4a39d7873b3efb1b4508befa780dad63d94234da937532f905f99c7a079de25b5a979f891dbc4ffe11e8a650d677de9b7f941fdc6b3a5c561ab733be55084314c589931d0fbd27621f046;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1968c31fbf5d2a6c40c9f5b5ffb6863a7e7d6fa097fe67835afb337a58d73ede74aec3310539c5b333afede5b437e10ecfaf0f1a70db051f9113c90f5b0cd76d0250bf408bf3dd75689e82b5b7e6e1bf08c23db8ea712c75efc154b9bd52155f0c94f95d60620a00325f6b3213fd61008b6dd917d457272b1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3db52b50decde31e7c46ff2fdcb96a3c93856fd0a4d0f52136e527f788ebd35487da925c90bc20748824e7599de06d6cebdf12900edf9e6a2797208994ea760e7b1f5fe282c6023827ffe4a891e3524ce75e409b4bf6a8d5dfa27c5d0236cfb4b975b2341cd945b12eb353ba6dc7d8d93e4b3200f92e8051;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c8dd1d4249c31a6cf949e7a9faf84a92d6b90b086de74cec86726c396947f2c157b4df8cf52bf52f1fd59f4afe73e82a45197e78b8001ab8451abce41154bfa6d4b41fdeb5a349b0da2e0aeda45efd66c49ab00cca6cd3486dcdfd3f0d66ba69161ab1a2cd6c13aadb625f71bcf557a144e601ae3986fdf0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h41c90355bf6c1495caf49e5fb0ead759709f16094a9e631388fc580b0ce164e42769ab21662892f0e99c2db7eb35a56f979d929e5fc4df05f15449e60e86099609bb711ce28611d7c612eee0781e96151c83a9aca7b30e4be2f44ae24b758ffd5ea005201ee49eeecfe081f81084ea02a4bf874c7930593c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19fb851abf2e70e9bf6e5191a4ce4b5fed95c3d474ccdc747d2c245fcc23f983c3e9d3335a8b7ef974e1b08319aee4d392d45c329687ad14e991ade7811926e127ff954a74c98990dbf174fbceb0a7569fbb14340331c29ef7a960aef1fd1f505dbd32d9003191c822f9c681beb31006830a6e19886f408aa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h529860af49c38a7e8780abfe3dd8ff649f1528a22b126c2c48163bbdfac2d8fec74cd174701072f6717c41b8023001338b9486e7b97fe67aa4221125b790503d90d96ee2108d3cb046c8650aed0f62c219185f892013b2b96e0e514b03be520f0f1c26930a62675a9b4ad508ef249cab3c68e0fec2232732;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1163b552b6b908e6fabaa03e46f788df126b496c523e4a7d1d725bdb4ff86ec1806d2793edbef14dda6273f11f8e770dd797f24095c85ffdf5f8337a56a052c90b4d19c41ee9f474acefc471fe216d0ee98e05fd48b94ec983d6570e9455337421984f822193c3d9661a9a181e5a5177ea532835d8585b7ae;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ee655c78134d6f5a970d38154bddf8240c6ff435d62196246f5131d981500326dbf32d0c211ecf93570ec8bdde27b155b53746f6139df23692821cbd12d997c7341685f1077aa226e3ded82e7f44f5854b30f90c20cec7a6613be6fe40c2ac39545d37e33dca484d372111a05a1b34bde031ccc16e1ae250;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1afa46e263dccf31ab137f7a1748a242a17ee41f479b6a5faf6afb6d72fde30c1c0b7520ff0f0ef8445a94f56393e05abc39616b214e13ccd3d4ee8308272b98c46b5377d8ffbdb250d4bf5c6536d64b734df57ebd55be5307ab21c129e8f44378c229f2af9f5273e979676f6bf764a617ffbba35ee340790;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h117cf94dfea4374aad264edf64d5cdfc6a243f6a04ccc6d2345d8874c67c8e6b9855e97ec6303724f42c522bea18273de12d67820b74412ce43be1f218eb841f627acc0d46e02b45ceb98e7938708af1f3fe2efe4d4eb391ad5a05f6cd3bc81a6645595a15df74f3d4c81f37a3bbc96b1c57155b598606571;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bb108b9f4dd27b6d79b82d31ea70828efdf2ca76a65b88054990e3e4ea758fc3e8dda1b72fdec08f82e8af84878d124f307d2b8f2be883c17e0cc7aa5a8a3aca5facc206e1b92450eb4f0cdab0b3dd4f7911796a5b398b3ecb4340c7e8e786342940efe745c617b8c752f69c4ae0396952d8955ff5b48039;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15f636fc39171e3c32a25e886989a29af059b47a721b50098d1e39cb87df99bf073798f87f572e637f760fa60f1d8880f7fc7b906890dfcc0971c8b2288662e0adc1e85cf56956f3ee29fcd7d15db492e2478ee20c458628f26b478d2bc4f558f5e3afca56a3ed7705a58dff8be8e07966d005225d81b1ba9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a563dcd8e5a2304c24123f1a077c70e24a1a8c80e81fbcbe2a39ff50765ef6e1ce7c5c5f937045db0e742740260d9fc57f879e00d6eff2a3138635b10752e44083237804909a4366994d38627fe8041c6171caa46ecbe5d38aacdd5e8295df8052a2990b3ec6aa93864da159c344cd50728746fc5c331a58;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b088f6c50c402672e5ef014fef6aca7318c4e89dc6104e9a540a44e16e410a5b3aaeaf04e74bca6ecf07493ad2f6456b87f41854f834da9df4bc91d2902cd2d22d17379918fc41c9040503014053e84d70680ea671e1bf676d7f16707efc0564a08b243fcaff4e7af9aec610b3388253367f0b416c38b0a8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1518e79b65b4f8a6f2d6e69b70213c0a25d61a3909fc2744fbe9cfc751b704544b22ffdd8c6f91f5510d938ad6e73a520bce9acef2e120795f59c684e312b6e81be163be6c4b0a4085fff7abd0b258bca47b258914fb73e93140539a2446d4f3b5c15a3e34f7110e818a13b9d8b77e6fd94574476528c797;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11522b267a3857699c654d3ef54a6cc8e850531534886696cab27947e77fc078eec4fc3494bcd9956b3f2834433476271d1bb28d4151d17ea25713c9d7e540f4ecc642a104bec41129888dffe188a5e1818ce2cbbb9e175354c5bd8aebf51f3395bac09e5809808da882ac8c9a13c61528a1bb6fb3014a3ef;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15e1320977e985aaf72f08f5ad2006998ac8c2903ed3324e9cdd42e8c39a5a4b7cccba6d8af0e2bf436a6fa9766dcf037cc9c11d78d286f59efa96064b472dde71b19e13e5be543fb51fc5af064ca3ffcb926ab6aae28b086231a53ca252994a97899742c99e0a4ede1bf9580700d4ff877512a41d0d977b3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbcc469e4b492587ad7f78f149ff07230fe9fd4dbb3ae4babc4ce0831aba1f56fab6374b66e3c3b633d1b72b874e7953f1cecdde2e22ccef1173caa82b2259a51a7512e79e99f67a10978d613116fe8446caee3ae4575f6e02fa99ed3ecce4ec003c8545a2e1125ae1315e0f6e67918ca314147d9cb464d2a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h60bc843397137b9d5bfa1137557262bc3aafadd38f0f8f7db48993a32c3632206a981f7b33f3d5d6456d442cbf4918bc51f8e0ddf0bcf93312ff045d4d59c25dca71c3ef7e94cc0bbf07e3578e49e7a6aed4948d6f42e5044720a7659a89908b9910949cd2d1d4939e8f672d62138edc5ca3c35587f6a6f0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cb7c69e02c93a4c69ba12dbb008e2f162c3639af55eab165bfa3c428999aaec2a03fbe8cbc8a27e0f8c8e51b8e0f1ce5a0244088635339ccfc95d50d8fe156587f9b25caac6d1bde574fe688cc2d2622a350c6076c54840ec3700c1d65503de75c5add442dc9f9a5b7bb7e0f7af128e570f61be3c5b47ee2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10c71881f69c9ea23497f83bedf5111983ce8f11aa510cd3690c6cdcfa1ca8f65b6fc675656f1c7be4b3bcc8fa1718c0de6681fecaae57040009f28ee1133fd5587da487751caca04683206f43cae7568509b821012d5721cb11ca513c1300123e5ac65548fccca1318068f8280b534b54dac9339d1910e0d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f2d659466aa9400afafe503cdedc4a8dd2048cc872f251ab37dd2a3351594e88b82406fae47b042283659f32cf3a33b98f608f546121398620320ec2f4f4e48ca7cc3630b3db945bdcd6b8654b59c165e1c9874106d5abcf03d2b0fa870bfe8fc176d0a00c864ec122ff79acf15e75e15440f3fe982538d1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h27cb4807a1b73cfbfa9141332d06f6ea4488b830327907b63ac7b4e10fdbece817dd7d088b56e5af702330e27013a95616cfd96af643bcb220b1d85b26cfe24c5e6af3549a94aa7e01d0860b39d0f14cb552d7192dc5fd2667c35357f20196eca535bc6a0a583726d828c05ad390f449df45215b32628f40;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13c29ee8092a9f83959793dcf6814b5684178a7c081f7ae9da5d7e236a45ec658b3ea8ab217cb0e69390794c6750ddee9fe6384ee760197f02e341e1c295e3d374520cd119ad2c1ec78481ef2262fc2258684464f6c9c732ca4019f4ff6d73b64d2494836c9e8a9294e32f74aca498d91e8a6155f02734b3b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e8ded002114b9fefedeb58ea2def7093b9ea008f5b7f5dc7c63d7f0f885b48dc46b1445f0f1248c7d49df8d16a92fc767af6b9790c394125ffabbcb76ea9205b8ceff312dee2ab721a18f251c3f3d9d7c653ba3f2c755b4633dd33fe80094106c4e929f698244047de19d517d73ec2ec2a7dfd96f795d289;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3022f5281bc7ec4261398c25a8c9f58fa17bad8ab1dc5fbf536207c9427aae04de12c5cd8e99059b9c22ff035f52006cb8d27345faf1ce2b9c600f18b760d7586ff68fc23900390923c05be57042c0a2ecf227282204ce3c5b65e35b57cf3b8da1d8d20b81ce2ed5f9b54f29fefe96fb3960ce4617e9b5d2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10473bd77e2e60004a865889de2922c587069bd7878f1e6095e8413984c1a0c7981497918531f5fe8c70055ad52828b97ee7eea67e537a54b9743b997d322df12fbdfdaef004a4334f952533c2a3f037b2792d8e06b423d78192984d7ad1ab3994fd45c611a061c29afe491470884c2a426c1c48196fe919c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7d6e83ffc8ae98b986bf6432012dc1a61c34a2649d0d56d023b84f7e9805723e47e06abb80e54fe9e113d02c70c047462ad68361b94dcf1010dae943f2adc03caf2669779e25ecc93266b079f2daa8980ecde3f363e9dd5e2157874c80409935e6c0ec92c31b119deda6b4a18c41cebc44aba220157588f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18d18499b76cb5291eda3ccf8c3cabd503343fd70d88fe9ee04c551fad1223d8541d65a8c5a047ff25a2bf172629b6f44a9d055df1968b906b718f59f23ab9a572c3e1a1df70b62cca0c20ee928471d2345e7c1e48b7eb3ab07215ffc7fd0426ba7c41e6f3d451bbae7b519ad05d821a22510ab083b7eeb3e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13d5362596896b50809c4c6e42ab34c2dc4c323647fb8f4f7a095e5be60da80f3d00e98e05e6489b4bccc1af971e56f19006a051438e3d7dde5710c7386afbdf4f538001a6e6ee513eb3c8787ef39a490657b88d5a4a8a86ca6c3646066f268533c6655496c6aa747e1358366fd9a5576fda1373903a9c0d7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h20449e0158fd8d1ad0b9f04ad29c2a8df3b7c4fa73c391b6555739436088479730883d76d29ba4a1a731c5dac4d04789c444343dca174c5e1ccdc09c95b91846e1d6dc6217655ab18a4dbe4d7be28201247aa00a83fb814cd7795371d8d741b9f1e6a9cb79183395d327690e3b98c5d5e9edf1ab1144488a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he842d855ecdb421cb3612b265cd8e38cba248adbb1e928aa956a30c5855a1189413ffa9e2c5d55746d1ee0194c931fba2eca1865019b4c0418c3b30f27bb8fb48d119facf82aadb98e5ad60d898f06fd0f3b0b4d5d59c18caa3c970acad0ee27214c1bac02306ca4e38871ddc4c19625339b854fad251195;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a1db610f7dd3d056b2c0bd99a5345fe1b08e8d0a5e786f03ba123324f3c93a12246c82033a9c02a8bab434be204f898b716eb3d438f39fc46de549213e2226f692837ebe970dc13caddf6a635402c52ffd3f07d37f7c56ce42be9b953f376dfdf4a2893573deffccb716b9bf6e89225383b61363f17e61c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha8d03236b92ee79587fcffbc0c56865f37d10ac47d2238addad9602a96c118f6d6bf4e1d1d76d9efb8657bc26df3cd144e84061bb224b3fd89d7b66e1ba5143e15567ff6265c37ad201c4f454d3f8500a0dfbf7fa938ca4471edf1862a99a1eaf84d492f9e65744b4166a8f3a637d4cc6456ae0aa43756d6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1722ebf6014bd03ea2f23fcef83924a2a9ff7e1c9de77ed746cfa6cfe617884519a2a294f334bc8ace05e7c00897311e66e5d03b29d73e2bd4577b613bab58d637041f4c5325a4c372bb75fb11640b58f34407a5900983a2e41737a9eb9384d5d0ede10a7ef8abdf8859fd8bf368b61aa4a110546af0ee7ed;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h41c7a5690c856ff3e28eb4677842b79ec758ee3c358b54aebc19a13c8e96b4de62b74be17bdc70e698e7572c2b56b9d822c70d9353cfff7e2c29b116c17be4a2b82703b4962d8aa94681f488ad75874195b1f8644ecdcb0bab9608b08834c617f0b3995e22167d53d781e1962f95320dcee9ceee9c4ecd5b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10d043e0de91f4443e56136bcfe0de2a9ce36a1454a95610330665e94c1fb8fc42466657bd64dd2979ce8e76ff818c0f62dbfa4c2a7d78ab2777edcf19fe30b021f867477f22961ce87cd6c587482aed2c1c11363d0a0e6c8a15eccc96f88614c49e82cdfcc77fb525e0753737bbd2d3c8ac9d61cd4c9e056;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c6def02596ead3615fcc6be48ccdeaa03f58a11d260325cbff30f357dce2cb0540a36314d9ddd3fd6dfdb744980b8d79d9c1f00c4694554c9396cc0df5f0ab85d8f35f105b506ebcc766755886b00dc71a810ec879a85e41260938160aa11adcb7d5441be252363c5ef07dfdbb24a5aa7a9d105d6c6b71b6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16f10d013746c3c3dbd57ced566447632fddbcbb1a3c3a70ed8326a5a2a32617e0f0fbb18c037fc2e29159c32a4d7049f19a08970e754fc7863e6cc032a0d2b67a7402b66c4ec2ef915d0f93d6ae1841ab9fe02fa4120d755d78a8b89f4bf07dc2e694e172c6d5b40dcc9b6f3a2d5f85d587cd8fca87693c2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc74a0d4ce6a595c62c58ab0a3ab50ec83c52d3e7f3a8698af0c3af4e455b0f5814b262d47c12333cbdb911a8a6d857db5df0cff773aae1fd613674216f85ece64f69f7704072963e5c0787dd41cb0915b34ee8c2c907a3480572687b43937289a0162ae83f170d9b191553cbd7b734fd320896cb5f0a9e5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6bc08c78a66691c0f9772798f010050588a93be2817538c6397d3f714dc6b3533373e2b8779527752249407927346c723f6f3ce8fd1aa39cc5310af0ca19118d3caa295e9155464e7b293589c3432f7f606a9a0a079b3588a918adc9e105fdda6417064114808317b226dd2bc7c8805ab107217b066d234c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h34fa7c6b116322e3ba9913298a8a469d57d7673a3def4c93ae8e7342fcd1cb19dacb3befbdcc1f0b7f6b10878c671414354320e29cedd091fc49d696d8f3965d54339e627d31ff9e4ef3dba8b6f23b6e1d148779699f3c639a9f5c14d5dc002e14b8b7eb0ee18bdc75fb444c24079c2d0aabaa771bf0466a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he354d2e147e8551d2960391e7c539d5c738d6cce6f94ec7ce85cd24972ef98eb8a93559956b3b8e3c829ed21035404a285c9c0ea43e7e63e77370b098d253faddb3b58ffbdfe7c5a227bd2e1fd83da9698b1fbd82d79c56423fc66af6e36b3c0650f33f1ea5dde4d940b477fd3d2b2489920673e94c26830;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dc574acfa6387e6d7d1e34e47b5fabdebe2ed4022b35a9dd170f51f384f9677ce690e5de87570743006b4de313be7ad9124f604d4b1f70ac9f7bb2c64da87e599132e00e03012d5ac13fc4937c17340707963b862f563f031afb1b800d42441a38ed0e76a08455353d95d882904610d812aecc3b92e652e0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fa41352a38be027147eac97c9a389ac422115b8e10d227beb8fc8fa78cdbc42fa1be152629586c9fd7a2da2d4152613e090b0ddf7aebcac9e3ba777227a77e2327a62d14dd2fe983f8725e8c503c04313dbdbb17da75dfdf4974e8eeaea3aba4f38fa4287ef56893cb633d0e85d6d7b25c369a00888c5542;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h22f10fc4342a72e04077884e49725ba7379613abc2c31adf3a0713aa86beef3a79443ec94fca7b737c044ca900fd74d676793e34644ac3a7feef217e76f3a855a098a7731418d0ed577d396610805c45d1aa3235f687249eb877c316d1d5758901559692e34391b67fa6cf26783c8e5eb506d059cbb4ad92;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1664c26b6e425ff42b3a71097251ae1552417fdf546eff5f9104cac23d800b8ef8d69c1e3a1bfd2c10acd6bc14fd5d088dacc8f9d3515abdfbce44fd3b22d72c59d96961695afd81ad5d76116bc0393237cb1c9cb3cdc09ad2d2e74a8177ef5d59f3f70b79ef154ba8e6169fb1baa6f649a749685df031954;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf280020590a2f633e4fb58faff0aa0e66dcfe87f5d4954d0afba8867855059a43c35b8a96ddc7baaa18cb2634a87da292f63695211f3ca34467d3b39d218a7874f9f3430cafaf33ec8697eb35e8c3635468f9498cc83cf06d6a771e0711864b0f2e173d9e9a09992d15ea535bd60b70a9437ea980ebff67b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h793ed1dca73b195fcf5f36435ddb544f70f741a6ef944d7670d58fa017dadcf293844147bb5bf5f75f46e210f5a3148caedcdb2bd35fa6ab46fac8b0ede2fe5d448b6bf3c4a20aa58ba37540ab16eb10969af567bb35a8697b3f52a17e209328658946025f9d618defe70d4c8ffe5b6b5fe7cb54b01b9b37;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h123e8b380d730f9aefd75e41620ae7c52dd1265b92d9c85669feefd9be0bf8ef9b84640a8a331f88165eb31a924e880e4cbedabb3546f9f60f715952740c57db0f4ebf61a1d7454d46ece1a5a1fa834d4f24437060fe81662bf2263bcd477da11d49cf624a990e383fcbae0ee971d411499ad16d078394bb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h561920136f2862d652f18da51f4db91ab3d5e10ee95c7e4b68fc5b9bb8de347339ffb64fa077c06bfe311c2abc559267496f649212b6f143e13e24dafbc5b087e234e145528a9804f4dd47fd94c8f6916c96b604d7d825d797eabb648692fae30178b1ddf1f6e62a3d09ac61a43a157eb8ec02b19c2047ba;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h385c0fafe35c2c8df0214944fd5929de1e4b0ec12955eae48681cc3b55db40f135b8f37e085c4ef035a0d62763a353d88f4c2d88c372463ae16936da091830862fa5b388a0120deab420e1989cdcae6afa03a88f7d79d413db47dffe1e3740294904bcbc80adadef1e00b878167ccc265f60a6075ab957b6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b696cb6572e928d62ebfe1a8099bc87045e9b604cc1a4e35ec6ba58503a47ddc778e2e5578efcaf422d4f763502418f1a66449dcedc84dbef40fe7af33664a42941c7272e36630cad033782e6d7aec8dafb157cc405324da148778f879ebe71ca9e6f2bee3cdd357fe2b8a2ac97fed7704ad5b29c72002db;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf9718297d162a5f6ba38c4967ac0c36c2ed37936929565f85846c9597b5e95a8477ba1cc71bc3cbc3343a922b88876024d0067b827c5ba814529d5ac67c2dec6ec6f106718e92479207b6826d30e59c6412aa9300db84e7d9087dbb6050f699c6eaf001bb96b83f366c97e8212acd75fb3a03f5c84272b88;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb0b74da6ebb9991331fa97ad5d61c7a697d24d9cdeb9a29a67f31756de91e8f61bbf2dadc11e3ef575d3d7c73bff9e7702ddb3c10a56379076f2410cdc28a0e97656a225516df81309369c7963039ac711ab74b9b2705ecbec55be5bdba971c2163bf133532cf89bf5c81c67141be6618a85518a4f44ed45;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h183cc736f8570522b96c0285c80fd3781c882b1f33dd282f0eea73641b1698b318334dc37afb5cde5c4fce0d39ece8151ba0ab91969330d2cb60dfba6e64f212895dbac221756099bda37fc49a17b095a04d1ce54c507a743e3fe002c6df2a460efbdbed19e346509238e840636de51fbf08176834cdc9e16;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3189f090edeb054da01b34402db5df771d31aec5caa9f226b32f5e0298b9560e532d8d757f45b5393a9c8fd4f619f8f9f0c4cfbe170aef7188643dd2bd2f72ff1c5271d3b2c5aa6dbeeeaa9f69a59d49ff77ccc323ebbdddf8de88c74ee1de82116d666da17b7d1a9b44f135d5554b5c2011f64f3e694d1a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h71f5cdf24dce5ede6ce178a51a97185f35ba5fcd07804dfc8cb88e8b62aa3e8a9b45a832667bd5adef91a8e9b672a9253498d939e246098f0d48513d243b2b3f955cf11aa3e1861317bef4f7cfad4e4a74f142577b40720cac3dfe6156b098f76ca7a9eb9aff343ce5075ee6c2b6ebdb3bad9330ccdc4371;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he09b2bbef6e596610528a1121f76c2291b93ef9ee032e912262cd389399acd881d9fafe97b2be831bde95c074acaeb683c14e5c4230e3db764e1df994eeb3f0a63b0a4173a4f8ef513fbad1da82741f130b518b6f2a974cdefa8e2e53c23ae02ce07d615d7565966a3629463559fddbc57bf44c48e0d4371;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17a72918c6435f66c163ded39dc3cceef56574de13a956aa4c85f4e1b0ff40a6eba4ef8b92b758c3782927560ccafdf82cff694613b0f6469281092ae72efe1398ed8184234f35729154f16bd6a7b5fbd0801664ab68bceaf182e94dc41def2a436119fcc1d77a496824283d4473a7d73545e925967aec608;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1003888a9fcc864c538fe39de977c81d485b60fb4646eddb4adf84aba6fc8a6229abb6aa3d7bccef387964dce8331b6a2c0eedef8135a12cb17881751231cea78b588733ce016ab5fcb56a1b5fdffcde6ec4e4762a7ea18406360ab4d28787a4080b9234534aa472f7642148cfece104c5dfeb80d26f8f2aa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h100d3c4a3e16ae1c83b9dda075cf4b2929c366551f468ba1cd01d8be075ab35ae966f7906fca80f745a94cf276510341461e38c0c150597f75c0118c07e15133e8c1b93046d9f54e55adc91ff40b055a2f2d172e54f2697b026d5cfb30b01efd2968a4b77cd7eec53296284f39af238dffc05d0860b5d09c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e88f467728aaf9d2cd61a9e5a67ce23fd9f77e4e734fa9df880f93fd48bd310fe2d6364fb32c11726f97ca95c25183d8c378a6e516bf1abe2aee2b435e5a088d5b7248798ae2f46f7a11157ee8ef64d8071be6cbd7e715175035011caba86f544fef1061708a430e7250a8608d0c6782cb080fc09e3521ec;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17de87314d14942e9b2933515c8ba94fc85ae494dbf6e5ff7be350e736e4d1d968aa95389b05130937e32c774d65a86e8875a6b620b19d820ffaad3778b9e027e678d9494a69f0f879d39f093d2942e4a72c14d085be96398eba573c74626a2d233b61b2ac6e3fe6738d6b0a158b8103b7f96f77ebb77b9a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6d118d608234522f9be6a1d30f082aff7895c1cae9c20f63a0a8bd4373f273f2d6146057f5e2a0e5d0b098618360e8d5f66d1ee0c816dc2ba4942ff02cf037e0d8acda0dc3604c2481717ef0e87d702ae481458cdcdc115b6e93fe28f5292f26e478c25afc626709d7372952c2ea6fed434e1b4cda71196a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he17cb6411e9708818d5bb1a452873ca991456fc232c9f9e9deb92c95733f692f73ac2154b3f5cdda9e55d339287ca771cb5b4808dcd96d64de37d5c7d897214d3c5bded05005099e0149eaabac2cfa58c4ea7f564e375d9d5b83eb7728b516620ab8264390da3da7a3ef157293e7bf88fcd566e013ba3fbd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11dd7ccbc352201057f74cae6571b68e75024434097a2bdf936222bf25a04f39105bdbd72f41300133a6ec5682a4a8a451d3e744413162430c41cc04343b3b65dd42f47c033aa27c03f168648e642e7ea6bcef2f1733682ba3c506d02a03daa739d6ea58024fa22a3c5cc412fb4f746fc69bba409f57af63f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he5ab99dfadea57268f3c777951880c102a0c630b5f994c7c9a5e479b176c9eeaa2450c49d4e2f87746a7036d6a779d52670719a79f491d234fc209ccc2168fd02662543892c7b0b9cc8bdd1705e177736e4ab6c5424ed70e34119d53060f52837a7b94765425ee76a001b5b1747b9273d3a9511f0a44d756;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1356725b9834ea4b52dda2fa1f28cc990d642d682cb834fc0c6c2f9f8ffdd354d056e65dba9290128e2922ed9bd8fc867e216fe64facbed1ebfc33cd109ff50cfbd63c8e223151f4b6c7e127c60b23eb1711969e83c1e5984f1e8c1cd7b2e29886725b30ffe4b620be6b26b45b7239dc6f1a8cd777a6d7bc6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h146a1db128f526ad003541848cadac4eec7fec7a79472ce1976b165708db4ff7b208f1089713fecce31d0ee4016a5bc49c8e9c6b33daf6918a33ce5e4db2c8578953beae030896757c17cd09f5e8070e3cfcfb264444561fb36de9e6bc4f15b42d78c3346282dfdedeba22f6b3909182628ad2d2977586553;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1851aa55a0db26672a2e96e6ff85e73e6d7cd33596e16c9111ced67df4c7ff61615ff8567974c857fd7f4fe6a3caf51b6c85ba9be42e2881c9d5449812ffceb2a0b3f088e89705e75c5a285ddcd1a96477eb2a313ea93ec7202a6e1668a5612cecdbc11685f90424d8aa9c1180e7e0a161d4736abacdbe39e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1773971410791a9234215321d56203b489b70473ebcf453156d2eb89a326a98d66b7c368cae7cd0d6d27d035d2b629c13a6862adc8210e522bab62006cc46ad99ad04e543ce419e5541509b02557ab6c24408d27adfea7172d3336971bde182a46f78d33076646f1a5d706d5d523a33df4d80f0b777b8771e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17ccc4803835326d9d81e7e8b71c12e819b6b224273d1c8128ff85d17b036e8d54923141c2d6f7060102bc80d43fda7d9f52b134919caa85284df95b7e8f18e99315f979e5dcd994bfebab8f2c0e43b26b3dceb3c39efbb0ae341e820e6d2d4880cd1014fd88b802811371b671024a6a58be1b38918371d6f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1293edb60d893d605358344553d97e6ce1bdf5bd3b8c0f776eba87f8b338dfd360bc9c2b048c95fd27c026f0044760a445ff6a732afcb0e9a563e594f180871177954a9be1da12bfbe75af465412ba7ee453e6555bc785f33416e9072cc81fe2e81f7d85c10a74ee384c3984bcabba2e2de047fb4d6394ad5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h185aec03f7826a0573963dccdca04e7b3d04ce1aec7b944920c12b281c6397cd8eec545230d1a7b1f7a824c8434baddef00e0498ec13fe1556b21eab2f6775c9a6cb1a5a87e738cdf7fbc0a24bf4975b05d489870a1db216e6e80f409594b086596b0956bb204c0c7d4e8f5d060e241e5f34b648551462b2f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14d856a36518a3feb34ee8936364e6700621f035836ba76c03154d2e513523b75e2cf33a629f914ebf350a56300bf4f7c5ed766ba8da3edc3fb781755919be26ad0b20a45563aebbd2ac600579cef09b20bf2765c9c76207a898cf1ebb0bef187285e74edd30cafd5fe1dff068d3c697b5ae044fb3ddbe9dd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6e499a738b9c1d90d423c244443dfe0a9c122cc3d453deb743abc72aff66313a4471fb7b1ee01d89da976f447b3a4b1d5c763d929955fc3c64b0ab537171a8ada5b3f5e22474d166dcd064c6ca036f87bb4a8778c5ec190b01b753bdaefc67aa6f669f94d5c5c947f246ec347442477739c60fc7f9378738;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h942b6986beda980f3c8a0c1b1aa920ed17eae481482b33d684c61cdd85c64e7fc3c1c0fc4a0ad891669f06c59b8b627bbb592b92571ccfe0e5f11ea16a1dd90419ef4ba5a16fd2b2f74f535d55a33a0a07166c69dbaf2412438306906c93858ee3c69321b1f0ac3bb8ffef658b368e93d3beac9565aca3da;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1842c3bdc6f782255fb44789a87178058d6e9b7b2a51866ade28958207e2ca88ad9c531cfc824b51a2bf2c00daad8b6651e14086d483556948759abf1c81454c0a8e846ad2f39dde3bc8dcca972d5e615b8465e004bd5fe9e7d43e7191871dce3f8e9f55a6c5e9c06d57c81ce0742e718900813782b2c8e13;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b571ce0b540e90cd46f9cc72a86b5ee0e7bf9f1e6b31c8d8954ee90e8af8f2b96dc559972c5f95812892defd772c985a78c94ee30398b3a9b42c3a3f4d972c05b7f258151aad5321376e51ce069c3c41c2ebf4e52dc90c1f1e857501a65a742b845f90d1f2806200e819afaac0c2db63034771ad9b2117fa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h137da76164badc49f5469abc47e6c114271f20411d3739353d42dccf2ef42e5cd69097267fa376f36cac863335a207d00d1547e3628e2c06f3a9ff4bd06c523dba4d4b2017d145d3819f35629ead3184acb0078fb18964502e161b3c0ff50ac5290e3dc59601c1e53e257f044abc8e232da48f74005b82abe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2c4d5754fa9b2531d37d8c9dd08a5e46ba6ff381868d41c3a8bfd668504f870b89ab6fe260adaf11c178c5c62d100c3dcc30ca6ea8ba641f4d0a72f56ae65bf533ad57af3179b048b1cd8df75539db47bf4d9449ad312f53e4c07f49b3d9645eda18be97590c9a8a37ad5fb3371fcaf6075820d202a35f7e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dc22eb7a60c9bceb9d9501f87ccfb130e3fe63b67302cd0396a6700f612401975639c982ab387e9c8df2ce06b4d6de1cd6d0a69c0be6030ebaa2ba76858a081d530bc396264ca3d3884991e9200781ab6336a4bb49887760060fd478aacaeccad4450393e574fa1d4d603f15d8de54e12a546a9552057b93;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h194238914312c76b0ac137664b48d711164a224293fe7057d2bb6cb708bd3f57e4309d76f9fa7bf1131fac1bcd94fc94e9e41165152887c73896f47f909f8a4aaa6b1224ab0814a6aa11f02da98ca04a1cb79823df49250beee0bac8ee2a468cd7a2e05507959304c1c436386eccc663ea3503ee3651867b0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h174dc738b28f835caa5ccb8293ce73518581ebff1ce2aa83f06f58c5430eff0e2cc2ecbee056713f2756783b64d3d1a778a57452c0c0cd0e96f1c62fb853e3f8f498611e5b877950c350dfcca2ed306689296f17c7ec30f75a2b0461d787d1255d59206cb29f75b74c3874208f03508a34fe354af7ba8f589;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1451c0a6020f923ab99dfd74d5f279e3ffe2fafdaa8ec0b879931009811e0ab4ff6dde53fcfd42bb8d7f517673a5a766895400e467ec0629f59a9ba1493bf20c0a758e3e28b73ef880a32032d7cf2c569423a12a526d3394507b21581eea6c2faf4dc40686493b69ec6eaa6a18b2934a6dee02a1cbff159b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c3e1bfd8068ead0f8021406973e5dbba4595e2160e2a5383301a2e1428d4962892bafa6d6911a4d0e53832cf4f23c0f41cb4f137fcd4c2fdac3d6003a158f385c1078590ac166ae2804b0ab4a329563be384feb3bfd1d3eaa0686a0c3a89dd6097de03bde4fd646d6dd95b1f10053aa576cfd26e042e044f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9f80946a8f469a0eda93df8bd97581b7634545c448be44dc7064461e2b7e4839d3e93650b05d77f7798d5f9ad8349443f234e44b222b2e842e41a37a3f5a87f12bc1c2f6898e7640835fc128871c372b97ed9f5bbd2dfbb2a04edf4c0858725de394e0203afaf78f7e777685ff9d45a5976ff1cd30a736ae;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h69a9255db9975893ef9acbce961b2c66d947912b2da1b21c1f3353b610bcd3ebf9ab47b13e86cf88fefe48a8ff9ae6b6bf8b80e01d22fc235ffd982ccff684953d1cf58a1f9322b3c2c4911911eaada5413e2e6a2c5f2e8795ae216ca65209caeaa7ded6b537f276534500c974fe4ca6478dc890cf4554d2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16ce0dd46fcad6580aee1cd2140ce718fef58d22bbf7073423eab83db170e6c085466eb4b5e10e73c31c0452bcfb605bedeab97a4f20cf287893b13db5b5cfd7b7e183a9ea020a08018bcdd9d2e4a40cc324344e6eb0729c7f779722545832273ffe48e355cdacbd2172cc10c4635e72407cf60d8b0c62f3a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18b7f543704bc8a20c08049fc5e5c09c38134335afb1b05775d2b7c010d98fee45d358b1c8d99e7f84e78b4a8f015b72f58f220d156fec04f7fff014310f2c08ba849cdeb22c2196969b7d7866d71e53ab36a62edcace3c8988ddbc20c1be52014f54e75b8a0538a9bfa3da3e11f7ebf2a7c0ec509b97e69a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16b6f25db138c049b2d3a745efd33cbcaf78c244b5a3a1c1adce6b422ee7714360ccc22eaef02d63a6f8e5090132cfa105f75b1276f2dcfcf445d480a144bb95a943a1842397e9c5c7ee5f21fe1fdc60847bcaf560835724e4589d82a63ec3444fe2baa38effca15dfda2ebe8090b4ed877f2a655b2b6959;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3af7de5ba9dedf9d392549afa1b0d8128ddeb68ed4675b38f80c2986ff6aed2b502896667eeefc34e5878237f799e98d8834da70e99da47a824477ba79ba410185bd1479089cf850f36fab36c93b78b79f50f593f071862b14c7388fc9cf4dd9d2963a9b4284e897dcf791ae4cdddf8925e4f8d200d154a2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1610ac80d0c463d3c780628184a101df503f5d4bd913de381c205c948f37336b83cb1b81f9d8c44992ffe527eda0158309f76eb6f3f57cc79fd5d1515a9346066ef2a2ea4966bfed6cae7227180f24dad3e48bafa71063d5d69100c6a8d3730c8bfe29ee2ed8860561c35d8062b630816d7b15bb5a9f4a5b3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c2c42750dd31d3099b04beadbc5e383f78ed0b422a54b3f6045dff6f045ba0086e47c8c874cd9d6daafe267465b2a10aa79ed399e29b2091706d0e7992e8c8acb5c5ff441f796c75257edc029691c8dbe2a00c5433cf14b8ff3366035c50efa627bb70e11bfa556cc50c55e146337de56d42028407630f89;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h178b8359f03ecad8b363db77891daa0908f84052181f545f53129b611408ca6efc54ef4d4c2b70c99a236a9a0765b05f653fae77cadb1567e8e7502b3bcfeaf17d672b7b8ef4a1ec32d172f3684ba61fea5b64f2cb344c1efe2520943f29291f79967e57c93d33688eba5d5c3c1eea1c74c6fcd935f3b2a9c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12b11a30e3c860beed4e34168ad20be253f3d48d9ecf17a954a64b44a9cbf00bb9089ca972c37f1367bffab16e571bb6b8da6b26f16dce750f4cc4d55a352e0b177d316d0dfb4235ed4d5a2a0e0cc0d656ce2f5293b2f42eda3a69cf15a8fd4ed4976b372190519e801e5b1ac53e6b332df1fec79fa2b160a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15ea04b39bfeca74732710037e4a9368c77cbeb9cf8ab75fd52833f7527ec6355ff1de36006b7fa762ac7491ba790f0591486e6fecab7ebbdf6fc9c6ff2a5f6148c4ef6303f3169e156d4a3982b690b23d10427da8e833022603dfe10e2658810fd49d5622452a4ca3f747f6c2736104cb9e2df78a5f4150c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha8e9c69292295376191b91a106c20bcc9973b3e2d5ebf8090d527bf613d8f9ceeab5bd8636550468d868eb293a25f64812676641e234cf0f829c2cdc05e129e02d2c25f849e9e032176d5fd1bf8e959ccc1952f07bf835fe5b65b378f0e887cb8bbb693abec4d85bfe8520c0ce76256656c471ccc2b1a2e8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcd024f7fe9ed8b7f7a4528b726430459a9f3168417bd99a49240c487f17c1e854f69ec44b72ddcb78802c4b20c9c9f3cfc65724a49f6c1fa45a8697469be293dc706a9bba710f05d2db2cb2e2ef5d9eaa8663af689f65f001cf232d99823dbc89e479b7de729373a1bf473225bf1b42a0557e5505b21a373;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13227e8fe5ac746e210a15d4bbdcf00342ad46297f8323732807cc185c4da92429592ed1eebb3a681d667e1402d12002b0a10f6badaf656779f18bcc426b932a6e8257ca04a7d0b86a3232dd361b8eb57f9bbe83807f73012a93810fb48624a67b759a9de7cfa2623b75386863d34b4e9842b509c8b9246d0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcafa4f1e34cabd4b9f7a91d528a2c30ade6403663880390b851e203d3d9dbf24323404ef5e2b27c4ffd0a4dd19499c0dc0c8848f0a84f710311786a3320ee8abaa3a55d54dc241529834b0b7f1fe9b89cd68eca40acd8c94e9034f3b32448e98a4a39b1a60330c853ff856667b53a506c815150ff35bfcd7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ba67bfc78bfb5df01f7ca540f1893624d50a89c16fc83a51a42a77a3ec6cee26c8d84069bd55f41d045b6b9f48e823764142a3006cbc395941236db6095bea46c4e35a512a2e7a54ada7d3d326b674fd3c02bed1534759b15e620dae29a17127d20518ca371d42cfde10b74fe4a8fe9b1ee831374e512de7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd50f93e9015cd8bbe7e75fd0a19df48304ca2c150a2a1b707e7b48602e12360897e64e04544aa104a57638d68fef6626dcf952ecf8aa078e71fe170a39ae1a9a86ba9bfcb5008812221ef9529482eceef74cde62e3cef8d5ba171167dbabb5fe853badb422b9f205264752dd1501771303e6d5625026f36f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9608bb6210886de34ab03f268ad46b3f202d2e5124ec8be2edf8ff20e9d520b73522ec967f54aa9915f439a6a927cb27197b23cb55d7674b04407a2abe5ae33622dcb654cbd97f7116ceb8344ce17c176bcd127fa98606c16047abd1eac99e650204b27c5609bbd532e2801b52483cb8d5d1eed901336df8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h41710a3b72357988fc4f30dd0d3ccb4f762514a2b4a0508fae8e29fdf0abbb510e050b355b6b22d4e21256c3003930a8df2fb52669ae6e7bd20a141046a3737695cc4f61688829168507974e8c854603959be194a3ca753865f04683b78caa960c68f53e8cb3dccdadd44d2038e74b6bc99dab3cbef3aa1e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17a317e523ab2cd21d4dc68f0f0e2f117b54396a2b6931086c09bb19f07e4d859f558db81cf4d110f859d5f8feeb1fe73c30e3ea1dab815eef37f5295008b6e20494120aad34f0c3d415443d80f327c1e2ff861236345e40b8d3e26940515504928e5048f2b7554d86ee14216a055d7cc3e5fc05c974398fc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h169a9e3967ac7365916640079acb9e71ef55e2c5d343541f7c5a1d98a94462f464fde5bee520791e800b70b8b505c26654d17a605d9bec8b727e90cb5fa7e56574534370caadc835d878f4986f65f8979126dd8dc4792fb5d6775922c3a169df3d24f3e15713346b9dba4b75e214b3cfb41ddf79603d43c84;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13fc5c39b5a3ea32586bd3e61e85ce95da2c8f1086820d390dc01a53c215f4a720eb64efd1767c8037ad482b2e0081b5c5104d74d647e167b248e9072e4e632fc58424d43ccb55fa511ba28cc2b78c52b7064556b4cc55d3ac338bdcf20b2a4144f7c488ba010384c6de697ca11fc2a2561932b7cae4b45d0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h72445c1641433af10a45157f0f8a342941e68834d4bb2778cc14db96807e36be9d54265e4303aa92487ed25ffffc0d10a4eb95727f75682a119fc43d89e09e40d31016d6f76ce68513db3a27b85d0483a89d28605ce9524df7eafd4229e174535987f391115fa41cc23086f725b18c5fb2f3488625a3c29f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb0acfe9a5163be0fe9cf0875b66608d233198e3a18d17a45fc5b544e3bad3dec3c572edc844fdbcb101fd50c447a9e95769a74ebf12cada7ab45e2d46b663963744ed5c9298dc6a19f8e3b8b17d72aedf7dc429e08b0c0042db2c93edaaccdb77c7aa08448eb0ce242422d5b94eceea1e13931305e2772a7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h51416951dfa2c59421db66de454292db19821c4f93c264e068333cf7c87c376949b0137c02078bb35bfbe933974be3f1985bd0c7f313c8ae989b4902ac85217e935f0407ba877dc17f415dd39c2838b2d893c59d25c3441e4c6c169469a45fe45b9d3a416cc03c58a3cc525b99b23cf6d6544a86a374b7ad;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fae6c9387b20abee85214bac1b7c3b8a992829546a8a138391be798880b9b4334fd071ccad31c57bc0de292d9fa2bd8481ecfe627c19044121350a7aa49754b59bfdda8da1ad0b69d623380147a91726970d7aeb88aac630841742f15b758cc3cecdc57fab09c61df1f0e911776647af36b2a16233b17d0d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h494f091280a3e5f3f8473a482b0028e399d02fe5e958ceb26fd8d73bbc68001b528eb08dad1c741d1a5bd50ab665bbf17070181f42d716886594288e25c544b6d70ef3eb269bda53cc72b275338a32bf87b24de89b869a6bb93a08424aaf7057045aba43a98c135ca679b131d09ab30b1359d05d4e9c44a6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11437aa7b2eb0daa1fff162f40770a9afaf96f403a09d3d32e4de8c7b180ee9aff8485143aa1a8da17c51634543c7f531388964a50cb08e8baaef3979ac147b3d8f69553ed11072bfb07009df63513427d7ade391fbad3d3f57553d0e6cdf497832f407e9a2c0955509f91e6f7db1ada1e68f5d85c458866e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7e56b2989863d0a461878b59713112c7f11d5f157d5c89e0f5babd907bf4645d27e0cf858e1314139b84a63b3827d13dc6c73d4b64d284902dc2899f1f71192d87b9a353f2799e79f36a8fbfea35e08af48edce9b74fa2f86420b40ab7140db882cc1e4b406dc289fa7d901f20e487de546a00f9cb9e29e2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dd84eb023f25e2dfc475310fa2ac805274f9969b38b8da6c78b2f0d191d688d79a59f9472bcfe360dee4dd322f4d58bbccbc1443ef2d4ccbc2e0b65593bbeedcf420b99b2aefe215640c1d8d638b29683ba40ec1eb02709bc3d03655d932e76d18e4f70eed49ce850e1313324df1b4009645392819d0ba86;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf87c8651e7f878c5df44468276f3b850de36a96b30fd3183753d08ab505bd65daccb24d059dd72aa5597a2945ee261f49ea1d5e4261f842882fc59ba16638b2e9f488a8dee79eba6e955abd806c4d5fabffb21af5643db7f98875b8f405a0a193bb4bf042f8109315f8570fdbbcbdc67ca4798d8d407ddda;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13e7615196e58f27639fc43ed5bd7c6e4596fe37c45a2914db06da2949923c9ff41631b7469526825b89c5f464e943a5d9f25e4f65ed3844791ea0a7f2d0ce9a14970747c4dd637aaed4db2af79147da3c034375e7b4dab5dc7d4b14db89ba4f3c5219300806a85e74c2ab18b24b597cd6ff1ca1e6cc26cd0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h189019cab86cce0961b22ff270eaf0dfc86c42b94ad2312745321676702d469b9789ce3c9b90a7a7153e24e56ccedff941ed0c727297497a2721889b1adf20736cd57a0ab14dae86b495c8594af46bc58ca469e1a067d94a301400398330e561b43ed858ec7fdb74be42bd4091fc20ac7ed500dc9e824ac29;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h27563fd8d1c90d73843f00c0809e45a330bd764b1da5f77b3c6c443a4a1ec4ba4f3c08e21a6e8e55925cb13ddefaedd7b7cc72a3f170e660ac1c35050a6be75223d23ace8c18960b11949cc4f3868b42a0006bab35ebe86623107474f439ed8a169dfaf7c5516d292cdebecce6e0cb23a7d957a34f204228;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1701169f3e93d96009ef5d65099ee7fefd754959e7fdb66a4e4720f275f269d8788cf09a5ca859148e32c39db8cbfae7aca0ad9a26a8a17a774d51f57e4889edd677e0697f37babbf0243289785e6ac360a28e2c52aeb1cbf5061cfe8d5a4268d17c89db07f7bf39c815014a684e0669c227a692734bd7c72;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd76d2572876bf54b2218978f308744018b23133278e38096e2f337afa247f536fc64aea320afc5e626489e2b6e33f7674ba04277aa2109edff9b962ee5e11e19348dc20e1cbbb84014681750b936adf155106afa4ba479cd95b2cea67bdc04a787a2e8551d5e846b8b680de894f170d08d9bbc4760154831;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hddd3aa8d25526024b988ae2ff32cd81eca53be184caaaa5f1e37cfc9f77695cc50c09bb1d17c7578f1c2957d3deffac0a94d5dc807ace02a3af9184c19e39b7157709d3384685db1b9e8815dffde5a11965a9445014749f61117a30cc5c6adf3b47809009b5f055c318be010e0ea0af0d1b9e108bd018d12;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7da82fc6818fe5d23f327987162c1216e530365b0d5e92c3ff15ede2ea52544962a80c7742f4f3160a42e8903171daeab67fc58ce6c9827a2e242f65d9c7bd763c89efe65d450baa6a47a45575863e4ba757e456873b4b9a625d916110a5ffc2b9a9fb8f8bed0794592f8d6f4043936ad5b9cdd3afdb1a91;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h390de5e7e585d9ae817a7d2ba4c24eed1eb706fdb30886b6f9dce9c4de48b89d140d36c006bf5d942d48e2550dedc62a3a8fdc21f8d54a2fc02d20a2a911927eda9f497b49755eff94c6f3c2f3b95fb62d431ad47ac49613db3425df92ebd4655e6ea8b9c25f3e07798b10a7d7a5264a48f69c8048b0a87b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17067b0c9bb3abb872c4a835484a8159cb0efdbff8c952da55e5e7816f5b10557efbaa7db410a7fb8ab0c673561085d7f4709343d2a00a389acbd5ffc301607eb918326e6facc52b1971b85f99382f4d6e493eaf1233e7667f497fcf72e5999c4c4f97fb0913a70a900dbba3f7196eaa48705581eb61b9db9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hebc7eb7d19419790eac5ad307dcb18fecfb47d1e81e5ce9bd6d7f9e660fca34ee2e58f1b95dbcdba1e66d5295d3c1c062a3e549b560a3040ef484d20452a6ab6f78d729646de9a0e0e0601d436dd6faf7f128b985e69452ca3fad340e8eef69fd5df5c5fcb73937b481847a800c8c91f660f0690509f457b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc22b0c5b92706ce7b726c27614c33619ba9ad0cd066368941f9850af00ee44c2295eae70b7062576a7de1cf448d852f1efb0e4b87899cfbb0c4e88666f02dea528249c7c678edaf48b9e541ce146af6fe1f25d0067fd3889df6a5f542e17b5627b348b64318e5a0ac3aa76b52a530a6a360170fcd6698d05;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h162053ec9b627686c68804e28bdbc522075f556c3cff5746cceacd6178c9caa65bc3bf936b0e65605586d9be8eecab2ed8f04368f009a1594e7303ecfe8c373e83853080a71923d3e044e42e94c2d4e307e6e0c9c096600a4eb16b7c99e876bfd4ce08f3d1b5cfb5fd10ae4365e43e3ee45ecedf3680a7da5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h187ab1aa709db12686451bc1965e1bfd2ca87bd2502e7929aa10ae14090543f8c307b185547c27215400bd39d398c8a12ee082afa62331622f970c9b26ed938172479185eb06ff34bf04cbfd4ee1c78035d2b1fc9e16bbf0c256422b236cdedb9d6859c2e2422cd58bc6cfd9f888fad348d45b4875a11dbe0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h383961823937ba67292924417c76f39e4f10907aad94f789e6e4e6cb260b67750b8e542dc641296093cc5569121f56ed69818b966651299fcbc4635c240896cbfd8022b4e0d542830121ec321616ad8ab5f770656b829907e4d0f9b9fa6c269d4957c1438dde2548b1135b9bd28c694bcab9e06a4b00ba4c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1798d387454df59bfcaede6768306291d7cf7f9a49d0d33fac6e66b185aad339a132d512b2b062faf48a0de7e26716baea4d7aa7980d71f62666c3898adf9a93141aa1da1a0167ad82d8ce56b5a61ed1c44dff815fbd93965866f3b6dc9292e636b913d39fb44d360feab93b20f77212fccf328c24f04ad41;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5eff1da88dadb1b9afb45c7baf8bf9b736302eb7bf7da2a9de9e80ed6944811c39d564a9d7fd907838a728a1988b551c6e6de2b69fdb03b533ba18b809170973dde02ad27415558265e384ee472733e0bc91922bc735985b342228d4114c34e40ec6dc2b7e763556f86ca05c1d83c3814afb5ccd20c08e04;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h117eb7a4b42aea63100e31e07b7fae0f901a4d264d6977ecb9733aadae34eaa0486565975fc79d8124e7e9179c9e7b5fe621e07a583c1f63723d674b0146c4a5a366b442e7b67d5e9cd5c9131c7d2c27dbdbbc99b7533e0842ee1c6e9d51f4298f31fc80fdd56df49c08e1690885aa912d71e4b11c0de7f44;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8405846e2cea263f0972a194e467d0b841f6295a13f0428c08a0c4d1ee77d6232aebb0403dfe0c3fa1533e6a3e96cbf5fda85e0a266dad40ddc4230ab7a9059bfa0961db257af8b3cac09dd124103243c55759c0dfa81e1abe45e7a6f117de4b885cfc6d8a18e2505f2fc282bba9e74aaa20936be1b68c2a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f697399ff8a8f058930a2f1e8121326c7de598d62c4d3e07a51d0bb44b9ab8d13e93ca7f57fc57bfcde03768802cf2647af83429f1240ecf2fbebe6ef50f3cc0b8b757e3988ce9fa278600d2d5867b45202b68fc81445490643f2a757f7907563d8da916e1b404e6bab023cbcb0ee35f066ba9ebc3088d60;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12f419a233594283131e86b7f0c61de9f3a5a4c5c85610b42e15de95b8d97092ff77384b8175c10a376fa5d3256746e1df1acb2acbdd368d1b87bb6c8a60d394e591663c6d6f3c1d9c28c861cd6419b3adca476f839c1587737c89c03f587db9771be9b8f217c52cd5ab0f9fcb99c1a2f1325a04ca900c38e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1289ffe4065ad67fa7ddf57239ec5c24f89bb21d9e7ddb91824ea25bf8ce5b444da832573b3d0bf4f15cb5b42da777f8a3a700920d6e0398de38d89b9f72fea23427e43ebf3375d455c1e71e29d30dc70c1437395c36ae61fb1890b7e41dd686ac9fde0dd8bb53c03270a3a704e04b8705fb17b47b136f0d2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h88c613538c047ac46b0e1218ca12503100aeb36c7a2409fd2a5c3423134b5655a777f7b2021cebc2d68f4b50f5a71b2ffe4d5e85112761d36900a18e161ffd58f6149b5e7709959bf4328bc9d857ba6994ea11103072ce88bd1cdbad9e6e2b02876e9e06cff4916455dd5f2379b97754ec7bf005b0c66042;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha2b11144149ba224b03fa0622281fe14a64a4643283a89e4498973292de9d4ae5896935048386e64d7be87840b69ed9f8b9dc3575b78bbf69a919f8af396364ba7519aca9a465bcbfa6b9f8f17d68e685dc77854df99d6ef0248cd9bc3913e48b9e2ae3a20a2ace0f3f9161bc8b3b8bb069b486e3421e761;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2964f69126a5f95e3dab884d3937acf6c0083d87a434657d6ac0633730d3108e534229295ab3d1a3b814d57c5aa5d128670cd378ee752ffa0e6e2ac46a26e2cad7b090a51f36eb271db67141ffb034186e97393e95dcc45a28f1c9345e3493a19df9fef3b8bc208b0bc2f57fa14d9ac51476a3f0c26d8e90;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e6c30b91ea8032c2fc9b68a6ce1a5a19e8016b5571e94fd96a24e9d1bb9969f5fa0ebd3be9bf7a7c278e0ddb4751e953fb0729464604789e8e1de76b1381f64fcc1a75e389dd9322c6ee312f77730eed0a574c6f833a93fe620e7fa348840f53c4b35440008a63395afc9353291b3f4e4fa88a92f9d05387;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h540eb9fad9c38d39d04a7c7ac3c6022929fd3853ff091624198ec777d9efc6d1cf97d26af5052365f1cc27b39d853fdea3bf5eac88633212de6b21df82a41fcab33b8a57e5f1be7cf46878e5360f0651304897270e8ed6321181f68071024f2be77b593c2677d61406b5b7c9a59df53cd0bce8af7f2bd95a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cda2c2fab9bbebb6641c1fb2bcffa457bae1d91b0d726677e6eb30674a8fe8103ff1c1b0ba0d524441974fa04e21fcef48ba083d783d205662665efb0bacdff60445e96ecf207674505f1e64ee42a81362746b2923f4ab5d03894e4605bab319fdf476da45ed0c1a67500c36a288290fb30d8d294fe73407;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb82967a7d608debdf1ab6b7356faddfc0cae04639d0262cf793a4b0c209294d248846dacba7e773ad2b861ad7c94471d7590afd73f504ffdb378ca4121828e28a085b79a32aa289a75ffe40a838a63b224cdad358e08e479738227db8fa0dbbc40a26a146a142a31baea549bd9a36b9afff4414208f4586a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f1247172b57e4fe7bf3687716c799b7ecca0e8fc5d4e2169b234871f395b3906ea13ab9c5c439b506e891f14b67e7fa92917da2e9a292d08202f74ef3258da174389f8bd9b51607fa7be1791ffd803a6df8dc744d811750781614b221352e3e7eaefdfad24e25a74773097f37efb34f16792cd4c320c1e30;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h556a736f3bb734f92d5b5337ae2ccc3f9fb30d20f6a022a00454a15a94a268240b0f22831ab75f223cb07a4b0ec1b01e9c11b546fd2f819d0b74dd9eb2bca3ecfa56d37e729e2f749291674a1e58100968b1a6ab686b34c9fec261ff9f2e2df3a10528539e64677dd1a98e03a12295132a352fe6ffc71f07;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf59e1a29a8558094c7baabda64ea6de9c1fbcc5dc351d86da129a41b3e127cae4071235f56c4bb73b80a2e5f869185b8aad6fb34648742071a209a33336f96924a5debe2fd64aaa494da6ed7ac45d4452c29fd32fad2d46c51b1078b19b79c0eb9b23c9d7c1c63078adfc9478d16b5eb0be8c216a1aeea97;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h49f1813878d185980515e5adb2d9296d53f4610b3315c31b4c492272a8fc1e27aa1bce46683de6a04fb9ea2dc014eb3bb270962b9b8003f84835e77a06f5a22d67c5ad6688d87127b4e0d8e4b0ee5ce1ecf70bb665bdba6b9b6a4d4bdf8b7573356c8fd2b1b957db43dff2d6b947b89f451513c0a1b3d856;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h70c30a799446b581c56a33b07a3e033a63d690f9be77ea85500c44e83256cba4656217a371177c4df22977cc9b97e7e343e1af4da90be1e5e567eb298ce985d1f48f498e5af625451c0cc6c562b1ba585d02ac137083fefeaa97623f9ae40679d838bf8d5c5655598b581172deb28d858745bfbe59df83e8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h788e14c6110d37c2d1ecf79272c73378c6ec44478373b28de68a20362f45939d6100642e140cb84b871ad322dacf72501bd1358b3ff28de56fe9736f01b453c38f7da018e337a9023af00d0989acfe2a942fdd6cb3f71bf683ff9f42216e392069ad3d06f3d4f69c231555d86177c20d74fbd1f0b85dc229;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11fdf9a1e1d26c50d83a7ab3dfb5db45f89269a22a0ac444429b789f2898b9c7440a9d5b80bced46ed329699ebaa62a89e74021f964659fcc8590a90234721dac65a12ed08301e2b4b50ad47e654955fca319030ed9eb3d5c5dcc0ede368b27b2ce419db2ccfa64ceb1a6dd1e72bb73a6de50346c6cbcbc49;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d22a60edf091e1443b91f0a050da2b4fda9cf179b2ee0ed4c91399b5294a8d9f6479a090fafb402d9258c727247bb5382824e35683f1548fc97945ce8f252ec1f5e9b9715a65fc64614163a0a6057a7efcf886380ad15a27ae47c3d9084370decff69d92a238f41e5f58a14e8dd978c64a90a88ecbbf4209;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcb140f808f769e717f4bcd7de73e3c508aa269057ba053ce15635f6ba61bbc10fb094d71085ea8818e22a7e70bc23f1015e524d1bb81185089a2b28c5eb8e1c261265b96d847576896e3db5805695d0ba44d431687629a9d43b21cd32833b724219e11da71279e4c558534d4f374512d306f835dad396ff7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5a49438c789076dae7b08d3679e0c38676a41f975619c8a318c7f7d3e22e1e0467c908c4a5cda05ccad554901124daa03694249adcf68e11b25b30f1c48342e07f6b31d8966eff841c4d6fe21e75ab1d2512fb1a9e485c457a6c502ef3e38de70533accb5098e88336cd880094fba91aed4680c4453fe7f2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1622cd174eacb062a3faa911658c82d8d2ee6c4008b85a29ae594265435dcaaf091031d2fb34748d2d6deec625a780cc1c11eaffadfd2ed45c31c6a749f54d95cb4c80c37640f79d39ff3f73be21e26975cbc998b53e64d5b12480b2acdf466e57486e96580969413d1daf55d92d7946f386852f7caa7989a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h161714240d1a1a250f9163ccbc2cd8aee924d828aa2798b8a9b5f86dee4e1c8d4e6cb1c480e2f5c8c6ac3ef38f3ebb29c534c9fd1effff2349aebbd62167e571daa9ea1936c9d82d9066ae1d88ea105b2d279bf2bcf92f39804e3913fe011efcc96916097278fd4a46561233aef7c2359b917d4faa9da3abf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18ef6759594459f0d77813b28bee0129bc7ee225efe0c1f43968eb0e6ba7ada62869e434603585d4be2b2c991ad74d870a6e143558098b3ac5c8e469ecc3d2b7daa95f588774d7413b4705a9a88f29117491d2b9222d853d1e50da321370561e75d879db038fb188938e572a5623bdc642a2b6d0122bbbb10;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h86d9146cfe14ad3c377f0ba5c2c2dd72133da3d082f7a81b830c7fc6c79573fb6efb4817ff973cf2e1db1defee52d2d6eef20386ae7e985b6fd2773de2a46c5546708bde57968942076e9e387967d1b424c6d010d4dedb976e823916c300fb56b0b5e54261119aa60ab88b3121ac1de5064bb1a970eb7d2e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f286142202f70387b13384cd41eccc4f249ce5a85c2d21908afd0c51abed067b8239067d906c49cf072b9b86e82d2705052917f2349b1b1f285f5ed69adf6d4d515fbf900994cd59e6f49a373d982c64bd9eec63f388dc18b60d014a4c42d77714f9f608d5e671e6b61098f5920cca2ed98b3c78373be920;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h151d7af9ce056d2fd946fa9dfdc69f3df7977979966b8787ed16c1bebd38f146f0e827f3f10a7148b2ce84a449f8aa2bc51089c65b4ea0eb1b883275fd8ec04485dc8f1844314d48d88695f6609c1cded51b7b1d374bcec8ea608231b6a71d65775c37a6bbebb25550cc5d0ba7eb5e3d33d6c15abe514b3d3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12eddc7fe50788ed24a70f0296a268f1a7be05480ae0a968715de94ee6bc1ecfc13f97bdb7be44dc53c74c86d86ee0c876e09605ca6d1004646ff7d4ce80f054fb400fa07d113ef940d5b08ff33c047f27e9ad7ab810683d563b3be142d1062311386e37ada896a7bc35c73e89e4bd1a6bd4d394bdb8ce273;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcf241619459958591d21bfb79d5b98c69ff1ab2117ea0e451b9fb0f4f28f0281ee0ba2bb9d116b31563b765eeb346ead826c00ed709d136bc0e1779f837680c5fbbc04a8892e479cc1a7dced09b1a4b90bf5d312ff0b21f666213099c64f2c92c8e858fadbe1c05fa384ab7818052af1750234e02f6b103a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h130303cdb2edad271e26caf06b598dcc8ef49727e1bcc9ab2952b6f9f1bc62489390cd0b6a2313196c94bfc537e6c1ae65a415fe9568d09b48cfb030bc5fafbe07b7e1867e5c89ae065ade33fe1533708a038829e268c092370efac203cba41d063a964bf0e9c83e2e2215e64f75886ebf5c6d977419b6ec7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2f920d95c2ff0c3e251c3b3a870a56d927cc7a8e4d1cd42defaf789fb16b46acd6a5fb6c6d0b2c0becdcfc98926b71001e6d6f34341fb5e3b96485be9ed73f773be092521c07ba7433f1efa7c412904db5b7ac556979a60ac542076162d46daeb2ef6f3e82405a3c898dbae4a4edb7150480c60a49cc0e88;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e798947e3ad78c2777c80e991f17a244ded86d019c5c8b286e14a2c097f598d9440f89ca6fe83b67ed9e57504c0ffa6f1925d2afc494b57ff2bab9a8ca39f558066008a04d5d06afbce87b532a067b253cbeeae622b2a9c6ec1f90631860aef583cbb18797c53c147e6b6aacb283333350165b6b9e3db98f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16b14f044b6f7300b10624da68ac9d167a6646030db5794dcb84d3ad553b3c047a3e26cad7808339d8edbc1277d61aa1cf31907cfd9fe5556a26d2daa1663a9730b2a9321219cb1eefa798acc0de8bff1c34e76c88ee94420dc59dc729b9cc548068d7121c1dda420fde0c2d98e879b311d8493f11c344930;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h146c708c3932b3986b60ecfabfdac2dff430e44d00b6765332b1b6e94a616d4261d084e48b685fecba18cd8e49bb4bf3b204a0dd29f29a412765e190969093dfdaf5bda309ebc6f937d39865f247a35c1096d06660941c98ed1aebb19d87b3519fd07ccb1115f2bdf5ba5a6dd108839d1998b9710b96853e8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3fb33b7e9d14a4bedf6379beb0ac811f31691855999967613b61c7e5c41dfb96e97e6de30a67870089604fc1da43ee090edc18a4335b93670e5534d1e6a259c5eb4060841b4da74370aa62b52b3e102b4b6deb68de8ccc3268d77aa554dabb8117c0bec958ddc6a670f48fb7a2c977f48c8e05aa5dba84e2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16d95274daae2e8486e04e6d31048e3907d8a5d2ea26b0a3b9203bf79d8ad1a79311cb5884591b71740c994e339dd5bcdfca7eb49b81df728cafff2ebfc7a0a11377da6a888ce53f2f798e3904bb0327994924e94c2605dcb0d59684ce811002c8ebdb85921c34c3b24b1379f98e72bf11b754847dc25940a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h106554c74a98490d6eec4be2dcfee35c85f7f5eebc7344bc8adceb4e8c882d6219480dec21331a2cb661cd6ca7372abc38d36af9d009129890eece3d5b2cb7dc16d76dde915cae1b6ad6e3d4cb62694dc319d8671cc2d44fd66b828a0dfe6aa0154f958e5bcb5925971209e825cbd1b022ac7284734e79162;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15b5c86de720d74cb311617b115fddbe2a1aac9ec9ed2d15ea9ee2bc84f78eff6c0d60d9e26dab4950a4b3af9d059a007748b8f019c84730b8a9c15114f26180cbe85aabe596427b7868f523d9639d86235bc5c8517eacbc52c075ab93cab914eeb1e1ea5af199be4efb23ccdd84faa733d203323922875d4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdf65dd89fc22b99c51b5881280b9d38187eda377abc1bf2320fa383339e06f18df12db82e754c1b23d40670f2efe59b6ecd1d16bd59423ae6fdfe72acd93a06d366cf5021bd36f42dbe82f33442b42c125c08e99b272c827d22a90ab3ca544c36c981c6ab45245cb1f09667c0fb9127a62ced10fb7c6d362;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5c234f27b34906d7db6b1099c6e3de0c688149fb817065dca6fbbaf740e695c264cf56267c171d4f9ab9ba9c8c8624f7f5b3cd70aba4eb16129b62914bc243cc4f3f3db4e634788f827db2fb0c480f0e05fd548188dc8acddfa4b6f91e81ce4a7dd60ead8431313c298032803219bfd5769c8254a59759f5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h143df6efe7d0305dba7dd2c4a82482088d2668dc74b827b874fa0c2587b29a8b01c1f6d53e1f67b0d68a4190e2fc90017c3b8b2f65026b2fa4245271298b25b93f159037ae542e57e7aef9ed3dc0abd2a0ce1f0c3eec2a48546cacfca52b6ee19377fd8ef843b6cade5aca450057e3ce7b943bf216c4193c8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ea1dc2d4ef66164773fe0d12c649f04f4232d3f0c41110c39b3bad6a80c23c729f962ce205c0f7c82902985b970a0b4449c01fd3bc747f1d42f85a952f99d6eee3a88659468bc9700c0019de0d3c13222265adea955df762b458683c91d1acc0ab9f7fc3b613fc96f4480898b82daad4d98a42d7aa5cb330;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1089db048e3bae801ee75928b54c6bda13b5164d052f03c125307af73e5ccf7c37856a3c6807c60647d20abd0e91bf84ad7090dd29b9e0b1f43a297705185212e9294d629623808725ebbe0efae154d83d42fb965951483139faaddedfe22bd0fe4ae07da6235540fd3f18e4743005bb5401e21e78d63ab13;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h25096b082976c067a991cb56b3f65ca2b96b82c6ef59ac4d0ca6f1615d7c1455968185508a1437ae4c6658daa1e48d51dd482f0fde9b1e1eb5d4faa77ec0ed329ea4101680fa27910ab0e2c9f4dd8b5c2f89177dc13ffc3a034e1977e69a236414a7503a85fbe86bf983c243f972083203e1254ae7d440f2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7a767585dbdec3f1fe93f9727d2de9e247b6b89eadd84732449a1ea09f148694798d3dd633a16e652a72cf4aae87de5bbbb9b5db74bd14e84d41ba23ebb9433420923601ee861020d9fa07ed16f2526b7beb35c3604f36aba4891134c12ae0edc1f5a7173a4f33f450c7fa4673711982c3665c1e73a34ada;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h65ed596b98daeff1333b7c310ce5c214dd08e91f4d53fd945d38c29a0e14346376c5e90feae03bab58049180f4513884d228f2370b3746590c8d7e17d0c9d9381484fc8847b5d371d65bb4af47f1435ac84b3e5b379c0ff3be936dae99dcc9b18f90a8d9db1a0a46ab0d666502d8fd349c7e822f4e90b34a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fdf651b6df9b6e26ae4d45ccf1baf52cfc68117d7e18c18923fb0b80dc09008d7447ebbf94030f33d1bca28cd3d527539390e7b5226126cf126ca2229e7e4c8b294f98cd27df992b0f00546035b61f1d75bb143441185d49fb1d8884a01199c472fac7e5065348fe6ae48437b0ad2b56e6787b18add9c9fb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfc455b0b68cc5681e4d93d29ebba185b77aa4d3151cae381a1d2384108d7137c4efccd95ecd8ff356b750e9d7ca76fa272e7d16401ac54f3cccb25434099f7f84627c440df4c147ffa050801bdc10f7080a459c0c55526a9ea6c072a1ff7a209d5bee0252a0422d8a9ac4399eb8186cdc046e49f48cecb33;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18742901c987f33672e6d61d8f24066755fe3157810b9d5aa0f3cb1ca52d15810bc4b12a7f89ab713753adf31896b644f534366bd49c815c23e45b0f5ef24b7f459c1f8794949fa83b2392e2407bc47a4bc43536f3665980c240a0742b5be8597c5c29cf68cb32227de35d963069663f448a3e2f9a8d7730a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h75ddc4078ee1cd33230889530ca4949ae44454dcf6014117db8c35d89172a3500829f68816d2eaca48342668ac072d9c83f6266904581b2bf4b88674e2d374a53cc792b18e36f38f1fd7f8c76527ff4ce0c5f427f3b2001098ce6bec36c9593d4d0aaa4f209f100a68a3bde9fa4ae60de398ee2860de5f8a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcbfade5217f79788ea9908d2d5819c0209ca4d7bce22acbda19a4d92c0690f09d3d327363eac796443aa61deeb028fe9bba140fee6fcda17537bf5fc079e6047d4f6420b6e9e7cbb5bd06231e17194afd65fd4bce997ccd627eea07aec645c9be6c19096469cab4f245c00947e48f7c2efb7e24de82f4227;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13d02d57fd8e24a7b93b1a8fad70165b368b62023d9c0c36d350b3e539097a3df49dea19c103a5932976fc3f0a6e3ba94f23e27366891ef64dd16f7ebfc1eee2851cab79ab7863c01e8c3840dc6b5c21e3852507c6ba939b73f008af05c54883e19d595aa5234096779e5f260837d2322643935e2f72b62d1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d1b04dc6e0ef591d6cbeac9f1f36bb60bff0b8d601b6dc8a443430f0bae3ac8f9a7fda28e86e1d9262980bd24271c3e5426aaf1f2e0116c9e6994e17e95403588700b30cd218d333969941209147bc1a622dc5e16bbda7d51726710f7325a9f771ebc8c9e2489acde7c33810331912bc2deecc1e3b3c4763;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19bdaaa9dbf0596c4507c2420b89d180d93d5dfce6a3db119e0a4a94536a6067757e714135cb31fbb2bfcffc6f6d3c802a610c0faca44b9252b66cc1ba5b6389fb406391861207457f266cdbb5345921341ad2e30d2d85f1345507c4d0c7a8045ce4c9f6efbd3f93ec80e8f1a5af58ab77d6d933780cc8edc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h717e6e4a1f71195c3541eb6177ec1d1606d5ec23248ba6eb887f383dfbff556403837a0ac6d88850fe8c60944a9958a70a298718ff3077c33692bacdd4697b696ae1d8600f75839080299adc1e7705755ec535a773b86a9496d46c5ca4aa301d82a8f17b737d04bb66248515b3522cc7e28b4282ff3a711a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7b741ca10db16de3b6ebfac23207120de2ed81d3194fdac635deec0006f9eceed4ea6b1256c85e887756c5de8393ad1b90398a5660f3d4b1eb2d90864887dd8c58ebd0eb32b42c4669541d7cf9c301c5efc26747da3ecc254e076b2680011374a72ad9158f5f36303138b06106f266ed1fcf458e89a75b76;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1abcb8723d109648bb8664497145ae4f3af1ed5d509bc39215d0a29a58409cc27bb8728cdbf1b7e8835203e77ca567b4523041ac865e46c6e7a55a53cd77aed4d15697cd0509fbe15820592ce36ddb8e8be350564bac0503379c92808e78dc1b4adeb5b55b737f615c78d0818ef443518b73fd3f7d758bfd4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12900dc9ab235bca4ec7356bcb853d2b33bbee6a91a804bdce370cf09b9fcf98e9e091a21aaa482e5d70fac309d9e8a7131dd30c52e86b108439398fb09ec0fedf8631f2038d570d91e451906e7b41b0a8b81f35c029782c2a334573f8afa2d89172aa5441e0b104f087ad9c7dbcb3a4089d2d78995cc6c4f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h91c71dbe0870720e128c4712fbc171bdb5973085624d6e749aa15e68d67491a0506c53f49f280a1d245696a8ffbac0c8d9d6f678b58440f7e69d1176638c9a3d0ae6257dd656fd96a1a07a2f4cfad6b7c284dba928c4ed34d1181613d3cdff843409af6e4038e9f0c41c08ea3f3235acd04450c88bc6c91e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e32e9861964d28576a4db8d1bd9f4bc69af1ed7ad2791478d64018d86d45a7bfc7a114fcab3563e40197d71f76b330ce2e799cd4038d03b18734422d196338d8e77ff3c54cccb617e368ba70a56124dfa2a59b369f556e97cd90ce8efd5ad2e20c1fd30ec17856005c62853ae07b7bb7024bb99777d36f86;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6ea826a440c9e88b65245a2945078da21ab6a55bbfe4c436e580176e9d213607094969f920171605178df7174268980ad198ea8cbc9d415bb30685cc8d89a81f22619f7c11cdb40bc1509fb7b5535636e1c8d0ad44a38eaa8eefe9203d1468bcd3d7f457c33804dae6c4f6c046a29c640109d4205bc9bc9d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ed166887bc009624438682012371e0dba694f07926a70e82b44efaed595f9c0f13e6d3fe872d9742e957d49a2caa1a92cef55f5879b100776f8a48e8d77b24cbc597b1fcb18257c2b8cc6d577f9e88bca4cd4bf0b787094e906a7cde650bb90cbc1d5aa55abe7fd92866b9fba471376b8f9941acc63c2cd3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd2c9bb0c42812c263a163f8763f14436fe896c8298c564f44055a040a1fb8f6c96ef1f50cd1873f640af0e4200633bc924aff509eed3058ee634d4b0424e6fb17b80316402b0f8b4137ba9302ebc99f3dd07cee02459deb05922bf63d72733105605d86bbb2bf7bf68d26c96c5844e7640efd2af2731a40c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b26d23a10a511d3103bc8e4e106b3aa5348ace8225cab95266c60f506fc0aa771ae3d5fc8a2f1f5f6dce314ae25abcb7f346f68e25212c7ad9e0312e07a1b0e4e0323e35a5b70e268d1a2af8115dd5b8ce20445a957279688d887251f453329e19c835ec189ffddef3383c29f36396a93cd60c9d1c1ae4ec;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h52fe66ad2737eb3f20c1b513bfae36dd4f6432bd0faab6ed362a0b59e72f5002edaa0d6b2cd9cdb4b268cd08803ca04e2583d4c9a05060c81bdac5244f48d765a201440f4e68db8172501192090111a9c7de80bc9946faaaaed6de7526b0818f5afad1172cbde60e09e3c09d32e7619994b01651853903fb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h72f5993c6a68dd7008d31e36a4d86dd8b597a679cdf7b60a6a74ca5c45ffb5ef7f944f2351ce4e13dac9b6548fcce904859bf6ea39614a2ab287f37eae8c3c3ae6b14b75ceb920b28b4655f162256fdb9c3aa317cf770aefc865df109cc9083756d36436e64f838a93e94d150791636a7685ab098a9e2894;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb2536288485091dbc595fd83c3514093e2a17065a0fe048312389823312cd9478cb49b430aab70240903b548a57b3dc63851bb3bdfe195d397a7745a480b079c222d5ed0e3d78256fbc9155dca035a15a207a37ff6cc2e0ea36163ca8dccec82a1cdfc5023e350807fb5924bf4939f0582f83da4802c435f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h142b2393ac02b42dbef868644eb5b93846ee763b1a979342ce05ea84c501b31d377a3f70c791f8eeefa851a38cc8d3a761a8cf636d491584ccc96913328913c771c4af038958c6fdf019d110d0e14114cfccbae074de454f1c2da0d4f15aca496c775bd6efa009ec56afd744d494647c863dcc76f0b5c760e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8e789bf1ee6684cf1147b12820d475b3f2c5f65b1f4bd7e75b0ed582e17de2d8d3f293473dbab2467558d08ed2e8dcb59caa4882e44d036ce006e9f1ae1604f3900c31b4894c5be2bb271c30a82083f16410babc27d07941c160c550dec0883e5edce8c16c41069ad35e08ad697ab583ac8e2d86347540c2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he11f63c54e98d2cd08c6766bfb7a30a692bcd5c3c29d239a4491b17f305773335054026bddc26af56f5c7fb5c76b719853428b1914f96c90ff2236ba9c51a3e07a301b6a1ff0f6d37740da8c07bb252eeba3afc564798afb00f732e6c4e4653c6e240c047b990b548623dd5855592c1015aee75e13c57223;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c9d58685e762d47216f894b61bfd671ac8f94fa370d5f4be8a3b2e9c538bbf72e174a6f36885254115c1f1f902fc26c40b92f10874e5603a4798d4b0e4016e49c0c658a61428c684d7738787d68db77a22847fc7bb3fb9bd92cdaf69cc4e94d88e2157e7823681dfdef2e0fe2e7929664698d545353d2495;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1026e90356d3928549b1ef0927701e683247777219763b636fa3bef4397707455d9e022d96de03095d1278567a3607542d55fe41614b4288b3089c4eb65e47ca561d5b8f565c015a4269d0897bdb8837db11e56924277b2d0e7b2f2fc51dd7f929eeb5dd2d020f8b2e3ad14a34ad9fa6a33e7a5047e1735ba;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19ae317c5b4317e603143d01be2611fdce2622621ebe5bc0de88e711d8d2085cd7015846580542a8adb23945f48b1450b8a91792ddaeb5e87d3b53a34e896c3363adb2e4b7c1f7bf6dfa16ee73a3a84883b7a8fd789cf8a07d62d66bd57883f6b71e392e3832ae78b3e98dee383c59199fc7d60fa90a24f0a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c7e1bc5391a5aa411e978caff3356c7186504aff20b91b5a46fd8ada9def682de24d092f95a0038fc00544c4e7400ccff0de581c27e8e7385510dcb1bbd0d77e4529a5db75171d0d7a695fff64d2a2ae3ad0cba341028152968bfa6f0e2d1d1bf67b22c6ce2ec424542c54c1611a5658ac3b37e3e53817f1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5cb673752c42826b53b97079651d0e545fae092b99e3b4a22be1e12a52ac11b58a72a713bc928e6e3ca2e470bf29345ff9a475beeee20db54c0a06dc1a6c7381412eadcd3e3b12cba2ac6ed5fe9c185fa354c43c39d08a380777e7ca06060bda85820c9d45299f82948441b11338b4d17dfb7ff305775961;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc5a514a627aa06acee2af192d37cb0bd36f598f2575333cdcec1da227a8d80a5aae3bdaba340fa7b72f265802e1bfe4360d92a0dd4e5c55161b8e4311c2755e2772e87546b8b912d00485ad0d9109654fd06948a345bf27b52db4e5cf969d3a8c72f285db93ad6b964be1a213253943cadb94dda9ff85a81;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1981b0f506bfcb2eb73ce9d16a9870b529e1da26e4a1e16f83c957c0df4f413e945e7076afb79fb1e1651bed9eca6c1c4931efa440cd7049854dd61f959eecc5700040c51e76adde420bb1c53a762ab4cbb79f0f1a4156e37520b2e818310f57e19b5ed143e27ba6789bcca7efc8b1572c259ddce91b3d0be;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10afc41de4dfd8d6ff09f72d8802dd27ef2b38d8b6cecdc727e0e663e43b38399140ba101bb2a63c8415ba301d4fde60bf83ea1f588db045dae4de7c1a8f86c406825a01e71b03a6339aed16fd100dc51e6f49f5227fc290974f31bebf7db511e66f61a288373ead976691b7af7ced2e1dd68698ad44f4030;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a8d174268789bd492287d0d2efc7421298decb3b83b9635ade6258eb18bb60db38fa468eb36a52bc8426ae498cdcc034c57063ec42174591a2793c1a19a72a05202870d73920e945e37f0690039214360757545440967f6cd48d09756cb51b5d0c934a6599103a180bd5ab05efb8cd0f955d0befe937a775;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc08033b776e935e9ad437fbc1a4339d9b015dc150d78c132ed23cc4a6a9f0865acdb4744909084b773a1aa4d96e88dbfa33a7053a68c6af79507586d8d43637d622225581e527aebe8b467d74a469820b665fb527f3f0e7813c469b002d444bbe4148c19ab7d1d523d79d511a27e126a954aeb40a193a1f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8db91d580959637c1e5e281a5c5788d8e8524b8bbab7bf8ab8fed89e31c2bb68e6ef79bb5607657092d5fd098f352256742c5c328e29bf22e5bedcd973311a51a5c35d59176117a92ceab58c2ab78b4fb75c04c195fca91d87aac323fb8dec6b22733d88626114cfb8ca92928fccee9340cc882e2378cf19;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19f4eee45a2dc15776367233b390d19fce12e034778ba629c7d72c128748cb995b075bde0b30a86bd40ff43b51fc407f78e2a89b4cb8f0cbe889c99a2c5d3e8e1d8c7c60ecb101186b5e78eee99e04bd80e5e1d8870cb9cde4c574bac6965980d8f788456f6b67a3821f8676f07809913805dd2b509db7b78;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f9aec2db6f740eea720238f655827a08de23fd4ee490516a92dfe1bd9a78dd7487bd81eed0008fb978da54a7e888a41709a9888292474b30109cfeb69d56dc1f2751c6dba3a98d7222a3c447b0386dd30ca8637a4b934016271ad4caefb519195df84ca3acb7c6572f275908edd63c03cb11b585d68bd3cc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1adcef85c9bef2871789fe00d5cff0438b86cefe59dc57f9c797459599de4f0b92b14717d9dc2eb878ed56166f013c193ac37d83fd06ee9289fb517b102ff00d44609574d383cc18d7e8a71606e47899ca6913329b8c7b5a5870d4f66d37557915150e187549dc3d5ec606395e886391be6b7a3ed2cd6b106;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h28e6d5e7ca0e8be9773e6437f1c44a00b8556e9bd3fa54997af6c13967f58a27c1a8703a0485820f1329f49380faa184abfead36d58de5f18523d18fbe23592c8726cab18efaa9c3069efa7c10daf6c80d95e78800f99ef0cfe84a1be125ea063dd2a40600d21f7a51f32d4495812ccc56f97a193958e960;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h83d529b5735b1b0396df15cdc2d2673e1c8b28fb953b5e01b66af58855a38874acb8663e7e5d2a8c00bcde9a6103f0e30b085f93b4ddb35b6f3d44c85ba7c6994fb8bc9ecf3abd12461de8dcb3b826cc26147bb3bb3a939889463137e893ba1a5260271ca8005e0c8f3a4c3b5b010a8963796ce16466da73;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf3466f5f7648c04a6f0e7b8f19f1a92c7b49c474baf67bcea26ffd8823c3066c9e07e489a8775037253ec813d3d86490c6775000adb0beb822b8d5f7c442025ab2230b1697b2427331f3fc68d94184e6ff1c4a3e04ad6b27e1cfae11c0d2673fbfab767013a03e815d199e9926e8632ef85edc6842e8009f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h68b4e07772743b9a90e73854e49b986c43c4e8ef68d76d388c2c48aa68623d09f97f903b12f2a9753c0a9fef76fcf28984204e6010f5a4ac3dcaa1ebe27c035092b811bdb65f29c17a85d3757792380cc4b4fae1943a7fdd0aba7a1a646fb7795da3500ef97e5d0d2b47499c04402ad70461e1cbc0523d14;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3885ef4befc5de5133a098c5fdaa4b2fb0d0bd404441403c97f67dcdd8a2103e734a96da151bc4c55c2058101ba16a8f6a5688825d483dd6f6cc714f5221f00d265560e5da2da0d9427a52c23753a900c6d793d2dbd2f4292ca8306685f9e31f287fcdddb85cd8e93f354412ce8604987474f29ed9d480a8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1201c4b053bdc74149fdb605c797b2d31397891d8056fb9826989a9617ed6858e1450b1917e3f4b71f2418c50f1c3433a2b878a8ff982c9517dbb2317140b92a1e9468b6480de4f142caef3b4a709773f89fdbd65a4d431752e5e8c140cd01776eaa079d3b8aa07fb7a7a23adb80cdf678f8be9c875709604;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7ad3b6f86d7fe90d266705bc4bd3173e1d5c9486eeb16db11d68db61f144bf02f13e3dec7243eb3368a901e6e3f0d9bf8817739c42f4d528d46d75a36f3021eac98af73518537e136b03e77b2f8b136f46d6597e35fba73902e5090df72bc18dd548dcdd903a6293b1ef0c656ce5aad225f8a2a710a0baa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he7062303cfcf994d84177174ae1580db35cf18c749c6af1a53c224c00d83670ac3f321f8e3f6a5b7c7cdb9f386d27842accd1232ec1b73aa40bb060fe4b45a2f2b0408a972ab2085f41a89da789bef41415f8690fdd258379344c2ab7ad42a45289d94a9f013c4289faa80a8c6d4c578c09d06b203a15e24;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h869b60cb357a3e2e486f40f136292eb3efe7fd85d1387d4b2b4d200866c80a451ea8bbf6ba21cfe490c402592b250837854d9bd29081f68947d0360cf7a250f2d45ae64abe454de41cf6fa08245a034382ae216f8a62b6fe8daf590f1b74c5437a3b0bc95a7c4340db432ee616cef4aca8509f84bedeba8b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdd80e6deeceaff1b2863ec15e038b4d369169c7cd859a7da0ee2cef01ad7c470b38caab2c5d60c3497d161c7b85726dac6158cc79e987793bddb5dccd9696736ef211d2fe96f5c69e2e88988d999e19f4c13ab77fb9fce7e668458047d8fa0178b47bd2b4e02579939a59e0e218f19448994bada471b445a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12b96d6487446f381d21cf8c3477b1a053d4b1e9009062306a572ede0707b4297fd1362cb65de799dbd0aa2a0119f3e000ed0c2e9216dd893555130d9ef7f74e39dfeb2c041e6876355e27bfe442e3802e37068b4856dc0f9d6529d9a641c64703a9ae8e5b2a131753fc4160a5621f68739d23846431c6698;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc59f7180e4f586859b5cba7ffc5b1219bb65b4543dc8c4dd7ca85b5bb6fdfd78554dd3aeacb3dd22d469fb4eef2d38a66d05255bd5ad03026c521e2145bd0d6e75e9b26056849d98da23c0b5a9c562ecb3e755ba99121e2ed99e4d518ddf0a84672c065e67bff829c16b300f3d28a15c5dfb8e28353d072b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h792460782272cff2037ee2b13295a5b11b815a7d2eded4e532454476acb5929cbfbb356abe675e3519e73df493fc3812814457438aa0eef5a0b1abf77bded63f4e76676eff554d67ed4384f663dc3ad9443b4b94de899edea7fbd6d9f2de6549c3a2025191ef359dfe054231b765fa826b80e2071504e36e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h71a48f44761460d0c18cc1f2691ab5229f041ee539e76d62310e12768e2c16dfe2ebe078d903ce00beac3b39c8a02d6277ffe6653e1e8b360d84ff682604ef4841bfe305082d31fa5325c2099d1348a105b2b0d484c936ce27c3e50b71152b56e4b08115a6409878777c7b8b4c6fda27eda149ae23052777;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h29bff8b3167995244a715e733527f6d180fc426ef8f7b066c7cfeebc9d4ba4eef787dd7660ed86ce5641ed1cc6a6039a607e52eff8ab101b4ab6600fc6aec7557ec70713c4ec6680fcb977f3fefddb4d3b5f7be5431914f65c4fbef1eaf206be07d6317dd65987d333897bd2c7c702f71432506c3ed41696;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6f0607cf01ef874c9b250e403d2568eeea118f9d482ee2ab5eabb7b1f68f16939507d9ab9abe51515866ff6677e24535fe63aff317e7be6ea6c0dd0b109f28de2d1bea9629f00022c08063dda3d808a670fca7e5ff9e197953ba4a1e2b36166fa03867f697b805cc5ca570ee98be370a192f316cebb8297b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ff968a46d4818b7f3fe099d613036e4ad54c08f741642310afc7efeadeb993343159653445ef3ecc3baa0b40374a8bb16ad184e12d246187a8a03b6e2bd7d3fd044a442f1b31b980073f5f501b218798d91a03dbeacb30577c8dd28d081665ec57daecd2e9a55a6918815676fd7016bdee10dc30f5eea014;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdf0d19e06c55e372ec3ccd39738e4682fe508e35fb0bac88fc8cd28fe9b45a348410381c72e78d930b15b917a351b2c2a153d073c2c92c9bb116b9c8c0a87d2ae4475e338eb806b5519b91107f45c3fdc83baaf14c3bf2e6ec89e31eef9bcbac6806e9cad5bdfcae7403e4967fe914eaed4db402e7db9f66;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f7b4934e4d3b9a7db53471e62a89d2de7f34974c883ecf03ba3dd408d087654d99d917da6992f88675a2cd9e92c2d709a1efed445638ee532ccf1d037bdb423d79fc9842a6efa6ef9fbe375a53e7cc5b11d5cbac18b4eacfbf5bb5535e79d476f2e373b8d650b64ec0625d0a0ed918a991ab95ac9ad1c5f8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h153b058324c8a5a8177b75b60349d0d6b71cc9604637276b6e8155c727e63fd396048b561c9cbd91a91124c7c5a5437994669ac66b243fa4610529d67e094e803c0760d29c1f5d4399c8fbdecf9ae11eec6aaae4138de0e0e64ef8e768ab69f1f079db57038ada7247751a837e82a819aada35fe4038c23d1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h73530284ef2208ac99221f874d7a5b9b43138d5761b200aceb3a1f0e4d24294ac566fdceb8e99572ed76330f47a59fa0f17aec02bdf255a7dace3980d5071eb952c623d254b6b660387f02e7f10029817748295b945ee33357a5e40517e0a8b8728ed6d091ca1e8f4ed29a2186154fcac51c7fb1c9ba843d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a9b7491e10e46142a8af19e01ca52226fe71fbf9f5250e2c9132d1a095c3c54d85831acb897737380d4c543a559ef5aa15e3a39d58215773c134170705cfc656f1bc1e19fefd62bd98a3b6cc438eb030fc5ac51c0164d7056812ec7368f542a65f02172ea02fbc6746bf300b9c339f7b184c75dc460760b9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5f67372e1723a5c479124c73ac4897f5402d80183170135591a178875811677c43dd4578f40d9dbccf13f5c89d0996bf975e6ee07cbe884478188334e2a0f354861706451b0bba47b773d240af08b92a4bbc1bb98cb49e00983cadbe779a095cee8f6fdc18691b99715e6e8f151de76dbf90105c50cc4177;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9d9131bbf5f63c150c419abd1edcfaded0b49e07007b8352ffd3f74c450eeca66059132033780d4f1dd03ca95af98a70f75a1f1769d469251cb944ada3d736f38b30b2cf30116955cd5e5837dd11d1009b57756e4564bff75143fdaaa4a742f0584f5f90455734309cd9ce306892c4063090a8207393d92e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h106a5c62933735fe2ab08ef84b3200aa32a96b5bb500e9e2410f119513b8c35d1385b3811a4ce930a5c8a312bb9583bb6ad39d13c768b829c1ad03d550b202010754c567a0546cfff1c9ffc9a785812837e2d29079625bf62228ce72394c92faad6afd24d46319e6df988f26cb1b5858a5614952e72f70b2a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fe51f13154ecf09e8cf9a37fecb23179ec0cb097b5d11fda89c5d23d3549585f4eb363d8138068028f9162b6d7402614b11f4986edf3127f739fae5dacdbdb3d6a85f5fc96dfbe907fc4e226726d149b0738e4147778fe84c082ffe96437f0aa6bf1d78fe5c7f635b2155c919c094c7f02e9efb898cc7bd9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h118b3a834a4fb176be5f07259bcd39aa9942e450c9a29d4bd43205ad022abd2e70a0b12138fd9ea9108a65575bf7dd85223124dba010724460d631134ffa0654b7b6d6375bbbaaf42cc5e0b21289640b85f3eb0479b3133a97ee10fb4ad07c4ddf1d2cc2321b753ed4ae3ef8f7bde103bd2c69f07f4dfc6e3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdf1d17a6f942f5272cb86467f5ff366d51c3694ab6a6d9cda80577100d3eab62c6b16016082439d31c6946783fb24d19cbf28f8c5a7af68ea98800121a47805fe552620dbf2193caa42df840d598e8b300dad7c7d904edc7b507c3c81e776cd2a80bc5ac09c255a2e454d177ca2c4bc67daaad709f31026c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c9a414bcfc4ff4761508508f66b2f86c9ccc20ea7c6707678d48f93fee3563393492e15c9be655638848a1332645dd7b9cf932555c8e46047aa3d14d68355804f51f3836dc82c129d1c6f910fd6e3207114dd03a912e64bdfe0d4b1d8ce7654a379e0fcbcfa480763bc31f19fa7cf3c27a15774fe3a5a2bd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8403c0e9440e55d8d94926f89a5658d8980ce9e5f36dcfe4aeb0371efd95ad8eac1910acdcebfd4f2a370f28d320c01e535c007374e379d1b6b8a83c113b6b5b5a380c8760bd66b0406a8a314ae29abc41785b75629b40278fc238afc6712361b4b191806f66fa130041883a08a0118dfb4d94f44b616537;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h118e70b07cc1987402f929712f45e5339a162431be3d8924642c87574bb0e1c0000d90000b374d7c950ecadf2bc0022ab162b48c56d992e771c1d06db45fb53fb3eb8ccb72a1ad6b1caef3356b24d53c66cc2e500f1666d6133fade4581d9a831f5a5ec86adb447cd2933ab723d9f0a986675305a012d8857;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haa2481f7acdfba4bf7617979e2bda08319155d865c92e619ea72942098698638ed36e676ae38fc3c221473ee542f6fc900ae5ab5f8316536accb2904c103ddf8b2a8b0b0bd0afc351191eab4ec61a33f1f768e0f95f2e9a363fc00be08c141e2bc19c5ef130bc496af312b344a26c6f57a43cbfb45969bca;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dd2ff3d9bfb8c284c8c49dd7a2b21b7561b73334073d7d88155cddb9aaba3ea16e47534eaa99bae8ff750d88b2dbbb10e75255b480c350ea9d072f26160df99b49c8a7a609724b6351744a41272a4f4ff70e6fb55f50a034578e42cd84a781b9bc478e8015f8fafabc2a50e59eef9c3e22e6a70ad322a1fb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8a68d98351132fd47ba0669ffe1f79d1f9a73fab91c7f1a72f7eb5c3bbf7b66ff2f6d466f7978111a445356cced12e85e7f9d284274283b0df4610e3b629a9977d4a9472511868ec938a8e39302d6c2470b97c06736abee6b2601634b785a1586bb987bd416c8dfc2831f3667de165bad9bd5072258d2597;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7d64c8c544080d19be7009bc5a14de41a85e8c7cc80fedda4798a0c2c37b0f86ea2123e337a6c5e6d65ea620bacb4b4f40c20e21422748c3822500b253a34754083915343dc68af21103c4caf0f7fd9c53dc55b5b661997b92b462944de0a10006586c0d9cadf0170a773b7d9452313d2558cd34ece231c4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8f85d69dcca5dc7c4e29190da327fb72ebd8bc5be1f3f237539b1965363c0cca7fb7a52cc5956f4af79499d4be4dc77f1dfb78139f7f107c042d612046783da5a52ebb0168e2914d70ab838a8beee9fe1268dcad095b7688dedee08fa45e69fa6dcd06c0dd762e1343c5aa14623145a2b76267214f7e1563;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb5e9207540afe93b1bfd0fe1803ba5dd664f660ccc90b2c7a1451955d5b07b98c75c69ece88568b0b65ec4891585252c0f39cc06d4635283bfde0523b08282059451a445cf2e3438977668811dfeeae06f4de66c5c574c6e77196d8d496d76f703bfcd56c91989ad785742ad9fa829c8ddb7159847fc8385;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7dad7a53b87234ed171919993f73f2b70b011fbd38db3319d042cf37f0199a0ba7cf8a6959b9dfd3897e5b29e00e90ac9b2c031484eeed73c3a826910d9f5705b8817a26a05f97c87dab59d0e6f81d4f4ea2d492c5aa78a1380d4d718e28691b0a0187a25d67ecbf0738f18e81d35b553329fb6b1356aad0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4e8282f598b3810430fe3f3c144c6ae33436e9914ce05473ebef35b027c7c1f398464fca220fcc58ecbd30502ce943063439a8fce89621ae0c1942d46d010eac8ba68a75bd86adac71a2fbaec3aa0effd76a715a440eeaed0b5dc983963d1ad83a08e389f2da800914ca5ababb734630623d64f3d06643ea;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h111b39a8376144f5ddd2340ac9cf9333676083704f98e47f5fe8f3b3b77df2bf1e67cf97819c3aac7be9601d80d8a4ca2312214faac66d324db399615c166f1a74a665ce4fd2a4c0c517044337ad06cbe231f08d7eb619ca7e04c2131479d0229ec3f39117039a91edadfdd5e715d818137692caeb81bf18f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h56a4e191bd6faf0b46b49899e3aadac08dd6bdccacf3e53c1d9ec896a4492465a9bea7a3ffe8e707fa76034fb6fbe5a3e950f9d87754f1a79dc468cf64a68a9566515a5791b953dcd10e5ef461125b3233ff7886d366e8e9734d49e25f6ad9d3e8a941a101af47acf6b0b1d4891e5719055e859c3d37e4f0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h156814776012ffa086c6df96e01cb489188d11af2b77f0d186c4bcf01f661216ec5fa7b5da477aa1f5154f5b2729881e1fd1b5e0c9bde5bd062b5c81d4359ba79478b36e2b6a7b8e598829b471d85376c5710c975bdb33cebd0cbb8be53308ae6265bb4ba5474e2187208457a248507cb94450de1a75fb955;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13e8a4843ebea027d9b49af1c13eb8bd1cfc72c2b252105f889044ecded2b88316b5ec7319326d75f6ce5f782890e4b2ff6d60b8cdacfaca70aebc4436a26ed900286ef42fc04373813994292e5e027a980e4bb0ba5f48d70486c68830e0998e4b1788d608b03522666d09398d320f6456881cdb22b71b5f6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19f7f4f6fb2248f615856bb7c3eb9f24e4aff96adf9ec59b2e8693c1ee1c49e9145414110ae7296ebb7a9307fa4b79c8947a6554fbe3226986d15b78676794fd587ccd052f13fec79a4b1ba1fdefe06171bbcb99288e47e8fe8f0057ae38d4d4a93c2c6adad84faab1e625aba3538560a228d0d0367975c72;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1221b4c7c78ea1c22bb974f03ff6651b6a8255e12949797e3340aacd53ace30ee6c38be564b64316b09d0d89d19725847133e67d78d4fe4dc910a74dd5bb346396bcb9281d249aeea070da6dc921346d3f63e6b4584241728a817f772235d45d1d876e6698ad18531c9f1d2226d5aefe4aef6280409eca57a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'had2135734369c11631210627815cce4df528fcca864527ef5b257a3650d71a2647e83ab8449ad78a4198c0819232a2707028ebe02dd9d12e4061221d5b4413e5d4f9ab9a695a6e4dab92af10c9d3862788aa1f942b55228e48435ca56701a9385a183c5352be6ab14d736bdd86666930d1c3ec6b90cf5672;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h68686fa462b85382ac5eb8cc6c600a43b3d0f2e76de16cca510c0b67773accd69138644007fc9c67c1221c765816ee23fb1983bff8125bf4cda376212f5aa2037dceebac64b1876975ffebcc3ad273fc899806992e436cc91412b339a6a910aa4234cc03bf18bd7f0c05c0e79c966155c064f7fc75908fce;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12d212c8fea32e9a510a653860ea70e0b7e12050250fa775b48235d8680d0a9d9c7984b5e29fd93c9576551529aa80a891c508b94673bdde0f388feffd120579ed830ac758f4ef749065abea9b816566687d61956417d42e0494043d73bcff598ceeb05eaf6bb3fc235cf0dc5ca014f72be0cef42bfa79b89;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e40129a3fc070a644b1fcd2e1ecc92b14ec22c67c06b5ec1bf5028816a17858380cea4bbed91bb4e90c3d7d6e41082c72ccbbe659f37498f846862e7149d4ad92e46e79f5c453ca673d2bf7cdf82b575dd4ecd8acc1da7dab33f312168e24314980cc121531a21ac1fd70834135267ebb1c7be789eab8780;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf18882f9ca5b604e86069f26c0b636f61853911690c245372b31efc1e4030eaf39f07fc154b8bb9963853c8ea3e2643f8621e9d3b046c77e657ee028e1492fefbacf160ca8c63cfe2fe5fb02fa47a0a69cc4cdcf01e6e25163ab4904397ccd78a15086fa035ba3f43f9e9094720b06f54254b791ecb47a42;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he6bc57236f1f116131d9122782b7ad8cefe7f6388adb08fa315e6c8aa0ada492746f7e3acc1303a346567dbf330b3168e926d4acfd05626a84bca099eac73ebd291bf11dadb34d06ea9da5849dd4b0382afaf0d62adea641ab2f80aa8d26f93e66ed56c33eb75f7dbed3d270cb3cdf8105d4818628483850;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ce1afb30e15dd3d89e1ad6c14fcc59d0afe99e14b1d03e769e086e6d1781db2f3e34ccebf79fb70f595206d957cf306c1a33bc86faa15e6b1a646237c96b04264a1109f9a43db08ac6f727e8750cc0ce71b58e5d6a454e5c7a1ae6cfa1fc918703d43c1cd02b34449055adc59f56654c6f64e91ebc4cf073;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha162d789d523320b252cfcbade86d9e59119221676790c8f32014966f4345ef69d0d093ccf4cd8689625b8390a96cd02c2cfdc77edf8d5e9505a6b84523fd4ab5acdd8623b6bda0133c94def4250c28049e3b430341ef8df4a8dee52f1c856ed08b5dff5930fd76d7bd0b307bdb708dea865466d45270f40;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h139925efb62e5e97ad7d5647a8e3f9f52b748ee3091c261261a63b1074a122c2c92b15afd9939aa0db5983e0be35ee84d468db4b626a538ed53aebbc3b03c1bde931d199c32f6d39d95098049be918a0859170091a95dde35f8a770dc5cff30d605fc121c0a97fc5cb0872a8ac65c239c47d4d042e9eaa5f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13e9407d5896aaf7ba2d1cbf6dc05d2ebdbf1e637db03147a78a5aebe82d07b4064c97282da24bb1657e0757ff4e62cde4df339572daed07d615e9a6a50ea3d840ef1f3d4cd4ad66da202f8774b840a30300fb8fc8670e5620bff8d862a188f707cfee39e6fcf592f4df688cc15946a4450af2cd0aeda00ed;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1401a6dac9712c727fdfcc5f627ad9c1ed252a1ed9729543f25bdd70c6a075cf39fdea478a4f97f0852219d0d347b4d39c9f58ee26a0cd8c6624899367d57667ece6503ee2ab11acea2d94381a970a781802ffc35bb1f8ef0826c087df8117e7ca89ca5fdd4616a48568e3b139a1d074c6b8ec0c5398c4e8d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17ff79a454420b162d1ec2573cf0e6444456aabdf2269d51833efbb4b30888dd7e7a1a838db9ffffb5841a5704ac8f1c25a4f9ac9b8e12c3c39ac677b766b1659902996126ee30ce3631a2c77e0ad831bbf14518ab81b144b2e659a115b95289d9a17d38a51812600692600193e181e8325d287de233f0fdf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h751039cdfb21020bc40910d829f3d63d778d6a689fea89f1f96b7110b3cbe17f78ca4a6b9e820a1a943fff033ab3dff4a18864b9c5808b78546a74c88bea84f023c4c15428dfaf5a622aa61abc3c7112da625d6699d7b277ede52827fd875192ac7490a9aaba77f288e869df3556b4adf05bc0806bc02e99;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a376844e76da7b3eb4466e77d18eada1bb75c1c78d5e46349757625f16b215bcc9d6ad999a57ea378d7451e4f31b299a7460fc5ecbfb22e45bf49abee3b87f06b252f3c41f6bfe70151a2cea831ec4c10c47d0c9cd10d21c80badf52eb5e9e653efef27cfbd0aa869153dfde091c22c0403b3829214d38bf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ff89a4587475583ba51006053521e5c4f820ccfb38be89abc4a6640da16b55767c4db1043db79b1afacb3fb17817f230ba0b9df259040889e09d41e842327241e18661c76fcc813b3ffa9a9a7c8eccc3f624a95ee305a7c2951835882be3295e8a42c8fa207d5f6208aeff9648b47a075e1d92cf9135a34c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16ef040db52cff979dc949186a698a4f53f59cc92d4e1eb19e307a70602722aa2dd56a7d4ea44b7c2e3fd8205cce379792be0fb35a3e99bf8b53cbab405e4a98007c1456ba76cd46ace213e4546d80c049497c794ee049e3127f79688783e4625d8e01a0501077631ac02f82198e19ab0d6ae92b3667cb852;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h128601ed9aa83c359ac897fbdfde68e0efbc49327b0e7ee50dd9604df4ed23d4996dce3fea1c209a5cd223ddf4bd44fc3b4d066a18362d27a471811525276b339e6d1b355cbbc4c77c2af160dc09c87f33f015b60adbda4c68de024890d6b9e89754967fcb13205f804d2f50f6be809f05650e85d7705eeb9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf7cb58e6334547c514c8b53799dd70e290147a51beeac8853dde5ff5126f838f1d1819495a682271891028a265d72c1f2fa4e7423bd63bd85eeb259780e185be4410dd1c2ca6b61834ef894145e625aba87175e09574aa4a3cfb7fa573380e6ddd215bf21119b406e966186c0033ca6ae3bc1777ec91fe60;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hccf45d2d2909fdc59ed37bd5146e7960441281445c23a771c363f3f10f37ea5df37fc499de042b1b94d6c6b0a3abe95aa544159aa620f6dc2f91aa4d214e902ad06ef86569574debf4c4e5cf1b900fada98f9bce23a427cfca67f7d88c3290e2a248ffaef67d55831fba05924a500f5ad0ed7198c136d8a3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h45d2cddc0030c79c8c1a1217f313751d1e794936acc080cd134145af3cabb738cbaad7c6ac4920f43b18a21fd8f93cc6cad734a51b726252a203410e2a0b8c3ea5f44377cc04fa8df49927d1fa6b721c291529c862953bfca5408a26707e7dc04b68b635b16a4e7868746f9d506867578fd18a5251ea88b0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13768e808e1b8c5d47178c1f4224044b3ed249f5ce6ff062784fca1170c16605c14c8085038f52fe6efd583bdea015c7c1fed1b99a0a6b44b5a0fedfba9740a58d63267dfa79dc21d03646fd2eb03d1cf606a464edc105d182b9a321ab62f67ddbadcaa1c4ea79c1980807e17a83b58907457214c58aed57f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a8a875835144925609d7c844d8a73a4fe66b254946fa5388daee049989e580b04078eaf7e0a6ebb3b04765f8b210de73eaa9fd82d77fd4fc1c27a9da0cdd68e062f91bdfb7ab1ddc8709d67c196b2d6de98d5ceda71bedc981f54017ac1ca3b7e1d5d270c3fb212e21ae16e1e9d9b2f27748b16ee1ce0054;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1298a71baeda74b273660ac367b42121c1d310577e5eee4cbf81b018702303dfa928cb97371e53858b9d5897485f32d246008b8134bb2527bd01331b996cd2b0bc53ea742af71ce6c22526ef71e4ee360a970861f239b029d1ea9864fad66eee4ad16ba0bcb81178b67b24a903f6c49b67a6e7820f5d0d0bd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h196a8ac2ccc9dae953fad682816436d1cc9d08e67541de4dff689851b8bc021b78d03034fef51e030df61d33eb9fba499dab026cc8f0a4d2068e532681f5479d1b95d68fa8299338fcc7bdadb74145d2f2a7a200236f24568f7a70f1d4c81c405c5d02c5dc6466b4da8e10ffbcb851d47c56ec1cdfbca1860;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dad491458f4fd22ee5479dcd0d1590ee8975ec5519e29ea8524304c76d37eb8e90748246d8469d73bd6c8093fc445821c5ca14c8138748acafb624f45fe90e90616567973721e3b36a45acff21ca9ddeeb89a95bca46b912b8547775239c283457cc9c3d1d6f999978d38c39824bcf2dd0507358d6078572;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5141ec61426c7435d5045b439582a7791bf9b636f1366e415d5dae93c0400c5a81040f260eff74328fd5c5912d02834737b4a5b98bf74295b4c67aad6aecff5a1ff8431a4610625d4a9467f16de5e5eec682809174b3954b998b0d26262732f4a3df8d08ac021db1b5ca6463e8bce8bc936b150ab40d3325;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8e75581d7d128858ff64eae826a0a3e1c1d186381f61f1469732c18dbd9c2be5966d920cc115e79dba8e046541c1c342820108d6021ffbf38a75fa00e6572aaad9239fd26a066f1dc3c177dd32155311b8b8cda18687763bf24039eababafa544ed503afc77e79432698d230f4d1e16dde38893a0a1c43fd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf4d3bf4ee0d1c24eb6db54d3611af8c5f7dd32749783783c4ded1595e0980a54e5e73c01b319a8bfb409d090aabdd0d7580bad35110c1ccec3e6bafb09b8489f8e7e8b409a5b37e2232d34ade1935f5c15ecca9cb2f0328b306af3c7005a9cfaa284b88bbb511ca3cb44d55bd1bb20ac6d4938a16442b0d5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5dd933ac0d252d2adfa99b8d40af97c8e6879d827c786eee5c9fd17a126e092e5f7140f59c4153927b56c0c07e0e76169899ba19f38ce552b5ca0efa78cc17bcba5ff93b4f8dbacf9defcc33a8c4c29d15ee69d654a54a74e920ae07cf8f7b73ff653c3d9c2960026833ad3eaabd913b26bffbb05dc4f754;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14d806fb3bd8d09b4b9698644c9bf4b50b739bbba764ec1320a35f8c58d67f0d8995729dcf0cca34ce9fa103b5a9b5479f502ca638e47edc914196f8489bbdae15d5833346de33fa719515b4064d9ce36ae5a10c53c22322583e31925c861aadee8608049c1958da1179b2e9461ef3d2b34eee9fa5e290e67;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hee6e4a7927a43c619e4fa86b244ab770f48d86a41c3cdb8de11e2ecbf1ad1258fd2b857f6d467d4fa2e28269234fc1ae8ce8b8754ccd12eeff526ea6f2c384b3aca78c253007e7aa7cb46ab3bb2deb86013b768fd01a73b303835caed42f4337942c35612a1e079dc28c52592a45edafa86b03762ed15b9b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17e0fe9c526d948f5e3016a584e8f22545362906526efa1338f6deed1bc8a8a860be2648fbcc4be09ac8eb9bfa034ed81af2d25db49e2779fd8b52a4ee13574bfa7df053a9a76b3c9cc9adca3c2df5a64faa414e203b3bac867dfdb4c50bbe289c992fd6170a3d011e6c0e3ecbfac6f52be0a113f67a4f4c3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1116de43e6b7de59ab2c163b9085a748e6e46f90a8e4245817c977d080d3979b761682e2f68e8c6207b0900dca8052ca220cd284d56ceb76339397adf2558e7126c692127634c7e76336c0d92337fc98cdbc121b601f60ca49046b9a831192354e095da9f9d93fdf754bb5d0fdaa040f22e7871ec7f57aad;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1faedde909b9c753397d7476884ede43e0137455284e5fc0e82a75fa1979632fa23e119ddff4151090364ee4932505dc1f19a80035d4b989e0334853c7a40509c0f714c34ea7d9a2f56902a46d6e4186a1990081b4fde6e2fb2ccf68cbc44a8cac0d77901fc150766a6e51582e01cffa680d36e33c6832ac1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1717e849cbe3ca345eb88bd90bebd54bff401bab67f9c89c66eedd163d1ef934a6775518fe0ee7f83d7f5931ab1217b5fe965fda3c18015dbfaa147e7adb869990de26b6edd4cf70ec7b967e575d3b4ed6ef188fd960c4d469fa32d5c560beec4b3f588e9a9d17b27d2c6ce97cf2b2b68f954a2bbc0f0e8ca;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bea6d7f68d1daeeca0c36cca097e06931fbaaf613c6d2d45a452b7d08408cadc71a5dff39aa31faa95c0f60ff2f1032405950139ac51cb3b12e2001a234edb1fc4dd423d54047717d29a859b9a7084dfa9e7340d46947231205ba200515a77df398a17894dad8447f716c23f4a7c1931f47baa1c5265bc42;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16c43d851bb6c46926c3373d331923a1e409aa5fe725cbba73ddd8d1a790affb33287a957300f6ef66fe46a9826ae0d27534961a484833b24081d7c3781eab503d8810e9ec945a2c5817db4aa7f38c3676dfac177129172fa80f8a208b919c3fc4743f0028d14372d522aa6e31797d2b84ae2a49102c94fe3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hda4c251a65bc3be790d58704f816e60929fefebd3f7b24c17d163eb9dd4550a8e53b7c1acbce267daae49794b7fef417b6693b14a9fdc7f6c66c35632f7fd01855bcece53b64cbfcfbeb0546179c9c7d64972a37341ae4896a5d018ae07b7d52ca67d8e327711d73b94f0ec6476059d2baef471f8239300e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h569a975d1e4a9509b412af1733b0a6e47ca91d3dcf75056225a0b170c1668dfbae367a43b1ff334a3316bd873bd85920e131a1243c461373a9a29a33868fb1302855e54f00038625b3d78f1fd1fcc51faca4363e6127d6a2f1752d2addc8e06f7d2d32410f97829af704ae623948eeb9f0f4b661464f0713;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bf5741cfb267dab6e4787382db5ac680c0059f7936225c2822cc585445a7a7c27d6b2b65c0343073cc77cc5ef797572fbb56fa48bd23426b7d0e1d0eb77a3d40abcf32d1f2484458ac94f0e1be2cf13ca2d78383d8a3b658ae1adb6aead093c5a78fc7038ded99ba0a365f36a398c19dac0ff6f859f3eaea;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h88576a5bf4d52d350f854745a42cca03797a51666dfe0b671095edee979fd8f2ffbd2a11d643740ccaa0d90db3c13ea0ff5ed0c67af4ffe2cdf06248a4e81bb2c6e0465d9d3013f4e72e7427971b23b3753d069061fd784e03386f80b5753d36d1fcf7a5c324bef9de57f8e625473a978cfd8cfa156bacb5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2a066a9cac61aaf4488ced5b50f93031e216f417ab867df693d32c98ddfa4070576f029e29023d386031f6376449423803e439409db32f8932ae73476620737d9fc7ca9be72465020676fc17e711e6ea11064a9d01d5afdd376d80b14649aed307faca13da8e7508d4d31ed44c0a340f1b3f551ce47cee76;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b75957eb35e4552194134d70c55051b0aea5beed45d9eb346751db0c4258b60f42327e69d0ac41c69ab13b730c5df13ffbb7d0d01f3fce5647f55d7a55172a967ba0c79f4770e6f8c58cb7d2a75d0f68d4396c18d88cee32ec1c282b80edaf9dac6b3ff62d93ae67872e95f7fa1cea620170f686ae1eb035;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h122100c0a09d8432315489c0e4b61b2f8463f032031fa6c6d4723f0c6af58f32ab485f5783b20f4fe1b1deea964aaabdb6d2a2ea1c0a178e138ac54f4f3b25b18cb6792eddfb7fa8c637d2586f5a3029c4d3a62127cf8c94c124fd67514257bd52316689c3b295a78e6105274fc85ec93e24e08daa7fdafd2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18a74bea2393d0ef19c2e083fe7b38c4b0d6f853273e646827a1ab58f494d48649afe8bf55019a31cd06543b7ffc8e18790302297ff8bf2ddc771299a7be4f22dfdb62d0a7486971f197d4a372ec95f0d968801c0193548c1dc2aed5630da30bc3dcec067c04fb87cdfc1ccb49ce719effd3e5b832b47cab5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1945778a0011ba8db8344389428329ef2bb38aba691e3708c4299772bd47495a2884d6c8d0228d82b08169e34be3cd530b865531ff2732fa0ba16d8230f2c6039ddb7082b349e453b94c97e2d26ecd8e80560f600b1274d22b5b87f3030484bb1421518b7fe526d6a2f3b77b7779fe490abb8f1c865b205d7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dc61022793cd636fe62e77349452f897088029fa4e8f1f140089f4c3d611a38093e16697bbc4e4124abd054d66fce6f058f6507eb206b11d8b028c8c383c4d1397cd615d712ef7d9d309215a58bfd8bd57c478ac3a9c7a965c0fe0aaf242375469882a1ece840c2db2381e6e302e8c46e08ba182ee9ca493;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd513ee4c4f2b21f559ce727ee384db03dae76c0917b3321c5763bca43e3ad6908cac30f77d6cb581d47b9d95f771c17fff61f5d8a48c7bb3d64161424546a5747b5014c536f14c3414beb4e5aa377c2b2aa88b97ebe9c1bb7513c78a0856691c3b8ad7185ee7dcb5abad10046c3cd1dcb62dd7b3067e199f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h104ceed06b1f619f4a136d4c48d135f3292565e7631fe359f246c1739aedac3c8ca004f954666f2be2bd4179950f3881d47396ec0f585307fdd77ee1bf5e58b5edc64aa4239d9f71108a211fb68acf706fbe2f48e77759d3a835273b5817a0d3fc290db23fef65e46a70f4f71427b3bcf61e4896af9debd72;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10542ceb1bef7bb29c9c511ec0f227640a7700b6fb5e43607d8a00f8866507135c79fbc32b084d259396c9cbd74376dfd73467aae37462d1e875de511ab9a871e2759dadf4368f3057777995f97e1d81bc2d0148bf53d7b6c9cd73f52693ece0bacad68014ebc75b3d24bb63fdf808c9ce76c59eddfb0cdc0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1237b14a2feaab497ef250519561a8bff08e817844849fdcecf483b074af55280734019a4c4c1a19e4781f0099a9dfe68e133a69bc71cd5493e3a38a78569dad1de6abe1a419a825a2a6efb41a25dc15772aeb25aa13fb73c689c72af52ec3a9e50d81c6dee32edcbd171c567042551f23adcc84d08874b66;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3ae2257afcc7e3f2b5385db00d0720bd46cada5db08a4fab195ca3ce6dd98acdd7b517e14783816a8eba0472924255470ac186fe1f582d4bbab9662bf11e299e2b5cc57a8dd2d28b7001b6ec5a561f5abfddac6ac9d5e7d52c90fda3885dddb9e75c78b004ad4d467660af462b6c26d542643510863bb136;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b85db718e952ad6be1852b24730b3f3ea329e7d2787a880de7dcf628c62599da2bcdf35887a9b1cd75bf993d919b6ff42a57e91f6580c59254b92fc140d384ce102255d45352d3618dd745150b2ea9a58de6f958d5d4110663b40f86448c07373e822a7f70c369cd868d23ee4763997b7ff5859084f97106;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h84f7d2274d41bb84326e979f8573aafbbefc221e94ab64749298fe1839b642da7f455f80ffa8d41ab7bccab4f16f40c00abb3bf98cad11f9989dfa00f002aaa56046c01252312d8e4b6562352a508be18af53b462ea1f7b228a4fbcd8d38cb6315b8151f55806436fd3d97285098572e7fe49fc3ca618e1a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h558fcaaf0439a5d2f6751f296e507f4827b2ac2ec4659ae1b58a54a322b6e2216a4243405657db271e29299c304615f29b0f0c4813216ae7e4b0bf09f80cd65774c6e9cb8e7ab7011c995976f1bafcc2616afaebc772cb3b5ba099bb671620c3ae9e584b237deb54734d950c36ee139384edf597c0592a36;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b07287106593e475d73315ddd8ee6a3dfb0689451088651807726124faaab9926b2bc7f5227f2cdd07b74c85fb33855249afd069ff58a187f8cd6e2b3c11fbf49cb3edc2a5f1ff45e6fdc2ead834eb05fd7243b434d48f9e1c7a8bf0cebaeebb91b9bb278784cbd7829d0561ff6032952d8874ee112945fa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h33597ad95e22cc074357f101855896d16126b2c3cd860708feb6dfab31f6d607eb00e49e8c6f67c2ce7006ea5047b7089ba83766213cea82b921e5c779040d6df644284f5e9e3209af52aeedf0fba23b4fae80c691bcb44e9ff8e33d74de0518b10a5bf0042336ebaa350d015a2430b3bc81919ec7dbe3f7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1443339c3fe7d949ac0fd43e56b0ce2cab1381e5438420f7c133b51a716b923ee180ebcf98892f5487d3f58ae75ee414cffed1007b3761641fdafb7b423bbe08ba1819c0e0ffcbedbad1cab1c0c50c51d33a646b5d7bb95831973eb9da85c4be149ddd7c8f6d678067ab131d3c44b754300dda90008c81a60;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1561d63d46f2d7ddff569b19575b3551e02fcee831e36726a9cd578b0bb4ab6d86770cbe680cb896b9dfa32137e89aaaa12b346418ff3bdaf84575b38f52595f3717b7ee939b480054596806f9764daa5affe5c0f7a1c431792e5d87981e529b160f2e9037874c26d6169c64534554526f27a3e8bff0e06a2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8e51c84b23bc5732df26112e0949da69449ce634460655a9555df13e4ebf6d3d76fa6c6554262b46ec73c1a981ec970308b22ba2a1f96586db60d3e3def0cc9a0f55aa71a2e967dbaf212b2bed0914f47982dc5e0e6fef49cf62229365891647170200eb8b79fbad30e159da09b3ff79e051e950de3f0ddc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d897374fc17ad12944db793bd6438a4e4fab5e05a88352374cb6bdda7a9f8c4c52713f7ed67db2ee2ea4ccb0955ef82a845ce5353d4ea83fe585ad9ce29c04db87893ab91f4ee180608f3f7920dfd0440d31a88a29ac78350ab781dbf87c5353bdc7ce141a3ecb2a071219a3c6e4eb2b7e247aacfb11313;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ba382d896f0b0909ce7ba056f98ec14be5aa6aabcdd199c6621af259cd2b035c43875dad99f871fc0c3a3d834d907c49cb448adf0a5eb221908884e0ef5dab3b647d22c318543a7dbf2176ee62a36d71431de84e2c9764c5cb3eab3d33351a380b7736452d66187c81bd5056127c6276f9830752d2dfc44b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17c6f3a8a61e9e548e3ac79c6279448337d421b059611c228ed292bf484a432def73e001799072c77985bddfd1fbddb24a0afcd906a2fc566fd2a7b6311942117f42dec25871e90ddce5a38dcfe2718d722ea2a2cd0292d42614af3f47076127bd20a7caf93d7c3efd26386e192372c2d6b20586c9a827ea7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e09e2929b115ace3fc5cfb045843aada0e71acc2ae2f38381c156b311e8210357a67fff0d18ca03b9d1871eee87a2cbbadada1a877a7d7ebdeabc46ec6a87f2ca002a3f486f8946a1f36a223eaae60e90ebfca0bfd67f4ab59352988d8ed929184509446de1de59fcaaf08bb893b737760e557f168b10ab5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h71db04491dd477ba93ed4648f99dadcca4a4a5bff1629a8afa372278a0c2c33b5bad02bb60dc43a0e62caf6baf7e629a2362c2795dc8d6eaa30c1303db709e1c1d95e9e5eab66e35fcd54eea69b6de3afe1031b0b97cc3beba985d3613a252148124bab3e2a1b9835a875725b8454f91a9b10efc0ce8d4be;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha9c7273dcfccd548f8d2bf6846e75552ded41b688ccc5b0e51359e20c78f3ee7d98398065cff85d54dff9c0cd338c4b7b16c283e19e643b6ecad9390543e6f362022e5ec8dae3afa01c88e5ca7312376114c2e2b2e13881e6dfc08da463fa411211b11584c15a2bd41fb6be3c6ba4dde76099074e2cb3e37;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fd7fe0fec3695d82306df4291598ab7ffda2514b80590d38ad1024ebf56c110f5b4e71f8dc7548f2d561a3c4b0ebe0c254ba27c585a186a088073d92bdfd3ef7395b8febf4f30dc6eba484b9d897d64171e0f2606f37fef01e9589ab1afe79a211f587f145fb7c421f6b9a868f28634654d8ac85c13d01d8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19c8304c32b5b0a501f9e76c374ad04ad06a14df514dd53ac638023e63329546aa34615b7a6ec646d87aeba8d49fc4fdc0f557e246d07b40401a158ebb70c130cb92ddad2c1d859227b62e8e6272447513b02161d0dda6a2576198fcf689cd301dbf798f123b05a8b0da7761f651ce8ac5fb70a9b449b5d12;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3c94656df632fe3a0cdf47a0501def522f6ef918d6d45b5c635e2cc92f387784ba4af4b8c7ce2ca6a51f55bb0c59539d374b59112413b4a6b006de2814216662baa30c98718aae586c97ea2ec613c7c9f2a808dcccd05555280cc1b08c12e7a786c087d472a2818899a300e4881112dbce5fcea7442ded36;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1506ff6985d799d399b8e41b521b7a320e5e2dd465a6ddc762a6692d878ca745553ac004125d1bbf871d418addf24f54c4a30f9f4dae0eaf44c74807ecc3e8ab2ed76627e64e922b26921dd76032c1d67b11887b86e4f16f3afd829015ba16bdd5d6ed9604904ba9dec77f93f2f81036ad63794c17c760b94;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19f33e3a05c331bf0414e922fdd19feec40c17630119923265a56ee3164668e363ca986e83b3cda7fb56c3056f94071c7cdf5d9e6970e0087fa152cf114e3e3f0e2b63700a626134a8fc73aa10cafdbd000e98367aa61b68e991cb26ef4faa950df656d2ae0ed644cdf3f4d935a823b63860308fa30ecc160;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbd33c8d0805a4efd1dd99d584839e4231bf17947266c35293a4ce2eb77d950de4316a6073b2d84c0e5030a8854c74a9bc796e915efb8d474cf1f796be3f7c5093770c5a6253cb94b265586fec3169c36a39fbef6466ba729254cc16312ac0d7a466555e9608dcd749f9593b1fa7af512f6fbd014cd23978b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18f119e03505dd400c4a75814d87f7f50d15380210d96644d7962a0acee37d43fba902494e7f785625829d91880c223d2aff59f49f7e8018c447c710fba2dedec9de2671d8a8d0952c35182a8508f8fced1259ef6c112575aefba9a1c365aac7d4fb444e8a248074a0856613f83bf1fdf31c358dbdcd95c7f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cc24bcb7fbcc7a784da7c4df613c9a62ac295fff846373a804495cd182c2a4203bb8f9d5e793a3f72ac3fabe886fe8a18a80ac1f5c4b8dd0d3253a58bfae876cbd8fb6f1cea8a63b51dc44703aa07b57070696d976038025ce9ef533dfef7749e813a2dadcddb52e8483d96de89d94c7518eee2be9f1d409;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha5ab1a68196ae8744306bd2a80ca4b607e77503f118e79c0e20638c5b628fcc35ed40432b1cc633b608e0c59589c0c9531bae08218b0de5ce2e219d7d61e1eb95984ddaa2221b35fbec459942bfa39bcf4b77b09a7fd43f5a339504615fad7054a029c6d8d87cc9964aeef3bbde78805092b853018bf6e7e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3e077483f983dc7a1a259fe83ba1c6370155c87b0139f1ed7aac782a3849936dc73bd8488b09d65a2547f45849324e325678116356a78f4b039487a3819cb66910da476893e5fb21d223d984124939b18e84d091f125af0777479a9fb70460e022d5e15517fec8bc33967825dfce9c85a2262deb736ae3ee;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haf8d993e54c22951fdfb8067369ba44f8d0ba9e285254295b5698d2bf7ad2bd621f607bd8535e0aefc7fadc2e3dfe3a4337175c5d064ea8849058d34100de9328e3c1579baea3a655e5fd48d84d40d7754aa222f61881024bf2676d6e8017fea4340dab35d8ab16b63b60e0f54f7642df57fd64356e581cb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5b3db6212c870bedda0b46211041c410fbaf4d30eb98e27b7945afc12c134ec5c57e12161528a5d59fb82b3f569d7f6d582ba6a4c5c89f6b4552db90b2c74dfecfb8f919d81f000beb891e4df391c2768e69fea575e6e6a366db16c843937244006d01479baae22aeb3f51368b06ea19e57400e321124268;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1429b18ce6aa2bf8a5a175d5ff682f6144a16bab3dd6546658f897c5d49484e88edbad9af51fde68a2c86d26696aa49eb6e7da4b598b84e7397abc325298fe8af9571a3a9b76f8db5e78f04e16450a950f951638859d924efcbe12e58fd3a540ec5283508552940dc92d67c1f7fc497ca80db3b00c7bca117;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hef622b929065eb0934fd7306b6b33e04dd22345ea4f4f8000154c52980463eb344a79a3427d5d66e5cb442ff4c10f98247354d6d218ebb4ea72ea181db25585c672a6e46a0774f0cfb92aea63bc9ddeb6619632595f3c078ee6c100ff600775090146f6285f468ad5ac31540bf03ebe326ee6cc65c380015;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ead09283530ed4df680e569b74de1a07c26b23e477fe8b2c524126216ec91bd2810264ed9828246d6d22b9512eacc100c3dcfb5e2b75f965a4b400fcda4f5c4c5d9a1b4925d5e9d22ed1ecba8204a35f81ef117a7c433359e35f65d8f2a7bf68f129316602b10baa0729bd5bef46add4a013f49f3150662f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h157a2a52f036ffac812bcd403630d8e7811e9bbebeaef713cf387c84f796171ca0226b0ce6bcec98c2d5592b25ce29cbdf7afa232e4780b25686ac1b64bf4543f84db6385d32a40f8125912e278b3db6df039d0f32d436d653ff6d701016f6b68855c0147d36bc39c1d52a1e06258889d50b36e7768ab7a64;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11cc99e939a5a4e9a3996e130dfcd0eea78407d2649f68574203e59a9cbc9235fa8a6782599a1933d4447edc6b3fd44d0660c7ef3e614bf563573112e180b168875d2a07933c37c52918e72fd44f7316034b80dc57bdb65cd25d18c46fa1a8f958392e2c3e00a7008d2ad2737059fe7cb46127f3b99a4cafc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h67f03332f74066023911db2df01176ce478e645a11304eb35240f83c43078dee4b11f31675a08246db69d6473b29226fd570a85aa353c42572288cfda6cfc7fe11f94eba0dbac5016abf9276b9880b9d02a6d3b27956a79a1477d74d62160fd72155ea369eec33aa153264bb9e5b3a5a22d38fe966f5105f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cceecbf56fa48a746b0d26421cfa242730c11a31fd60e4d0772f28dcafa949656a612d35e0edb20c59c85ffeafe324ba45a144c2be60a4c75b946b970100e55486f01b608b9a18ffcc1ffcd9f11dc04d526c71daf7748cc9c7036f74a24a41f5faa92b5c4b4569bfc6ac12a9f192d5be743ccc274c872424;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h911f816d20ea8d45382478deea9c500c7427726c9ed595965818133af9ee47be301816b84bd63f2d8c9c48c47566d49893f93b14d6ee771a2b95022411463c1f008d151e7dcc56540302ae9537f0a8268614a1d27c2ac7f1b8ad156d2ee237b0ca30038cd9a6fb609266a58859a48788dde1f1f697cc5d66;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12deedeaf2402c8881834274cf6ed6d820c9161f336e8821382203fc3e5d7387bc6933c9874d31c5542e365a6bceb17deeddd2840f00286a0c1db48137641921621bcb251c39f7b3d53714fa52b5fd90add40445b5e658edfa398c7c3d520e6e891c84d071f1ac0e6b17b4208eef20fb7ce02ee0329caab47;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2b1fae99d8ea68a79369b7f3ef48770b9d6cf0c18b4a416e906f71826337fc9a502d1943b3dac312c6494630d91af4842004d190c7847eb80639e9b044bf4dfee456113eb327507246acc8d7a53134c77651f240e635724d5bec926ec6b18a1f1488407873125306d6c19caac743b4a7b2f31790ed6e4240;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f597d2aade8c0e31a779b009ad91d195d0200114b57989ce1f6e505fc025dbd67fe2fc5dffa3c1a176f6fb6ac0863c861f40485a3f3ef3b8e2ec7d145f9cb78970b3935c179dc92c1a26a82783399bf567ae539b7717a230ba6ebaaeda214f1e8e8e234ade6767387ca471be64c6b02c8e447023312ac0e4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he3f81c4451c0ef00f1979d92ccf6e9b979e23bf1141675083f4a674182dfd82f4e3eafacf79c818b27da91f737e7fb5ada6484efdd96689490d5894e23ff869b5556a3215cd3ee732ae8a07d04f9fd4c9bc74007ad0f4b8a23d0a471630e0d73ec599d70b7a89ff954865678ccabb772775fb04b3fa167da;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hed986fa346c8844d6aa7f324ecef2add306090200466ebb252670e1dbee25a7aa9db3dc3b7d1770a8b885da5e5f8a6acb2a05d21e9ddc19f4982a4dace976647105b9bf9e022ab22ec4e318cbe0e94db81f65e66c7fa907dc252936e23ec92a8d213fdfa2cd1bdf8851aecf7b594e6837b757f117b3046f6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h636231e35d84d5b978bf4c2e7cfcd75d53018448bd416ba792d309eb505f55cc78214195965870e9f0594b07258912cc826f85a798810b3fd4ccbe1eba964e80cd50cf42addf4f8a24e91d8385a82e5bd6f11c62ef0758343af88536e46415b6680666d010689c3a272339aa6ec198170cd19f0e21ec44c1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h157c8ceba8b2ec5572b324a3b20fa7c3b3a9357b23ce1f13f09140fe3e5b214975e39a96d423487a14bca82b103b3894b123c7a896ac564f0f660e04001399b1a5590e7d1068ed64e7d2cd7b8d083490e24f4051e783f7c7680354ea938883092e5820f5baa1d23cce59d9a85555dc7819ce328389d9236fc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11fd2a24f1d4eaccdf704314e1cc08c09b6f67b97a7e6d068c36722120b208a691f96ca3f9006cdae74998be68be2f2475efc81e995d1a17b40d9fdc0c948d30e8e61927d3ed361fd903d365aaa076e7d68b49ae18bb08f4d84b6f50fabcbb15f877e2c04f54d307fd150fff4a0212450d7ec2c3c77dc3791;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14d1492f5e9f675a4cac1aa9e84b3a4d1c996eccf1c0d5373799100b1fe5848a30ec2458057c5a0d0a945989501f6129fedd7e18c27db8fc270303ec5cdb0fb4ea69818f502754f130950cead7581235f2e6b48c511b74455ca3a0ad039f63fd583bd14edf871f6d074c995ceab0da0449cb1f27e31718768;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h313ecfa6e659c55942fdd2a27d85b1f4717a8df91f17dee1faeaa423722eb52b879579dffbf6f0efe2f621525ee3d42c8786f185dd8ee7fbf09c2b709a70d3fb483b25cc2114aee6bd39ff50877b62111781b04479ef9fba98035858e6829d34fce8aa92d37ae64d6655b8fe9ab11733ecaf4592bd76cbef;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h327b961bfd5dbbdda79b333f65438493ea05b81b51df7257d140862315f452330a433dc251a79d3656814d4242535a58b9357cff11e4c0d62d69b8be5ebff1a958bf7f79259f2d78999cda1d504bd0a7df1f33efaf4889b028ecdb1e74e6312c57b541ea85ed5d7ef9168f2a872d386eb82b77676a2012d2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h604873444e35c543b7f226e19cdca854dea44d5f64718680be3fccf9444d97d456f0778f0dc9004211308e06a27e4efa595588c96965afc79be0981eeb18db7dd230ee938db68c06f22996979f3f21282e70f0d37c4393ef555852e525bf1af527e36e21bc2059d11a4e49590f999c2ccf6754800aaa024;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d75524639536aa41a343955512bf5b41e760020822ffb4702b9d3b4ba06f2f46d81d93d8fe7991dbf061c141e941e54b1525c0f51df8aa08c65da01e474e5bd8f5c618cedc35989c445cf225e9792bf611d310c495cebb3982c1c7e9e09920adef4a68036531a161201431a56ebd6dac9fd723ae9ff21985;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcb43b419a93d6094d7a73f7eecc85872d909cd02c2bc1fada687c7ba822eed5bb3bdf175f1e8a9aef890733dd9c58d2631906b7f4c26a6fb37278d7faedf6bc13e09d97a071557f0a7c6b14ed1bb40f15b936c99d35a2e40784901ca1ec79ab5834ed23dfb6727eaffd716c24ef683c908e51c6dc2becd8d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h142ac02a8f83f69df2257f950ce537972357b2126cfea70586d3454b8ce5e4d37f5f8b9100511c54a1df99fea9bd029100df4d311509bd2f6f2f80fcc948ac912b87cfbfe76111dd23d57bf4c212dc2b510e162835ee9c8a45cd9a57e9e2ebc087ee919dc57fe9e41e15e8208732f94db014bb999b2aa3ed6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h192a891216471a4b3400995ba7b6966dd733ca02a343c4f08fe189562535655b056ff000420a0838d35214c5c8fad6852db7357c3e6c7dcf087fde3a79194e0b8ec0d1997d5244c49536d930a8a1a43f7c84b5714058b2c6f402c18b1f62c7b143477fba082f61de12d12a92bb64ec387139a792b204dc8b6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1388976d21a64425fdaabab4f44dab6f912b8b01893c61717f2706606d5d78135c84be0e2df3cf88e71875bb45a048e9e6af6928cf65757272b6be3677dfd4b9e51a0be10abe3cd66207e350fe7793a9f4cfc5ce2203bec8cdbcdde317f9ab969ce246b9934c8e8352f6841055158a4f3a63283ab230a6d38;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdf0218d407cfbceeb9fd45ea91e0d2b0fc6132a7735d1a4a8c8bf922d03bb55ad556fa41e6eb8fb3794002c926ad2297539db01696cb6cc775243507bb44731d5099d22a7b544f8b37633ef64a94a27aa41108ed08c9666f5761ab666ea66d061d23b8e3e2f2047cc356a652e54357e7acfd36e2a51bd04b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b55f9729791190c6cf3bb9055c9184d7ea204c0e5ab885055ed0355935e226e8162a275fb20bb35fac37bf2e9ae4190d982d21081ed664108dec6683c1aad87a42ce7c465a350737599e2eb77074458f08ac2973302d4bc28c43ec960fc0dd6166b4f0c134061b1d862f5b495bf422e9a0db7356bdbe2e09;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13af8c8d9eb93139ed5a3b4ab5a99fd6845d55007625a038a5a933bd599b8a0eee918bbdf86fb66f7b244a964795e407ad39ae19ce22d05a9aaadfcef3249b2cfea0b62da0d9417fed6849041c118da1ee89e83184cab2e9d096a316dd72039a9e9b53da098e8e192bf204304504c8c8eab8e98dcc469e055;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e2253fa3fed17785daee50ef8febaa4965d17cdce9e82c1baaae4d9ae1aad05ef05cbdff885019d6eb3e472773d1c2ced7ec3e6b91a906c930271961cb48c35095c12df0c9d76e0a9d043296efe7f5630c49069129650bd0f847597914f8e8a8245ab6e0b17aa2b9ef20bfb15feae139c049d5631092a3a7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h823f9259d700b1f42e41c0252b5cc99eae78ac8bbdf97427495f99a037a1e8bfe733aa3d16593ca23ae1f08451a5374e0fc9be8edd84219e241ce0d9c84c7a4571b6b95097a90e2ad906325b5291ed0f38583d890d5e3d45cc2e1ec620df0eb8698698b2e108257808589f28e33fccea275f8ee6bebdd86d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2526a355f7c5672df3af4d9c5bfdaf929cf3e9e9cddd47d7310198896f5c527968837e39f846fdf691bb31fe553d507deabf73e62ab11a690eeacecac33cad7ccf101424341c72790adb7d31d84daa0079fd8411b98393d7f54ecf83dd0228bb1b5fd75da80e390b2bc21c584c9e2ae4b3730b25229605b4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b5542757872d2efb47c578ab600a1e5e13d0ee62314d2f6a45e2cce2b81fab4c5e836e5fd51d3c45e898afa0c080d71bbced123ea9dfc08442319b661729a42282006011f4f3833c9d80e0f80ae1020c36bc1f31dd0646dfb3a5dbff5f18886d1ac2e0a39ef7fff47694dedc3035089f2434b1ed76213d3b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1941376c0956623cdc7bb37dda7cf950944059fff8bee41477a85828a73e905b8acc4d92708ee409dc01d669b142e26bf61d55c1e2df16d4c438f954c23dff97dee8e88e2e502efd5ad2e953f3f3fe876b4db9821f7dd8d289e191013c7028401e9d50fc833c515ada997138956665d58a954cdc7aad4eaa5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4300639a584a7f76b6f43dd821282d7b3f3e7d91fa276cdac94e954371783c3a467337b1d915186bb28462ce11d4a2c27cfc52d33954e21aaad21bb99463e2ef512a7f84c8b9eb7ee35d034887d9b3c1fb5748148152ca4d59e347f4e3e3210ccc65ae60ee2b648269e650e28725038c4f5d3ae79ac202a9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h118552e5e7dbc80e91f7d750408e430598cbe3c1f9007eb7863268edfb120582db75f77c9c699929a01cb38d674ef7ee416d4f8f40c4e8fca0305c4d352cde1d91bd47b1fa96a78277052c480d8f94610eea363fd55abbaa1047abc79f6de2f331f6ac0e1b0eeff7e8e18c3d2c86c96e633a5aac77cbe6171;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aac899c8b475d5bb0fc92626b0d38ce41e35a7c2b9db0014d13cc72abc3a1c97c4c315e282c8ce3b4cf48f21ff33128e430a88eee07b315ed7578189d065da7290b83b87ebb7aa7c4364a3697450e9eca80bfc120515e9f4169ef9b692fa2645c2c9713fae5717393853264e68edc4adce5b0538b5e03466;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h152a80e7b65dad7aafbcb480f7716f7414cb7918c4c6e07f3dfbd6a0348628bf83cbf464e2a1e3f55713c149cf412dc78039cddffbaaf61f3759afb2f22e2abe323b2241e2f0ec3864b3c88cd00d7ce8486a784dd8732b61d89fd21edd110630f4e4c5a30b5f716b9a0599c88a3a435e8d4f383339efbeb56;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h186403eb65c15be8d36c8008889cbebb1449d5691bad551c1fd776f9bd276de0bf16229970f6b401c2e8dbc95847a01b1317d949b9eb37594dc909732f1dad9667646fc8239f52c68605f558a6f0fc7bec4b53addacfe6ec7b19ade40da02e27ca7ac3af6f7b75b5ee1950f6233b14b541e4c0f5c0933b9d0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'had9e9557a2c40f067b71e48d265cc8ddb693b054c48bb6cddd5e899064ae563c8fc390449549bbf7aac1ff80fa73752339a3d835c5834ab20329d5bfd8bc7198516f5dbab43d5768df3c304bf7af6c7d0877f62c11c6d17b0db18fa914b6475950d6a20e105c67f49cf173719e8b2d50a4c31c0dfeff5f89;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5d71e3aa2c8b9cd5087ad9c7f812bc2ed1e8a384dc4600b1ebebc21ca5e99630812ed1692910e9fd3bfe0d6c583888c98ae307d5e6e4cc616d283beb04faceb17d30650c38ab02063c8bc78f948c0248c04794a3f79cdec2fe48f960c7c96539494a6bc1de2a33bcd382bed8978be924e3388504bc823e66;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h58f01f19fedddd7fdd1eae7e72a5c896d88f26fe0bdde8b64dad432506cba6bb5ebe038c2581cb90e246435af9cf883e556a4c0ae12a118be3384857102610cd8a9097feb72a67b97875db17b89d64338444b2d203436bb7b1735ba06a2877c97488ebfc13523685f6e5abd4e781917378565924c03a55ad;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d612d0415306f87791510e53f827dec531586ac41d138f1596db27066009ee13da17c5691e6988e0bbbfb2355d6366a449e36ee946a540b34cb9383ef9ab0cf6cbcb0c497199d5087511e3072ec361e83cda66b52d4f41dc7248224e46831f851d62c880e48ed14d7a543fc934de197d812c01c8f59b75b8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d41e0cf7552faea8f23e9e48ccdb5402a035a1ddb8f8adf0666173c5eb6b74dd2f799d0e10d50beb75fd6841b53db96af8d7c528718e85ccd7510c59907ef0492f7ee8ed04eea6b9adef6c6d8877bfce98dea7771da0ec697c2bedcb633bacd58e64f312c869bac2b197bdfe0d37c7e7bb8121fd83894fb5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h114524db78525c6643c46e87c32db1327babfd38421d3926787aa83cfc0509961c10cff66bd1c9eb6377336733bb1a2ea83c16950c094ad3c005adbb077bf698263ee5d79da08bba227a47a06beca955623c09017e2e708cb3c64ed80cca8fdb4125b4648dad6e067b6f30fbe0577fc0b7b1c170b567fd62d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aca74e70b8fbd261a39c2d8ad223344c85615d1892b5f22140d976befbf19c39551d1ff74d9638b6a3685e5e5a49eaec3bab97192f8fb83088f7b123993963df65b8799cf38296141f611a53b24da7af0f4c14c61d4ae7c319592542356b1a4a1f20cc0d6c59de53a5ee762c9094f7a28312700125505f3f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8402ad6f4c81e2f9df53be59194841aae4853b7778f006f83ad1d64e8bc4e0af8105075ff2020932c8c473e85885485870fec498e8a952ac82cb74e7f2f9d8a449349a3387be0d8564f8e54a838d5a82792ebea1909af044e3d8b4a0d2dcbf318be9ceaa6f1519d75b098ebed22bb198054d794b0b3b8af7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb8a6576fff18f4d35c518ecd626cb00a420a788af56b2ecaa72ca33739959d9c02ec271a1b8f3aeda9f344e22eb2de93888891fdaf45b0d186de64bded37727ff30ca7ef2955fd3e0c44e540186853a8da2dfdac4a4bfd9266f4505e2dab2efd37a4d8056a0e636abb90b93759dc1a3704af80578dab9edc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5de254b121abc793fb82229f702792c55d9da891966e11b9c46fb75497947bdda80e33ef9ce226a93a0edf06527b4d206a1908d778ec51601bd880fb44f4a6d44e5dc655857682025a0413cf147197ca64a3ffbc897b2c19501dda09814b87f3efc5b1ee77581da7d4432beacf3f3a9aa6c99110a875f6ae;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b303181424edc3ab5022955ce77dd4c0d7a5cca4a73226506fa3262ce3857ad4dd74c1376242729be55b4bc1623183e4fd15ff0628f08ff94428d8d21446539a9ce29a309e142083959fb0aa2c77593011c9c27b0ea24962d5aa7c4d6ee302d2e178b04a9b73748b0ed28a9f4ddb9a9ec34084d9513272af;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10de73551dcbd76bb21761e5f7e9643281133edc110c5e19c85d0eb74caefbd3c0e862b9eb9bf4cd79c5483b71c2268a981933a51c4b2aa0210527f67f911139085cb834e3e620b96a401c6eec13adc9afe949e09e58e4fe5223879bed791199ebdbf3853dc43517de5d89be19e0949d887bd6d8c3b4472a3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he4a350023d40cfb708c7fbba6809954ce5fafda790198154eb960c9f98573e35eaa2f684fb1b44a5eef357c636688a0f19c3981f6382a74304192ea79e806e134a630bd15963dd80b9274d6e4ebb490069633ef0d6a0d13c9322a3527bfb2fedcd21377515380199b6832650075ced3a8e0b8be143b6fa6e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7440a148589f0e2c56875974a2c3918fbad3a538fc8db90818420f12e315e26d4caf913138ff3cd5eea35c7de318f6356526fa08cbd8206f8fa692549b780698c228920ef5e93edc63c9bc5331ae54f3521d6452b6812bfcca24e12ff6d602d8064faa73f3a3529c2ee1d438a875169809e8519a2c301616;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5d7324da8b6731e7101f72435a33ac9bb111a203f047a3ad7701a799bdaa45574a63e2c3241f363a925495fe9d405cae1db5a3336899a7c3f5a3e2a926736e71614f96d351844530dcbeedfdab3d93e75239655690762aeb1e3ecd4879b4beb524ac95df09b8db6b55830d3a7d82f10f20bd2d6166bcf0d8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd1fcc29f76af0c933fb662518edad2e9358c0027877e878a80f2401e4338d7b47812ee8729bcc41755d52434683f9be0bd0dd7cc654be7ff01e0f416eca8f874ecb14e47ca41557d1996089418ac3ab9df4b81493f658ae9f0673d82f0d597e51196862182c4f9049e0e14d461d1aee354a572feedfe5bff;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2d85b7ac46db6b2b9a62d448e0751b487507db307e11a33dd220465625f192a1814b17bd588adcab274a4bf531c58a1f16ce5b589d88a869fb2cbe4ed83fafad6098e03cb92b3b176f33c4e725b296be4920663b8ebc34da8f4f14b1a3f02661cbe32a78e1e30e6476d99d96deccbc8b3c873ed49b86fc9e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1512f25e7154a753d67a226536632847c3153b276c009ac111ad0ddbc7d82906b5a643839aad388c38966e2c0e2f207984cbdc2ba7ba9c6765e0a05b1504f16b18fcc159af98e113afc7f93848eb217fabf99d1dec51b1624228a9da578615eb2607a0ff36c9bc15c866eb14dd27e4783fd51542fb518ba8b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf23927bb98942ea4b463648731efcb92ded4c93b4c47881906a175f0d772979448ca19474292db379bae89f685c7e0df2c139ebe8b89f227609920d36e030ebe884194aae3e14096c192b4ce9da14a27cab185a076a6d30f9642fe01a80a6d3a683b7d51587f2a6641ce31e6e7615fe0be19d29870baa92;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he38bd9145cf1c958bcaf949ec8b16347af4b3675ee97317b4def25b89bd1581aaa79acb2f6b89e09c2e59fdd27389e098bbf5d6bdae4574f19540a2a0af93698917a7fd3191b367c6fdf8bdf30936fb2562d6fa92e8a6b9b0861889a697fa525cdfc42ce20cac7627b8adfb83dc0e1d88ecb5df7cc7bdff1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha8d80eb94732a3ed92685dc93e547d5d227f67b73098a38f49e76c9d96edada68c535f3d6b66b291170a4d50deb04d4ead7ef618a5ff23059fdfc943e2e022e93436579deadcdcf301fabf7e4845a1183c74659f1412b494b4713c741ea8f4366dd64e592f10dd730c49d9f59464f28001b31a40e1e62d30;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h71936b2374ce113a982bbc4b65290805dbb09b91bcf55a9f2bcdbf145c86190e7e335180c1d1094e19ad761b357798811623fadf80069555ffddffb074825f3388bc912eae1d5e545b1664f7f2e811693f822430f8e04cb40a138d519f13a89c6ad3c91ecf81c7e3da2e8286fd431bbd32b5e5363863a1a3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1685546209578cca74bd752f44faa5b1ae591cdaa16cd03e4d00086c8f4ab00f2cc3b3feb4e8ff7c1c56ef8940b1e6b7ea2e8a093d02cf1d756a8c929c48085ff49d2637863c4e7774aa219373da2408de7769e5472f85f9736a91db8c5735c3e6fe73ce178dec6745f747974b906449dcc18d1055df51465;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3d603002a4ab3b60d8963022f8a51b7ff3252e561edffd2a85ebefa92f9c0838c17490b39dcc4e8b42ab3354bc7f4a8ff8b757cb653062738df79a6e868701c2096f3a22b4a361f1fb2bcc413ca430d094dffe335820b623835c4569b463ecf498090f345182c59085b822fcb9bd2193ed93571d3560ad6c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1713730f164b1de926221b0020fdeb1e9ac67e4236ab8c8ef8dc27df0e53b935f8be89d2d01de08a0874b3637073ad476940b8497a6976774a38c999890270aed9b32633414f06d7303927f6bcf45292c6f22ab017e9984474e08da4dda5874db1a0c38deadb4da3b3d09a554da6521fad4c80833135af4dd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15d3ff08dc36af7691c4f3f29bbb8d425f3ffa4a08deb10fb51d9eb2f18b215ec87b38be182dff1783cd67bb289d1da09e9b1587b4a1a4bd476a4fca62440d350902f1a9f6c07bbe4ca028c48f35542b3f35df95e4578f4eb6d0eea5cc129da22dfad7632278d0b149fccdb1213c971eaa019cea566b1bd92;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h121dbd9e9ff641d392043ba62ae337b494ed2de3b91311955df0acc1978cb598aadfe35ec2753ef8bf229874654a24a4bf4e46695da5ff48e569a49a80fb60c1b55bdbef8adfd2181441cfdc4851df3e1c8b3ca3ce29b61d1a7e4443d95e9e6811b94792a8548a7a6c01db69ff94f4d0b2c559b6da13347a3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he0b3f2b79e01391f7d89db3ea775db9e1498d3bbc46caf8a524690305ccdb784ad299cf1a0c8256f1bb1b5fdc0da29275c97f44122f1d6c8788d0436182b4d81bcf2e30e95b2360d73dcbbc991a96ef2b5fdd550d7354195b6b393d0b1ff7c19c12c2ce4cd566cc87f894f85e11ef66b5ea5605d65aeb94b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h310e5365891a77142b75562408bd1990ac65efb9166d1d1305fd1aa53a990c8bfc08dc3f5580f0732405d6548c0c3b767921d7dd05446f6e160b50ea023b012fab129735f5049da938893de9abc35367feb2f030c5ebafb19089a8d6099c270467f0eaabda116b611bc7658ff6b41b81a34c78639c68498b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1833975a314f7e2229a2833951501677a463b1e5ec5504ddbc7ecf98f558605c58cf9d40854e7e80a0d60a3b0a2ecc219714d8c46b2821bf40d43ba12155ab1bd95ca5ec1366e665e197cfa0ed049efca55069f4600d05654ab482cc6aca9e4b3d306cdc3eaa3eb13f6b41a123c3cd958c79d6c301024a294;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h545307672578841d3e858d813c4daf98ad5a780f04ae83aae33dca36ef7c9b111ab09145e50d192c4dc01c2d47e597f13eb6c6f6be5caa623f0d453178298ab9a2a9bbc3faf255e380fbb50d957ff8c0d180cf791828f2e2ccb3990297b811b5ae7614a1dded31d4285e50de20dc95e32baf6a624a65ee24;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf8368820f09ce225b4237e83ff71bf405b915f4f62a94c7ebfeffbda06e39c6bdc098a1ffcddab6dade29e2c385f94f9d719cd60c9f10e9c406d982956865f61f3ba6d8baecd8547acf395ddde5ba73e94b52411753a114671a037f6e278ba0653b21f2c5a59546ad4ddabd2e6b40c9e477d8cea18093529;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7e39003f77816555413d072eb096870b1ab3565d186ab9d3174213e554f5ced9823e22133c0730107aa6bfb904d2ac4905d637d1e39dc5c6fd9e6892d71f294fdff5b7d5202d449806224b9c4218f9e483f0c4ec270c67b8d5fe19ac6e1163895ab6ef6feb4df6b2c405481592abab7808308cf890746abd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcc37f5419bb3e1ea0c1fa3dceafa8bd50ddb27c2c55a0d02d7addf32018e4561f4e103e692a692b1d5809f736c51c59d29d6574dc6251f777579ec97ecd2549f09397d7ee3bdda0871ef2e2bda3d972a74856c8e9cb1c13d1dea3344d40bc29f94f8221872bf68716dab6b6a1f9a8e6e056a567555bec19d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2513b1d469f2ee70a7760f23330587b841a043c61073fa8c677588df2f0a552089d273f0af904921ab826240d441d8b8dc4d7ea81d4e6405e6380b86878a651fb941a2141d9017fe1be112fbcd3c195b7b855be746ee4c58c708ed385ffd741213991f372a9e4a8fb00c244e67370ca5474e4d8875e9bac3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha70e31f157609fa2e158f43e54591453b257b4bc870e36c28bb964296922fa3d55b9080b37d67508ee7b1ac2e205ac34eed26d1c061f3cc879a08a1cf18643e8bf5d435995d387e780b27fa3c932ee475c283f0c0fd653cd215978b080432ef83c9114bee31aba48f1e4eca56554e1ba53694cfd295f2745;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15796617df52f4c8141214a64a57ba4d14723c78a25b31dabbbc34563cfdfa79a3ddbd1a8cfc44d7681d84ecff3051e93b650f76186c110e33def00edf0b424680545554d892c7690a5eaaa854e40aa80a39d547654fb4e58320dde853c1df32330b965c8572b868b9727fc69239d2b3b8d5280f67ab43541;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h39a554ea87e0dcc9292e6383d5c831d4f364ac386a8acdc4d31e9e3ad9f8aa116ba1420f5403eac7529220278a1aae6e3b1966eb9e16cf1f9f4ebbfcc0d422871827f130b2623590685f6c71d6a7f3003174d21ff085e6f1addb05dbbded68a650beed56e552cd091275a06e959ceea424503418c8c8b02a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h584f9588a71920d4947ca8c90a2b836e5dd10580b5f2e33cde2c3e78dce6d52cf586e8d04a11447b2bd5ae760c943998167dfa60bd8789442f129b8307e106435adcea164ff6760e180caba4369f9392d9bafdc6c89768832826cdfdb9d32eaf130b7c29d3e340527ce3a7d1faee6e49e842c011dce47b14;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he5dd0d7d673f472a9a410935d100252b9f6aceb1ce38859091668bd7fbfe06864eab7d5fa82282c0a95acdc6fb439c5c10ecbc4dd8dbef2fee9c9d00ca3e792419f22fab3c82f501795e99d53e0cd9eba4229d66175d61f8baed63d504cec7259fbd21f794b35117a40d2075fb3ef9cb9b1d547cc276541c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18a7d0154043f75150849d63589c490321f655ebcc65ca840be0b2ed834a5164d68ab17b817734951ead6fae482591502439e2a2c58d9387c8cafb703a50783203d2d8f841e467da986914cffcff7e5dceac094003e4e8bf7e8bc5794bd8fb66f56bed2ad633fcb14524f2c01309dfa6a1807cf15f035399d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19099bf7db95916501b762c39f4ada895d1521c5dfc58b6be67fd81bef129e63f3a7dc17995109f5971f47fa07ed50f1d52a19a2bd7b02145e3118811ece3a67461fed0ecb55db066c5e9733c16d3ab6091f7c4c63ba70e6628ba4c5e1ad3f761926aae283114597b84510f430cdb6b5258501f229ba5ef9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e449ed24fb82af454dcdfa8788cff757b37fea5eb2f9f23dd9075065153af93e90498cfa35553c01a117254223a004796315bf741140602c8d899e38be45ddf286e0f9fc42d89812b4eb4141fbb6ed5609f7114817de8a0d600a1a29b4fe8c2afaa80c2744de79b9d57d2106ce7b86d49065e6277dd63dc3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1abdfed1233131112a1ce9b2fcc84de5ddd8bf3c40aae36a6d80d40d819348da59d644fdf0d71b7a8524f0a02e666205bf27e0ee443dbf031ef32d567c5571d0ff012ace0690d2c50f1fe4cc5efd99da102f17dc689070fa6d4a6e6c03eba25bc02efdcffc8e3e4d29bece2e6c7160b36629dca758fdbce64;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18da727e821475e3960c23f94a713dc500a8644f24d70f9106a747b91215c61d3d8ab90a6fd8f2673c081790f72191c0ccc3e55f39673c142c249f07b88868402e93d9c837b31cca8352fe1e3b862757fa5f736fdd02643c23dcc55aa40206ae5b1a8c2a6d3e9e1ecd25e158c134355a5079bc501939e81cf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d7a75853e52a3df8b5f15462d08b4e072fc3b4febb9a7d974a953f441ee259fae0eda1bd3360e32c49fd5b816001bfd33721cb0241057359ee61d5985e32338d51832685b6112607e784f6d8e5a1765b6d7e0ec91a02f6a19c2a926a5fcb009909efc5a3962864c33d59a0a6068048f2fff39397b0193fe7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a639b0181f07e5a27e4eb64b65c408bfd66c2846fbe21d040983ac07f3d731fa4f38e6ddefeeed96b5c5bc628d98398322e7e632869271f1c805d0e80f4c1c4f41eaccef66794c2c633b3e2fc3a435f8d66be472197e1f1a4630ec8022dc659317abe1291b0ef913b8989c537b0fb757f8e41799279ff8b2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h349e6cb02669a54f2fd10de87db2e565fdab6b7e1f80a626d1128775114e9311a727c7b9e0806daa5ebad1bf5ba34bfb3fcbcd3c65a1034daef8e4277ab897ddf0bf8e6b39db3be3ba17c314501dfff7ef1f11f9047f1edf8a5c487c38e4f1147633805678f57b3ec25260f8eaaa1f5144c451dcb98c5bc9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13076c4cb9067e3d5cf24ddb264f822a85dd054619e77833768fc81f970587247a91098e54e2a4595922f582e90a7cf3a43b472c5f77d7c542053fb5e58562bc70a5d230ca86fb9de14f5b8775dd6ed78aa213c41145e016ad64b2c94922318dc39181bba26ad107ec2af4aa26f4ddd7322116e3539694d2b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d92723f7804f40de5fb76ef877a5c1f34b8a6b6a3bfe6b172480c4899f2c7afca981e79e2d3bf61cd4ed41fb72aa6396446007f3569535386798c30b1ffe8d10a19f4794b83eff76d7c759069d39b85c4477387983c9f2399b19ca6b05555fb39e7439aecef012f273a368369061d15730d59cc250a289fe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e478af6219dfb4d2d31bd8cb72760532fbf2bd885ac17cda04c9f629001c46fb711c40f9dbffc03d65bcfa0e7782270c73307b9e73faa60171427490ca00ad52a11182f10c31d7fa47ff1cbada1a1872305b35a8624d4964662c7f15ec71a87f8a03d148e9fc69911f0b402cb87bebb6ac6cd3e955fed4d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17f72d77c1a3d021e9afd3494cb84eeb40bfd0e7af52fa1e2c383a814a776643a27aad3090e207d3b1db6015fdb22723e16fc2a4cf9966c3757db50259c68902b3acfcbd10b85e0e81790578abb0f1c2aff2f89e448ea733aeeeb2e33b515a33155e254bb7cdaff02c572b2a8e69ef5c0c9ec1fe665b43d6a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c5b524290989e9ca0ed578b6c1bca5c92c9df9961df5d8e6515792c8d2a8f307bfe46d79976c073a100f956f14a9c3434272e4ea52fcf94c39a52a8913a3df5024fcb066a9a442d89a08ce481cdeeb1252fcbfb2df3931d4f3c197327eb072f644ece6c6b1b98f81f7417697c271d6db73166d867221ecc7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf820645c472acbc58ef2ce45ed4ce710932e3f5a3011c1916d6748d8175fc9f8ac96a0726ea8d171d2d8060dc3d70fd215a415cfb69db567c82b67042975f9324be11ae182bafad223f2fcd445044ea4f765c87999b06566193cd2a3d3255c804e5a018aa7eb3f2f485f9936efbf5c1a6d916159f1d33058;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h85a43352061248f10846fb7ba58fb3ec862c4c17e95f8985f4af4a3b086634236ba6a15fd5b735e7f355efc6d9f4bbd2455b3c0a491e3183049ca70f68d464cf2ca45aeaa30f39566e73655f5fe876b08159ef56cc207d3e06184e861db62d342f5278e02b7b94621287d94e87eb8b09164bb6b0065195bf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h78c87a2c57b36a481e8cc17aed3a02ea539eb84b6ea632b0f22f742680b6666e261c796bfc159cd8fc230313c922a2da138df0759a207989a79975f9403816fb1e2ee238f56b97aaa871fcaaa836a75da2b23d9222463b1f5dab6ba6947686f81effe191e3f18ee8333853e3f867a0b3f005f3e6c1068cdf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15f85a6d48078ee3350ed4df48c4f1d92110b58fd45c54878e0fe43d55f193f824cf4df078aa4c825227bbf1019d2c8b97062273a1912d6aa189b993b6cb03e33d890c89463be31fabb6109c22f971e167419e580c4a013c35c91f59498528636a295b7de8a1c3eb0b67d2f52194683d0f684b8b38c288dc8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19da516dc1b95ef1397d6397b3d5861da9351f5848ca997aed10083d8324accd111ac5eb4cd3c8e636cf57283330ae7d2ab5cc9e57b11589e4356b069ce077e55d6ec61a2a58defa37f38de994ea86b6bc1aea8e918caf17f58e35fab99c3837e8eee21cada8d3cb4260bac5976454aa638d5ccd496aec7a1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h179c8219aaad5c27ba97d534ee1802bc6a57e68509988a014543d2a1785a3a3b63dfa578d8ca1eb48ad3dd8f83a8e2d74c13e02fd81561b979d19d635041563b36cbc4b444a4e1f2fbc4e83fc8fa56f0c1da1aec6141144550ac7d294425512a7542d03a0b519e5cd521ec0d699e831fb9c482077809ddb19;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dac89cfc88f27bd097f77ccdcb6ab3b13ce552a0a11adf591ff7360f8bfee78ed921f9aa8fcbfef7cb8f0153cdd242c11b0d3d2c91f4bd1e0e526685781a9dbc12645b57da26192099883d8285253b9dd70de5a130a4da1af03cc9efdc1df10cd7175ff8d9245981070a0497f459096f8345c48d09bf0501;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdf9edb03da077f4ea7e80185e34c194771dbfc58ce20b66f6e6903fa6ca93da6208ae58a068f5f69950ee06ced263ac2ee99eeced25afbccc1e8ab0cdc851ba1f95abdafd2b796b2c6fe1164e46a88157b622cb0d4f3e60ad5f786eaad25bec681be4038649e4a80285939d278f3b7b3b6d3b8e18700c188;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2e6ce4b8743ce347bcdb8ed3c162a1d7b46b773290c4c069b54076d3d8e34fc4d2685bd7900bf7e3fb5155d4bdfc56a057378d99f93c7d36734024fe76d7fbbafda608133ee925201cd341b4f65df9ed88e16b73dcce52fd0fb87808a24b7cb6f287b40b3e1942a19a24bef4a90e9adccdbd823250ce5e01;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h38fbd856705aa6ec50457cf0931a9520119b8535d03b0d7f9cee2d60d0f1a0044d5cedf3c2b3f3c379d16e4f767e8ca0078b0a8b137d2febdaf7e621d5bb0bcbdfd8f02b0217658184de2ae0eef27ec14fb479ba9667e7470cace5f7593774dc46c37f6c2f225276fe345ef169052606857a71625f938dab;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12ca6e93ff6ac4a7a2ed49e4440856ab2f38d86c1b6b350139371d421ff1a39d2dc9fd56a2f9c87bc02f2645ecd0e2f09a830e3e890b2f427ed939c62fc53925e962d23ab70ffd9d80155a3b12eae6f9e727970da91886c3ce600a6bbfc6449c3ecf063ad0ce31958a6d2f1471acb836141830369360ad7a9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10aeee52d4bf453612459b4ac09df46d79712dfb8f19712b68003fe7d688b557b3ff8f075d87982ab0083007da772cd8535c12463b7f74ccf60fe6a211da635c242d68363e7ebf9e1198fcd10e144a72e835d19d9e0eb7e5f428e3eb4dd16d843963a96d580b830adef961efae2fb70c6dd23654a2da3eae;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2ec0a285615d95db3bcd4e1d7e391fc6a3808ba658f0a2d6487da79455480694f00b09516406808a56b311a6505ffa141792e50dae24d1a2ac3009ef731c6deee17453a3e505f172b20eb93577fd264fce0411f168653f5b1c6342bf1606c3dc5827d339b340970e7df40b7080c60e27bba6ca4c77c30d6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h958e9e421f6d65b5e3e1280f0797ff67967b298e39c4c980eb00b856b1f24683f34e523f4fa0ce660c9a9923f4c9bff5149a3181ae4cdbb2c4df13977b22177a53ae943384edf1a883b5b078db789f6b41cd71c51a723e7fe3b2df144f6f6267273f18f30f72faf73fa5bca37a721e2bd6e23e88ab1ce904;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h33eb966e60005143a6aecc964df5cc7bc389c2addfc90ee22881e84a8fd0d4d11bfe2c896cc0cbc7a507a2de50150bcb6d8e35f86b1827b3753a9acb25319015624b488e5380b7f1d684d43541f9cdeda1c4d4cd746eb7cc44fd08dfb2aa6e41b4cc1e56b90982105049f8669ce4a8f1534d8fe9d41a8c99;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8c472d055420288d37b02dd57350b119a5f68d6fdebfdc5d74d3b9b80c69ba146b2c8af99962bcdf5ab21cbe527262ad901a5aee3bffe06487c5cc2d2b114a074c81ed8a7311ab019d49156338b9d49326bca2aacda5b90aee933f18c82f82ed4a703b4f5f636f0a2169890f3450c44adb197be68c428c84;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ebd15466833a6e7a8535712d11f42384276a058361f06bc92f4fb404d9891b8397682d55c4e8fd1e6f7cee5953447c5546f6a5a227c63c298e501001427e584c71962bfd6c7e2a07cc3d48c1b24489968422dd3124720787a56b9a013e3a99ad51fc692c1330c50b9755dc49aaa1702029ef6bb4f31557fd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13e85a5ed0c66c846cd939d11e6db995bc4188912d10e91e94b1905bb8df5aa97c49e1aa3e927456881ae83377645227ea8c7107d48e973f62c758c5450d981f2c1179cc0725adc22a331dc82f3877f2a0aaac51978d8a7d8d74cdad01c34ba6c405f63da761609b8f0c1489f89e64e25a3a4c2335de7c8ce;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h113ace5318effe6b34882b9a723abbb5ad40a682dfa7436ab7cb222de18052b649f989da87a9e7592ac4a08f908a5b079caffdb715150b8998184b03ba31b4b17fb19a9fa4bdd14b041515e5ac27389fa42d4fdc124a880c37cc8407efe3b6cda8b7b00b7f034b06a8439403d5456aff916213ecee25d61d5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19d3df1d9fdc62c40759e3c18e0dfcdcbff8fdfa52c1680150fba308e76a30302214abc19fff3ce838f79d740e54b90872134510e358278f459664412ef1afe1fbb0d632b1f48bff315b79ee5e046aee42428466f405cae27d6841b063120b4ca414ea2ad44b6a29ef3482f433a8ac7498e43a375b2045d13;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1423388147ebae10642bcd637338c90112941ecd56f5a980fcad59c4e273a618a74b73f7663f367ae8bef29c78238bc5f59e3c0abfc16598e5d392ec1cab81ec10d8df35762b1e639bec95cbe79ea1f0e9116580dfb13c88e06b3fd07ec24a4f1fd50f26e6b9493112479a7e40c983e2d2bacd16750427eed;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h216c442d1119dcf781db04f90c1e8d63484e61cad3b7c86c7455a3af0f99a629e5adf8e2913cc2e514a5722d4d514ea3486bcc2a9813432ed3e13c12c5560eb5207589bd31f600ebdf8322cfe0f3c95e288c32573f07d9c2290218a4c6c5f25590b61c7781fc0c7bdf391e08bfb8bf4091f3b69d591a6135;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h102702bc33bf825237e55ac27a8c8ee2415607fac398910847a965c0a1cbed34c1b0598a330ea895cb82e313eaf8b2c82dee37146fef4261aeefbb08050616aa1b1fb2675a5013df08298a4f2d8c69d166e2acbebb4502c188cd542eb105ca197d8b886ef0b5baed991b4f2b7d558488e51b42e4ad873c401;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f306585a8db9349a24eec4e1d07a59d4159feb2860507dfa8c4967e0e2fdd5b3b2b05684679416739e4cac07374995c6cf93da5fe51aac839347173aa6ad49159eda9c2fb34a5cdb81064bc42c7280b00d963fe64aa88db8c3f0662e25165f2e02dd6043e3ac744a828243b8308c253ad2de1fcd9432ecb9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15f6b28c53bce5c16f024f5df291f16259791e4067b1ca88e660ee8fad3a7e2cf9335ba6b04d6de005d2225c50e1a04705273df60fa2bd962c11f7d697654822c8ec6ce33465af9de7369e1b3cf82ea4aa4824e9bcd2b063b77f2d7b912d95da61753b3cfd053ab138e632012bba3a0db031b16b5b2432ec;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbe030f3a638ce9ce59d3d0c0d9c65c79c5adaabc1784b18a6db8be06e078efb6ce53bdfd4a2d55931214276373a3001e7f442c93517cb06b1a57823aed371f342336239c00e59b8df54e91eb1aca87a5faec92ecbe4a33cec34141f5cf9aa4bbacdb56b68baad90b7cf0fcb17a6139397628125e731cb5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5644190b71b0037d547a4ab40bee9736e76e9d533a4a666406f7bd0ab2b906fb5d74730973451ad155379a88f5699db7db4b7ad8062e49a636d14a2c7d2423e506ad9a0635fd04b6430c36becc2923e00e1cc10fd3ed530314a38fd96ee1420e8bb56f124e941b3a9537bb9154246631c6d03153019490d6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e50c2889919651f6ca13ebfa4e736e2bc1689dc0030846c08e0d8b0282c8ceab43fbfcb70587dc432e32723e033bd63b4f14fff2d770510079db28431a8d0780d5701ec191c8e09645935b7908d6a8eec59b06214f05c8f06feb88dd429093db5f841719ca7fe213329e9c49b36960184fbb16a9c454d9b8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd09e54f16b34bec8b7715f276f2441ab1413b58741812b7fa2f919a91b015c050f56ba09bde498a6bc838425c66a85d0cbc0fe53ecdd20e673e70b470dc228fa97e230dbf9cc68839eaeed240124b6e7ace80807d2dcf26106fe6cc6edead044bbc421d99887b2a0a5314aee2642a2b2e41fec2d1ee2a5cc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2f2e6cb6dc1ba77902771a87d23e06f2d9993a1da4aeb13fa51607c973279d5e4dc586d0205a1be1f2c1c695e4bc9b995a3c8726f0cfc1934492cca51ac60df635c2d3b3d641f826578670ff9f31f24705899c974b5d23e672fa58ad8a964219384fdeff39e39c28dd27b9dab4a7b746b03bdae5a62075df;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1457f0247e916528e4e31cbb5ef19ba0f86680e599e5c599f2538475b0f822f9047480d64eaf96a8db068a24de697dfa96c0263507bdbf2026b43e4fa45d7946743f63eea50c88bacd4726b0da84e8f9f82e69211919e88d9e00f3daf93b6b38044184af363478acd554021e9433334b4661b93200afff0bc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he9d2699c7c824cfe054c609a229dccb606fa7ef6a7dc58afb2b74486c7c2507b5f3337a96b6390668318615e9d78d2f060ba2c677c923cb66bd5b676a62d2f73e9b9f294466f4cb3c17569320bd4d96b6bf44189edcd22ece055f7c7740a73b7301ab27391d0ef93e914f9d91f59fc095570266291240d96;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10817b09d50dc77cf5d8ab1b4384d662ea30a1718d5941eab3d313ae7cb12d31003da1cab3a861279a58465966a62fdcf676fe79a10db30b2cc626fbb1bd1dafeb6961310e7a5e1c2d95f2067297fc15278824019a204b8851a22194af13ac84aec30d65b6ca871187e07854ead3493fb5409fe15236a1b04;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbd1bf6ba304c9f126b7e1699ccf9e3524d76f4880fda58d847c5effb4fb48d837e2b5a64cf9eafa9da1b263efeb4f135e3f17a72761103a0b91c0e2c5465ac5719d6ed2483c470be0e663d162ff68a5578df4870291e41c39f6dcda5e9248fdd1dd3cba7223aced91d65e03fab131cedbc9a0bc28488e7d1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h182f251e28cb0397f47eaab1abf24f4fdf01762a30a00a9430f8353bfe70a0ef64e5985b3beb2193f36586a7656404d1dce74c537bdbce7031cd4215bcd649717b731d627de71798082cfc8d05087ad4d54690c04e39485d775c9ae75af9ebc7fd93ed8b36efdaf45e75790fa4fb5d9596a8ea82afa89d02a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haa47f150e1ebec84fbeb916d54381620a53897fd8e4ab3114a916b971d8b11c9cc54cd6deb5a95b926d4bd3a70c28d21774190a29969dcb5858637a4ece5bf16e7741e0ffed1b6f1fd6c22642d135578417827a7d2344700cdf497234305f91cd042d2d62e903aabbc88cb451f5d6afbe891340d9daba90;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1358fd6f79291427c6c8e55d0c38e0a2ce027169bbe37ecbb6b5b0d13a05b7ce0a652d85b0a948f7ec323f907354257bd60e6edc6f4f5071c7f1b02d39671bc8c4907fcc358d1403649081677bd6495d50309979fee70818401a3780702b9737b65a0ddc87799d5ddfbc0a1b3d0af440034bd5a299b4d2505;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h149facc294393ac38d3a4aad53fadc254e15fb856c35d7bfacfe38ee0ab4339740f4c2123c081170dee4b608341529c1cf8cce31b67eefdb0280712767f3e22afde9eb57dd4829704a748c2caa9c0e0f205adb2483425ddb60aac4abff01a259ba94ece68ba928d4e467a99482215d6c14d6145edc247ec06;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14608ff319f05a7a85f19188b8329fd06f1d44c57aa067646e3d343de15dcb87c19107959d600b7bba6eae861fe3bff97a23404e1a8d474b4cdecf2ca14b47cc92228a4d31ea5d3142edb985fa8bfb60cd7ebf5ab13ad7390e1c3e370c6c9009f0f7c958356219e00cf8afc4152a79e72f0662195cce699bc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbc9bc166c807ba4fe34c671571acdf2d134b66abc596cae877144c6e8ce5b8c50644b02e6e311679285d1244a2d24bed4a76bb5d287d9f49d66ec0e45d7bbbadd4fc81f241f4a7b5ecd15efa4a13a07b14b80ee75f6f83dbc95a9e8eeee97951ab4d0d0de4d8b5b1df746d98d2dd0826b818db3575943121;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5a4ea7ab8e0f9e8ee658ef727639773bdad03e250588eb241ce6073db381a5a54cd970e2a6502936833a107551392c8ea50af14e4e9330103b59eabb528b9bc17a2638c72c5e3c07a5381969e32556197e3c67dedfb2bb2528beb6753701d30abad25b57dab6c7d9af6ce37a52811f9620fe8bff9b070905;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d3374130820125c997461c566691e3a466b604fbb4281948eda6b96961f0aaa7c0079edf923a3913680523cb700eae1bb43ab782cdc4fa65cbba01a17e74e00dac5e9a86ef97557555bb729d34c1946d5dd1ac72a2cf59b6a741c7775bea85a896f27ee10f16c6cd3ee2422b1ec110a303061a8bf820146d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3b8f32cfc963a2e2af40e60700e56aeac2404611f5109f89404f2e30c3d2f629948503a36a8a289a102c5c99b92e47f7540b34fdfe3ba9c4e0ee0602ec08a902ee1f49162773afaeca3c837e7d5ddbac2b4ee01be6a7fe04b9cc1634cbfd0bd6a8e5b57034219bc94a2b3c6e61510ec12c0a8f99946fedff;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c94636c28dbaae80f2c85acecda12cb1cec375484312cfdd97146d90f1fca5a4d05848553940b85bd2a9fc4e2ed6265dc9b4e4bc3809391f435d78f7696bb939cc627afac138f99a3e0ce2c3423297c84560e40043e396cdc9381cda8f54278427a145d10f089c0ee3abc18e08189eeae8ac60b887d54b19;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h22b6e8895eeb166b1ed431226a57dc6a437ab46a241b0af828cd7cc6dc4a39ec53a9472f08f06917c12eeb54fed5a57a5d5f717837a3497b865d0402d3100bdf55dcf1eb0ae77e0dac106842e832959e16b1f3fa14012b2127ad7c3b5e5d2b5b3e3120a5f1dfdee565530779ca39258ef42cf0143eef058b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd4c28c02c24c515fbbe221bbd247fd1c441cd6ac676156166334989b9f36ea04aa8de98fd5b10fe86f97ce87d320a4ea82cc0739d4aa543d728e688d5f39f4619967b1ca20590eb76048380c7c6c7e69115e0490913f233bb399d10feddae103837814f165268102d58f93145952a4759b02c7d70fce0c4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1123222481e398e72ea3902ee2164049f11feda946c92a45c5fd14afa8d4799a2b63fca5ae201daefde599fbbb87b58489a468d2f06f99833c805f55acfbb94a3f11e822bf6604f15b4454c153fb9334924e7a74c9b8afb33086632eef16174195a361f2a1758636bf0ff32c504c37b0dc7cae98766897ec9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h43a8625fb0816b5b3f58615e2d0270d1030047ae5569874e7d65e189f0efbea4a5f3dfbf95b08c983348e952fa55642a8420099f4a0de76260dc6776acdf0e2ddcd9eb2f620e9e4162cb0a4f159e2948ba48da7348efebe9b93e509ea378dadf12a104265b4e6d285d960742f45461a9ecdd116a8fa07404;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ac9bcb4d3774e835c1d122d62ba57ab07ddbe472a3b98e664c8acdc5524fb2c3c2b69992fb1c6e36676609b274e7b5bcb6b96e6bd6d4785d0cd5cb096a0c944866f76fe87d18dcbeff9ac3bf2a1a85115e03e5dc153a8d06a2fbf304d85c446f9c9dc8015068388bfae5a217108a91c90a937011d9dffaab;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h136bc07d27a567c1a4a4323ea101765f126cb39ff5f138173297220658f5837c9e2445950808ac1fdf5cb612ca535fe2b56ddca4ddf7147219a1e74b75328df2daefcc6b42d7f5e2a2c4cc3f7901effe6653d6ad4999261a13a9b05b34645598702edfd8c05f86a15894e0d88616eef4cab0fcca3f56119de;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h25b0f2579309a1517d39a307df401d83dd33f2f78aaf410c563a2f7539a9c28630603d8be608cb34e51e20261692ccfc302cfd146e1b6717113471abed8dddd22c7488868810479ed70308f9f2d2471db6a60d5434415b398f7661a543765093363c4653433c9abff9ea6567386444384d9c320c4714e306;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15741367649fd152a4194c53b5f0e454fc192603b1c8963d5cf6894c39212e20f3bd3c4fe0cfa16a20192cf04153efe5b651fb787c46f4d194b61124e8a64694b634ad0cf77c231f76ebbb68412aca6a72beb94dd7e61b2632b42f25020a50dbab723aa028d6f102f51c2daaab3d7c7d4fe31a819a38c17d3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h194e5b073d6de7be30418d09d8d42e95d1431ab374c726043efe5fac4d76c5235e57a34377f5adf24d13ad2d8725f561c8f99b72bec9952dbc0908e609412af08da45bb678057fee60756195a85c19e86daa6d1a990e03287f119b0d211e285fade00f863d86ce1ba650d2ff3015aca6659294aee98eac5de;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h118658b248b39869a0fe1d1402b082c713b34eb28aeabe516d6ed921b04eacd93eea9c4a6cf570ae172f61248c8c8a7785fd3fada4511e892923fb34130618922e638ba2e09ea89d753f242cef1a248f54ef434f935628d7985c17d1932ba4d2f0e001502aa74e610f14df3db44b6a01fd980a6dbd5809005;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5e9cf0a23f2b03295c907bdd2834f6058295d12d4d7a9c4cd7db704a54b3fd7e59baaa6759fa328298261eb52cb4f86e5b49b8929cab740bc5014f363189c19beb41f2a0a3420c2fee40a4d465a6e4133505759810ba00c1322a5cd02594c6339e54c646924ae266835eca688e87b80da6e5c5563c5cc14c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e163c1728296c2f4b6e28eba8cd03593bb1f4ce0cdceaace7c5b40bd7248c40bb102293675537291f64f349246829ded3d0771ce9c54b248eb51a967a051f6a0ccb890d345f804b5584a0e3ee981f4fbc157e1f5688a993bc5e5d6f81b0f1ea85aa896de6df17f6da5a91953b56dd7eaa16fcb5df541a611;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdd7c417a292316ecb33f27c62f18d6d6cb7c3dcb44bc37b31531e124d2c5b322539c5c272991ddf16f06c57d3ecfa3bf3404681772caa439b0eeb7fe3fd152cf40a8cbaf130d5ada93a3618bb418e4535b14f9224a73936be65f3aef21341c7701b7db6d1ccb01049d507190eb02ab79395ad21e4621a7b5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11e32db3921d0eeca7e31d2755944e62e3f92d018c5c92d0533d0e039aeccef7cb585c0d29bb986d8fc05e7994b14732ee3d47886937ab726ef2ca1fc0a1f5ae1ccc5c582891d01a5f176148bba3beb1d00bb98a19c677d5f63a9ed491953a5bdd7d185c3cdc288e767f0abd74a02c240f9a832c6e1b29603;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f2c71767de3c470df43279f649ba5c7525a059515f3e6c4e0bca357aeb18a94893344bcb88aa5558951bf4436a972b4edf164902bc4ae5ab03735ab12f38770160967af73b6e9538243161fe3d11d46de4c418047a2f164cf173c12d6d1af3eeba08910748f71adc5d44700f03158baf036df9351809a9c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1072b0502706c457651444f8f19a62dd4782e0afc6d39c45424f526b32978b977284ec5a4e2e95694269b2a9ef409cdb6d38f0f6b0fb76892b4bf335d6dc9752cef38b0ec1ebea8758c7489a87a4104baeca5ed5a3a6d788a2d8f9ed6a1ee76002026151761b6d24d20fee3ce135c24292892c257724f299f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6f21112e215a790cc363a67e6802d8b3d00fccf9fcd20322bddeeb3044cfa75572983a0cde657a2e0b9ac6e7a264e949150f3acb1af2eb97423bd8fc61123489b70018f5c20f3e5a4b15517ff11ea640ff0f42fa184a0f0337bf109a1f07b51fbe58c91b88a8804e97608e81c9f204651af6cf79cccab04d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d2087528da369ade392746b838d96566145112b652e0e512f7cc7012b6e78469d667961460fe020875f7f2ed3b47ed74557fb8e1ff4f8ffd7b457691efdee2c79faf604eb2d59b017d2a5953de405775225e5caebf20080cfa5ac2d0a492faf3b721224cc42ef67b591298b9b17644ddbb8de4517d4adddf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bcbb133afe7cc033390ee2e90455597c7d099c84c3ba7216057481e8923680c7c65f915b67a68395d19557d8175006e0980dd1f5ab0a7b88c9477a4639345a471aa5dd6e30d8494d07ef55bfb2176055dddc8d7b82e5456444fe9533af822d7d0bc79f7c32c4dca98d9809c4b66f915ea6941e0d9caffc14;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2d7337fd0a82d9a6c25dc14109d9d2d9a65059f21839039f761c473f6b62af38ebef5f227f5bbaeb6f6244c0f53424723a44c070d87594ff4458009e340435f19192f09b7bb8a9fbe09b9805023a76bf4b1d5d58f0c3b405f9ca827cae78695ced2493b12dd65eebe39525e67d02d965a034c659aacb7e68;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he62e52d3976c55b1afdd5d4f6402d7c357ae442df67935a2d5ad8a396e17d3abfbcd6ac165805d3ef922d2b6ced0e2884f46fb4bd0f58f3102d96aa0cb1047f2bb0e1f608bf6df98181767d1bb3c30d1a56ade34d56f5985ad179214eaa38b9f3f1d79187f6e3de2627a295b752c51346a376b604a707fce;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc9fa9889acd4591f806e7efcb0c9e98c7cbc94d4ce3c4eec0c14c6dd35518dc00b8024c693130881ca692f9dd4488b7d7ab50c923f62e89ec6fff9f4d5c61b07779b2bca7a463fc92595b11fdb20fc234fb0d28ada912dd78433069b5e05da08f5996d968506fc983783f1a4877bfbee1ae201743104bfb8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5fa49f0e4bf557510d5c0e3fd3d1b6decf27f34add3ec122ef200f7988633a950d221bd6e24d972a1980df7e33b558b2669e73cf7c25e76817865440750c203cea82e4ef116b43b01e83d014c317deb08230c0d3420c14b248078542465a21c8d6602379bf358733f17e19b3bf59fc691962f18261c41f8e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11a9a393fee047cf33d7bb9884bbd45f3e569c684b5dd36b995fc0f48a6cf06c42d9856024d64fc32bd172992ce643769f451a04b03c9a035ca40215387adcb343a4e725a0ac8aadb282e57d238cd292b82c5bc1a4ecdec8c710596e7153838a13e8cfcc4106f1fa4e08cfff6c64279cff3213d3d479fe41f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h127071afe5b69856c8bb22971495d436ff66805cc6cf47a6bcfd3acddfffa80c51cdbb1e4da635f8d90cd8fd8e59b491a2a2ea4ced17b7ca26195e5f676e830bb85590179406aa71f59542fcabd444af61852b24b76d30a31d58ee2ec12d5225644bf3746151c86f117cf746d453a3174ab4eb763a1a92e42;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9d97e55dd464b4fde3f7d59eba533e150448ccecd55b1a068e6ad9e9608b2c798a49a435ff5b1c9fa84f3c0df98b439be61c29e287e207612063c996b8a3d5358c63fdb83524509bf8f723892366a25021c7fbc0d7b3ab6f9c4a4f7345551638f5147eaf3f497142445377df06314b494fa0c9947ee7ecd9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h115310b32c9bde4418dc0ac93dc8d149078834af76f6c6f9c00210e5fcfc898227a0989be2f6cc28fae85651bb679d3be20d39f45b69fad315c1885e071598e416e1f199ae719fc3f4a25914ad6f78126900376aa9a79af8f3762623d9fb28c7298c5ce8f45613a91325e60e75cedc85490e471d91c05f8cd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h49ca793c63addce657ff932b96c7d6958551256d1d0e0300e503ae92273a36ae861068b50ff8db22dbc961458ab9f0616fb043255a3a89f27cb2aa2e6f16186edcf89c2840438a93b40d997774df1b35839c7834ad5604d80b981e713e3d3455a9c750caa405902e99d07dc022e1673c00886567c291b780;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf56566dbbb4e4b77151dea39bb07498f3fb849535eb1ad7ff458d8003bcfc3f44269d2f42ff445fcf4ad34ecff7cbe9c4d857589023429d0593d5eb1e8a2f08f6491bc59d853d922bb93d8fd42b6ebb2130731a0b039f555f7af452137ea345b31339a593ee939bd667eb71ea6133f82ce2ca00f607efc1f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ec8ca76e8ea41b404743d2cd3e5798f2d8eea2b105667d8ed69ce6be8651bb88512ee230943822cf4e5d82513ca360fcc574e4d0f5283738d9a9d0ad573df91ec9191ebeee0912dd5076336ce07bb815cb5ec9926a73d66ede0001795df6fd86075360947ba46a67c8de8edc38d86b0190b7d55566716cd1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12e3d500283f2687a81a904ee94d752e5711fa20fb21004662e77e7d8da54a58f82ed6637138e1ba1fb3bfaeea5c5a401dc1ac472344ce4d675b49f688f40cf066d0beb9fe56d2037f741ceb5447420ac1a9a22d6e6372e170a6cb5acd10c750c3cee6d509a29bd15aa220edfa25aaadfefa439bdc342e8e8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h175e1b657c3dd3d9e24b6e6db70136b39075271f46a8fa3d44d048193600dbcca45591798804c5e88845e88f0b80a47d22c7a04cf118d6dd3aafc6e11abd00c50423861c9adc8ca0acfebf6d8964b697a0d3f6ee5d031f1ed468ee8f238fc1400f71ed51c50fbf1b11b6860b0c986191b13a8086577fba7a1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b3b93882a070daf5fd4948df815b4cf8a52e390f1dd60ba8ca1c3449fd85843777e7bfa3b1072d8e0906903a0406256649547b62c1b5dc49951dbe4454df6ac785b725016f86e73dedfe7e7a852127b758d61afdcd2b7b9381150ffe7de5115a66849961f0d51a8a5ce550efde4b5422c3d9491431103bd6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1617c06c6832c836bd028a7f6e3b9f139411413c89cb4d16fc10bbbd884f9326bd2bea06061ebe9e74e891f8dbc79e240202c344969b26281f263cc3d949f445d918330776579455a12a904abde8594e77fa15be5ed0590a60e53f92708255e12ae581a21c8aefffbfdd8f6ad82296c087e2f01c2f5f7e9a0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19baf5dbe55e0345a30e0869d3bb922be56e1d8b953f04a427d638662d21b2d36404fbd4cb98c8887b4972d635944880c1e0a5f72458af96fe827fc215d489657306548cc5a652355bd9247415dab25233452e101106fd1e1974915051cb918616c28c4ce2751786a4bc55bd21638ff50164c9ef11b37545d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11d39862b68b0008d4ea4f31ef08f5580af969d57f3f1bbcc26c7d0ef0a368acda00091616d2de09d3f3a86064a46b363a47b6c334bec03251b28e9bca5c67716d31b6f5c5c5d5f1d9a17623a14744e4395e10f2c0d5f59ae6f5d1176be18b9e5d7152db493b55ca54e149ddf12662d5278b9428de0114e5c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd1e9b982bd45123dadf143e2a88ec6aba89f39173835bd98d5f38034cea30e447d0a8f65d7efce113cd310878622fa0bd63823bf19f17d5c0a8ba39234dce4fbf47ecfb37913090360d6a01043d96e480c89a60ca43e2639e849b4b5847c1c1a1a99c36022addcd846a37fdac1f288447b3f1d02352f9590;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9dc5c510c5a5812a1e8b43b2a94c201c2dbc9f4dcb929e1f9d02b19c60cf2d957d54471103d66c815657986ef79e71e25a5c9f9af15359acedfe5ea05da36cd3937175b000bccd4874361e02610ac637d64b9b5c83989b802c129e888a6669267fda893ef3d8e7c73dc270af590e0c51f62750267173b436;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3ed51af67ceea78105a4d10b4174b5199635c3d0753335a36f49cde88938492f69399c009f3d8992217a77feeda6729a855b336c665bec26296ad2094f0978706849c817c2970b2ef2a85cba18ad380c506894b95808287a1da1895f34205eda00057a8e38660792d411a5afcbd088d1645c18af6041ee9d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha3c17bac86ca1b7747950e9497a2111ffa219d86790ccd4aa15bd06279e4e378e85a746f340300bf387a5708504a8d571798fa1d32c9b71b41951b4f34d41e4f2b3f57622b6166ec4f63c15a558ff55bbaab7f2de5977a444bac6fe215dfe61b009008e60b918feb0770555f71a66d5a2886d25d67fdba72;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3f56f379d13c164a043945e3af1ea943280138f76b384446036f51ab1079be7ca2ceff76b59933fd850b662f8d1d08df7887cf4d4c9810db71d04ac9eb7556d0d0d7793d16120be75cb3f80eda7af4361f01b13de4209e6a7c47247761f427407a59c308cdaa4c45e6aaf66d4c85d6bfa8707e650c8ecf12;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc783355b1cbdce87e12d2b8be5c3fe9e075839ef340982b8bbaa62fe9421f0a5572cc2deee4dbe7dc01219e1a24fbc7c2425fe02e79d1d3dc8201df24c74b5816e4874a985bae6a84b4f6c05cfed46cc617f10044b5696d878897e0804aa9b16a61bb46ad040330a5f22c4413d3342799c81b338939d3f43;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h107a334d6b2b87c7f4017111167b30bf20d5886679c895c74482b1128b27fb7a089e5bcd36edfa982d01e9eff76fc8e86fdf7a7fbb87ae6fa32413d71e910700dcbe43ced14965c2d74e879e7273af11728d5a93fc90075080b3df95a4f94819ebccdf8a401a5857395f1238796beaa9d1edb5b0e9f3f5436;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1265f7713568ad2c4252d29d66fcabf35d49bfa046733c9769900f640923872ebc04de1e28d4e461c5d194a5b29f56564e41c78efb93ad61169106c4ed1022e084ef8bc1a5222dfbee872387960cb5b74bdca583d740139e93befc8b9dd7dc741e5ba1bf8223aff9c40ea7f634c108e1d92a63060b9b3f05a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cd7ca5429a6cac191c839a535c4ccb0986eaa02b5a302f022426ac5e894c84b6f1b0fbdee0bbb4f52158d4a70c82643d827bb8f4f2039800086aa810fa4b224f4cdc2001ed8c11f7ab1a626cb262744dc674d395af66386649ab4ee1ce8cdf6a119159386dee70a6fe6eb450558f73b38b9a478973ad1660;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11f994bcd242755efcf78dee2bcca26aab8c6e9a6f5d8e1e46c531fe46cd687bdd40423fe6427c336af9c8d0fdf356de16d55964db816a4c5d50f39370f7beea3d36c35b24de79ab66ffa3c122b03726eabe2ef23b29aff87562ba8ce64f2fcd04f4398931c0f8d43d94715dfc96ff478f5da3173c8ec782f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16873a6aff84b139aeb8ce4ff90b97756b286a9f821b32f064f84977f94cf74388536246a844992dbf0cf85800c9495aa0557e343034bd43399871b84c26f7287a9c01753df71996b4a96d716e2bc181623c8960d0525cd4a9da1fa9f102078742eba0a750e0a7ac684ecef883f2e80a50f58d4a8396b1c86;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10abd8a6292889283e0304737eb8f191b20ea0c27878e2d5ad76aba291bd10f998d7a8056ac08f008fc539df8ab0be73fddae027f2393ff1d4b052c350bf0747a46616f74df2a382a7de4d44bb6a49d3ffddd7eab53b103a6ef53b8b75a65f691a98e2fbf848982dcb29dd3524d2c1e4b9ffab8eb5b78fa87;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha848e5f6d23b37f584fcf31b2ed1d46fe31ffbdfea18e74c1957dbbe4044cae87f576cbc660b0dc6c4193203ada12ea9f70e2a6bafb5f9048afce146598adb4da9fa52dca0e12870089b120fe173d66e2dcb03ca9391fcabf0decaca736d42a429f006f6f1e024c7598efa4a6932e4bf33c5d2835e1288a4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h89646e7ab83ba2da0ab311156bdda284656f53c7e83a3326cceaf2db6005f138e90b5537f9ee56ce4d11be4df2e76c3a37f18f2f67d4dc7261b0b7fdf441b1ebde2e1f9833d9b8f9131d83bc6e4e1397fda84fa850024a8a32b2661bbac59462c3985c30ec7abed62951a0cc5b0bb52251c14e4f993f3d6e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h694973da34cfd933e46553f6e0cc18f831cc50f17b8109df7ff660bb6d5b69260bc0915efeac052c36cd22020d4e8e99875c4c0416d9da9bc3010c00a08f3c49dd00e24378af44953c04402584a2c5c4354da0bec40f31875cdb94bd8ad73fe636ba6167d7c9e02e24ec1dedffd1fdd61957da3de5d6ca4e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h128d3202639d431d2672d2f1713ebf29d0d89fb2004dea9d08453eec81a226945d7472a19f2937106d6fbd0dd8c14eb4624df6cbed5a93b7288b13912733a2fff64ed121561465a18676fdde449fea7e96b53a5e6e64e49b91a6b1924ac738263408f6c718fe77cf93ec952a1e3ff7d5874cfa9840ea4c048;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbc2f86b2c3bcf68f8cd7012d5a5a4d91f428e393b1c2d7b96721621f7bc2ed69e65f899073c563bfc6ed733315cd012c6b24191e6c32cce9fcf8c2effbecc451501a25675ca1ba84ab7f42d536ea952ac64d9c4a743b12d568b885577cd56971a0014d3153421d429d4d59236a7b420d672b03fcef8de214;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc1a7914f865c30828c014be08ed67c667fbc026b70cce0d3417c10963eec83e9f2e89be124f562b236e0c141ca1b46762e6901be88e7e91e0a75465e08499da05b6167362e7142484fd0fc5d6818b9877ee1ce1977efbdb5d216b543f11846806708927e431a03a3a81e6346564cc4699abcc16998b48b61;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6c9ac0970dd9c47d7df79c1bd139ba75329dce66307e2c488719d7c956ac711b453d14381356779be32709f3de95eaf1b7ad41090644824882c480900ebee89078ed1f396ab2125959920dc528f71ac345a389ccc2a115e9f07e2798fb9ef3c7a06872ce86715fc263745dce3506ec51ae876301b9c4dc59;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf4f5a881370f7a0e590f4bc5a7aff755e8d4bd1bb7c365c642c7c0ee0a695ee39290cd28eb146d4b0bfdd581e7b7c51ded234b3cb741c43c51bf0749f6fe916ed5c93768d9c8407c535995cc90668649ecc8bdd3af99a9d4cc5a8824f70890afa3b4b8dcb6975974e5701a6a9babd472bde595a96da35123;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hac77596503c65b70fa3392575c9ad1c7900af01207c04a4b6e6259a727e3a6d30f85a56678ff4df278c8066f2d96601664ba8a99b568edff10091fbd58af97667c61fa1085676e9b25cddca9d8ff03a54010159b93c70323b257c163e789bc3e7099a9c69b393efc4258486d446ef4cefa2ca60deed633e4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13851982bf4c84f2510adc9574667dea267ace99d996dd8385f1cf8cacc910be29e10f742732f1734065fe27cc537a4592110472b87be60db9d337d60485d4ff2d1a7ce1c61dfc5452d3ced7ca65dafd820f8d1734a57da22a7c4a2c7d9e6d543fc5a4eebc254815b47815d9cdfadbca04e465105c3daa471;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hafad476313cf9cc9cac1ccde338864775401800418d9a1916e829686898e45cec31b72de3212e27d873e5943a9e257400a571585e2b3b05b4a146c2621d56391c3e4de788b4149d7c3dbe7177ea5b4b200f317513debeb3f5dad813997fb4def49f41e040d03a3edacf8ec0c2a06693208123c1d78dd67dd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5d50c10f5cb8d73d4f18c574a7c4853cd417f7f58b57b5caf3efff94eb65512ff928a5b18d7ea5f05cd438323f1601b351a245e3ba27fd7a7ccf95095f31cc36e22571f71f86510220ad457ae9eb432f8654f49808dc73a45a637ffd5e1a9f58fb10849cc432b08aadcd85187bd5e41c6aef75d3d3c9273e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6d657f254c5f8fb6d31758c80fbc01f58f816aebfdd50b14c6f5be475e5d34c0fd4894352a261fb912c0f19610519f4b3598d97030634669743f06b1cd51b014e0af2eeba93107cdfe93af97e75c2ade038f4f11fe6a44b829029aa48859b4c0079a4763d82eaca62acc1cf35f12f66b0f6cf631f922448;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14cd97672c0528b0e7796881c403aa8eca283f09def6baffafa3dc00b9f90633cae675a2214d1da7d71c122c5576d6b9a053370d5290bf885dd55735e096b6c3d53c01caf7951285e99b8dd24591978b71ef4bf367a61ea558cd33ed191e3ce5d303aaada2f4bb43caa92f279299bbca8820a844830e76d5c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3cab0c8f260f1b791ea4838032b241364d043f4b6dd557fc2ced11bdc82f23309ceda3eb7c92382ddcf4794a9b3ea5620640e1d2cb2a9bacdb7c3e0550f98b07e2fcee0d1bf910945b933c13129899661f783181dd20237f6d17cedc5dc7a5a321429afe8d7aee44e8eb422d0fd5a0e3759c58840d6b60a1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14eccfe6b838af1cacf94cbf513a10af4cf62fed77e72d1a08b59f4a6089a37b391f0ab558defff14516099ea43caa172e1921329db2deed1203a5d98a665f95bcccd0d393f267b59ff4f9d22080a00d75073f5a15e49966b14a2d15a169ae18a522c3e3be7fd1a05b786fc2a3832102ec6c269ac47fb29ff;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fe290acd818fcdc6f5deb4287dd6baccc8e050fe8e726e261cadfc76031dfa8ab9964deb54008cdb2f4a81d69fd426949566946f3458d809a18cb8e521d05b03ee68bdc05cb8f3379b8b84689e181a4fd8bfb595b20b73381d551dc78b807d57a5893fe404654436c7379290f2747830e966a7376e48d2d2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdd4639cfea68e79c0c1b6a7cfcad58699de6e760969415008cc9cb0b3bfae86372600286e3390abaeccb8f1a964c64f60070e1ed19cfa7f64ffe156ebc40c12097facb0fc675651a948fe318778e0a41f5f0af5010f253d35ae41b95c8d2a2767799d6fd80ff12b713b157e96499788e4e980859f01e379;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha4b9138b3e65d9b59d1766f86bbe43da82d8dedbdaf69247c679b6f40e36c144601b1262dd5e6690a28d3745682217a5cd9cacbaec2d5435e2321ac2288eaaa995181622a33da5fb6cfd3d4614825bd4bbd31271d8287e75fecc045965a035cf2d991f357843503f4b3e2b38bed2697a28ffddcbc0613555;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h336e895a637971e0c2376ed9ea6e756d6a46b2cad4e1f0cee8a4ffb4de7c9b6dfecba3317cb977ead1c2d43888023bacc247a5985d230dae855372a5c07d013a507e24f3afc93f538c0e59a86a1f8146055c44242236bd59163316c21651d805e9e188ca9ac177309b809892a707e9db9c7a818810b81259;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e9993dcbe8d8be3d0ed01d2d0e6309785146661f02b8f92a9e1c9395402c510922482648d528da134d6e3994e3afdfb90d93c252efbf9bdbbf38fa6a8e5e2fced7ef2c3b199a4cd2300629e908aecec1555baad5607cc1ab5edcea972acd4bdde4ae3f5949bf667d04005b659fc7cd2e69fce807687d97a3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1716f8b955fd97a7108f7fc6171f37bc26cf2ac25ac50a510dbf08501fa03215d956a730b3ad4bbf2979bc38ead59932107940ca97d5bd0d09e2c83cc0d2981c91e7ef285b9d172dd1a0733e20b40eec74f1fddd4a5550e8b3f7f4845bd9b2e8caa93c474da4e430cca8f2516a18810f4fb15a64f52994a6b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6cc05934e77a67a7df6d510629f4c66ba53f9061c94778d996c3e177374563522e44850e598d2f883f2a2b7e00b21bbda227b547ba7796bf3117721d246fd8986f5c6088c0a6a3ad120d30e231b0b052cd13045492aead2df18c9971be5ec24d54357396aa9a6367a1044549129026ceda1112fd789e7f57;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b6d14536b6f80920ae434ca2872df8758564c5e9493ce87e7aa1a1e58530a44a8d100e3a7561645a2bb26d153a2332987c0194b54aff1408088542af4b063b21705678904326d4f9ffae3f013a6a2daac48d26e46216fdd3413a5b7d431a02102c7605a9f9f0ec169f37da4f57f145af9edd6acd2e86354a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd4e6058de1c83349dab135a7d011ec84ac8ff2eb216262c66c703630b3b59172c5d584339e4fd73c099e25c700b7953b9799c14a92e242f3cbbe8604fa3ff336bb9e743376e74f142a34b26afebf08e6319b84a89141a8b3732fc16a777dab72b0b2b146bd570fc40c5e99fa0cbc86396ed0922497246ba7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he2f6b28d9e89ebbdf2cf7355e31f3d58ac5b675558715546808d65c8e873fea6aefea758fcbb6ff9e775b5bb1771f7de5a2f82677f93198f986b5ed9eb1b2afd20795f72181194669115cc10f4bbf48b7d3a4069f2d5dc42aec68c3bae20c3c3a8e672fdead1c4c22b8be727463b436db52f263638b5fb1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14bebd5c8b527291598cf21fc718cbd1e0eec51eebeb4fc5f957fcc5b81f88fa3cff63942fa67abc243bb8751393d9235bcaf39a0879beb0fd33cce91605fb64b6927b45cefaed0e65d589b3643cf15c8b259f13e1777092ea91b17ae4cf0f009641b2ea16844427a83d5efe20f0c30f64d8769e7e8eec278;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aae5c3d11f2fe23e41c5d877b6f308796971b140a9fcbcf98e61cfae11de3d672a5d16e96c46008a6b41dfc27eb22baa5be7b0af949305c29b442360022e6fb8f08a1033dc21fe5570a7af4d6bce737f335a07e7613a33be934ee635861bed67d860f6c6e3905a448cfdc67f79fba5cec4d981cf0dc39539;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcbdf067f84e29dcf6460553adbc3f69bd77baf0d5cfea423460f7f239b01d450be46f32a1b4b29781f58c5dd36aeeb60d783d27f0e3ca28d5d8439cc656a6dd6424bb3b76a783455139cf46288da1fa94a2aaa461a495fc767b890ff5738af8dab21a6807016a40ff8d21a08dc182b6b6ad4ab19fc64b5ac;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h90bd4b5ea936443f5f3a6738d5d952e0034f634dda6b95c3882b15ee53d47aaabe4e39e18a5c8a2fbde96ce20850779c6e24809eefb34ebed323a8bdb3395282473ae8c1b2878c35b9c1064eb328dbf28e335bd50a2b03597a865d881607b65acc2fb3bce8ded0dc680afca24eda0ab0ff6aca590a7c46d2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb30daa1f6ee481d66c7038143e81b5567eb52eed7cc7ee4e452be530ef59dad2a4f811ead61f5cd43ca2dbc130322ba4ebe38af2e73d12ac1d5c602050e2567b96247cc02efc0bce296e8ee24eb1054c2a5c3a7c9496f951b520d8bfba9c1074704834a264b61cba744312c0f77256eee4ea82169bd36151;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h101b8c7db818dc24a3cd1fa36b3dd4f105676b22cc5172fbf02ed0d9e3518d00873d429fb4502d65cf4b4029ad0675f2ba4f19dbc3b96e2d6e12fb5634469680c34ef52938b0645fe3d1804ce71ba49d49f408fae5fc93c17fd779ff2bb3d3015becefff732b4447a6ffe9f7d7e70fbbf05c06bd4ef8ad266;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h868631833484188033ac29098db201190b59123dc86037dfa11d9c8c6ea8e59b8c41a773528b34164c2fc01a3d758a3524379dfeecf322e0e59493429dc4de044a44705df385eefa7b73ba383c4ed31d017905fdf37147121f8f0e0c64b09577f547e9c79d096825a3433ba1718625025239b047595262e3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1617080b13049c81d4fa74bd83052fe4914966bd0bfb886445efd1c5a622929e480215d5cc14e274410bbdfc0e1ba846c3fd0dd4b54b0b6222cbb6c1c1a0a35a602c53388340c561d88e76d584d3e51ceadfd6224603d7b8496c61194bb21596bb834211a2363ca85956f956b72a9ab36215965a125a699d6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc49b1d87a8621980de18e9e0501f6677d20c52108817ca7aa820dc06873b66cdc290676f9e33ed1cfa3a45d31ad0b31d8d41118eaf97942d946b75b0317b395878f66b6c4908d22a1015035c75ecd3594adbb9459377200028c0425f2c33389478664435f8ae755fdef74228677ea3194fd9faf832ae9d43;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h693d3b96d8a2950a167c579ad84e56e42bf8d2e41b8fe11752642e9f6f8fdcc2e3b20d7e58c2946dd7c415db006484045e932387405f94a0ca3869b8856055fa7b9dca4c665cc597499cd9a23bc8251b802f8fea62857949848d8f8f4207cb3aa950a7740e3cf3c0289581ba97f1b3de90fd8326f1e2ddc4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1632d079ac6b8282294f67448e0c87e78fb96da8432d0abab21254e5b7465619b9ec50c5e4014c214c9c03436006639627b9168def7d0a9c5a01a89cf66c7c62c82130d587790d160d5db4f0e7cc8185cc6329567c5d9d9abf72df4ec4fdfc114ccea1feaee84325476a27ebe5f648151ef46de6aefe38320;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18cd86bec231f4ebf2e11067dea3f7dca24c29a08fea143168e8b2781ab617b4116377320027c330abde06997e43890e2217204d79a5930a2fb7fc464355bad4d41d10b869fa6f60380293dddf13e4faba4b57f1d306a49fe912e28900b729c19cd608c3accb29915fff6381a6855f2c40b66c9b23464356e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17f7d7269d4471036dce66f2461d05c27260a01a0f91298fdef330790e04b8b3a618d04b9f16de19be8fced7645668e55971936f059e017a8a859e1d4e15cf391ee2cce91f7d23ba388faa2c8e6c8f0a97afb568c920de9817536155b54763ac51fa691258d615cd8a6e17b7674ac6d961bb74dd31037ee77;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bba387a16cc5e780982ae82c22ac7e1aa0ae1098b031f31947e96a7a8c401f36be6769b32dcd1c91a64bdb20a71a0ce1f55b69bd6354c8d260412fc75de15daae7e559d945031363911c4242f262f30748c35c345ce7fb7b7d1fd1d0d066e8050ae82f4e120233d290b8d0bcc1e936cfc6d04cd162046ea8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hda9f1b935af617767ad69fcca630ce6e142c074e2e62f40fc64bddf9cdd2df249a7b7d02582c701bbfaa97519b51cb2fbf8f9a83e7f600e62efd6170fb2b3b3960d9e932154c2c3d4d41d7b3806ff06a28e86c7246e157686a3e057071b783b75b0ff2b7291d6d1b38ff4cbb8f0bdae7e22065f32a24e616;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12be8716fd81055395807a97791ab08c527171910486f3c4e94ed1847610c4efb44c4f5ff295e83f32590058d9bc838cb1c4df2c3d830ba540eb137d8e00cf7fe585082e77792bc8a05a106b1be891b0b66fcb6ea4b6ca1e12f0af6ac20d93b82959039ff9cc20a4aea968878e4f177f74f694c7f0e5b89c7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7703eea5dd69a543290ce61b5fa7aeff625d05307aa1d113d813b8075d81e2d725cbb85fdc20413840c5cd4685153690ffb8fbaa5d0f2065050ad7c8dfcf6aa3b00b97bdb0157247d6cadba80b5ee286fdfa471e535e5f9bf049f6f5cd9213b4c9b469f1c6cd4ad91c2986c3d6ed367689a05d6bf04646a1;
        #1
        $finish();
    end
endmodule
