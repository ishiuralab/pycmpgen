module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [23:0] src25;
    reg [22:0] src26;
    reg [21:0] src27;
    reg [20:0] src28;
    reg [19:0] src29;
    reg [18:0] src30;
    reg [17:0] src31;
    reg [16:0] src32;
    reg [15:0] src33;
    reg [14:0] src34;
    reg [13:0] src35;
    reg [12:0] src36;
    reg [11:0] src37;
    reg [10:0] src38;
    reg [9:0] src39;
    reg [8:0] src40;
    reg [7:0] src41;
    reg [6:0] src42;
    reg [5:0] src43;
    reg [4:0] src44;
    reg [3:0] src45;
    reg [2:0] src46;
    reg [1:0] src47;
    reg [0:0] src48;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [49:0] srcsum;
    wire [49:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3])<<45) + ((src46[0] + src46[1] + src46[2])<<46) + ((src47[0] + src47[1])<<47) + ((src48[0])<<48);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hde58f5ec9a2adf6b57591b2ab32be369f380d29be0a66677cf4c0e294a617d46856b90d757241c863b7af2e5620ae4ba08f461d1e2bd92334b9a83b429c71701fb3d281caeea28652766dc3c5416;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h142f1e3b9efe8b8a78426c7d6a55f0bbcd1fe4da64380f986f51a783a59fd2ff64e003bd35078484af040bd80db8263d4b258fae136491044845a928394d1c731aaddf86741789be9f088e2e6cca9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d461184b855a4d4d5dfbd8bb836744c7998d2d77ef28a73bc1b7a7aae071b710c31dceffaf2801910557ce8e28f1d3cf21fad3d64a1a3ec2cf74edab5caec4edabba620bb37b4fd8207238e112bc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h50912473a36358f9caca133fba98cfc072a9ce99a4c9f87ca2040cb11067d5a4599b0c75f265382b7fc05c8097eb180cce72d873fdaa64523dfd077dd28d14df7025c986accccefff4dd573a22e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5c3895b916f6b89e9f19db579fc84d97c35ab6f4293a3e1e01a50ea05d09262f83742d21739fb02a534b0d2235d2228e7f4ced8f9b9f015457868c667111e733daf7401aa938b2d71a9a9124cbff;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ac8825e100c2aafb8caf1cd42867dd1098480d89a2af8dadc3866bcabac68764a0dd4f34f7bae493ba47ef79827a36f8943958097438f63c34cfa0d1f02a93ba81e0053c6093fa562adf2712fd9b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h91a9651d9ff1021b776af5d5a5a0c53ebc9ee79631b2e2ec78388186e8fa7b9552fdb033e5d8ab8f0a3b27b0a9d2717c5552cc9ceaf96d30ec27c66a22298301c44857625546a52e1cb53baef6dc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dacba1bb2839c378782a7ffcae3b1f86b120a2fb0bff717ed49148fd2423f7380b1a09ad695a3d71bee928843f9995549e2790cb6e37e0852a1d3605b82348bea08a6788aeb48649192404803068;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a375b249ae0d3e16dfbe8251d5d6869f02945933df80487732c07fd31064462c45fd5711d480521d25feea871e50dc5bd71f2f501236a82d164a378c7e2203281c92c465866f6c0de1abb01b7a3f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1af03e3f824cf03a7cb9b61cd45fafc568bd7c1c539e74d7624ca28cabc3e2baeb94a7ff7fd56189d9b7694c84ce989359f973f84dc23cc25fb3e747ae61d3fc209a3183acee974f182fd5cceb6af;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1572df3eab2bb025e11119007e72644d3e7e6cd6d3b7be723e4a8bbe85f7d3c1cb906364410067c136830e00896e1cecfd8ab0c6e69ba0447348a83b37427700d5a8742415ebb8ba0e431bb8c15d4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aef16fc0497f9a7dde5cc913427f0158df57aebc3a1f3b7a65108a5925927e0bc844f108a3f670a150ce44b51696505d3a12a43afa2a4d716c057222d5f7c009db5fd26b350202a44ad475184e32;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf0f4a5dfeb53024c748d9124d35d65f66b2de6c5ed985242335bd442b58db6aa1035066729494dfb577503c77385110c40fe2319f923abbe6f74e09e10bce63aed8b5ecefd4730ca6527f84c64db;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aec078a986b4407c8ded2d1289eb7c56932c549b17e6e609c245a8f81338753388cc58283a0fa4e98b68a70557779d1e33c4b2b9fc391b9d537dc66d1d46a8783ab68114a24adad1652328ee9109;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d18a3367797855692b8ca5d7d8e22b1459db16cce23ec5974514d8491018c9779e36ea59daa99c4fe7205a8b7207f9739b593e09c53a99a58688f53fbee516a6ead5386b9bfdb2a47ea1d7f396ef;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a29d60924ade141975dfabf6affe61cf1cca53639d801e0b3a501d5845707d04290382cd7bf3c69747cd286139561c041cb0353f4b4c6a797c3a57b1a8a5b2ad137eaec6fa0123baeabcc7c76bcb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1def5016fcb47ba99b99c659982c80517232fd4e79fa2254d80f98f6c9674e7727d5af167bc506bf982da640af1d2baa201fc7ba6b8aa05bc0b8f8cea3288e429c0c8271b32ffad6b27d0454bbae;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1999a34b4609fe01da42931dbc1be8f8fa1bbedaac53d48c1a0552ed6848045bdc4e5be2ced245828eea0f7a4102a052539b47fc74d20f73e2f910f07c6767ccd60e65ec890e1b3dfcbc988124b09;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bd7e2b60866abf9aed3619c3681a56364f85bc412a3086f60d90e423567e8b92a9e6dd045a607c3c18dfb8936073a043eb841cbc69b26bcf034a0587c7942196f8dbebe79a074661b68e89b619d7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5e60591d9d8a941a885a1c78ee8018ab4120c983c599ba3cbc77e2cbf42904a5b045450e4b41397b117072d10d008d7b9589a91e8f68de87bd86ff6b80d86b4a333c11056dbbbf3b60b11595cbad;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a613f4b84fd2238bea846267c1df42efa82c7e6bc459d71aada37f426a67440a33b3a0f196d89a8831d9f0e325b2db86842dc18a0227ec66867d406226f222af2cc63c3e4b3fddb3f864b5354c23;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9e9374ac307a1963ff32baaf5562e51c183767bb009e46c8cdbd56823dbae91580e0febac358d6beb896767ab978c55b65477dc72e1228764e90bcff0c6304c2cb24fc0a16be131a62bbc4d50f3b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd939a60d8dfdc86c9acd54b346bf06de9226a555c3c33fe0aef2dc35ad13e7720012abe375a620f99f0e7b69c78d937389c21faafdd25fc3d18317b523f682da45a8c25f2a70c7cb8a619ea4fd0b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1701a915f1f2580a63665c3c821742d9304368ba74115abdb63035549bec133dd32505ecd4a515a0dfc931b9d9336022ea461e695c333f2d5e40aed16434deb6e815019bef09b2f1c9c9c7e384145;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc53e6660bf5f17a404b2d612fbad2aff5e9dc466c04ec9d812772ae605a4bf35c2732ed462a515d01a7bf5420b98c6ac7aed043938fb0dd4091c0795c93a0f33392e7c4891922f1cb9b86174cc40;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h91ba31038112795b92c513f14799cba02f01d4233ec4feca25b4f2e42ae1c687e583d39c760f60bee3bcd4989068d236b4640bd150e3baf6a5cb8094e7af4174c9ec38c7ffd413271531eec31f72;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4f097c1f1ab7f4d8a5e97a76eace9f45de3433c527691ac80093d4f961532112b9c35badd67ea30becf5c62f4cf266cca493d24ef953d91a7d3044def3339c8ea0c5420385c1cc11cb0600ff75af;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hedba6791459283368e83fe6af52cd7ed0ebf8e4d23623eb46321b8a2dda3d7d1f67f482c1812bef48c6148cf2b5da0d701b4f545a7bc3557a60fc035d8c6206d1ce8b130c7c689b8d2d134373632;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ed15c69349a7d81848ccc690683c0171e28fedef5bd9bd92b3799b2f861ceeb6d0a329da195f5e00591108a46771f2c68f0949e89c35f5b002c6c1874384a3f598e621abab0d95336169788f2874;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h640d85dbb912fa54a9d8d0b667efdecf22568980364b042a10ff3a51a8bc6f2b445a37d6ea643a99615d9d6d9dba90720f05273a5c30eee647e796b06f0e9a84d03fedcccc0f78854ed57fdb6e73;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fb4f781ab9fb3da54892578fe24a9114f9228f08226cf646d570af4e18fda647b0d5faaaaeac7023ac1366be0fda95f9557c3d1657f475788cf0da295c87ee98a04928e2976e9a6c7a9d64ef520a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6837e057e81a19f83a062212d1f9d3fc2f1d9594fcdc5c2a9ffc08d3d49895782861a05b991c27ae08d2def1aac82f6ec0bb46883a4e097086a9c4afdfb73b83d6243f62938c7f60e4aa78c37796;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f1ab2eb35085e3645dc72f9514d7c684993667e1187af912473999c49e1e218ae243c1b5fe03e89806285b9383b501b5c651f9be169d6d7788fb3122878165205cbe90a51fef344801396a80d3ca;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b024563dd959aa91bc980c19d0fe9a74bd1e452873b794ed684da46c93fedd533afa7cbd5ae073dea9e66f73173950fbec9c1d0e55d1caaf0349e14f92cc2a74f60eec45466ce35f79c92a81b0cb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3bc450e23c66b35b4c5be36146ef367fbd34e6fbd3be21c85f36f3f8651a593638da23825babf60719413a3477f194e13f16bb1a7025b816a50b5d1e59479164e538721079ae990e60ce2044cbb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c8741ed855f551cad9bb0f60df85a781cf21e555066209d5b47a1aa16b0821afc6bc8d3987d2cc6dacc4745ec677314d2bda7aaff9684cc9001069fe95a1ac6c1584b04d01caec098a9738ae7a85;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9a137bee317739deb0a3331a602ce3f2dd730fcfe867ce8667fb91cf993a79e987956b55b4b2a22bc1a23f35bf0946f6fa03efdf05700d5a5c8594d73489e64103c070fa969baa927bbe91f004af;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6efa7000ba992179c3c1f5089bc2c48b61b757a3d28fc7245ac0e19e811d0ec6e38b4101dbfe5f96cc520a5df8f3bae5f6345bdbaddbe4e590e8f96fd9145b335136b641f0f1ef36744145f3a5a9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h137bb9d6eaafb51aa4c93d93ee5a1128cc8010e4061460d75461619c7c6fad189f845f42274ba29e5272677ec0dc743d0601bea4d722d817fefc5af47d7c6a48573c2f2159945b9a14d021551d81c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf9cdd6975c4413100566acc50d1ec459f5002cd571c95dbc1b3e01ebcd8f07858bf84493c7b25ded175e9b4ba29f9fce371bebe1b68e143dba5c554d0d4b8b1e10b6b9abd629d7562a934a10783e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6bfd88c05db198ee135a2d7561e4ba73f8104e597e55dde79d563e19f952d447518b05f0d6bb39c8f59b0a64b1ccfbbf46c3ca12ed2f49c757a81e3e7692ac8a85a2f122892e863769a7b9b8a3a1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb273b8c5cfb3a8b2e57c9523f6b14cf36bdc5914cb32ba2098c95aa74c52634d5eb188813fedb599eab22d46f622c45cfa6d75cb522b48fd75e9da120254956eb16490fc06b5f86995e0ebaea782;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h59bba71418ed98eb52c00340ed22a0a4325f1a5b4f695c01f105146a7cfe49fcd669130df3377598243d125a0692f543bd1aaae6cf05632ed31f53a5a843b7ca657f5cc4c13779697362145523ec;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16507317749d50d4aec6906e2f15f2f2062dad0a5f5a7771843e11d12b4072bfe2f4c567f44f59f7b391642fbf24096ba3430c110d76d6b3e5ec5d872b83275888df1fbd01c45f62767d04d0399cf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2ea98e7c231a86bf216cff9405fcc46d182223f70c5e8f4d4a21fc18d472bceb161a1c44897201bc719950e4f67ece8edf07787bdd6c00d2b3e8acf0953cc4c467eeae4c9f49e08fc4d533073e67;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c12b6a9bec2f4284ec22211ad8fa051d706d0442b212e11816a15d55bf836970e551a948c957a631a8ebdbd52765e870a17a66612e199350a424e8465b53cb438fa1be3e42205c481336f79aeb43;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h77ec7476e6830f3ca0d34d654823feb85c9d1ed16aea882a29cf0a09f4688fee6c51a36e4b7d4a7fdba01699e4a5ce31b4d360aebea1359f82474dbd1a736807bf698df1f72a518ad713215aa0be;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h251d7e17277cd9bb6f6a0932c41ebd289c780011a3665e8ddc0620f1cc55412ad5f7f712052318967ffdb3daee3565a92ecd8b0430214b081bb92ba487017c1133309912c51441c784848f72486c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h140f9b7c24bf9830bc552b93c4035ceed4e38b2f2cf4ed7d0cddf78f5d9af28ee90e715ec6db8ba69e2283febdb6b5b45a13328772576947053e801db0215d889012bee6646943344b6fd3734a831;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6b668af9bd36a9116110e6af1213f0426dcc134d05fbc2995c2c19c66252c7e757e6d61cc48001c91c2b563a00ac67d877cc842d02a7f89d77a688ef8717b832b0307645e8e54565a0a47ccb98f3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18138e6e1f9524dfb026c3db0aa6d0290b7312bbd727fb51d540bc2f01d53e2fb4324ff4720a6db70e3d10a1817640d28f37822c3ad5e19e9661e8d80e13844784d19b280aae33980824b79795a1d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf2bf2a5b1c16ebc36f6d5e22e825f130fcbd3abcdd59962ee1fb1b1248bdb8519dd8ff290a2a1cfc1c40c6eddbfe067bf5486e86dfd423d2fdddd6fa74f74f0d6cdd89138ca2ae57fcb4fec90836;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hac5fd60339911561f2e09c611bf58d7f06fe0ebb588bd4a89590bd037b5648686e65bc0af30bab0cabc910e54f6925fde7c0d4d06bb5472acfddb5bc596e07d00a330f62ebd76596ac054ed492ab;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2a738ce44a11756f6f15e5371b693ebc62ca89f99a30488a0478ac51c3d33524a7e3c6e8c5e95b39b2b69e72438edb4c74e1f14f58b725828e8fb9ef6ef01da42a90c3432abed7c739008b91a42d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a31bd037b1326076ce081b52e04a7440d6e245475889253b08e5b5ecfed5587a8682f42ba5fbacc27d65ebd69f505b7c7638496f76450ac2a6154b0a6ad8911d8ca3d8b26d1ccdd4c88515f7ff1b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he8c7efff0eb4ea0a211e71821b082cb42b03708f23c2f93cd3f884db77745ce40536ca769a646e56c140f66ee7b498a26ce93bd601b938e33945ab05d441db0cf0c291c423439f28addc8b334c81;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b912817b7616d76a0bcb68cd948990d0ad9a965c8eace9c637abcbf4ebeacaf726a374c0a7c4c8f4abe865cea4e5bc88254a9800928c03d6ced253688fc719d84605fca2df52fb07bdc8abe1b6c1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11091f8077787d5c9478a8c77832e60986b2bd0f650856882a0aea63f00e6bdf49ab163f0270300df1385af618a2282c4b5519278d6d508334eff73f7ad0d8cb266c6f9686eb4fddd5dab91cf39d1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1778717cfc751c29b71b4f98cc577b12171f3ec6e495049de18f7afc0c6d76db7b466b8028bc0a99e12a56aae5bf815c93bec1702d0449082c6341aac75eaa4694e2f61d245debf661ea09da565f3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1397fe04f143de7888a9be07acbfa76342edafc860529e2278e5215359fa9bbd9f8657eb78f3d363ec22c86c577cde490fc9a034ba51454947f3e9f312c5e7d3fff05ee03dea00a02af82c9aa8bb6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15385553ed4eae6c6b23b0975ea2137e4cca8991d2858899b4c978294c7a385d08e5e9c45b6c8304e51869ccf1aa856d514f273d12cc10934df18e02306e60bba2e5bc92ab6a9c2fb90a11f1cd48f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a23a768c16742ebc68aeb2c629a5b417b8a6caa3898aeee354cbeb9d8110ecbfc93d0f7afc6a926f237109790a7da46685e2e190f76603b33a19b2dc003e6fcba719d765f36c6465c080b443ca5a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17161c91f47f9dc6bb497f698a65969447261bc00924a709b786bef53f41afb425cf19e873bebdccf6642cd9eecd67cc62c89bad1fadaf22d2eaed814317394355f3c1e6e23a2815226845bbe12cc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd81dbb53114ea2fadf9f2109cfa7c1ca17ae395d90065119b1b263c7bfbe4616afe6b0c0b563fd9a5024bad4884d426921d73b35423859cd029ffc0a15501690cb052bde78a897c2a8f4daed23cd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h918db621c983329e7a1b578c57cc37ac84df5884d7c66285bcefc0289217dfb64038948b71625b2df8787ebbe0dfc08d197252b18bcc638c87f66eb8de6948d6774f9be74c1bce0fd829e1834576;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b24be3dc80e883f2f6628d41afe71098d134c4dfe157342b1968f7828f698ac4b594f355c5523e095fd83ae0d3a3c25ef1cc79c0fcbfe8f14699132c03c8eb473a5a9b55d99a379705235cde3854;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5918cfce2dea500bc97a0c642c505899d2ebc7ffaaa109e2e1afbf9398f703d616a8c1cd85a9ca1f9c8d3d131b405b43421795befd4a2d32f8dc372e19b0f02426945108bf039e259774e52d1118;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb750d396855f04165c847605db5734800453988dc1d835920fd5ee2b2f639e6efc615b3122f2928479fea7b0ee23e3a4e29636d315debcdada068f00a2fd19084dfb64ae9d01299d1c6d8a587c1c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bea1ea2a0f0e5dfdcf8357cbb092c603c8a40895484c93067d95da909ae65516584522f0b31a5530086613b73d974518a01b4ed36a4cfb366fac6825ae9aefd74a6978d18a6c91ca186be4a50b01;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dbcb599412f8d32c492c15829195e72107e0d903d0c892a7293220a7ea7ff4eb9281cee54289752ef9fcc5167f1377e1b0a2602b1dce20f67c5f9f84f23f80288db100d9cc70ef361cd48adfb039;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf106d8b22d1fe05ca516146ee708895055e4e8b523fefea2eeb94238f16dcae8d164ffa3af67ff16f68edd6fd4d8b27d85c4aba8ad54bf6c159c901b65f343c56b30c05607dcab0005c10996b993;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8ccb33f6c2bb2c48315cf02da315f8df331ae49e0c62f5ed2141e41538ef20f6730df0f4378d33b5e5cc089e941421fabeabb64fbbf3e1cfdc45f1ec0e778d0ddad3a3b0bb33744de820475e1c01;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h157d22c4c83e522fb1713baa6f072532dcc239fb94c599441d965eada393dac92e5cc7ad7287f085e19c62ba4b47becab962bef280f93043ac5deedde258a28fdd6d579daefdadf633d12611022a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f115ad2274916bded431ac8cf9e1b3763e05c8c9a1366644f7b5e5788e7ffef1fc3880182efb5e7790acb5ac4d97d2bc1fd7eb522ad468bea5770be16b3329fee5f5833d754faac2db0b85ab8a7d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c3b7a7ecea65e906866213239e9e495d17e7a9304a03237767d029a057ab545c48b6fae1fe956e78c65662679fad1c2046c813ac19a06ab8dc9db965dfd80751cf98e9895845bf42674969fe013f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d9f8213a9fb6f46e2d66e4a4f49e715e1e0ab4e031a9b9c695d3d520be64b34a7bf838d8ff9d35546ae5473b4c858caeabd7920d1ffbce2f17d2b2a20d2c29c884161aea783904440b7a765d3b4e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h138297715e7610741586d3e7db9bafcc3d5e107f110a4dbca16774cf0bccbb79fd7a989ca3db978655e446aaf1323da561323ca843ca64f9004389e16bd063ec2efd197e191659e403c550d8187be;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h817cd2e712139beecd280da5c580340c87630e5fb8e9ffa70ebc17b5120e79a50c8bf86b0606ca059c544e8114b96c25c2bb093f2c7fe8969a576e209fd685c4463ebd8dc294d1bfea336e0e3629;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d4846abede061224075a2ae34a1de2804c8635778048c27508646637a32259e79fcf5ec12655ad0631db4330d8aa213eb707c1feb3d77158ca8ca07bbb23083b21df6963c849645ed629c43e647b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc0cb531f2ce28ff7e3f4f9de34eb22628ff8ebf2780f996154dadf16125f9fb760ac9740d541f14d537130de5790871bd719e3d43165bf4b263889ff1b6aa0beb9a0bc2e30ac6f74c44c524e90fa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3d7fac5925d3924a1f4e7be221c745fa0e13d393067d0b8241fd508ebe21698c0ab9008c0d821cefddacf27e1baa45870e8cf1977eee39cbbae186abcd9006b4c3831c90ca90a7792119332b0d9d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1afbfb77228e04d074c9bfd08e89439e980590ac99e76335acd7d68e146efc565774bef4dad2af6494cbe89a3022898709a66b39931c0b97c2aa8a8e6511c0ca66bd3fb8aba87fe454ca7f3622bb2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h923bef913715d2beb06a0d4a50ed71d4a3a0d8ab77ec73ffe2c9350cb4322bf241d101d2883ab349f87b273e9302e62bf7b05495ea3152d1e59d1c964759da3585fe2270db8234ac8d1dc1c2a590;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1365bff3c4df90455ea2e3b3fdf82e2cd166baeb95b591fb4bd723210e60b9052ab0828236b52dd7276978c8cb08973eca5d22871889d75ab24feb0f2163f45c306f1769b5afc9d1a4dbfe8ca1784;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd4c10b8846e04f0a85f06663f9cd6232289615afdec8a454cc3ddc450f1c0539c0c38ed52632c0c5483a6574946c2de1664225d4f38b6e8ca9bbed71ee1fd66c58c5632e305056a6c27f91f97d9e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h118a2c481b31723d0b802b60860c7c21aab3a5630f40e2c59928eff957356249fa1831077b483d04a143a160efd97d5ab49236b8982a2c4e3a06b2dd8cb10419c558f07b046408fba6de03f92a443;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc99d5988645ba3238da0c18e3255983cb2fe88ab48518f83eccad8db0518faaaaf80fae2a15056d5edf76f334029c350c3f7c14c827a2ccefaf2abad9c5300272738be35e920ae71dbd045e48a35;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c100efcd4a3da5a1e88deee717851a9d5bf324f17283a0600a7d94ab67896ac32a22e7c80d56c91dabd44d780dfe5ff476b8e4b57f40ea1fe022f22986a06942605d85110d50bd643aacb2c919d0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h34cecd2f85fcb350b2b035b05c0bb6068a7a4b2418878391fd5455041777f99724f055df14c633e1936fa27d8f081169d97cd6dfc1869cd5954218ace72e357d1e34f8898507ee1455e0c4560e4c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5392db3324021356094f96585ebbb320967c87dbfa6e2630f206d0303a2b3a07d3e663701e6bc60856b2ac15fde18c524695dd55064af3db0a5d52a999c57e09d0010346cef8299592858cfdf620;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1661519cac09b799d7a13852b154e5e20d634dc966a5808e25de38e14fcc18b27c10dd134e3d4f8231eeb55ab98873c7b736149c3b2dad25e18dbf6778beba3f94d23be74a08f4b72d3bcea32611e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc97ccbd5c3b20be5f57781312b4cda2942265703b98632a62727de06d6be5b73afec26ea2e4792bfe187f4924fe2422d902fd3954103bd814ff3cde00ea1966247cfe52b71926bdf8e499903dd4d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h169cc57fc87c43d3601783bf2ac49a4e3fc106b4e17028952068523130547d2f4464b2d7bd5d579a85fbf8a3f465325f26f945db0d3b6671d41ead840367b97a4639ef1f4dc2d456758526d3ea300;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h82ddb16d637f22d956c3bc149b644c499eeb1ed09429de8b7d3d8904a557f148fb5e91de7c2e2a683f9ca7e938d009d12c0f8d39d135febef1dc8a076268d77b94ccd117cbf1473886efaa36bfb2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heb2b41ac4e1fb6bb8df4eadfbafa4d6f8c236c31df06fb1c8ac87449b273bfb19efbbc1e64718f54102cd77c6319158ed623e0c4043dafaaa7dc7e7b35e394574137f6f0d0897307c274ead78eab;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e8deb2cff31f289336cb338fbacd8d6795e42ff3c3eea884aeafce7cde47b0837655963865cf55bd4d122ebd7ff2bbe0f2ec73761e4ca65c4dc1c5d76571e47924892dd9e5318b94864e522a4a90;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eea18efda30dfd6e97bf0564e4163a5f5315d1c8f963b1548eb0ee1a58c7cedf06cbd7f9a49000e981faa1eacb918678783b5a7646d5f4249272e7fdc365627c57ee146fb70ce81dd8c9b743a46f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13c253a679d6948fd296918ed1396edbc957e9830cf96f289c4831fe3aabff1c01f4a657e5f300ec85cc63b7f1fbca30410cd544a2f24c94dcb3b9e72ab5400be664e33442079bb2d77f9709b352c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19ed8a7423a249b255f936d39e4b8fc2a591f80be4cade5c761245b676f16584cac5ae491ba19f20e2e7e455cab5ec669e844e802cd3656bcc72cfe8b0f3acf128928ab3f865efe234be4063c37b8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15b10b7c81cbb902283caf266c112c228917dd910d258b52fc1a3b41b5af6332b0396c23ed28151ad12e29e70ff9b217ea4fd985523822e1b5b04d152c5bdcbc94e73ce3a6343e524668dfae45dfa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6a0a3440e166868df5e64b6ae36a147e78c84d3ac7c580345cc61ddbccd0530f463f637d1fc633146bfa68ea934b956f18f11e908ec94effd53b1217e3c4f61ac1c625bf8f11b0883bb14b871846;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18088839a400ba4d8435c875784f443badf18a49187f0b24b2c7608fe42b64586c5457a2741a369c9e66f62d076edd04deb9233208aab277b801cd1e54951f41e5afe549619134717da03236e8e3a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19f57d2320b5a2bd29fb035e97e219b5ae5c58f9de3dd027c0570400f8825937657283d007ee5f88de3f72855780fe1958ce44acec5ff381d28edf5a04c1c3bf68a23fe304865ff586d13e7e1661b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f15a82b9bb2e2c774ed232fa700f3919f478cd8907b7c9e28b289334c552d174bda9681e580b5bfb49d4743ec95cf791820981765c36486c6584cfc2676164615245a76ea86305b1830c8782d027;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he0da24369f0a7c9e81a5d72dfeb6ed167c597b967d1fc7caa0f186e3b56d35c29432ee8e9b9bef8108c8ea098cdef1b5068908af6cd19c6449d2f48f45c4e9c4170387a4247fc6ac1fdfa6490c7a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dc9d1ec97badcf7ac4d8b1356300a64f0973acfaaa5de34d82ece2a8a36e4d0e061bf8e98398f37bf59ffd8319a846661be29679f69a44d0663e5b2a33fb63ddf20498cd2749164f219a071e679b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19735e1bcdf418e9799b473b648550b17c692594d7af19d1ee8cb1f56d2adaa024de88fb751f1282e5eb908658042e84d0cb67a647363a3377069678cc3d4e6487687924a2e8d0ab51f417cf5da44;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h162e34af292b36e9efc1835a4ae9fac4eb2d064e21bf6c0d22a57973e61f6a592c73e16e30a4cc13a3459a1ac5368a549fdde10eb5908590b932faba735691ca16d8a7661616c0b730275999889b8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c7259bd2b60d8d97ee4ab898950fc871acf726daa9bea3cd6c8a269e6457818649993a72f98eb426bb12285e447971222004e9d7a0806793569220d48e1577270cfdb7077c7ec0682898cbbf95a8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h200eddae4e7e8a75ef4090063143f11d1ecfce09d2c04f2f9bf35166e8f932cb216c1f3c2fc0d883ac0c79ce0de206eef0ceb1cab61cde0531ea0da47a34e50f6ef80fcd1b17bfaae768ccd36cf0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd9b61cfaec386c447d3155d463ec7e52c4d91c21993e8ed1f8cf384de37b3d76b4d4bff7f67f0931c2ad4cb7232d6e594a738924dbd60ca5a104bdc04b0f621339c7ef3fe988b3ff3998f36d126b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h35d9521792615f8148c7bc1348cbcc0a6f73cf5451ac0c3e7d791fc9e00dadfd14add4a2e67bb3a43295f8ea84e154230e636c750fae8af1b54bd12668e9c9104457a6b67db8436652fcd5dd956e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11fd95b728bce34bd12962754d992653910675a7a4a46ae956c60b770da0b89c8cd83b8bf8cc2018b6c0d4ce7b724e0a434da2daa0ed8590bf1ecfcbc06ab3d568929e8497f73150299ad7a42db24;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h190e2d9bc80951e60eea1a12ca954cefca2fb2a0f3426784e3bfa39d26cfe534795e108b238100c3cdbe750a24d2d17e44633006bafd62260fe0ebf5a2269881db8ecf77df1255645a2a712ebd6f2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h85d385b6f1cfdcb2842b34c6363c890e4b5935ec1da9888e3c7017f52cc6cc9cbae9bdc12d2fca4cdd228309f7e7f151444d182b07ba059ca6cd645d9bc3ddb17bf4b3b2f6e820fd81998d795d4e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1259a5365a483c8f8beaeb69deb2cbe85bf174b8192faaab9a5fc51c9ba46529d2424c5adecb5a3bcb2abd5167224e0c8d74d413c8d85f3d02e073e5972e6bd77a953db4f7750437ee552ae29feda;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16c204c926c3e6055cad2dbbda55cd22888aa9b46e845d1a66da73c55e28801978283149828813bb64acf2e38aec9127de9f86010ce184eb33823ea0f890880fccd15f58980e9dde49377be32b4f0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbc35fa43a46631ffbf6ae660285f448c927e14f3a8d746c88b618af0d83f18e43098eade3f4bef75b3fd1cd5450384b17fc0e41b670935104f1da2d8993bc27426751ed413e56ce764ca7579ff22;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hed649ac0b55726277cb7730d56d9c910ef0066b7d02b9a4c8b049b2154d5f0b8b417fa693d55803b619a14101428173767f64a2d4f67b655a645e333e5b0addd27d55536872f310fef11c4001904;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1597ff4f4934f31db2bcefef58e0e9ea744728ce9b0c3f927375719ea4a896f253d0edf9db1e2505222a6839826e715f2aca73bbe42208c04d80d7c7cb9928a7943c488627444121aaa876a4e21a3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd9b39e0b063c53442eff1802cc278f46c816fd5219e135926fcced1cdd44f1bbc8971dc3a75c6220bf475352333eb4eff8ba30372711ed2f12dafd3ed20a948c5755263ecdda1bf3d095fc9be9bf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4085f2640eb88ffeb5b90ab89e2cce9697314659955dda72175818bcc74c601f909a38efcf6e698cc4d4d646454ec988a7e949c87c41e2d31d9060d35cc5a6988c570ea63ba64a584cc2395dff4e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8a863f8ae8e356797b0825c8ef6ddf73d807cdc7c9ad882765d4d8c158be4312394a5fac70717edf6b8077da7cd232dc96e8e388b338ce1c6e9e93a1fda5bffbfe49e27b874a61b4afabdfb00c5d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h135a02f8b131a79d8561fddf667236c5bf010a94a3a959dff9017891782adf78b521f47847c095df607cb0ad105cc4ba8a2aa5e53e4ab1ef1197472eafa8f57e510fce998898c305b225905f2a258;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h103ee4b27a58a49c534783c5f57a4cedeca6f073b0823224721bcb6b7cd0a2c1c32780b11e064fdfb4f2311c373428c46ad486e37c370acc3e7f58979cc169efb14167327b291028872998419ddf6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha452d309250e8485aa2375ab34fcf51d07c3b6eab8d4e4fbd80746b7880aa30119d60ac1678590fd7affd104a55d54e92a0f58e50e7a5993ab08b221ecef474a1d2dd9ea9b367b1be03faa62191c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h863fdebf8203b7438bb2bee8a7159848743bc173f17719414b2167df9722a73412517ef21c8cee06bf1f1704d9b19b43c86323782378ce1b7330a0fff1916b5459c88e83a1043d392f094791f1a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5b908e30c50dfe6592c90a7f52a2557c49c3faf0d51d581df53bc165debf0385a409124f83902dff9cfa4a51878f90aaf4e3540c248f0cb5775cd3e11b12cc2776f654a9e2b599ffec18aaa7dc7c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb3628d7b186551714b579e0293ad12017cdf2730a5f5e7e375974465bbdc02f867a511d8f5770b608152d26568a0d1a8cdc2d2382f86c7d556c61d0e0a6520010ca7ed88183d755f14d9ab198e3d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16a7683bb5fa6ce8fd11a0540a344dd4beb7bf4214e9dcad7734cd79208978bc6ef9022be9488ce51f32e11e6307f9c5055059bf713e2b44afd36caa570e0183252b28eaad327fe85a0a6435c8f2d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h332d43c9ed0ffbf2189236e5cc84140585d8b6794b7aa8acf73f508ffd3ba9f3a7d9f4d860acc5d3ef97f2669cabd7204d53a520899391489ca5231d6d9c8605555f70c4f51a9b64253d33a83312;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11561668dc2f5aa359641952386bc14a8b66b57b699ac55a2ac3e911181910d33d29a34236406e336c07d32ee72ebdb52dc87141caf771c6c526461a7c39dd737d20432e8769db45e7038abaa8d01;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc152ff22130e0a051093627b818dcbcc7b74a39d9cafc02d7aea15d21940fb05055a1241c658686c6451019e5f4585ae725e01d2ba6b218af83815f4b94f9d14aa1f5c6381f9833822b3f6075c04;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h667c366c683bedf36ef2cfd885221c5dd0ed45707ac6a107781da8925b1a3c58096b9a4460f98ea6587744728282aa4a2c5988bcf03ead21d96b9b9889d91a6b50027edc2808b8407837ad9dd654;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3ded7dd802043fb9a53b711abe2ff6fa507210c15f8d1ae912ddf4f8dee1b47847ab3c1431b35e4ab35a25e950c88b69459fe5172b9a4f1019a64e8eac852fea80787721631aff6c5760d9551bc8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h857db685ab51cbe8a702ad452e071de9788bb5edea5571e327da8ec376bf60cadf806390190e1f07e59b643a5048e66548c19412cd96463a55a0c7a6afa8db0e798b6ba755d4f3efebd0b041503a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b2208df65792348d00b24b2c4c4186cef2eed422b970de2a6cd4b6fbaaf881c06ca2fc537bbfef90163d4cf5276c211698bc277f2419de9a360af6ea377561c5733c5ccb7be9e3f6e5880576cbb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd93b40d6e9587aabe069ff9bbea71d772f2726c894de1fe219d361c1082e3d2677326644918839da4de2e1a32713634e43f6e013630384f5d22d46b66baf2eea85ab868f397229cfa9ed85620b53;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha31c3f5ae75765753ad9024cbd1363e8421b6cd8354b335fde8e0305862a95ffa789c7fc3f3342802b83411929497e2f21f64107552ea05dc10040e87e5e3a107d0bc81b6cf1dd1a323214ba593;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1497c8b9b7ac7fe307c36261bb2799aee6df53fa4475046c5a984c08b0a345f8a90a7b9d8161ae35d0873de86da31a08cb067ddfb9f8780fcae301e9e0d29ba9a420cf6106127cf1399f66d72e786;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1892fd62eee53dfe5796e9a8175e1d4f85f33591b71f2fdabe162d4594a5b473a9ca1b969dee77ccf0cfb77b2bce96b1b00d1509154e9bf8015436c92c9a2e171633743a3888fa8ee2e0f0a5c814b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12e348e0d017ee0d8bec636c6a3d0a4d0d6c4d3b0e107bda8540a61296769a23853e68def41651492b6e811ff98ddc27ef97b5499660bf19ba8e42b80af903679a4d3cc7d87ecf032ed1a4fc8ef5a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h763f68f874b8802585992dd8c808089641718ed3bc80dcb71474a94c2fdfc17f9bf7b5bbc4eee9721ccc477e98dfe0f9767243a6eb11c925c83f0ab428724e4418833f4d9388282238170a121781;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h605fb41874c6c3d9ae46f78d78ef96287e38ffd2bf5e40dc64a14ee5d46d94adf4d8e57f12b3cb0833e0177f7ed171902bff8c9241b193456002db73a48fca00c890037b265da913552bb2d70832;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a4c780933b1067a1afe62c9e18adf536cc2aaad9223ec68a68f00dc355da16c3b2948c6104708fdf2404ac96d107ffc9b65722f91b204f04ce7f74ed9325430b24eef3fefaf5644e115dae2ff05;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h165c196afa8cf9c8b578e130bec8f7152f75b8c06c9c807e295d489393430eed98d5e8b66b686aaef10606466d61ecc5098256a94c677c6d5df4777cec3b187958e7991224a36977850682209d2db;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6a13d227520d090324232368e163e6f7663c93c98a470648828fd301a177303fe6246921399a210562c5b067781082a8d0965bbb9def3fb11d28fd66093cb76b1d67b7e54a56e58e7cc29c15fbc6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4e87be3893cf82f317dd8488f48db06fec655844a7d76963a1d37ae895cc8882b500f3b3901dfe49a72fd054788379fb6dd8b5ace9feafa28a6fe9020018f0af1c9b739d8b6675f002798dd34cc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14c4559dfbea057c8e2be4464a75136c786cf753e3a0ec4c5eadeb7808ea4e2c368772cbc4119d348d6e8b026fffa32acf4ae818e58be996d9aab22ae24ebb8aff1fda78c053d29b84ea2f221b65c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15b7a5656fe7d6c19de6368a40722dbe1d6ee37d906ebc1ccf8e80b1194ffc46b426040075c271f02c552dc9b1aa63b070f4035f0e51fe9a8510185cb824c859b08491dee20ba47be1f0d5964f39b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h85c667e83065dd57661d4d8a171cb5a692c6708e2b3f15fd4caac66beb8784c85c3f718bddf4ba7294170d9017d3f2fa815588b0b6aa7978b86db47c6a4ccf72f9f80d23318ceadbb51570860171;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aea0e4f1e399aab8ed49bf4ca955f87a152840bcfc3d31f9a002bec99a18f913e610ea1ffd25da1f4a1995815fa647a63629284def2b0f2b3f75853b7e8e873f7c0936e362e977202a3dd125df70;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb569f01592fab689797c5fbdecd99b066c415b7d764f8d533a485efacbbd7b32954f150322e9c620fa08a68134b2227c8915ca8b5caa6ca2ea61597a38e8dc883b9b83d94e3d5b262eec165d8c4c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h491326c70eec207cb96cd8c0d0b14d8e732184ecc711bb1fc392973ffff60006b1f7e369999eb195c398ea2487e5c1d0f1710ee70554c644566e2b969a2aa73e1e05519eb6e72cb6423b91e0178e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1afdcd23ba72bb3dee720657bb6ff925ee8492f8e58f00effe9dec807142e49a7c5c6c6374f2caf99f1355eea600ee7859d20f45448ec8cea0749c585acc058025463f3cafd5b65969628a52779c6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'head7bd914d8ba486ddb1c44911481e002a2bb3a111f62596a860d3fcc598dde64defa1532ef8ef1120cdc47be3c592284a2cbe76161605ebef68ffae0a89f8ba13ba1c3679ea3e54ac9d320fcd4c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha8a0a453513f627587836e0c6c47bbc35fb59deeebb57efd6d5441d23dbec987f3a6e6c7f8d3d8afc0a5f2b0d16ffcd1517dbcd3228219e0ce0e1c0f59827a289c75aa88388925ffb9a63e682df7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h40e16e7c5fe986bfdf96a3e4a3cfe22030e37d5c3a2fbe4ee8feb5710cce6280b1e6b7ae9c1e2c874da59cdcff5897a11ecb01df0d699a720523a04b64fd08d8ed60bbca50e21a5b34bab851c4c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dc7913699dd792268bfea11c4b124dfeff5320a49bd081defcf0cae746176357bb12069b036d7e1f44dc9b6172cda0603ec8dd82b7f141636162534f420e4220c0cfd5e14bbcdf9231564f9fdcdf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h67208b715351f95b0851d3036be23d318a71e9fe73b7374766faed7b094b724420d1142749d5223d7f21ac6854314702d4e608a9232f00d59b10f275f78a86557f8e174224d7779aad14ab94b088;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h139b5ce786a632f2556c9a4a6cd5ee69d13b752b555d8cddefc680657a395cb07a0169c9c76208f3f2b93d0b00f178148acdda32250b05c324bc346a21e34865bf33e2c918656c5a9efff73a8b151;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4ca7e37a2e7fff39f102075e4d5b5733f4c793f9634be91230529e7b8a40adca65d9bd8381928aceb9f3ac25baf456323aa2aa915b27041ef9ac93a5c2c113e23b1514c150d9bd19c63cc3a8880f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c643406905e626c0f87c8d5f6bcb8ffa1c5a230cf8119c5c1a7356adb1b3b5232ae19616d59b1359886c0cb5e98b3f7fdba27e5fa806039a3a9a756236e2569043f82bc3ca40b6ed3453b184821f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e17b5827831f63b0c45add0008875fb6422d17ddb6840205092a994a5c02a1159763e4d361be5259cfb1c122fe6bd925d5f4c71c788df15e1aa85fa21745a8e577fd31818aaa7fb717ffca555fbe;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16e4030ef883f078d7f46e5c7656abea28df04b44f9e8913a70165b50c8a79b280126b696eb0e9318a5c0bd9147f84e9ca211964f79ca9331e09f4508c0633ad46e1b0fc2d89829847074dd50e8e9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbd1cd28fe36deb79143110457ab23c3ad79000b5e3f6de233fbe381233613d29907a1af0bd7fb64c95e6ec649e7e0f5179e09cb89b3722e2537c831f79f6480395aec2fa16578a8e548f12ba7937;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha9b080bccc1fae2f8e2fb3e3c930087a27e9780c38a663a6f1fabb5cfa17b1021507f098e88c22fcf8171f0c25dd17d0199634fb7d0e46de439564ac882c2ab0d40d05811ce6b14b1cecd3f8b199;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1156d91047a6acf744b39b8c71aaea1f362ac06119a0f0f46e71c87690fbb7e2507ea087b9aabef822d77e53482e09e903c9c8c49dd72ebb72d94287e733c0e3cbae273e59efc543f4fe9713446b6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1779cfa4dbd9693f713b10ba7393f23026e41dd1611e195c5df3af2b1dd1646b8b1b36e030b4776e4fac5db047d068808a46c2f155919852f77e56746fdc3f3cc6e2147802d7a2c67f3d44f3b7d3e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h55f55d92a9969e3ebc1437fc528609b364dbd1b4f09a909d74dd2ae2675eb98c83dbf13e97c527e54d34fca8390d3311b9e325c771d3b3c0f3fe57443187ca804d5a4541dd0dc2927be035649f65;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd8e2eeaf87396cde14906d0f820ee2dd1fc86cad852c1249cb67503b54c44ac7aef7faa96d06d7e62dbf9415de9b2154fc0e4c27943e93079b73dac48e9d287ef1813e861d788158d7ad377d1d79;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d254f5e6902b70ca0ee263524c1cc57c440a1284a238709f0825f6ffc37780d7bbe9d0d97c27959aa18e4a74c428345286d6f22c91e79c8c31bd68fdb48b6aefb2191184008b43fba1e111b6a45b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf6819c79646c0a3cc80715ef79db88bf80135d5d648ddba47a318d09c205bf507f64a6484dacd91660aed40783a620e917911b8fa6c2284b0e17ec06ff9aa8c4d1678d3e96a7022ad9ecde4c05a4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15eaf45be47f134838ba606859916e26b71afd513a408f4c1375b5fac3d25c8c6328f6efc95385231efccec57940c0d0e2390110d73ac6d4cb24279aeaf8e65f4583d651b20b0ebf173a56efc934;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha97d730401e2b8e122c5d9ace972f53c1d6a6854d165f9601bac69a508d0a4ef4f58bd52b67c36a5ede12b598d9d68e9af53c462b694ebdc9822616673c98a1b501aef7126481ccca2f99c838841;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc77717f32ee26baa2960daa76a5da8e54380f71b2af634f117c7d5c5c69f049c73abe84a87c833c8735a96334031193bc7ab55b9c33d0ca77df14c87128b5fcd85a2020176e7b4e0fd72b087f213;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e30a320292420fa86670684867c280d6ae1bc714bbb2202b6c99df3f021811d6335747dae091809dfd4d9d3f48bebb084949d2887009d062f76c1539a6d958b338ee4e7b3e5c4e2857ef35ad6dba;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fbe36a4d2b1fcc98210fb4d0d38a3f4ec26662e9d8deb8654a974f02e5957e3f826bd3032983151ef163d57b83863eff9524724fda7962e7136219951d57d2e0c19e96245f6572f0fbb9b4cab33f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5b754b58540ff3c67e61a75e1b14b4f6ec062fccdeefb24434a2b870385e907e257ec09c9229f813adcb0e8e1d62b489da7669d960cb4a549bdbeb213492d87f66c735cc24428250a5e95a596900;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2d8461d50481c8902aa1bc5bc74247792adf07c9babb45d60597ee349e466387f16d9b637f57bba317f7120ad0d37d41e533f981cc56432bb8e0c2cebd6b78912bd907308f497e496209a2a03275;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hed324c3f61a399cd7dd08d5287b7a5b36e9e387fe5e3593353c4ec4b85575761a82310a5134a12df27b7cfbe5d7c3016c0a03afa84d936bd5ffc67b52a5324a919679902ceb7e842ddaf591c8970;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ed78e87a0d9ea914ac4cfe1995ec0746124a5f24f9b95ea62a0371627f20e490ad30a080312fb939a028c3aa417ce76d1cfdd10c3506ba6089d98cf7e052d38cc00efe3009055a4a117009083fbc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hda818707b5782f8f6324fcb0a5f4be45966c96398991457628792507f5a1d920490c4fa1ea5460477f1271f58d6f597dda9ac788fdba529ef3e161790a697d95dc67a8c61725fa99ffcf816eecc6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3cfdd69d2d575c01211a038c04375a2d589fa7ae4c2bc9f2a41ce9c1737dd6ddb23bc3a661c08eacbedb5c7f220f5d2286259ec72f48ee693934396c4bfb0eb4ddfe197bc48e2429bfd82da065d2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10526cdc10c68a6b321b04275a22fcde028ec3ae767d42c4ecb39b95e3d6f324533aa0158203a81abf2e8a685cfeb22df3348d02547085bfec830d9c091862555cc980e0f03179df8a8344dbaf957;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcce73316539171feb0189d0bfc7911ce78a60f9c1408d7453e1e4d007038f8e19ff427615247f1d3ab3f8c367a24ca84849c6bc691617f2fa12b02edd77bd281583e5305358c2b11ff7f5a04faa3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1894ceba36dffbae4088d011e78ecce077deade99f7193eccc8c0367fc3da465c63d533f75f1a33a6c3f4c5da62eae4d8f109e9c0060225d0044efef47f026317d9a510464882e0321fa9d8506f20;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb95b67ab638196a5d2654b02261c9ac8128894edcfbe75ee09a10b50b8362bba51ce4742abd087496c49a91f9efc7d4977baee2345650fd06c7492aa8d7dd5953055d3a2e98a24032a91c6809c7f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha96e9ef96bd8a25ed906934bad8351617aed14a3264db89f4b14308bec786cd9689de140bc968d9d20ca3c5416b7d1070e805c6dbc0f4e3006f388445812ff951df6cee0bd799a2c88bdf7a739a5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc2cdc2f6c999b6cba9fa858a50a560574bbd4aea01efc29dd258a1a139dcaaea598bcaa366ce793d62de6952c355d7f1f6851fcf5486dcef3af12e2a4f630db6f6d5b2c788cab8ad2b4c03f59a2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13641436f3cb957418f16d778d373b755ffa6eea271693089b081563eadca9dd9ff86f4e2d94a86fcf1c96493482570530e2a0cdfd4136a87ac9e9590242967f877256d033ace4ec53d05b55e3033;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1562d6b189018e8f6ae4223b0564c1f79d4359028213a01acc33dfc89b08598509935471369165e6951a9a3c78438b27c48b787eb170558c81edc9a6127136921f7a38c82f585184529e972f26cbe;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he45da339b633afbb12a690b4c9c01ef86418998ab7a5070d529aecd944be5f4ad267a39de372376318df84cd1070354951ff1bf8826195fb4141fb6ed6d45af4ca3ea90b55db6faf0b5bc87e5960;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h83b2561e17266d7b3d44124d867265ee3e55261c64aeff219e7fdb2f4f8bdcb29471708ebb2d841191003e7bebe98f5cbec6ccac0ca1ffdcccbfeb8c2f3e06307f63faf49ed9f9b48be5c358f279;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha6fe2de2b4a1d496f7d4609a919b4fc3f9fe775c1fd55273fd2cb0b15c044de8eece5648f54e1aa7aeb5ad8bab82c4472066de9c4b3717cc11f555e79c6811f6e6df39be813f49bcc8cc235c99f9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1607d31a0e4c0de00e93dee47f5d095804ee00aa7f1a536d21b82896c6a0e10549cead2fc4a7e7656bd9d2090f155c515a827fc960637e1a1e23c0cc5136c67e07da229cbaf7d554c618dedcbf66b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d8826326b8c360edbd6f9d8fb7c7e5a0a3bd068b5fd5609a011a859172500dddb0c3060a1ade5ac943cfa9e9014014effd592d7e31bc0340a3341f181543eb8d49bd5913e4434c8d44f82ca6289a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19fa52afaea8d103b99353a67ee88558818c4fe4b07ee07b53be4fc312384118b26c7d0d7d892bee75e891303229518c456aab5e163a1b15b446bb10db48cf61d9f01d94b427fd164e908186d3821;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17b5e70b05c1b1227fcea72ef097bfb372ef85cac2048f1a69c86694e12dd12d56e01a17e0ac2903ba7d77d90bb606fe9a4af5e1716a629c42243d2048b1971b5d55b42e3c3dbe5997680f9487bd9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdf95d40014cda02c377cebbb150cc7b8537ef771e949cba6bf2d7fb6dcd077b8537f05e9715c5999a84144648bf0b7a20cee0ae8e4b3728b051b40fc7fd8df7ebed25ab0fb4ea9b2f3e27d3aa2b9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcc3fca0c81562b532622309f78087704890c1c743f99db59e7cba6b0489dfb546a5c7208dbcfc4216086bc41bcbed1b562945412e1b4648b4c704ab8753f880863e05af8d35caeb333c22226628b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h61a2056c390d5b1c33479614c9730c2595433231b0a2c236b76b6ff3db6d10991b9bd872d3f0265b1ab67c70c8ff71ca83482a5a8002821943097156852aeca0ca9220a3dcf54347c80f7bd74fb5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e40f05794b03cd2c24f8c5897d814b28ae6ac6b069002853409106404d9135d58061c170e6c70cc1c8bf45b6b7b99fcd70985ddfcd0c48d8c1a351ddcbf402a06c4f3c57d9ad98a3d0c1c2eebdc4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2c54785217bad05d12f0c3d56e986050d783e764e5e7558f5c63f5a7561b9fdf846aaf3300fbcf0a514f3e5ffa7adc59dc2d849e47430d1d106c1d10b0cc5a01c5330059702e7b729d04cc5d0847;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h128e093fec6fecefa5b7da1d31db25bb7a2b614fa7f510860511681026d9a123177013605c9a5a45895c39cc6d46acc4e22a5cf8140a3d8f390d518401fa62ebcb3d42cdfca90c0acd1efb4beddd2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h85f282139fc9210acab6adaaab6b923cede9c69c8bc39e0d9d50d958be96ec5a9907e0cea0d35daab3d224b8655ea00ec927446b6868df1df3fa01f9f256da438133a9ad5ec3664f6797cfcd4c23;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fd5313edd247e6c73f694d8bfff7bb2ff5ba33a447f253483e91ee4532976236a6f8004c6720e3ee1ab91e6ba8f26aecf40e9f23b4aa1875f3b5a236e25c0eaecddecd09af7dadd992a46fc292b5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h31f39431e6c3c1aa424f6104ab8a835bc77c617d4688d094064bb8f4b9a04e56bc916fff8d414d40da39361b69cef3a591fef22ff70eb75b87fa1be04655ef9e1cabe0c8e9463f1022ee0adad440;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cae0e3463fb38b82849407833fdc6ea3bdaf19a81bfcf3d91e12bb5e61a6b282a3e48c629963e322cc37c44f6329a9df71ce00f70af0d1bde249b579d5604bebe3c7fc9c97c801bb4d64d26e3b01;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf55ef923b942607c08f30e78f2dad986752e6d2acc6fb5a81b47e4909b8a2c823faf374240d00db7d882e094072bd26cb1e7dc26584db6b4e2e20c46952e5e859d92fc7be7267e0596ae62d2dde3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c9756c96a39c28891331b93f8563d557c541c1855d1eb2d02764a5c8ca266d4bc5d73e47de01c32fcabf35e1f8f5daa98bd3da5a6915430122e9dee6c625e9db4cab43f6b5950a14e170e21c1afd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e0ba9c026043fcf91e1947871f372aab22a7b74f9a785577ff63cb0aed823f7cb40f158ec55a7243f05f3398345f7b3f1a0455b61c6a0bdb1d29de8989ceddff330d23e21ed8657e0e1000c09d24;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb7f42c6a99defc4a12ae7b3a44309f38f8cdb5e2d1533546653d78d8367a1da77693afff7b77d41b03e02725163205f730bbde5759913b8ca4edf75421a44641aa8932cb584ffb9ee62a1c8d50b4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1baee0e7913c21f1c4f191f12de659675d54662e3a5fcd379ee7b6fc8f2b2d77ca59029250f9d71a5a1f653f8b5b1432ad5669d088a0c2a4a7c6c70c2c97b58dc8438b23b5995e8f5b09526e5cb5b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cfcb406a765d31ff2db94e997a14c31e71f943da685fc7ea9a77053e3ea7b99b1dcf9486b70ea038eda09689aaf7f5f415767d2849b1173a8ad195eabb56fd5600b7d843d9d3470406fb150b15a9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17670fcbd3cb9c67c6e1c933b0914f122eaf144932596606039fbf251a13b94982a2b57a9055d7ae2744be0dbee6e6f26a181a8702cc70462952cf58154b592f3891d1167c266824752889f90c1da;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c17d681b5e9a44d3ea0c67a58bb16957d5d539bec6003eaba1a9472d4b283aa7cb9464d9eca60e3fe6af72a18d1e36c6f32a810db29ff5aa1bcfdb2369d5124053e2f241aeedaf032f55f0ace85d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfba6e9fadc610e5e0315343f1492eb4548976be75cdf92733316d871e4e53f1369ac397a4f24afa55a46c413426fbe5942751541e07e60cd4dabf18bf2ea9f259301355df2076113edc4d96ff9be;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h187ca025cf02496970be51001a11fe418bc8e6ba4fbfca3612a7348eca5778d250b12990616b2f78f87d8834fc0104bc4facc336943a5e3a401e803c3dfcc33ca27d1511274c612c7fcd2008b9d9e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h166cc1a2d34ffc112303bfc0f8b9e561eba5c0daed4a507f02fe6434f6ab1b36d59c6342407813b1696a2ff5fece76da2021ffcae62bdb3cd2be167d20dde1eb1a7b6f1dbdaf308fbb21ff29637a9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha75fb5550012ff2b5b2129e8f3baef800b7f9c5facc4c16f03be3a74832de4fe99533bf6601d35aa7f2eec37258f45f7e15626ea6f1bdcdc73bcbdc0cef17c6c2c6062e68f1b133da5c3f15a212f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha3dd22c4b146ee698ee2e3ee8f2e30ce8f60225dcd47321b79bca1c22aeaa98b535bf245804c7709752101cd6dde95479c1a84d3e60d2d0a52c2660bd4de000052c95120bab83593751341f2b072;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h408c1addf0aecd51e947d361652ec597435120d2da2b938c3e598fb74898c511ca8d9dccdfdcd591343b076709b117bab17da873c9ef1bfb8ffd00cc7e1ada5e0bae22dbd3f8cb8fe020eb7625cf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7fed00920a2f3174f3b2409442e696b6e12dfe353c0bcf5480aad53b464f88a9f6f87c44e18540a3788f08ade18669e5e9ad978871bda898d94ba7bfd2553cd86c661c197842c43b9821840b2b57;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h173ab30903438441c53c4bd8b88d42de6b2e737fd706945b487f6f2ea131c5893ce9d52aabb70cc1c14261b2e2605631a03126ee09cdee67b487e5bff72ebaf6ac51b15e114cbf8416f0f7c130486;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfbff66029bb3f6e52ad967524efac788d8fa935aea7638677fa2eb23bdbd82aa60aa5979033152588eadd1de01328a2552bdfee5da91314a8974223c330962d308f7f0abc15b8b0d2c45b275f731;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eb15bbefda733540766388a90e43e900370e051aa4e1ab24417e5998e8df96a75df4ff54eb8f056b6c1627bd5ae2305df4344976016c9c8bfca2e0aa253d8ad57b6b524fec88aa0b697ab03ea066;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f9a4b95c91d99f7a5703e5db56910cfc7855595994a01344507319cb5d117b4ac9b31bead76d8a8e468ec3394d7000bf4ccbe8344beb469becbb44a6f3271f538fd303c15d677e76b5e0f9898a4f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha9d4cbe7b1a75f64ccdc6de0c5ba4e801094d5685238f773d419bec18b58687e1c329eca4cce281a87e38e627f6bf8c6726c048fcb581f7bb2f755e3a31b8c3a79afac7da7fd54f0ff142a4192be;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h110f513ad1cae0f0c59e61a0fb3a93e666c665e95d18e3ec3921fe24c891d60b9e281634d90c7e7f1c8915819031b9f5554f162e36ca3ed4ecf4e25edb414b18e95c2f3f1499eb74834d6ce8afa5a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19b7823b419dfb85ace1f65ea92c1bf86007023c95e94fc39466d3b7ccb50c8ada5a05fd208237f184e0098159c09b1f6e128ab8300ab88cd3d99cfe90ecbb1a0b93fceabfe0cd114b29e61cca8e0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he387ccc861698b714d9b43f01c504903f26ca941e2be21bb0c0827dd9fe3c97ee446019972414ff8b9df76bf66137a9e61f6e4811a540613996c817f84454cf3344843ccf8f98ef3dfd9f4b624d9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17a8af5cc3a90c5262a5efb1a1f21e35e9f5f6865daea75a770440b0824a31d3033c2c8cbe8ba2c70c2dfdb1dc9ec1ddc75536d0da35ee019c3bf0b2ff132541aca192e6cc57eb2c24b574d0a45b3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19c8f13fdf55f6ea2b057005dd12e20a28b34fd0ad3f2dfe0f93a6d4a5fa6f90bbdc95a60c02ea519aa928b30b4240d1739f5a0c99b74e7aa43ec686c7b7e1501c9799094b213a449fd2b579b6185;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b1904ef2df033cc4bc9fe47dd713f64bf7528e6a6d329c35b2f3c368ee3c161fde6e888f2f86b4924fb217d031bd23c2aabea49dcafd70491d485a10a3d4fb75ce0b647f26eb78deb51c2258b25;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10df13b74ad653c3e7d55282973b6463fec7f8ce540d0f9d20b5a6c0842543ac316680883db23fe97d61b9c6c5b79bc7b2bbd0914db125f87d9ffd50d1258e9bed4fca35b8724128646b0ed084e5b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ebc082f359f9a7dccfc52f717c8b00be5a860cd3ad5371777b9f400b000860da13bba891a4e93125c83615e885e2828b3087c219d1554b80a84142b7f7fb392d60ff830a374382ab385b167742ed;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5e981e130021a1f4c6b6acebb0e42f8b79b3591615fba2ea90f9880a4208e79022b9103c4c4cbd3fc8fd1ce5a0e030c876f556c753f4715ef22be36eae3dc68d76061948e1ed9a64ef4cd93c61dc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18c73d027cf7f611da228ffb137c6d23c3f27fbe6976855b2af0ea5acca6809d4aee979ffd8a84056c5b015b781586e8f6298154dd2f31b166bb452a8f01617d51983bbbba330b2b3313b25cf39ce;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h480819bc675481f173408d5034e2d4be5d17f349441b056acafed242036a7999924a9d72396dd3a50f1a5dea52c4c9e5743824488bedd8211b2aa034230139e61d26ebd56f39e65aed0ad70a3104;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc7cddb2d1ef9cbc3042d1340ff684b3453b39352b190b7cca36355423c04e975bf09c9f035dd478d55e60d43f059d4012904c3d2e4dce42ab53694a100b3cb28566d25bf9dc50c3dc11ac82bccaf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6a31e161dfd3b39fac2883bbab1cfff1147e96c300c05b92d45a7a090aba27461a29b3173a9bb084f4dac336e8cc8c820613c7532732ed7f89b7a15b9743e1daac8b2e91025422d94ef435068807;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1443dc42da19e092cdc8aa669f6eaee27d2a756d2639aa7ae4d25f285b969adf081e8e1d19a9fe7c3090aa7f514577a44b8aa9b0f5831a1d4ba631ab038f881c15c0238f2902022036aa05c014163;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17158584c31b70792b6238b27defe2f81a18822f93d56b8865d074c9e85ad0f7f69630d66dac6efa6db797bec4030ade79b05aad123040faf41a61422ea99696d0e04e870a805fb5b67d4e371852e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a38b88a23e4f1f6503f4981a328f9c48342d06218f96e86acc5c7cd3dac1a55560454fef93940ab76142cf50292feb181654129b74fd967afa47c63666c3c9c709e3f4157f4aba252741aedd1f51;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h313345c48842aa7079cc7a45547142a01124ea14c92c9f8eca4291702d863a2e85e22e5e4daa8e6fa1fc31ab487f0abe3e7749aa53bbb0bbc2dae98dd619be840de97e6d2592fe0f9eb8b2f7ecae;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9ac82cf8c297df0e0def589cc1534c0f970ebd8a45a914fa2adcf8479d7fdb530137df21b4cc90573df1ab51ac8d1b6d46e1736324efae84c70ff1ef6f872181b5a117147f989c69fee069932637;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ce4f7dc6de591393542179cf788a0c324da8786ab18de22fc208bd86ab55634e2323cc7fe13ab50e0a9e3a2075abf5c51692182c3039b0d4fcfb4157d72efafaf3039347f75630844ebe37254fcc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d69628c83f685ec7171cac0f97e7009d7cde897545c241c153858ef08f6855b224e7a1ca1ef61368cfdb1e588c440c1075fcf1ec4e9e10cbc2c3edec6a84034efb32db7b9d7535f784dbe82b3c67;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c101e9189121977163c4f3ea39253343b789691553d5f4387a419cbe76b7b2b0621fbd0399473da2a7b5ed957030ab357897615f6ea40d9bc5c6dd16a79eb672913c5a65d5ab73abf4407f637964;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e7ee3bf7c870fbf7087d56aeafac3fe4e755124def9643bd503bb8c3fa7644f3e38e10b3e765bb268a5d783a75e5aedac189489e2f3672fd1c89360b9b436d1c8f8c51a1c21b12e75e856bce03bb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5af9499f92d68f7073cd78bf4333f1916573e9f82aaff9fadbbc940cf0e3e9c39b76b6e70ffe39cc1a8624256adc56910627f55d74389e72dded3425ba40d2a38ef562d8be82f8b500ec825f7d7b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1232282fa88679e1836bfe8bbe5a16b6fc8369fa8c0f7f3a7c75a6fcd523a72e2a10ddb8568960f06a9e1a07c9cf3241158a3131038531efbac7fe380e261fad7f38298855740e7561fda75a6f7d4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h340e30398f85b3158756b7a8790c3075208fb672f3c433e74aec643a072dcb9aa25a72fb0d3f227875792636e704a3513b08b5f7b4c70c1bd3833bede435a80454f383c9163658d20dfd8592d9d4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h42609224f2fa32bf0dae1b8e3be55ed5c24383a86b6c6909696f8e7b09662cc8585ba918422e77884ead10d31084b64bd008f905b3ae9d0038fc37aab941cdac0af06c223737c301cedadf861afd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12b63bf586c4811b2a0628899e92c231bac54837d49757fec1df9527f03a24321dd63ca66b43c0d6cfe16f6c7ec3281f1110f2eeb9a505b382059966e5f9f36941f8bb902fc60f44fb6a6eaa78334;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h179a34e324f579039b268e0dbe6b15e28b4d7ebf22de244e2de8d232ecff8b4cff2f66235d9155288a2c15f4bb8d4cb80ff8bc89b03c8332809bbafb3a2a669f4178cb59f44d3c91009fa5f491245;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e9a18b174093d26a5daaec6aadc5ce2d9e633943180b85e5a5f44ab7a76ebc060381f303e19c4f9716a1ba7057172dfaecb5bd016258724022b8830e5bc03225d438f77f8055d7d1af7a8b3b948b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9a350b19415f3cec72497a7f160563e2d7872c3facb9b22b120227f2074fcdd47951be75dc1da5fe250df9d3aea40bb84d2fc4b60cf5ca3844801a616cace4cd61ce55c0babb56b63b6069b33876;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f45624d1684bace0317c99ec387f14a6ec3384f7339c4a6fcddb2208d05424b7fa903071896dfd1d8ca23902b2d89f28ffee197bc4e5dc4f7338720c99d23ee016d11510a70c995cccdfa514725;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e95685086d555ab9275e48db0199e51723e143f8cd1ffc86d41441177668544a5370358e9b132496ef3e4bae9e3fdc653054cc2e3643fd3953c265f6a8142a50ac80a426157f2706eb34bc6aab6d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h102cd3593a9af0155fa3b1d7c3372069c33181ee688ae63999b6c9d99eaab7161810075590edc1f439ab6db4cd5963226368d144a7c68f3497fd586b014211b8fd10fd2d64f9058312fa969f2e938;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1046029017d92dcf4707e9668c87258b606212e094ed01dbf837dc29f1ae864560840a2f8706a1ed08ed298aa6ce7bd3a8487aee542bbb299b0b9b7609b56f25008d25910f5c6ee3ed28ce974ec0c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h176f5056626d4cdcaa872b9d04f04fd6df54cb3b9d4af9ccd6ca5740e2767c6854da62200d0763634842c3990eb7e2ea3950910d700358558f66aba6938ba7e41634d46b7182ef8e62bf34079a358;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f4a8f0ff9aaa203437bd6abbc064c11fc4c711c7d56869b384ecaff4704f9e20f9609537606e02b7de25584a292f1c1ac37a84da4b96b914dff488a959693d041c933291d5fec2c94899ee9533ce;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10b7bdf15328077a906104f090e464089aa6c3fc93a6c5d5d7164427c96cc269c5496e94387f70d96260f34f8a8cfbaece2072391ed06cd7c713c90d596e10937595ae54d76c07164709db8d64cfd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17293b2b040867a22678ed4acb5bd1858243a7f8126615526aa3299b301e8b400b0e675df4a32e271563d07445cdd6d6f09edf37804245e21f0b5316258ed70413485b705bc2ebdccac8f932a25a8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdde2120048b9db491a3f965555a90f033f76b17c7d90571d53596f5e266bc029ac357c5c709f8b80354d18c4840aa14159206d3759d3328b163396d0769b619c9743bf0409bbb63004b1c5623e08;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11ab995e4490406ce48aaaa798c2f0aa80746d5fc5cfea75c4b588b289c9ec3aedf39facac6171b12a30cf67e68afb8f8cc4a771bf284574f7e1fc501dd63a9ef6ad5a7c4aa11314183b97d8abff7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h28d913903631a4b378e44cf14e92c5009d53046fd18e72c0eae92f9b4d564144db9780fcf00065bd4a985dc7e0f96ad8f0e595ca32ea687094e64190b2a3e066c4f10a642290bcbb57c705870885;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11eebaa627255059a6d84a78229df3d0ab0efd4a661486cc9c56d30c6076484196275725a68d5d61b916500edf4f3d9202afeae704a7e522f179d9bc097b5040196442a3df7ef44c8102fdc8fe0b6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'had524106483cd5a00e91248fb460119c7dd88394ecb0215f9571e8a935c30cf398a287aac1b110bf7440b603511f8d6f5870e20a39d381a04af4c67174df6c3816294ac544de5dbd8df535476042;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13ebb3329bd55fc0662991a74d7d53185da1ea0284d57ba063a6679979456c7e18c641f9b166a6f7794f6ff4473bf7ce975e0e1f182f7a464c5fadf6de35c75d333f4f2f3bb8f2219deab99942a77;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12151a74065a3007264d6b8f9ac2420ee8a37ef3610eefaa7408cb09bb953e690394b7f57cd907fa2ba704a8fb63b5a5af6bbe098f14d98068be8110cb9cb03f44bfae010dbf93d3ab91bdcaeebe0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h135a9cc32ab5d95eff45495f75c02582922fce6cb07fd9ddb3bc0a8dbe0cc0eb2f6a5732b8880ed57df967202e16fd904142d146a7a9d64b07280967af8589a40453ec67c5edc4730f897dcff3e5e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1590e15c236f7b7090be8ef6173d539d6e87b5facf3ac1896a856afef1f1ea578ca3d37da1216c6c02e252db6c66c55385dc00d31c3fcca4fd0fcef0ea58e2c675d3027096e647f3eb0ec9865397d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h458f831b77e3b41cbdca31bc514d911c492269be5425b86cf5416abf650febf6b914b2b73d0418b1e8299987a6315f45dc819c804f5fee5f72f3f14838649dfd62a078ffbd5e876576734f36fc23;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bebc737c0454caaf6c45d393bb7f0f8a15c6dddd62fadfef174c43d3b90380660d4217c425e6b95e9f49fdb5773147d4be10a369149c1af72bf766b8aa71ce22b89ab95b02f510d4a755b45be606;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13924b270483e26d079c350d14ea257195c2b42b985e1bac1f39d2fdc71e6daf32ae534bb6a440a9b87ca3e300592c9500cc0fa99146bd729e68ebf2e9f8cd4f386f336dfa44bc2982e1ef62627ea;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12ad6b18cc272178738db0c76de7da51b7d225ddc8d78cd4da39df6d56567169f31463a42e4b9aac9b21f4cbb7c9d5eec441b08c61c594ce562567bcbf6ada5a92e9f93867f9e6fc2a1233edb235f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1449f694d0b5e61371022e0b8aed2ff9a0175d21aaae9fa18932c6a7f3c6d71097c616d1f599318170d765d6dbb3df4372560c31410e7b7dddf10c3f8ac1d934c2cd9b659333afa9736315d58d3d1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf35f73a34f8cb833e1f9b130c4c890dd3202e91acea1c8e028082cd8b7c14915e5b201119fb04c823bdeccca74a65c9e65d9021fe3918e8661e03982709f60e5edbaa7e331b14bc355b20a378ab2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4ca2386e82fb5ef88adb3bf20fb9c28424e15c578b315b4461b66c869d019b6d857a484d28f21da76c11f0fb5f0c3e202d0710b4b206bd88a52779051d2e2cef0bf763ca664247d8eecf0244f8f7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11541637f1c715e2247da05823cd8e9fbd17ffc183c0f189de2e48567bc3219240ea62319892a24b82c1a459217c18486b5a30e35335bf4690aa3b1bf87c1201220a302b1fb3ff46c3740c583713e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h125f40ae9858060125e43fbbdf5c4e83cf32b7a8faedc775d8132b80c1dfa23dd8d756d822d64596f1ca29bb6c07f50f27882e433c51cadb6407211d70ddc49e61b470dea4fd0a910ca1b7b5aa142;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcbf25795ca4dc4e880c9ab81ed1a7316cb0581f5be089c87e005e9ce9211cc716db662fcaa08874990afb8cbe4f5e5d1450f8a095fdbb06f0d52434f69c1d8c05d3eefb6c6ee63705884666e21b4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1116d178c31cb8c5d7bda8e1604dd50a9f61d9e415d5efbfad709314384a0a9fc9ee41b02d09802bb5096c719b28f75eebca6d73a74f9d5cce0cb4dc4ad5b2e082f17ff3885529716e34f8f7cf973;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14374e742ce958bd8d647b1fca25bd0e8b90ca3b65c488b2170aef4ce8b1d66a695e71b43031ac69917e4f67bdfdbb0df35f2c74ca728adec51960d704438a0abb6ca142dba476290d165cfc72730;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f6e31a5ed635ab6983afa460f8666a68bcdc7f3e89060e23f2b7cae3cb9d071d6967815e63f3f710e06b014a90936a7fc9ab7ae0dd08f659ab07d0f6f066ee3914cbad28448322ba71330318891c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h78ec844326e7d7a85c61bfe3c393c212594be211670dbc1a08891981d89b906449b03f0d0f1384ccfe22cd27dc3e0d34294ac728580d5e0000c70956e82b2b593d5e0580fe01e5d5a46e3c1550f3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18da69c6f4c8321428ff270ae7c03c71f628f0c5c4aea61dc1b743b1dc0f792e359e929fa029ccada92e1a6bb0a16563883c69eece7f7b1eb0fc3624a92e80fe1d57d61b98b432353858ebd25ccdb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14828fff1c3664c9f865b3a0d691cc36bde5c87d7eb28d9e20dce323a3113d299d85265bf4e3de14f31e8f9e614adf01f715de257c902992dece5cfafdd1ffd734697126309681db4b458274d6978;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h183aba6f4d0d920d42c28cbf4e8795602893c930551cb80c1ffd03620664b6536669f703f72c617b5e1ffc2beb800185a405fd96399af7681dc26eab633a8db6e0ed4b1f47f3fee497c0ea6af1914;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he8409bc7d86039336ad6929c8abcc80dea63c268a5447d0a8db30fd31b1ad048e740d46b1c98639505df0613ce7bd224080c5feec19d778ee8606b35bdf23aaed1cb06f19bf087e2bbb424976eed;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha7f4803849e464f0f9ee9b976dff07b06536e2a9b88165cf257923278b742222b93512ae6e8391f8ede715e8cdea455f4c64944ef2ef9a0031af5030b0f243674500133c05911446b96e6e25c859;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h145e5b1f35e189e7b5dde0dab096da11b8eece3d9d133b2ac6993784971edf101a3cc5a78b7e9ebe83c33f11f1c477565e0284f8d7874c0f2751b8cb66e011f08ddc27731f13717f3f8b1c8df1513;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a6eeb7d06feeafdb64bd6975cd6f90cf2635e00b0ee1ef38b7c82e0ff5af68d9e66af2799f3a40694057f117c055f6b56631a3087746d6beb8cb71e2f222957447e6c2e0b8e837a63f80a88cf5ab;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3bc62753ea6e716fde59f4f2227ad810cbb26396e8120f4f063a7157c08b0f4c69bf4273919288c7a24bc090d8ffcd9b2bf163bf5d23480587b63b31bdd8fee9b1faa5eeba3ed4581cabfeb390e8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd7a62ed38a4c49996b3d043efc2b120ddd93f0cda5a7aa06d93f05627dc588b57358c8452f350b77608416e5f742dcf4ebb2d6d36bc7838e53f5a79d0ab9953f7a02b8b7b7aee76949cd24667564;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h67ffe45db07bdbbfdeb502c1f470ccc74c52059083aeea43d9a7df9996cbd3b98726cc370aa543372eeada1d76b2e89cc35782db3e355c5f6db6379ca0c4b404622e77df49f4fece7861ad487d2d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h49f619b861209eff1f03011ab55e0aed25d738cda85bef6fa1f9e381faa5a3ee058ad80121e2216e818fb04b37a6be832d0a39aa91de51cab1edfc7c37d627591bc401423dddce31359bdf620984;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h26fc97a67f87902f0a3d56bec7454cfc661a5cdb49577282b0b6a28ad8155a01f5bca1fbaa916dca000522ac5c8af650ee12053e6bdfb6f195e917a22603e62669a6f2b55b6b2658eb7590529cdb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h500c77c30cac338336c21d5feaa98e4ff8c073c7192e51923c4d47d2ae1ded0dcbd4bccd2c6e97ba97f70957c52cadaf6bf0a5e64d5660e22b2d48e4c7a5b9ece3324c9c84cbe5cdaa054d6143b7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19e75cb61fd37074ecae1199d3dd3be8150271a2011829df5247ec8d56bfdb09db4bb81689b45ee132a7bb4fcf2f077fe5ed5749e6f06f8af3d76505c4fee6f2e6fc72949cf1551fb289932bf9e97;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11bc649e3b09cb2c4778a1545e6de93550d547c85455b75ca9cffbbf954959951a3038c7ca0e27d57a155867ae9f974e8341a5097c8b739dab00b8c70384916992c1d1af849b53bc8461814b10687;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hffb64e8fdf62f91ce0b7b4204c9b52a396845120995b66bb1a8225dc630ed752c35b2c588362855e2393c5e5a5beebd33b7be18ef785a2a3f6c9fa78f3cfa7a8f24716b37b73262077dbb2bdf6a6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb5060fca7a55a897e52fb2172c8099f44498f18050881478435b686c80b7904b27e9587defe226eb3bbaf7ae9723359376fd1c8e7a4cd08dff0558fee84d8aa8022d45d8778d6830d9c811d67153;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14f29931a3a1b936781d68cf7b3f4e1c73a3d894d2ba12720fc2b69fff4d1601ebb2ce35477d22fdd8ce94cb2c0c3cd7fce58178df9b6f18665dfcc4bd3da0d005b87d95316ca8d390ffc6fd3f2ec;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ea9bb76f916d9cd20347fecf637a79b340931df64c5deeb043d12b24e50514f3d567fa9cad417d5bea535d789a189e033683d6b706c13376faf7d08fc368b3632b77eaaaa4bb316d6d5035123ab6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hae3254b0f73b4ac69a82ba6bbb8b085a46750dbc296853c65d40232dbd97b37ea47645c9b0f06b66887b261b0e34a0715f80d79c2e26e98d6dcead15cb0d12bcf19b6d38c5e51125d0b54d77b69;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18f14d53717a655512596cb428932421957079b2a67dd5a24f2dec6bb5eacbd4c1beb383dc2b1f1f16cbcc6cc63e2a65dcb1c2e20ac05e5c75c52989c33c2c4739329a3d3f31dcee14f54171439e3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h217d4ab65995cfd3b577c53ebe3555e24629d96260ec9ec4bdcd844d02c2f539f3b6d3d857eadbe3e541473d9a36b16d04d58993f00588412a922ce3a4a13c082a78eb0becff1d4d6bef30610f78;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2bf8cfab7d04eac03955d99715d490d36f1ed6335e8e5d2cb81a9a38d96f8b4fba10e0463152bb406b9ebef266bffd784ba799b1ab0e9a2b7dc21cd0d7c2a1f1d802f88443f23a5e55e8f9c97998;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7efde6db70137e948bf21638e888d7eee01af98d47277825bbd6b76447a4c7faeb64720c8fd807f86217007ccb9a8055aed2a398a158481c3e49c17a6291745d9c06be30e248a1ab8c0ed737f113;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b95dd5ec4b4178939b5a27bafaf82da09aae705b673c48a7a8d497ba6ba47b47d057b78162e01be826b1922a9b45665da89e88f947115a89832b80e563029b039164c256d1003f451f9f636b2f3e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f00793f2230ff54889c01cdd3d47c33e6e79d6b5f338c292bdf28b02558a6ed0c69851f6c1bdcd613f7b021a926647e33b9f1b4caf85c42f470c8fd9ce603bca184cb6964a2f8b7df2cb42fa9e96;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f110a8cde8505b9b21aca09f4179e11ad99ffc5852b84d16d4fd1e3647741413aa5c498ce03d6e2d0a1b81f8f46542a6190a3e8b155929359e5111ecf61dd31eb2f1a15785bb1e36b7c77c9e24b8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2d646af384cdddd69bcdc823198f09c8aa961e9e991550e10d9f1cd56e837a7c3ed22b8f0799c9addd6a2c46e1256477b958fc13c22ab8b9c91dd8fe1d7d0e5b2f66e5918d33ac503e725b04065;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h67908dfb8b54a3d01bf03fab83d823228fec312a27fc9cd3815cc151d5863908e051cdc65b55f646e7a18390690b604e8b76aac0d09e12d6dbd1b368c93275a8afaf9a51dc2e54ef0d1f7ec926b2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h141a8c0df543382de85427a61b0b3294a388edeba4694ec9f751bab1ff915598679058818ce47f8cfaf3248e34f7e61ace88aee412c195e6faee372cec705e658ba340f4791c9c2002be34472d0d4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h22eb323091d82cf1060593d9827f4fb2d9b83268010d2b526205af2c1b703c2c9b29d26a8b7d0867f2c4cb951e881f527905f92bde8ef2b1ce52e3ad69dc9a2c6615ab18a19e1f76661b3d9c509f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1760836d599a0a2a1719408277abb364411aa694fbe3e7305b9e7dfac83f949e107e5b91abb36145fc82682dfb6d49aa8a41160f9f0611141e2e4f77590261ee6cd81b8deb7b6b4f1f2eebd150f7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4f27903fb0e08e0b1eae330237d47135eca9916a10fcb9dc033276f6a97bea2c73b355537c67101db1cd09018d570a8249fcbfe8750d371e8dc954374a1e9277891940cee95b2f2b8ec294bc21d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb64656ec9e2967a84ce00dcaa55d5970f9e0c3086c6b6eea630f74da464d7a45232889c881589487e8ef9391e13bb41f42ed15d42dec4c431e1dfc39dab4d3388755f5184cb9fa0a715e74573196;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbf911c83137fc990779a08f2cfe894bd9c630b5d9b274ccff9eecfbfc9c6e8c535b613706811376f4f7a5f4908b7cb465f55396c8404f119113a50505989b128079354a747ae9ad2801b49cbde5e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h323fb09aff3afa2277cba2abc2adc9427d28d74ce0689ce2d54fb4d0c2adb16a5972fbe4c83e06f758f777d7c590b5b35650525121e21c523d32d8c9cc8a42935583c552842e1b3783a941f17a7b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h623964fd31055ef7b788824de02695ab0c606d551c82baf83fd985de05412c8d8e038c7363ae13967abb020fd2a1abcb495d6706ebd6e78be8291b3c19e3233e1668ed79404362ac1c8277b1219c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h27e67095eff17e0bcdf56d38eaed7b04344a98c7840d01ab059424b56011b27a6a8a496a6fcc24ca42dc70aadb309ba4273d2bafb3893059d0d77d53a05e0dc3ec4091b25b2e29a8a412240f0d4f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2cb57bd0a4044bc378f6bb6006fba0be46cf5365c57d81348b5b33797119f0d535e7643a5375a280ce631deb267c2fe0a13d178ea5f6c1370934e825b8c8c6cea3eab1c45743587e76ab17abf7b8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e2e5c57cfdeb29481c1214b67e47277c26f71ec8b6cd910e1ccfb946119a65bbd3d7aa1d5e231e9a94a1b20ef268a41cd8312d534d2da3bd57d73e79a1c7e12ca9a2d4d33e7a898b560044675166;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h118b74c9d41df384754633b80cef8cb32b219fb0c8f38173d52741db9181aa51abaa5b61e956104cb996fd2a5ac325dc926d13148d72dc8ae7da2b6e1be92d6a2f0d2890b43b1fb581341a67e38a0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h163d4f0ce5ab8b0b47ec4c9d952b4a609d23dfea8ee4e414c14d9a9618c918ed1088eb0ee0401fc4f8d81f7173805e20b5b0119ccea0c13608f845b70dd1e61e7fe12b1f5b9ac5c94abfcdaefdb0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h31ddeb949ec569fcc2201c7c9aa2b328cab0f6b13e7aa8ba7bb8b36cdde5122a651f9732cfaf2b0d002522dc806e295c14adc2be94f64d6d5b22c9f122265f1e2f75b6e887667e46d64f32a0181b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h54be8474368ba71f73ca55a4c4bb9bd34545d4563d1fd0e064fe2447025f3010fffe97b37e6cccd6a6e67f3f728ee754f99269cb7529ba53fcd960aab06de7c3930186edf8a490abdec403a6d008;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h926c72a3fa7ffc943f9c41d5fc2536da9b7d84db6bfbfa753e842e6adc62b1db7d0c96e2d4617a4c0b10971ad118335899bb563324be2fadfbd0e9601b0fe681eccafce68e1a20d1378f248ce44b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1db57b965610ec515063bbd996357786979f1ac6e6f9a37a08e7f7244b83ab932dfa7e85c58fa5ed72d15842f67f5b488f911452f283ce145ce72f441d35fec4cbdb1d73b268880c1808757eda3ba;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b1e2f80290024e130aba81c71b8d0ee80f573b50c2b201ad686eaeedf4a52b6cadae64f3eefbf72c871b526befcb596f49fc64cb83edb1a4ef0ac8a35fc134a5ce6f30d7e1de53672e70df360653;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h849b21faa36b809c1e16ff264a340342b8c5b3552a91f048746f0ac3aca44e8a985e4054386ff9b342d574b7f93459b9a501de52eed082362c2e95cb72f3fc2a4da110a46c7ec306c717ae36101e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h95241e5b8fbd0a3cd528d5338cd52b7dc830bfd8e54dd8332b4814aee67ef7cadc610a7d4729ed62f418a2855d992b37dec8482c8ecaa1cf35b03061244f4cc1e6bdcbe6e3a6e829dc7bb9d9def2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e94d0e4fff03a2e4cfbc0c3f5ce16a080a74bf4dddbd7ff4dfe6f2a37a8e04d40016536e4b1d1c0a1834d1495c65552b270fc6a103a39e1ce5c0f0ade2c8db113b4b0b682413620bb712a0937ecf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8445ef2185620bdd41beef17135176fe4d221b219d7968cf72a68ae3fa8c48cdafd912772a57ea5c6a3baff7abe1a358d25531fc7d66266d0de2b0b47f3468aea93256a4c0a06e297d3bfd0ce84c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1167ba0addd4de9b6e4cf2de06c79f30f6ae37296009275aecb0ae54eb3fa1439e276e60a9a78a49c491e927fefe8115b42f3b41545fe01ccfcedf1d05305cf3188f36094301ba0f1cac05622183b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ad6e1e20359e1777972bfa4af8c8180f6bdfd84caac43d9b42a6185cf022e6694a76fe2ae9b47e0bb4243e39636b58a24e2b333f03a97b39d7e6b0ebd13cb2de9de5103969af9ce460a28d349f1d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h105f99fba4797783fd3581c9923b609949dbb000c4e2cae5c6fe192a896b69bfb152650d079a99b745019201f8f9527170f66ee219a53ecd04cd3a526e38a34e7e8871613035c4584d8d6b6936b48;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h797c5eedfe0db8c6828cd06916af0f8e6676517e92c9e84af934418c61969f2352806010833021eee71827c4e733d7ad4a4b548d686f5bdae2c1743316af99a1df62159cbaf5f150536692322a1a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ae9a7020d88fb848780c813b3606b61c49cd42c3b178f8953f4525a5b2c6d1f174cff43f68ac544b1e0e2164936fe6eb1979dc733b03f6d766a64de5e0cce233d337941597379d96fafe12e363bc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdf88c307a5faa99e0028584d5f5c801f743c228b22155d8fabba935debce3da19a91566df761b810ed29bca991fd8aaa90469179b4020d3942d0a648a52d52a385ea1b0ac7afbbf3ec8324797b84;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h917c2e4502f69fbd7caa0e9428aec04adeed8f451a13d56a59da25fbc764c8e205edbf114bd82440464ef06d06be4ef5065366f7cb91234ef7303f5f53793daa23efab4717c73c66fae3eecbdf61;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13000f5ab165d93d3966c86ac77bfd87ef90e6bbd78f4b8eec808de11cde332f450d98f6cdefa4f7b0c90b7fe09c0b30f6473c740444df6b5f2e00e6c0090af276903de5eb03ad12848499f23b62d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hca1b18297a4b4ab1eb1ddf2705f73cd78b012e733e105b3616722327002cef8ac822a0f0bc4e885d22efebb256cdcd27bc6b540226693ada81bb89b9fdb10a27c9c3308942ea5f435098b6e6caa1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d2bbac75468e0c2db0ba46d46234a50592717f953181f413e7fcfcdd3f1d484b74e93af2dde76f04f80ef8607033be21826b8c8d09fe1f916d56dc51f41eacc2957e61ef6b108aa18442fc52f84b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb17cc9ab4b62909ab4d90b61708c560fce030091ffc9bdd5fdd32e4f213731a08bb29506124f9d491e8a1f26fb86704675868f3d1512a7bd149a1fc1f045a80759ee7b3bbc6fcef5683a1aa1c288;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h95f36f7b3731576c1088345db29aee62fa706748c4432d173849b257889b19698a4d78b705b795bbdce97f252c60ebd09e7711a9ea7a1b4f5a0ff3d96b5bc6321c9f9f54835493c1ffbe7297bdf9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12aa415f98279ee3dbb619c54e8f41cd79c2fdce41a5ddfbc0b6e816966f0d7c1055fd54f8882fca13e71413b1ce48d0149b311faf258a42a832686226bf1829ea12c6a315e803ce7069c644c9a0d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd22a453491964a222da66cd9cc502538b9695c0ac34b90272e07594598fc799e5f1d794b61edd7d409f2b318ec29873f6ba1070a649dc67a69fa5e15fa295ab33b846083a4d8de2b392511d0188c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18b5a254ed7e4166e0d9b0ec49cd4f4510ee0709039d36c3df59ad4488f6851eaf7f8a41e385c00c3e9c2b972289df236e26e180b9c8a1b09a75ca5a5c0259b6862afa6d8fd83068fb396d1d3bc3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f21e9559b98860f52315f1b0499b0707ea9fdf53ca66da8dc8e0eb63ebbd3274236a5276fda71c337a43ca3c5f81714f3325cc298e0251ee79d12a762c8786d0fced708a455209fcb704b1756260;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16e8c2b3486a6681fe0fc5106ac6125a90fe4a02e750afe3a309353f80a14f8150e8a118af29a297ca1d9656ddca1c65052ef496d61d55bef8e3da3260221b9c4a865976cb34d9375add50c1f141;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1416074c07eef39b2d137849ec590e61eb836452422f75eed90f5d8d0aedeb8c0c387d1b14cac62fad2c07b110c6b36a87081643dc07be4928be24490ebac83fb3e49aa9ae398c7b17032ee3d1ca6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c4af6d6e0e8566ad4ec8d8a84eea07389390182a268ff1ff37fa58b94013d8941df6754cc19079613f4f9b9b1fdc4fda5aa06255c2bef4fe2d1d69f4c09a650dd5e3cb34f215244bbed831c1fdb8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d7377ecf97cd10ecc7e0b8ccf75799cd586a568eb5725153fe399c7e6473c47f59792bd479fb738a9d2931df4d59fce55e9f944765a01b99b21ba72041be3a3e94bb7795a4d967c511d8c6b10de;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he2cba176bb89f16011dbf20c8be562ae8f9a778c3153b0d53f59a494717606e55206fc61315bd8d6b9e99ac33d01316cf037a3c13fb6576d0fefb4b0c36d47f4e5b910d3bf59d4e71f5c011e0e4c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h387f8d1812ecce221694a549fdca45cdce661bf5d711cf28c50311a0655483ee0b2c51b286ef98ee3917b17558932b20d7abbf5e292347ad917175a89e803fb5d10c67d587b973d8b7279d886847;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he9d35aaf79a9721a9b3e8deed3104b2a762cc69c020512c0c3f6e72d09ce2d110b3ff3c0ab28a6c2bc0fa6ed07a88406a485d4d26e1ae6f79b179125c5ae1152f68c4b578316885dea47d3318f3e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18d1a2925db27d8b4fe6901f162f8bc0332c8ae299fb942c79e2b98fc3a6f9f9ac584a094174cfde1abe34fd2e958ea462e3a4efa68c61708ab91950d20419b953f69de4602aaf46eef97ceedada6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19399bde273e051d0fe7305cd3177a59f8791146fbb05423abfa31037ac2ec1d337521c868364e6b1f1ea2c09eea4684e01d270f642a66a329352ce74e08140da6f7eafd8d18af80f4a7144374b01;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8257c8b62b156e2bbd31978846dd111caf89ad20e82f9b29dae5e9af4274ed4e0c8374786a39494137c8c85d473ff80e4db2a14c37d509cbcb9e50891be2e002391a3f8f8dd329b55b320029ac24;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10b7256e40d6b4d5aa5c6be7e22828fb5b9c5883f814d59edca09f081551d4399a96b42d649a577cbd4abe397d60a486fd7f54c4015b9c0637adce061f998e96c672ddd21c66181b585d9b52f5979;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bbf784837079d1807e44eae34e7ebd129762c0ac2c90ef821c84bd4c4993736d492e6215bddc99c7cfaa72b53b3c22f464c59593ca19a9ec16bc577bfa7c8eaf69497ab1e1f27707a735ef8cdc9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfea7f4b75e40a7fdf4db0381739560d6d4bc518c0b1d44d71d8d44482ebae367eb244b68a526a8a2e49de30fda9e5847503dfaebe2e56766e8f76f91206f8a7752fe59c3ee866d6d225cf3a9e3bd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hca53b8814affdfa1d17a511a02f00de929b697ab66539d26f4a61752f756ffc75eb02b3067488dcc6e3384c53357adb3376bbb5b45227727948b01276823135a37c54d68b618f494ddcac1409ee7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5415d5942ea980b3ca052914d32d5bff820a8f80bd2afd23e888fc5ef3ad56161a0ad7cdc2c0de1691dfe22205949abb5d3c30b691df2ddd3a4f9279a50b28b1b854c439a669e6ffe131caaf0055;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h109cbe44d01bc7ed0deb3ebc42adb5232fa230ff740bc09147b379087a6a48407fd62f6061c05eeafaee369ad43944994224858a48b10f891276bd7b4813e8959f4e91cc367ea1379d800a9fbb578;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13221a8434fedb5b8643df9dc75dd0303e849838d1bfd72e61541683c1c8c3099a86ca32eb7234e5d0e78d78f990a2b939f85dc2f543d948f90815849e351ec813ed8b129e0e0c4ffe2255bb70efa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc97bede56a955428e9fc604940b9dde9a2bf210407b75ba883614ccb2e885232d0565fb9e539f1371655e40defeb0674ff19cc6c44dd6c3dbc9af19a65ba1536108d7129c0384a516250ce5fdc69;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc5eba74e8b7143b941d00e292bece955fcbf140d18babf9f906c2a8a14501d2fa70e90a7962a3ca4440737748dcdd5382efa57188563a96af1356f673f01763a9e6b3fa3c6883653807050951dc3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he03894c7095c20098c5c9413630fa9c8c95be1ad9b074360ad94c0e87a3051c916019cbef86844d98c84f656823cdc051052729e83a3bd553b413ba09a014d585a4a9fc1d21df7c701ec62c64e0e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e8b3f33601233d8c73e59398ad24070340b109088a2559af033eb5c25179dabb5b909968646247b7a433e3b40dda6de1c17cc92d3eafe1b6da25d00842436869e18b174d5697620eb69b20e81fef;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2b82aa7b046cd7f62e21b05bbca123a149fe820421fa4559eec781fade96bd735a17d2dc853e0dfd6ccf6cc847f62289d0c49662e48db8abb3b1c1f1bf391df99179fd7f8fe76588a479c6ffbe05;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h171e0b1a06f330dd8d6c1e1053393732ea899e6f1524ff479971956595edf30bb2edad5f41dda9d2845d99d623d397e8362913027db2ac3b71ccdaa257bef899cce73aed719803259265f4419783c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12197c4a8547b30ec4c94b462ab57f185f5e6b0a9600b65790f1e9549f9924269d5b5cfc06ec40d4bd5658b17e980a562ef0b4dcadce0630e10e8679b0fe60753ec8695d5bd975a99d636a8ea90db;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cdb883bbba090922513cf5abcef60dc0c65c304c6998c0a0a9dc9b61af09fcf589ad8e188126c449331b685c2cb724844d72c6c06f65e1bc3434acda8396bc580a10bc4a2133b1811ca3ec3a582;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14b997c8764c55f079ccb68e0fde443793c2bdba17e64ac76b032afd79aa33ab5750366fad6c9661975fc80a5471a850f3d5d592544a845a71fdfdfac8912198ae5b531e68dffbd7b7185ac37632c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d7740158b3d2fbc9d8d2183154b867ac40d78ca2909899d9157e6b852aff25b719ac2164054319f7312e1fad50268b2b9c2c14f70862171097c92508ef801de42fdbf3b245b032ae4110e1fe3cf9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3fb102ae518784ba5d9d9a0a9ee507d8c4fd3792ba6a8217b3c37737769ab15884ce884ac18d333d077de379cd7a15897d381b4d34f90bda9e8f51bd7ba0b19c2d7dda9f8ee41b9bac98dc98c876;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h57cf4645faaa2bec24fac0dc69a3ce5c32bff79c0a9a0b100a4aace1eda51734c24db88ffeef81e041958d3c7efc2ed4f59e431e3d13ec909c1bb465f75725e07388d9d4deed124b27133dafdd2b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15e3ca32be37f93bced243686b6c08a2e9f95d8f75263afadadeb5cd1cc53ad3efb55ed7a7de94514abcba700d4a695e362f648ad12137a00373ec6a9924f13805092ef1966b6dcb6241df489221f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1606f2390abcf30ded675d0099d20fd9656bdd0db9392c96bdb360c5fb46f7826192e137696d058d880727b443a1fdbdf845a1883860870114bed7da2e2d527be9856cac330529955e9255c12509b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f3c1e05041c93b68be48c89710f613d3fc536578960e5ba7d351a840630b3cad3f153b3134521363b7276d06444f3f911706544217113ac1f024c8b12b95c46fcf94b48e4951983177fb17012edf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha4739ac062dc7b0d9f38c60005e83e30bbf7a3df7b94868276e806dc655c3d8139810ddbdca5cc228e3c517ed051152b289d52ab5ab7921d27ef3fdf2334daf537cfa699da164a5826fc368d4bd8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h896e74b7824ca375040303684b4658d189099880e70738f8b991fd3eee5834041db7cf0a611879c5e8eff6096aca1337a5a4debb388498dd115ed2addc2dfd2fe3fc0affecf5bd6ae3f88ce3768f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha592a1b3b7d3470370ac0734c77f15cd3789147d21b714795d903bf2fc4dec6fda2b201738460f8018c55d9e13fafcb29d72947816264110183b6f84647a823aa43dedafaab2d9f18db8a6d03902;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h55a74d32f53fe4bfa0cb2ba10b5f137dd66f4dcbe88c32c4d2304658c9aa57247c3b9232ae9d8dc0d150508028d4cef2950275549bd309cda0d297f9455b0f41a93652b62e4b29675c2b1afb2f67;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4caed4b4a3991b9f614e7edb1e9819c0b2e127ddb36a11291868e68b36bffc03f11b70eedcee1c5ee8934035ca87421a1420c3a88449c4715c58a2d4cd66833a8009b444ddb8b949482aed4cebee;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h40a6b9d63200f938f9579d7a0cff058f6f299d6ded5b7e221ed4ff0e21a2c6647a96ba4b34b8a051819e968ac71d88a056047a1e473e2cf647ca36989af7a861c24b8483232b50930cb5655a601a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11e6aaebdc7b333044ac26849e533c0a9a6bbe00d218ca2b73cb4372d8c3e8e7b1336c4e2bc56a6e757da687191bd62f5a7017317137bfb0a12c76e041bf50c736f05bb373ed939d40f8da0c3953;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc26185385b7b9743da979bd711695f681d73d060a15ddaa4974f18748877032f7e1a6d54ebe2f05d166c6bae1639e0017486551536f218d513dbc8901f30140c023f9cb8d6742043f7c286726470;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6d271781f05ddccbccdca47f64091ee9c2cf2a4e619fe14afab5de9a0e5e077523700987fe2ce36bd35a6d6e88bd2fb73df177913a112cebbb0ae7bf8259b8366471dea24449ee986d7c81649ca5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hae3b886f32f2dc4a9d48f272e474fdda7464a8d866012b271754cdffd9c51bd258a06a1944c93175ec4b8cdf4bd0060ccbf7e9ab293d37254c7c826ffb50a742dc7c5dfce599f0dc83a0402b0a02;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cf4254b92af32e1cdbc0a5154a6e9b088bf75f54e00eb0cd1ac5c297510c910782e04681d5921488460561bbc17ef05fa56f53888f66ff92fd9498288d41ac80ce31fa20fa2af8a450f8df1bac70;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d3d8558b09cfdb5ce589fe071509a31785d0878eafb310fec1de1dc3d4e81ad6e9febb41d787914cc0d2e6512f5fa7c8933773c8159dadc727116dc62fc6b35a3cc4fd4cdc0d12bdc1f501686f42;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10d409b9c4851bfb09e824570170eaedf36d303e69f99690b3dff12a4458ee5aea73af9bf15f1394f7d97fdff8719a5de97a3e008bfc5f7f86bc35b182a926ecd2b1c59d63818c4ffd83cf05c408;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h519123f1281493083781498161c3a0327b81c192a37df0f6fa8ec70b68ab280a22665a332114f7d30ac98954d3ba34568287a948ab1f8207824b880f265bcd6f7b63331b0b64cdeaa259ca10101e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17921acfb1883ade99a6e2ce4dbed46b914b1f160cc91aa48796062db5db9ac2c1ac9e5f3d7c95fe55d992ea62d00a626afafeb80e1b28c0ed45e81b1b8557bb242fca97aa9549d882df85476302a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18839bdf3748930bdeb2a016e4f1fea4e8a6a4a4b0b8c96eee62b7d6d23719cb212f307c2a439764e5b3355a2df42abc2cb10c0c450bb2977a9a7badc24da9fbbb41479947330a4532513c2d0194d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1579d8f4b9afc3c974748031197d778c10cc28972c6aeaf92fa58e19b664fd8f526ca2306e6fc11f6158e545cacfa357cc31b8506d54c1fb15f54a19c964dac177e40d5d5c0228abe1aef85366a45;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfe68d74aa1dac57c7626e638b87455aa25e68d89fae92b745ed58b23906e173cf030177c6e1153e973c1d5568cc5d8dd23ee92a1cf3c5386a8b6dcd17f9f3675e3928180ca0c744a6ddec29495e3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb44a6926c1adb16140191ec5e7cc360654977817dceb5e65b0b5b3346fd088955b32916c5e845e6eb6463cab96a57c9efcc6c6dacbbe0996503dd44eed407b094a6b72fd9852b02d5bf6c322a52b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e111613d8ceeab2035427fbaf6cfea93cf9c1e1074abcbb7a2f19579a57d2b474c2e2fbb66549f9f8ad12e2b32413c23bce40418769e2e6b466b48aff0682366da014913de4d531728ee892a6e8c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h135afe0c04c286d957b887354b767c22d775cb949886e574cec073dacfada8fd3ab3f1b5899730c3ad13d2090ef4b2f2e5246e32f67cdddd0b775ee20917daf12249732a24addd56f0cfb78a4ad6e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5b81d25f8e14bd1219ff2aac1313797cda38cac1775b70fd670ec235045be2e96d46b0d98ebcd2eee5209eabca928cdff560c3382d66df54b260f22f55bd55a5d69def532a7109780bf7f8324d4d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8064d0b5c0ca4571c2e57867f3a07e65e87813c4c6bdc2d359d1413def0c0a6ecf68a0651e3866b1905c9cd194d16882925a9570f7db7d2b3eefbcda5b35731b6fcbbbe6bec23430100c05fb7c4a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h86d607b79f47e662598bbf6c8baf656a1453b90f48a7b708fa21b6dde4d5636ea11c497778807a113cd4f6e73d24c5867e0868c65c1ff884ada0ea683f65f308ced05ff09b7e30536f143b3da041;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h31c9063fa6d495989a9da6c3a0c0950863b6ece2595a562f6efd41c4168bcaf61ba1972f8d796e3f5433ae5b8d77d86b388e79bda060bd6e02f338121048874289f4384067a1818343155d6adc6c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fe20ca8b624bd85a2f3f5aa74251b3386a9c9171d3d8a46749a1629c8056829a5b0af058f3618883bffd17fc1d0af80724915b84980b3c1d7ba2fe19e061116b8aee36f8ccbbbfa43a740699445c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h193e653ea08a7435cf7b07abbe237031044652e2ea201893cf4e3aa8ae5b610d0579cf08a5bff89b19281c035dd39f01a0dcf26b04c980f6f2f4f78a40fabdb75c8baedb5e336cd49d013ed8f831a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb733623cbd01deb5e6f8be98aab7ee44e145bf8cdda8f0c3e680c0f7e93a9af7570c031f0f33a6f5266ac14719b3ca113e7e75e59a2d7bb10ef467cfc7299ef887edf30322e6efc711e06345945d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7f80ce5ad42f9975d085a30390d860b4b6ce9c83a961a5791885b524de83d81e9a3164d288787212831870efce9d2eab4cdb1ce7afbe16e2625b99c5f380cc366745bad3af9b59ebdcf18a663afe;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18203c5ddb36aa816babc63029c6bf914c64cd28da0da1bfaae49fc1e319c97945ddb76817f0e432fb08b132e1af3515b9fbde544cad64d227a8c60442d26bb9ca5b33a9d0dc071e155f5e6269477;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb8b1b1323f66cbba051c5fb330e14afbdebf5316d62e75beb9003c618d63b475068493095c769d65d7ba54e034094e12c052ed53d8c751dd8d3401959fcfa228417e51ef53c7656e808c6a15a3f8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ffdf802a154a998b392f3b7534f3bd6c3826ddb084265389bb31a6494c8d242d2d5952142584eebf7ded7ac838dc41e960d32d50c5b1d749b177c2e0085ccd4118f3c4dface903b95f1ebb24e259;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ab4e11c3e4b494fde3c4980e2c1c64b3a65b71ad5fbe291b5aff913e3f07657b7f58fd9197c7cf013d235ba89186ddaf52d8ec6fe2855d2f48fc3a399b63fbf58ad82832d9f7910a24649b21f7a3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb54552d1afab3ed9f80af21ae73447376425adb3f8d95ae67ff986617697dcbb9e70149a21d9917366883646f9f8c6938fa6655487cfc5b2d8aaa15638333a5aa4bf4d3750049811370869c37457;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dd26c0a95a3f7051f8639878167ef560845334fd23e30b5981c37e563c72d6f8e5841c996eaa04ad9d00fb2797c5f3f57787934a27ec1da3ace5180934c58437ed3361b9757e9b710c51d41967a9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc2fc344927fa47045240253f28eef137cfbc917979d046cca5dad3a5e75a68a1c2f60e335d58fddbdc962252644f54f3633200a8cf86f390e1efe5366fd4af747d3a0bf2981ce8ab3b00608a3b4e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18a415f27addf69323d9005042c7343851c2cdb894397a6c21bb7675607c8d9c745604c3f4789779ded4738999c1827bc05c5364348adcad30daab2451af2bbdb14bf440a7a88be60ec51c876ed0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1acc4c4e497b94580b2a42c2c5f23da55cdeaabd6d4cda3338e01ca0a80f5a6ed1914dc503bd4eb6c1a6a567604877a4683f99c8d6f5259462ff8b8ae7a410743af74827dfc4a5caeb74d862801e6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h76e7a881239fd276287a462b5ee87bf659a0686490c5801d94b520e2cb6bd7fd795d159be4e3f03c55c2b2cdb439858f926deb43d6a4e1b72ae0fa8ac366d5322d37b45be7620ae7d1500a18bebf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h531c0f1c5887b10ba8d5c8620ca4428349a7f89341945ccc9cca0df69ff40fade7ba7f6122d7957a562c6d5953f79e22436dd2e999b3e5f6bfbe713c790239643c3b5559e5f84d782513d08394aa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17f0182e44baac760dee5c11e18cc11b0bb5f41a7e1154c18bd7efaa05490b36a6dedef5aa6a63f9be454dbc39260680b13cb48245fefcbaf64d34c895ac407e10a84991055b6618cf2d0dceb815d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b1ba302ac91e1eeff72807d72c50cd1b535babe2b6281f555b43c09bcefd1b0e1035ee3b2d6a06d7d17b0c42cce565cb0b203dcff67ca4ed7069f4c2878adb8683e2020fd2cff8687f4392845322;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d3673648577cba36e03c810b5717557b10c691f361042f5e3ec553b25f7acba94a3d22fd5ae137a0ff979dff7df1b0a3386de358b87809b67d009753e278722376aa4367edc381d8a44be3ffe35d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h283674374d65798db24b27c74270d04e6833704e0583a4fcd37e99b111a5a9c31ed48705fad37bd9a2b7e0771fd21359ca89450acbc220369359cb8b402e93ceddbbc867457ee13c6f2094d75f9d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3404bcb4ae5f9ecf5f88e06280784c519fccbeeafb73330c4f7ee07b655dc9c6327e703580112071c6d5a4969ced98d88a63250816779308fc1214a4f04a98789706085620bbc6ac86fdd6054dcf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha183464cf1b6c728c4399e315acb6cb833f308ca02ad30aa623e30e93ff0101339322a32e73bece9f5d12c738fe7241e24ab7e3a102a94d4e2c66eba78ac0bbc332c198efbc2f38fc8bb3d3ce6eb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16e571f0c498a7b8bb852394ffdf1679ae7fe109290592b966cddbad5006ae20ba2d72e45074a2a2bad4360fdbab64de0e6cc4820c878307b45ba46aa0f05e861200807c61159914768a5427c5433;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1659206675cf04227224887fa60bccb6d630eaee0633a6f559790cabeddd2b375f687c05addd7b923724f4772a1e04e0e72db8bd960e152cc4af0153f027880be1ce064e67917bb0de7e7fc85fe33;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb6ea8aa42d407f14ac6a0de7e9f1cd8b983a4bccf36eed47fdb4c5278682db4344486517ba70fdcae6f26b7216c62f85b64ffaca0abd6d8b8bccd4b7da5df4610934582ebc2e430d430a63476eb6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h187170032d884b314e8db867371df38d945a4cf31dc1a8bc2ab6c31a1c39a6fcee9389eeb6bdf6448a6979e0a82c31692d6b773a68e566e04980a1538347d269fde48df46caec99c44aa997757896;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9d6e52ba20faddedc705ec3e972bbdca79f0548505024d0d9ec31c4179be96880c3a434854253ef6c89b0e3d9c08efe85c9014320a807e10d0232dba389ea19bd81358deb7c9c81acaf6017f524e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18746e480f20c4f9a030ed25bf0a058e6bfa93670b7df39bad980c47d3e0b69cc22a256eb4e48812cfb88d3426035406ed2f3dacde8bd996d3d54ec968765982c527ac8fb6a40f05ffc7e62685421;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12a4e3a886a60ee7b9b11fcd4b3619ae9f78f9f2a38f4e2659a05189794a5b8d2a9903bced95d5630db4a9b0c105f50844b990c0a428c2482707bbd7a1fafc05e5a98dc68dd715a9412c7b1636cff;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h57e778b0ba09df59de94478d8df66097a80d9391ac6f13f227c10bb63189339b045908b94dc6ab503cd3bfb6cb33cbbb6047c9f58aec9f3ed01cfc68e84840dd88e3b0970f44e5dc7c0cece7d5f4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd426571f7c5861b8f3b81ba49f4d923985ed45059599c3095875e7ba2fae92042dcbb72d955ed145dda1f4323dd50b57f450ff4fd5a291ba55366fb4d202f5a51c38374695f0691c724a7386365e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3fd0eaafbebfd1c223135bfe14e9e4bfe990653f84428d884bf409a8cd6e35a6dec9bfaccae27e96118c7955aa4d31ebdf34ff07c0d2daf7b8e48a34bdad1594f959e383f9acfc2508a0e7319d8c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h72ddbb9fe819ab592aca6d23bc976342e67e3abb896578083fe1900700364b4e87dae1e22e3219dde374e5c5a15327f800d20853e87f46d278456125409dc79e14f3f4b8ce37d3c7e82123e071a5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ef19d26f952f5bc07cdfbaf3785320f4f5058cd4cfdf01693d94f2cb7ec097370252bb0a43eb3f6fa8f098b7efacef90266c9105062afab016a9445dca38e8f1c135076511ef7c529427df3a8903;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ccac9aa951868417fae5195ed58089477d217d7b81083a9f0023f6c27c309381689ceb4e2d3217c50519fad6b504c0b5c53b718e5f63d8ea2d35549ae59747e001227407bd9769b50b74807e8c1d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10ed6af52963ed967f19b0cdbc41ef735af11f734cd4c5fecdb30c980d45263a6c06a900565b9f1114b964c740565703d5e4064dfd198289262ee46e07e0016c8a3ad243a43ee71bb960790466696;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b8f7ddf40af558efa89f7c8ffac4569195f40a9e4b30cc1eead5188ea09948edae90968b6260df21b87c38e4fa93ab01edc1e4fedd8165de7d6b46ae3fd506a259b2a13fdd32eebdad2566540467;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12d8ff8118e6fe57d49cacf83dc3e5c1b3bdc30e46ccafd532e0be70616ec175d2c5ded1fbc2989eeadc8c9f14d3c31a51d1ccc7d7bbd6e944cb6e39df9446b76eb516a913f04e4633f6dfc75c1bf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3c947184230e1b09f442026b7cef4c70253b09b59144b534a3764bde100b9258a3801e5d2dbf0df592d8877e0cd643956a08d7a3ad76c34f5dea968210ff0b2e6f39db40a2944c6a6d116da58c66;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h159cbb7d9200b64320cbd04c6aa138632bfbd9bc3f5807f813c0d5efbd439d11feb678f8ebc398cf19c6912dbf061c91fd0302dace49d6422f61a1b8d1782599b873029db406a5b62a4f2f4e49e1b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he430e6da68e669f9a3f052da1915d3c596f8b4942481de388fc45e9004ed5d70276afb27b3c30bd905c38f1a6239ce610c01aeccc29d1243957c21c0c45625c3b9f8e3cc005d3bbe5c9dc5cf13b6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h22fe3be2500ed56c0dce8749e95eede838d2a94fc7c57cefab8ced00d47a0462973c138cfd761fbdf91dba95caffb1006032cdd417f1901b7e55259492fdda656806332ead472c81590061a338ad;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18f2c4ddb6ec0f393df13d93be2f25338ec2bdc19001b0c716b21beb95131955b9240f08bfc3241bbcb1affee36f201af4603d77472af01316628a7bfc2c33ebe5d19f0818856b2588e0b2b541866;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13b78385cc40b5cda0ce4952ae76117c42ce4ab09b3e115f958032c485a8a27174744edecf90fe25a7edfb0016461e118209f2d9a2445082f0b92189b025a23210664bbb43a3e4d74578a64efda8d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hed8e4b81c546ed9a54be87e5ecb736e8f3c22169ecc053ed322363405dddc8f6143fce6e96d6cf2a5e145f94ddcab0c3134c19362a29a93ff22e480b14b2368c61560fe519926d6ea4a9c303406e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16aeabc2a0118e99103ce08f75d927dab65370566dfb96357aedd2a93b73d225e77aaad66de1ec6b5bd56b1bf425d2a5fc8622421b06cf1146d8cf64df2e044cb7ea782a12ff249a8876a2f2610e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd96b8a8bedcb8c9cfbb7990de88df0d7a4837651af858c64927cb631679e483e20f95de3d7f576cd42f568af7844e2827a1a7d50dfdb392c3b45756fed4b4f927921c499924d1a0fdb8e9748e81;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ffb702ae3423121e57b249d78130c4a752b294b8498202d2892aa2bfdc8ac5371ef05d4908728cd58fffe48ff306d7e9be23be1dd541c8c1f29c8488aff5b7c0c48416c93c04796271e4cfd90f0a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6fb12f223b483b852a27d0a1789ad81e7ac30c369064467e25f08d9571da3bdc204283925d4108c44ff4424aa54bbe8d57d0fd0805711b180583a2c18a5d5be8d6084246d9b9718420caf24704eb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15383e5145aaf685a032faf31e0523019a81eb46d067fba3d168b025fa3b683133cf5fbda414ec3b6c7308251db61b26329e1d607b7381952ca1a47c3cc4d3486feb4dfc90998e1ccb3167303d8df;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b0ee6699ed0f74dd28fed5a1e1b50d466fb22e49382db9e29c22343295959582ff75b65e12e7190ebeb4ff6782dcbd6f0ad9fd57b893e7b994866e8a7e3c9a003bb718b15c9ef0dfd4adb4e73238;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12a24cd61f28c4dbce107a796f2e29aa9930b02528fe2c1c38a37766c138fed471291a79f8f4c4ee781d8fea51c3c0687dc5a5bcb2f1cb180f0c7d7301cda2ad5b3fcc4e33191142d76a05f975f6f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h188c759777ed5b5b19775b9d2004c9a0db88a7e1236e44ba2838ed1e3683922a300971c81e0c69b74d785509dd4a95d59b869b2c980cc9a0ce9d06865ba73372535a0444e1ad4af7647b7c615d401;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ffd65c271193a9c34d50f871e473583ba3b21a7f348e2cace878aabaf02282216c2aeb0896183175d87cadc140292a18b8ef917cdf4d271784434ca60fd4dadd039178721cb477f36d6fc5eb553a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10abf9b925b03ea9b7ee55e8d2630439278b76b628c216a6d78725575f1811b388fbfbeb8d82a1db53c2e8086e8dc242174e7d4dfc35817dc1472e831b68287dba35b319f0fda995cb9c717a11f17;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1437b97e19134c471892af0c6d3cf4032d33050e4279076ebc370d26eeda8be258e8b836ade79e69af1d94915a8ca3f1f753b6fcb0b175877f56a61433cf7762f65ad2635dbf5cc4e993b1e2b7b1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h89cf1b7bc70ca3f50d061c26d3dbc7f0c0c5b5c66056068b4289f2b8047aaaf93979e18a6bc890a56e4150d21c9288a3ef4ca59272f55dc9615376e94541b8688c79c70273ec5b873993d2be09f2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10cd996309c666f863a95cb76460796836c5a93c5eee80faf8ca6465d7f0340f5d297433ea9408fddaecf9c69a9209cd1c22ad74045587ea59bb018732cbf64ab6ee7e4d785053f72167f1b5ed7f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h49ebd1e67d99397d3a0d2297202f04c65b6258b63a140676adc3a66d03ddbad2e0f73eab5d5ee8bb977f805478ae9cea7af511a1afe9672661ae4f98345b986e0abc2004340525696c513acfae0c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h998ecb1d16db31b842e604f411d614ea1d7486f4147e8d6003511a6e5a1fe9a13433e370995e7024bb5587b2a099f4a81b3ba887d74484c0eee26a5831ae440cef21e8afbbae0579cf4054146454;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc8da30e0b8b841f4ce60831a80472f2fe33f61fbb9a0373020c544736eb9c79fd3289ba019d3ee06da2f7bf5131fa047789fe906943b756a5315f07225593a162a430c811ca20e65ae75cd70a437;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a8b0569cccadb6e5d8cc6fd6a3c2653f7a344f0a5446299f592d94e4c36ff241394d4d8eb15e5896c17996a3dd5d1728a9afd64eadc59da4ecbfb4c1090ba83331a74435a86ac09884283c87ef46;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c720f3c3751e1b37433fe5bf4b5fe842322f6ae8953b96a9ecb16a35ad87e8549d082e85c1b0eff98d867369ae4732cb5304c0cf5754e457d9849b46395c825a2186c76918a60e6f5d6a5475d6ff;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12f4b3cb7b514548b04fd3e873975cabde4fa5004ff915986df061eee33d673a3844ebfe0cbbe6eae51bb2b0e19ab4308917fcdf871676c319b69d9881856724e525dd06523ff47a61b8203e19457;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8a8c5630f166291d964ce5166cf44996d226f745be5db30a284d8ee3167bc5ee8e06083d98746860e4fcad324138cf3f3311d2937d2354b8785e42814047886ca0cbcc2c5db6141feff3e002278d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16e1a085d06b2b5b69a7ae14b51cdd06d98221f6ad0a4337ff595219809e50edf80a937682f40b4d85ec38685ab783e482fb031d41edab422b9d8bc3820b3c5310cbe224ea2ca30fe074f1825dfec;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11afc6c049ff71d85cf0bebbba339c0dfd204d4ad9239543c4cdce3b178615bb16ea4d8de541ef96a2ee0d72f1b33fd32a617260d67782fcd6554ef45027ee89a4b114ab6b10c9b490bbf3cb3eb3f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbec73c89d77549457f619ba6c9feff2d076e32b788e4935b5f26818ec11f58679d9ba4a129f6d3207851852b98f3456ac39525acdd03a848e4474b3fcf26f26c069703ffd33457b2544d74934b95;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9eda93cee88d1b7638b0d9844f2b4ffd8358fb21260c06a7ec6bd3b5ee504fe560374f59c5519ff38a1da30cded22d4f1e3e8c34d9b9c42b94cf2a8641add68a1fc03051ee3a2c81a2dfb34cb94f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ce60b4328aac85d48fe0725a53d38de6f8427925a883febb9c87efcfe5648b874669f22852671fc7062075a19b3879c7bab84711e3e00aa512e6bee266b46a4c5d45d27da3675daf44a117e9371e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9c92831fe5c7bf56ea37bda92897ec7279d5c623d788d9923dc41371fd8f594c596e24ae28ddb2a6aeb1f5a180f3fc3c27627787ef2d6a16bef188837c01d1088056f1fa14bfa681170c80758440;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1940c8b92600404cde445d25858412d6edf2cbf15c2fdc954600a3f4a616620eeed233de649d0b273d2479fe1ce441278f9f3a3625add743811b1fd010acf533860f5ca24838b8dc746756265a67b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf59206f72ceb94590d7e67539042d667b15e3c2f652db26488e2f3330ed7c109521cde463494a10a7dbefc6998372a594496acae408e4be82a9ae0135b1adb101b5adaf7ab0705d0a8784503f4e9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf3197033ef6cadf32296b29ad7d2d7f3ef014b1d205d9c748be2d90baba3b6abd54b1d671c67318832792dbfba62e2966fc2e00d43e2c7fd2871216ef26bcf3b32d6357bdebbb36f522aa71bbee4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h948a804dddb4603e733bdf18781b86b742e0397fb7abf8194d33cd2ef629f1825da1a394207df65a8a6a2e93bfa74c0c81880a2339861b4947fa3ab7a0208b4a1540c0664ba4f1eb6cf4ab87a597;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f8ccb5d14d83b0cc6463d802bcf877586c79b2c642c7711cbdfb1f3331c0cd0fec88edd4fc5fd9edecb0b9683bf96f11e3ffa6cbbfe032a487ae2e1a9b87256ca66fbd3b615d9399eff394f73492;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'had9e382b5bc77b611a250d81d0e79a67941a6bb663826e0753dcbfee2b7c3896fa111e4469bf16c822039ba9d2958ed5cdbb11e6738960156673ee85fdc7b9b6fd77a907aa61b64f72c144c7cd73;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d92028ca0e450f191f78caba8cf836c527b9e8895b8b2569b3f35bba1d15ad40d82719261043b0d535a3e44f66a38d13fae0753323f11e85e6986b01bbb2ea73fcab8409733aae63b30321d72212;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15f707f863aedffb2a8e5b08834878b4220fea69f37e101c91b484ea83782341e369e80669e2c8553c332303a951710949c7de49da85471781d4dc1f204638cb4ce87d2ff12d032883606c29c9768;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10a780f8e9b447bbe69d20f1c8f15364056751468dfe03fa616111503f1c7b1e9632cb426b08b4a352efbea849c3c326bc25437196a0866679639fc4cbf39e03f2938cb6934fd8d862e63e245992b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h129970b7d2f534675aec7e96f689ad6f8157c29a819231d0b35c552e37c8d09144d2780711a604c9f53a3c376789f1393c247ac45fe07baf13ad90a940314102febef3a1dc088523ca31eea6bf73;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fdb8fc94911ef0303161c9d18c29f2245df66ae6754e05333113ccaa670449d7653ba2c4ec000f1e7ed85a6c660e92f1b261583694e8b97971afa7591454830c2b58e130f695efeb6d5cde43cfd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h164f381edbfb53b8af68b345f0cc8a2847d5cae502631e41c0bbdb32e1fb71f4359da0e971dda007773875a0901182f2c3834d97804c322f844e37c492150b7a3fdefc0566ea013a532bce987fd25;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h174cc33d091937493ac33ac500955fc0cb199db31a1ba84e33eccea37cfbd35850ad4cf2b080dd0b4921613b812ae7de9fa43f426ec7bfcf13c3a6569441aa2e1a4a12348ddc3c7ba27d6dc1050d6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1391f3a364bc0a981d20e490fd2701f20bd9859a7c4c020b049561a468f554980b6a7169a87e7c7e7ec1f1fd37b3c96c47b4b24753d6d51330894f3ce96b5db4db59920f019068957f74d2997e1a2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e92ff856290fe28fdda92bae7eadb6062f117c2d5938ea06bc0e4572b5695300faf61f76f49c87dc6ee09ec5f010341ca030c60773978a8d9d26cd223bc5fbf736d062a5ccd7f452ec3b0cbf793a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dbb9ca31ee9533836244104b318f8b8ddd4fdb3cca3d7fdc111db049bd6a6c2878d2137f2acf15819a5aae0e53b4f02cd2a228631741bdc326a9ec4da7047c92857e7f236345c0b2514c5cb0e9d7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e1585a4ded0a99c1a182fd4271d4c5a2dcf8a86de78c44fb7364943dbc74aa0c0d86c9b973c673e8c1cae271d46eb6f854e4e11e9fc861b22dbfc49d408e8ab4adec706d5ef6a5986f1966892ff9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cc8468f80f2e16f1539bfa27f97591b202575428ce531a17b61a9c70305d493035a3889ed1ec6de78caa2397ef8f6c2806db16d2ca6bf70da9109e6c425bbba34ef09abc9d2e4250e1b41e192cda;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d057b5745f0bdadefae3d1291c5c50067c2831e77797e1d9e305742f1104cfaa245892996e45023d973d054a9c1889f80b681b10956a595523aaa4a71fa04a951ffb86b590e4cb3dd7f3112a0805;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12a50b746524174214a406c4f6ddb61781da1d8d952533b74782037a785ede68b250358e8640640f78a054eab795c6e8df77dac157121912124dc272a51178dad50aa7ec07a6be9a2b1c9a48f87b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hec8eefcc40305e8f454024da258f484a101f33b24871011e438d0887ffeb98e1da758d9cf033f0402cfcb9c9a16dee757a079bee6397cbdc3d0f7c9485ed0925387e1acd6739b770ff5c574a6f14;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4485fd624364b901b0bf6fe2e64e386b2d0bdaf2fb031171d30febe9fe64058405df7e3f3b0de61bafbcb72f33e2460b9beaa3af386ae9e023e5575e56ffe44720575c3622cd368ce9803e3755fa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ddc536633eacab9c8f84b834898b8258bfee2d22f01c5489bb7fc54aeb4133f02f1aaac769bec68fe6012de44be565bcdf8069aed2dc668656a0e2b4c82fc6f3693e929096f5650df315f5502d24;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd12925e1641306fe5337c983d675b757079bbc7e5456527812fcedcce1476b308aba8854d24b1f1c801a90ecc8899170ed6e30a4f00bfd67a51f00c2fa969f58fd67d63a495e787bf8fc43d48928;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4b598e3db95ed143dc3b92f07eb3f9a17e38cd8ad3be790a6b682fb3e9986207a723d9656be2aa26d95e3049ac271cfa02ac37c037d53861a9ba7eab3c251302b1250ad42157e53cdb06457850f1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bffdadb1486c7e74d1ca2258efd8811a468ffc53e42933d1b11b009f632a0fe0637ff7f4330dc4cf9754a00bb7a7c1f3a1ef9c74088cd91d8984ca6ff7f427597277a237d38d02d11de18393dad9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h534d4807c3e854542284df5f11fd18a8472514c51da5bf6a160ec04c737f96ee07f8be22073e9bc5766c40ce6e00364cc2e94538fd2f43b526128e94f92c631ba3e83ed065e5a7cfdab5a144e61;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16270af3469f666aa6128e363e414786492ce07ff95c80dd458aec395bcc7a582dae6fd6398087b3966a866fc6d312edf7f366b5ea2e253a81b53696479235a7f7b7ca14fbb4364c30c174542eb7b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d383f9520358d5f9d49573a9fa4f9664b6d6692d34eb8ba73f5d139e59202640696646e4491cd5b53b537b6364ec6ed82fd595332966a8e78bd83a0c75ce38dd5413726b49b5205fbbde7e7d78d4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cab38cc20a44f0b5236f662d00e0efd6da35f15da960a2f981936a50eb62f16b0e0e5899099e98e42a7e557327b9dbb649c07c72c63dae5c2cb3d4370f35df126525ea6464cbbd0b9e4ae019b29e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfb3038c954f18213146dafe39fda47660fc224939b09c01642fced8bdcb6472edbee89478efa3b2d6af3b901c28c6c23bb24bae5ae7353450ea0b64039a60708949179b8b09dee2a7733cdf4653c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7310266a748b28e2c104a87901ec5f8753ef8dd36ab1951082cc89a4b8e86584879bc7d83aa849bfb7a3f4325e14f4f3637734643680354ed7057db51025616b96e55872f6cb6e37e1e2afb67ba5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e54234f49acd0ca807ec97a1cd994d753985b57bb40aff2c0c0b1ce3e1190fa71b28e5e7c178c719f93db46e343b84c12e85a5117d2d55b80ef9539764e26eb0c4178bc9feb26a6610e5cf5e003c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2903d9405f18b8895a968c32ae3ac95b3adb544a4f8787d8f8dffc537e58ff52d68357c5d6835c519dc848489b40a2d80f00e9aa615bbc6f136d5e758c56124dc5c9def423a79a5bbaa02f08adda;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12368d1c948d0d1637dc332a046a686affc58476697aaab924e36223adb7f44437478c56e3a74f4259d38900785be3686f1eec8d56e3d03a3fd43112447bf0d2811b5f8ab4a41b1ef7872c28134c3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1126f9da2e7d3bf2eb634717fc7f4da4104bbaacd8a5bf95444c5e3996df055de6e8e8f351771927c68271d0823377f2de960308b7d74a51d50fbc3ae7b84a4bda1ba0add98ed4855c557aa774403;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cca4af0d97f70e9cddf8d6842d127bcc592ffee3454df83b7b00b3e47e2efc294e297a05b37042db69d493ac7d3d34f01646c7edb32f0bce27c869bc5703113621b7cae711d1f7fa235321f51aa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1908906e670ffff317392bf0bc85ba0efb1e45ed3abaadc648f29d165530fb954ff2efcdce889425c72772b675c12011496c86c5f40a0aefa691705651bfa5a05a81d9f314ca88c6c51a57eaeba08;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h114170c13b65d6428923736a885f9d946b0c7cfaf30a4677eda26fcccbeb0ea67c1b91e0620321628047988d7139f48adce639864bb9e711fbc93b329e1d240fe3deffe3777c7e438e8db1c654c50;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2c7f3554d70eba8b1ab1ce82333a2caee4f073cf4c67a4457064e4f2879fe1d242921209432045fba7c3d3703d1903b400d6f354cd6d43173f1410c6351509922b64b2b4ef52415dba1d037c34e9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h127fe9d9e7a188e1a70d31b04fe08cb2c57a32f019b273666b4b508a11275dc6451887cc4b8222290fda568333d6bafbc5df09c4b793438f640756e7e0ea4d88c6bd24a35a3f3b83f18806812e016;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bbe0037e4693237756650d8e24651456a12593903c61418ea25ab43d3a570c3d13223382475f5cbf30cc93bc2a8ecf5facc3e2de26e44c76129cbe61758f535449bd94c6041573cd4a07d30cf456;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf231b7b70a1cef3cb8be699d9d188feaa15dc121a0f1ca0d97192ac925ca4ef86be07d50ec7affb8941ec68328950b23a682de9487f9e7890a1b966a549b53894b9e1d24890029a67d9ae058db66;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14cfdfb29631fce3f25e2d8c4da2090ea7ad3c1946c52071cafa2fce796a2775cf983bec184c92245de5fd98433a910dd4bed42242d337142651ab5dd57302100c93ebd97fc2fcc4d27bddbf28190;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16e406db085be986037393433500e790915bdd1411e742d10e68679f39654e981fe6244a8ccb012db53a7e0779aad0c5f7b56d8c81c0d5187f9f9e29850c82674015202897e142e70af4703e79965;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eb3f1af6f1605b57717b9a7bbc1dca30657e25ccc8a4d1930ab101825a1223382d58fb19a075a24858f622e3073f72fad7acfc1038e5e6c0f83591525cc0640f77f8f8357d07617138e4b12b971d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h140f77143e38fa9daef389c81db7e76b74cc6f8d0260ac247afdd05e2e3d33291a9611a17105c3a88d27001f81ad20c9853cc8d5439338c38bb3860bcbcc2ebe011d2b3f5700537b7c2dc20ba6c3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h705a72b4fb19408a4d9b7e64e6b1f8a0b04dc8d8db2cdbfac0b123a6716ca2972954603570d2a21055619184f9db0d012fa18050ae0dae2ce8aec503d8787136eb3c1ee7a0467a8278f57bc6ba3f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h292c65b2d302bc0c395ea7f0a1f5ce1d205ec9f0a8bed00018230b6dd8666f09ac40f5667e33958e27afdf193f03353b4870057548a888d0ee3d5048559404e9b1be4a6cc3294faed9a12007ee86;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10b9f8afdd56d6407b908f0bc9669d956941f4a06e4a0c00b2f1b66bd1450af2f1e3220cb637a222ccb9816d65d904a8f7e20c54c72a64ece64dfc537a62ef8723c4e188f55c4242f14d78fa22880;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc3fc92de056d92a98ca620ac79c14591655156bb6662c0278b9758f6e61e3f14839a82d985f784d188f1826b7b4d088d07f468607e510bbd14e0c5f97246368178c0c87e081dbf6f4bf88e1c1e19;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e838325ddd9a48a9ddcf3d88bf14c2c09ed7a31651b17c99f73ba219189bc47dc4fedf54bbcdf822cb6085068643d14fd7695aa73f70e0e6dffbe2f0e2bede2b549e1f14335291fe740ee7febdb1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h74b44a89e3371daae439b12280ae671e5f98e849e5e9817d0d2478eff46d4b21a9a6ebab09c03069dac6020ae3858a006ec68b3eb6fbe6e0e3f81e0c65a19fd252c7c24f466fb5c53ddcffbbd39b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h893e0c918c572627a76bb3b4c138b16f9e93560f8cf082fe574688cdaec0f3d7b857383d4ebb2defb6afef21af66c4db22e67e8059e4ad79fae9dd9669a965a6e2337198e171abeb48905b4c3958;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19abf3c91a5b54bea71c4a1c818312b208b89282b7ccadf1f3bfc64de8e39763639ac89be2a95d690f2189043ff1d15c0574188b75907aa8c554e587046c31ec53c6d61cea3386e985dd1e0e5bac3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8120fd99e52fdb2b66ce329121d63a82d9bc2ac0158660dc0063495467c32e0e0b00f42e4ece9d66da99ec650f41a42a1b3751abbb45e75d62c2d3287e6bfe46e076138c211767fad74c38c1961f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5e62ed3ce5f101384a56b7d7e8c3624071b00bab75e657e8ad8af702e7eec4d8e40c4bd2aecef37a85b3870020b6fc8717934a10a3f695a1818d5257261e73ccc1d9223856959b4f6aea73274ab2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12c7d6d6d65eb7b284a99eace6fce711464ebefd7acd05d0e83ccfb511227e334ddbfcf2bda540a3ad8b9ecfafe860316d9099e9b51c4c289c8ad3b71ec34e2fb6399a2b243372a5ad5053016ef6c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cfbe39b574ca40d2c0c83390e3782f621961a3fa3b7b4b6a08a80f7b509ab4152095d0536878f9bdfb4b6a6d355f38cc2e15f4d009fceeb2731c3dfd4ffb17e57ee09c332c24463e01cce348fd18;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hee3b32f9907d3e152c045e4c94dea8a8bc83e97269144a8a1c7c40a32a95b7f5391bd6ef190ceb2f67317be95b1cc11b7946dadbec6819af8b71ad751f0b87c2e4aca18b78024f7a4ec7b51bbd61;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha08583dd86e6dc9adfbe9569bd85f5cb028f42b6e09e1eea6a4043269b5f28e29ce4064e1b46e1e6d882937e96634b7c5c266bc353a4a13febe05709611efd7209d0780d6f6e1cd81f8b0a89ab96;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h575d7c0237343002ba8222c8a62daedb77c02c751725be55935d86395edf4b2ad306624436c7e9ec759d36333c44295622dedcc7c774d9b177f169ed54d14029d96431fd29baab5aa7f18855f479;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h55a8d16520248c4380dd673c02df73e1a6369374690644ba1946e24c35c5b8204860cd378084b8018ead65233f108ba674355b46c75458af761dc627da8b984cb921d2f796e39b6053b5208fb28b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2fb6c8b852dd6690b77aee8080c1c8c8e2b64a9f383c92040ad09ab55a2b75c6c8b1b708e2425b45ab239091ed776f72943a4ab6596aab9e7e390163fcb2fdec442fa7af5a89d95a44552039c801;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h195e3c4b6aae92c851dc8eb3d900e64b680ad7de97e3e3678d8c0c7dc45369a2416e0f7eafa7550704805e239fe792fdf8661960a7bd50a71344795bb650c8b03f64259ad0c2ea0840176d41b9946;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19562779e9934a09873f0d8eef39ea23aeab92304315c0476a0ed3438cfbb56798fe9312dace15c8dc564b6e6543bf140e15bf1e32599e683a13af8afbd468796502b53c122fbc7baa935b4e69432;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he306a3618bd40728cd0a37523eaa1d094beec4fb356d93c9abffbd22d5b2676ad5aec586e525f01cf5ea3b187aefb75f1d1b6877bb27594fd82d2b44b7efade2085ad54fdd54512187aec6e2a08;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2a63cd70b083122f3772f020cba193a845f3bdab740eeb9b68437ad2da8b972793483d0a110784c506909042d6b97722f3710779b9e13b20b5580ee571f06d10f8d480c159cd308c73795ece5f44;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b41929f5afb3454511a5b57eb2c619abc09970c21b92415b10c65b9ea8bf87540fddfa88437ad2cdd1f7672a1187f2d1bf8d056e446005dbdccc1e1dfc855f77e5e5a6947c2180e4c8ecb081a5f0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13f937319e6e63faa1f72985533b80413c6521d33daa595329d93aa773e21c03ea2a11b0759bb295ce435d3a918f5100e833c705866b8e6f6fd138940863a50e125194faba974e5a9a88817cdc453;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd76e9347cb4ac8521dd2fd5944c1eddff4a19afd6855c7cfc483a6a569afbc54d6949def65d203a1e6217c6eeaba09275702c7158a48cf2e5b110be6ff4ea1534c9f46c01e400514d78f6255f74a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c233554e6a8d9f0fd940f0dc44ad8aff8473fb540cc72aca2baed659769b68b2c0ce8b72564a10df1260cb5019f0bf3c7e2246692214bf14bd7d896bf552bb1dc4276be7d14d95320921406d7a63;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdcaabc21be6dfa879be9743fb79d92fe525850d480980f7ccbc968582a341d2bcb7781fa82a004d14062287fe86f0801a34666a89f8e73fa229efe3cfac9aa62dfa31e56953398d51be970c91494;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h422bcc6ca84f886f4583c176ca3c4bf6fe2bf6bb8382b86a2123f3d3c60775658a54ba7fbbb418bfa16ad96d2820fe4bfe4289d8e55d1b008ec72a214a2e85703ec686bc4ba916881dd39543c436;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h107d1aa0b1032a9fc061a2b4effb4f5d1e4fa804f4798532cbaf1dc5e2f04566efc4dd5cb6a37c4d7adedeed2c3bd8dc37a7a756573797bf1a3ef9515c819fb92b31857f99ef4e9a9d6dbb6b59b26;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h137948513c19174eee04088623b948ef27ab5e59445fbade7933beea7b326013eeec0e4bed211516c9b81c4348de4af984e4af35af7943d176c82a4cc40d993de28a42abeedd4de7da85b906add28;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5aaaf2f024e00b52f7d253db9d951c1c0c6862d837358fe9085ea5ac02270841a1468195f1b9b591177aa574ad27165335cb84d3a769e3d7c3d146113f5c2dad3c2f6d76d67bd7ca933ba0e3675f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h86739000aea264422fc69671b5387e2f73c5a69abd2804081facd487e7048e66bb777099c72dd926f9c384b19170c36c4090a85738faa198a9ea468cd9149fa9aff022b55fa198877d48994e1b5d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dbc71e61567d42da96938ffad25e7db415d8750e115f5fbf5a8c1fe1ab01dda6e056f07fe3799ffd9834e6e86ae12341a73bafcbad47acd91993d3079374665a8335cc86db733b3e731f6b8b7356;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heb78646401e31396f5124b1942a0c7e320dcfa369838207120aa881810ed8c3c5fbff52cac89596681ff6a59d5ec1358f5d1a44c302b40b9bbbb883f43220d8176a5c0c5a69a7d79d46d6b7cec18;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h43c2264570ffa8f2ea7980e0dbee6fb48c60bfd1a6cec56a8d1287db461a6ae8ba7e0bc0f340035ffb430708fd504973ea68b0b1760f44afe8c95ad55dd7a6439948ea42f4885247360a9fdca67c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd069518d001a0098154deba903190327dc5ca6aae39d2c4bcc403ecef8adcb2202d46ec3d3dffb3a99fed1dcbc67ebc97c6852438f4b421e8a7dbe04c38418d5ef8ae5767d380a1fafa936c08324;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a955db2d8fb8a4455ca0dd923b4fe1113b20791a0c66bcda33b8a22685d8be91b2671b8b9e76598b73fa580e23b91b679b8ca8c245430595aa85d3d577083d5469c2ad6cf305214270482b80f246;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5570fad1e178da1aa731a5e2950386b23073a75c651ccc875d93a1504afcf9b411035f6d90edc4a32febfefe643ba66a278f7a9b6130626e733c85e4c47b0c74d78ceca683a1a677a5f331206c23;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcb3a1d21b7af07e7a71d1059e2fcc8a720a1cda550c10cc2b231ed81e953dde0d29443c532ef7b4abea7fc15e682fdc2b9bcdcd937044844e492d5dfc0576191e18c2cedfc5622fa6945ceae840;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11d7c28a57c0088ab747e865ffb504e54bef45d0166caedb044a4163f545569d893ad2f68b38e42adda30938815ad2f19c5831935bf4da2dbbd6040a68250a5b3258eed43624e0339b074909acf61;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14f6a1b77ba377e6be849e7d26dfaca8c5a267633794957187f48e35077da0d81c94c512fef57ad13d79bff5b78fd8a7d9e3fba98d22999eda5943261bfbd73713d5fc4d87ad4e52c9d813a024cc1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13621120ea742a542ae02fb85fad4e40e0fe4a49103489a809c2de8ed90d54cfbf1c11105390ef650868ab9da9f2805633bfd73d9e92672362c56d62b87419b423480cfbd000275a9be1202a8e61f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f53766d0af5760c084c900bad24ce6f972f4d3b9993589acb0ab59119bc78c6355674c0e490dbaf1a31599054a0ca8bbd379d46aa6738b8c5d1bd313c76c06313c92c0c55ccb0e37afc52fa3c53e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f864b9d113c03568f0387490d518e788e12f84d5ea90d0f4ebe90fd2417691622b59ea58342d248cfb629bbf8befe1c48d0bf993236b70c67780bff9471275e694fe3a2726af02376ccf8c1c7609;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10cbdbea31ff6b37f2e04d07861f68763f374504fafc36f47fa2080aa271f154fe63a1f5592727cbdcc857c5ab9e784835530e9510c673dffa774f22c30422814913a5d8ad9105fee3fcab03e9ee0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h194fad21dd79d28b17af7ad40b88e0a48fc82781b64b341b77a877a470617a91f54c0dc1efa1365a270a9f27e471a4460bf3679672d35582400281a73cb2621ef159460fd4be6ffcb784f685c8e71;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he39c79f00ed45012e06636d31b920d0abfb99d29449dab43e04fb7cc045c8e7fed373721179eee8931b18961997ef04de5ea5b698e8d8c7256d3c9c7ad19e584bc3d5c493948df8ad6f0983fe6a0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd7dd2ef13afe2ae24cd8e4caa91354ba536809d0aa00fa8e2b12e3f74cd487310928556e1b117fc8aef93eee12040b3500812beb73ad0b4f0e7e11775d1fd6338c773de992d335409bc657360ead;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7fa82f35cdd629d3782cdeeb5359b63426f5490dbd33475ae75c68e9849e85610a0eee6b697cf9f65ea894f47244ffa887dc5ea98b4374e53c2590f5616a0070642927695b269daf3cc238c6cc11;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h136fe08e73e2ca1c2754903192dd74490be81d536e88e2608628b1f9b62d949f8e418af6a854859b41cbce45097e1635132cb72bd68204a119a056c87ebc543fbaec75643e0590d1fa748c91b0b1d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h324a64e73e79df8583786f9d3650952c8969fcdd854ae6254f66eddc801c4a6cbdca0e6c3cc1ee61e28e4e9ad3c3c7d914096fcd7dcacf8aa7df140e808aed01c402eb42820208e8d38ee23f4501;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a0e361f82d6fc856254f7e735a6b5205a683e8eff3ef5ff2c681d6ed74b01bc525b7292b5974c46e5688a4327775c84f528983fd2ef86cccedd88901f227412e79060efa37a35c774fdfc9f4de94;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1acbc21c30f884ae56677d4e33bfb70c480d93ae99b7c6b7ff95c063b10d9acfb61683cd09a4ea0f826a16141e05430b8d8a7f86f9f6e6faaacab5bdb0a88275f2a52d9555d9c5c5fc4339e8993ee;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19f22d506f201e3c49416451412225653963e5a3854eeb5afe5c79230d7f9efede45077f0f7731c4b6ae991341963f8dbd743b65396dd67239e7250ad1515cfe725635f752dd38d11a70884240973;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fa66208f21c680b72bb41422ec929b4e481434978ce575706ed273aa25f9056a9c6b4b62e2ff2881d634b0503b10421b1b03470bf0439a31dde1bca8362197f572c31ea5dc21305980c846ebf0e6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1167f1c0e55aac1824fdabb971051fd30f9a16d674b6b0024d781c4405686a0d1cbc6abf35d9dc3643f3c9939d419bfef2a9ccd143ce893737f0e14f25d8b9f69766391c509377382b23091881088;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc9bc8667261b6bb00ec0b6770b78ac37ea2a7461c42042f7956159fff5ef3179708f73353a63dbf10ebf0a40bcf827a540bc587fab9f037c637eddec792f5b07e93be4bc57db108d264948a82150;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he9890c840ae535c1b5e71ea679e380a430f765f4e0a84df557f64aa435464ff2eef4b81dbb78c9118e997efd23a46f3f112c84240ac3cc8d9f0784ce0193ccd263bd21315775b1977b847d67add1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c745e87140b407062381d5eaa6f74848ff80a4dfb197dd75140cf273f1a1cc9d1b912d01807c6234a40dd03f639ee626347ccc4175c2c4e0a917df6e3fd86cbb954aa3bffebf4f12eb585d7bbabb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16b00cc9e2278257b2b6bed0e851b07c1b9e544865fbf1e49d18cc15042e2cd5a3bca9a87d30c05f905a55bba7b98b49ea777d33e7b6db2795979a755c8acd35df393e5cce0890b72908398208e73;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h54586f3d3b5496ff77aa8826917c6b9a65caadd6a4dd897d6466654cae3cf18bcfe808df3e98f1d2fde848594195fe4b4507712c9b76a7e54408ab512897f97d18f9d30106dd64646234c99b5688;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h115edd8ed06879bb0ccd2655fb48e5c3d0f4ec0a00be07d44afa3ee0c3348c75faa2931048c3a75448fa947e2159ed288c929f4dd280aa54b17407a8fba134ad086b977261a921a7e72ea23cdfc3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10c8aeb773ffdcd46fbbf5bbded0a68fe25ee7f5d443db3b0092eb66ed8b147706f7b5395823e8cf11e88c65b007b7fcd6a594020686ff6e36be2169d308cecfaf8922a824750c3df8b0f2d4b787a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9ea1001bab1c729a854ca9cd4f6dc312d98ffe0b52b590e110ea068de507ccb30955c5a172a576cbb7000ae33c4a35ee45f82267381db3bdc22c2db718fd758096c9e4aaf8a01a09c90b4bbfc843;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfef5aac3b24a24d61b07605d9a079c76adc0d90458eca933d322fe8fd59895760168e73a36e067682163201f50ce96e04e46818d73e39452241472782cd0c5f25e1c2714fa95416c289abc7b4d30;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3b8bf6b10a591c8dc1441da0a7cabf887b73890790505a26450cfd6df309bf54d398dfbcbdbb432e81c2b28f57365d0888182ee0d97023fa979d9941867f630433b9d5d627e8fc15da3a51086f67;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfe4de60a24d82511eb2a3fd809b09e85d3fc8dbabb7735d4a47725c8fbbfe269b3e20cb9b822b6c22b0b37d0a7caf2b176101b3391533bf707c4a0a8142fd42193b0a09522b96da40107fe13ed59;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c1bc658e860b70660d9f8687c5f5693f2a2e98b4b6603b760c9d046bd5345a8663cbd26543612d98fe3e00252c3881611f976d3e48a25213ed8114371344d92c4c5188faaa57c635dfdf4195c244;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d7802467a814ecf8c83d5c0b8ac025d9ba78281713a1fba8372035fd6e36b274ce0034f4d609ac7c440d311dc3d48f354661b25e4c00d3c392ffcc0a0fdc75a02ee4501dc0f90748a3b095331082;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h190a9793a21bdc706cb336277ea4ecf2583c8850b94343c98b0f299dd8537cdbfdb842cb807e2fbe58d9a1a703a5fe4f1a00eb05c9335c68e100e09048da56302e1cd9624ad481054cb6e91c9cf91;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h159bbf9937fc4c1d1502358841d7b6642fe21d497e022a9cd899083d884763399cd3aecec62b35f9f6ee36aba4665a0118e7596e3618992c3f7fddd197f37aef3cf106ec586d5715a2626c294ae89;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18af30e923cd9c1a43036485b8bb2d8b44ea7091a42d9bcffe5434fc0e64cf0d13651f1803318483a9d2c76585d5895a70d4e1307908b76aafaf63790d85dcfea2d55e4f48ca5126d205b303b9362;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13a0560197cf292f9ec53385fb01b5b39f6ab59ba863df7069e7f52f5007c024380bd44b477e452958f3f44a823aa43b8bfab836b0ccc2c307c4952a63cc5a0efa5bf6ef7c8ad0b8249b5ebb4e90c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2b8a2af9088170f03ddbdf332404acb9c9510f4067f0f56ba4b55515489acba66cf736027434531bc1c21620fb0a96e0fc0adb2c4fc70774bc75edfc324b079db6a6f39f5397be5ddc8523f65c4b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d285fd56f39d79ffe959ca4b1c64bd1fee832f11ce13042ffb63ea637f154a81a7a92deca29044d084baeb7cc1ea4eb8d66f48663ee5fbd88d678432943448ebd83aa5b9bbfdcf21b4b904c7755c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hda2b61409224d6bf6c1b88a8ec0665eaa2ed5ed28756a76db247011bf598e70a654cab751c24df96af7239605ecc5d1dae77c5901aa9d58aff1aff6dd1eefa101a2e5cd11fc0dca9d06bbb2789c9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fa9f901b70756be3fb4ccb61e078ddac7872fdf897bc1afd741bff2710e8964682846356dd3d7efa2f715fa4e3be2d7a2d1aad71478dd0746353d49bd3e035808fbeca778b10e83bf0d06e3a30d3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ff4739a4e7faa0b8b2c3fe7eba6c459aea80b216abb3d554365fae78a77e46fa28d9288dd998f4d17951aebd9822f1b3c1186f2ff40089e7bd4ac4a2f089fec75a3b2cf5fcb48067a63c514fd195;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1180f0bdbf7e27840d4f6e83965fd3ffb0ba09a23ebf89c75ccf7c9c06b99deaaa59ec63c722c32d1af129920f0df15a8b8a66aecd6ab2894c0a651550338998e6578315d7e920b8b3f0cd3b7f07f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17a9079ffcc40deeabef89c67fffe06720f20218182957701c639f032be0144dbad210821c4bc898a0e37688adc27159bab7044880eb40cbc015221231209f64ed0082910f4debe407d3eecc4f1cc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd04d18bc9e2fcf8c1d336983a5046a2db5571722f9f540010b9a33521e348a6099010df5496447f5947f10cfdad47e56550a3f96c4378c1864863b25e3e3284a6fc413712d1324c1ce3a53d6de6d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15caebc465af64286a2a331de76e019db3a5ef86dc0e260bfbf84215000beb218617cca7a9f19bcb5fed65eac71537dcc0e57dcc58b8e7e8e934df16dcd915176bd620c9d1c10c54099521ed525f5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h62c401c15e2cc9e050a5c6026572b803e2762e42c8558eba50282fe155226a10c498d3fb573f119c62255319a48d52722cad9479a302819ec63c540d83febf2193382b05c979ed091d526858c495;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ec8ddd2129bfcdba804fae2af7d0ff3c8f616eec5f74d2f336e64968ea45aa11bcfa6dc1d9d04b043015b51fe9b0ad6c113b2c3e0a7f411e9bc6c369295e0623bbb46792533de019ba3fa37fc63e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ea3e3df4e23b4a17df77736f9e9a9850d64a1f449e47a72526dbf11dfb4d7266b3ec19edd1933639b2cd384e82587ca8ecdfeb472df0664ab6c1b299659f22b88db473a58669d6eb045275bb52f1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bcd5039907abbdf55e31328893f09be31aa17e2f00cac01c0b2b26e57bda7c2425e13041935812218a8ff4bea3fc831ed28002dcd7539e45a3e5d26e375c7d131ca70264921af4694d08f0fff6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16a857444a08dc8afc030d9af0d3679b9dbfe3e30577b3532ad26be0f5b4b64312f21ab58c529ba34ee02adf6433e16df7b321c34d988daae42c5c9718eb81e8ac00a89c799480717820097337602;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6836063b90af9d170ec6fe9516b5277883b80d12f6cf7060689519b120da75080656201e43af2cf3859c3378b591786b6dd0f6c7d05c6e855ff26d7a15fd5797cc86b59a0b86dba464872b719f4f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19ee930fd711c8aa49a8b8ecf07c6cc997a2100649a5c757bc95c738b5bf0c0d567915a8f8c82124072ad4875dce76c41bc71269cbfeea943009aaaaa8cee8b19743a519efd95e5404eb8ad95af75;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12b222beba20aa59be115a9a9984f444dc40565e43ff02695336bb2c44da04062bb3ab98f29a08c2c93acbd7ddbad4c699b2d3981005405234908996fe8d1cb459a79a6f355790e6f7ef79619d55e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17eaf09c8b4b1aec21301224f22e7c5249364b23320bf5fe951017b7e1a0ef2c32a482019580cd9bf042046dcc3c2b5422b55a74227eface70b3f877ffabee834e18ce5d5fc8aa25236688394df89;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18908afa8596c16855d759506d5b353e94a76e63028846f88c952df9f68ce2e7772ea13c6f1f992d461bb6a68519efe8e7af1e3a0ddd2959b44a85a86a3a1b7d82a5f99f0974abd21d32338e9a1c7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdc5a03a94e12d5d6525358a35bf5a8c9daaf9af95ebbbb558d6cb72df484bf5caae77ea611c0d168de4478cbd0f2cb5c0b7d824ea5b02d84daceaa448e23299ca2bab3018fb6a78ef23958a3d118;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3662c6e18d1203c39a16b0e1fe8da1d5499a0dd17af4c93ddd22ae886acab62a77672c55a8714a1044765312c37faff49841559ea565c09bf71d27d929682e150dc8f05caaeda3449eeab91cc710;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h214406dc65744a378fa3fb06885ef08f425954ffb77a9a6d65cabf1c96f8ecbb84fd512a752c37b118c332bf18d4720442b16eed7f3b1fe994e20493d9482a32a8dd04bf98c0fc45cb9caa9ec24c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7f49af8e881f7512e0356578d40b2d92354a00a3c70ebce38b58cb19a224c3d28ba8f8a70d565ae1c64e1b847dad58aee7efe5f797f10a6f8b485a7a6bed8a37bd545dd369030f42ca7bf4d71e0f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b65b0fd2ea1b574148a9f6b66b17c5eb5600f24714161dc8125e6db518019f0c6ba9d189e821f4e6928dd48ec2e8589754294a1d0693f1f5edf53b36651a99b895922b03206baa3b937b93a88f04;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a27a3f350dd8c014dd313c8b10ffc71525790a08dac6e3f2cd6a3055da6339da45a37fb3d28b8a15d8a7e9633a0d0f51ee3e9cc5583a65b8b5cdee1c08203c5e16a344c7af9b53a6bb722fa25764;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8bf7f94b21b93b79366f2d9fec66b5b6858bdd091251e9ee0450a8b69a225798af99ca6c3f659d95b68595bdbf2d0c9c9af2eea5e188feffec4174f67eb0a6e0a5f84e21237ab7b2b88bd7af19c4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb5c35ac013ac15fdbcc55fba17dda9629bb4e234a713216c52a4551470aa4c668b1268bfb52e482b880cd1c39f1ac8f4b85ae8f80280cffd6ee1e5e7d81a45a485861a530c381be5c0f91de41ad1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha4f22b7abf219236a91d73b4fc21396975500745e1bcc6738e64da7cd654d04a9722b77ba8394ab63be5db829f64a5b9c28f3edc7643f690dea928b97900553ad1925ab4554d8c820a675435a57a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h929de8ddb4a15f2d73870ac7c75b2072ef401e1228bcf338a695e3958218e9f7076eb84e9c57e9263ace7d62c06f7c5601bb8d43472ba226d8c076e900ce8412c18f4adf82215c664927c78ce234;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1901205d2df85933eaf9648775edd32cac3a598cccb1ee3d400733af2b2760f2ac31d08f72a814517515198ea98151d4fb97ae1eb5cf8ab39924209ccab0c375a7b1e2b4a082e42abcbf69055505b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1095e9a654bfa25e9f88a38c36fd1cd51730cd16af6114265c2dff3310d6c1b98ff4865d751d1d5f18cfbf4ac89da82423ac6887a738b77d4aaf8135298a3bbe64ec613e9aee8d1d65f8fd2e257c6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16e0655395c308270740fac7a2e42db5b3dbfbc6075960047d515e6a699c0de6dfe19dfbee16dc29609ed8ecbcb436755a6361edc1c85b6f9259e93630141fbd369f6ade39a6b918eb4fc0bc62f91;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb5953d88bf2ed657d29f471ac315b3361ac01ee9560c583911c42b3e275e789ffd6d31e7398aae840b5ced7edc48019263151da3788d80aeb3fb47703000717254c5b851dfcf3c23e791ee839ce1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d8cacf5c1d4294d1986204cc302acfc4a8134657545cca4d917d1e285c82d4ec278595de45c43b673763c2e435bbd8cc68bdbfef8b0e65e763ee1fe741ab7113f3949dd67938d2f0f74df0dea275;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16ffaf2571204aab740bd31ce0e2efe4534d48545bd77805cc04b7291588c60e5aba6bbbe53b7427bb60e840531d9b4edcab6b0944dc4318d535d3ffb2a6208052d83e4ca712b52fd9c51d8231677;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he5c3a5259d7babe34351e7a09b36c84ed3b204c810b9975625e7b0832840234fc4fce14514680eacfaddbb9f0ff506b9179dc93e34cac6d9af390d9aa670e27dcda3d3741a506cecaf63e648afe1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h58f77f0d25b3d77fd76823bfae11b1e7bd3053040639286b6ab940e972ccd714105d48afaebf161e8c9af82fc5d8a08edc6d81642f259d4c049ff86b0d6bfef8e7d7c045ce8963d523c2902cb9f8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf294930f3717e04b0e0a85f77eccf2694551d3563858955115a7efb0a544e92c71d18d27257b3a962e1ef9b5ca44dfdfdac5ed24e8ed8894b828f2973e65681b22456eb66598dbabab30456490d8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9156db973c343a0f0459baaa9613647e7bb4fdcaa6794753f05ddd52edd10d7d8d201346ee00d9466acc40e871cda97f18907201d7952d0f9c3ae1aaf4a628a4e097feb9e3751c7a76b3c60c81ec;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha7f01a72a1a9e5c0d8f61719be766ac83bfcd3ad6f5d8e5aa1eec2ea8c970379b63fb13dccabe34dd845aeb92d589272357da348390555df727aabc45aac90c23e1eaa059f9746d1b56b94c42061;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h158ffb22f8f13a760314984172e52091247d8a991d294c812badf6ba97b2b4bbdac822c447f9b5578d5f809d03d5afd624f5e749941edf6874cec5130701fa9fe2762a4a8931c2556ad3edeeb91b4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h140d81c728b15779e7a0ffc3ffa6a6d139456a6988f91c5175f2f88078b127c5b11defde99772f37c7eb8fcc7b00b16a6a01fad62dcc3eca6a9f9fadd1ff91268d90fa61a086408d776d26d3c468c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h42bac4e8aa67c10e1b92cad5ec7d7b358b64ed499484659566e9cdf4cf3e810939758879c28a36e307037a4298eb98bc36e8e9b5f170fd027497308e9cdc48ba2b36032209383bdf35d263df3767;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d31a694e897568b9d4c6a7056e2a2a0d0d2d3e95feed099b6f72aefb336b6ae622323f400983ef9a2dd0bb61b2f6f8138a789671b2d77d16c12e461954ed0104533f94167dd43c9f18f6befdceaa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2db9cb13a3d5736fc735dbc4cf1393bb28194af207ae35ec0eb39b152c16ce7e844738299ec5d98fa535f11b19b8994a3a97ec1cdab673ed3a5716f8e08c9e4132d5b9c7bf65b72698a438fa64a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h141abe99896d3b52a2b258503bfa8c0c4a172c5d66adda53ad60af6fb19618299999bd37560c77cbdce91fd86d51efb203c1f2b257435feaface5edfdedcd5de0c30bff8514a43f3137e8db08c07d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17ddb510a70b40f45e22ec2201b85f487da8fa3cb38116b5b27b5380451da6dbf6b876bd1aee5eaf1ee8d52b5081fe60628dff8cb7e4d67ba1c40ea585c2a52b6891ff41f294680ef8ad7eb3115d8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f103a1240e20b160096aab24e8ee59804ec7f464b0d4ddfa4aec01d1ffc00ab408856ac5ee11cdc6881458111fa1f9311a02b3027cf05ba2076f9436ccf0b7e0c64ba031fdb8933d424b244c7f69;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2b30785db19ed30bf45c508f7801081308c4a229a3c928ec76eef266b22a7fa15e1168325908b82d1646d8d3ac9613173cdb02367583e20a5249121e04d6d4a8d906a3c211338519fafe45c3b19b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdeb03540f07fe4f11fe100963baf609d826aa414a3b35e7b7d6ec9d4a126d914c019532f3ac0e5779642f5fbd4b4ab4fa4aa99e6bda514954b760a8c38adc88c015fbb14ec1a637e3259739fb6f4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2fca4314def013ab2ee1b3e5cec85b762b0a57fc70935aeeb1b18c1ccdda5c972444e73022c9693f817e7658dbf56ad9c910de3b24a8866291ef16e30fb708dbb9bdfe44984c683e8bba3c90c268;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h141d98939c146f7b561db427240c2fb31bec047b642fa3793403451dee27420bf13899dec0415ce77658ab363ada93cd92976c96eae7df95b67adeb45e01832e38f5defe05d6d6955d079fc9f8ca0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7bb29a92d96ced2cb0d52eeca02182feccdf944edb14d828ddfb5e09ecb2e78617e4a9d5a4b7830cf80f3514e13c672852ead9f2c36ad2626758592e58c3762bab7532d685b32a90a794394c24ff;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha4af821778d059157bdaf3fc960599c987fdc5e5712fa843f4e7dfe4abbafaa3b02c45560bd64b3f47974e913558b3b3003d75ccda5f07951119af28602a366addc2e7025fc704e3c6390a85ccf1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16e1dc3bca4c507fd6a6c334b5441741cca7a7908d84bd906764c3914543c739190b40dbc2f029a1b27c757ba7a4280454fe3db0959f951831eaad3f17bfdb4b1a085bfd2c907c9970ef0c480f783;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb9302ec8c992c5d5b8b1715f956b56de9e9a32d806dbdaa54c2693c56bac43435945b73a21281bda5a6ba9e1eb0ea720674de1a9cf3ca4e5d86b64beff74ff57ba42af02798da3d3e638f8af7091;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h82a0eefb59e675d6fefaaf991b7377a3571650e5175e6af9bcbafe890450c3bec37dd8a3bb9ea92dcc86804785a5b0d3b50287f1d295110fd46f223f27cef50422654080635c98ebf19e091ea3f3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h36c6d4f7b1a089b49688b667a24513a9d753a7a30a9b5a05f469c83224d2a7d37f940cbd5b6b2ce8b02757f27d6f624c1dd54470d1dea618387e47a6108fbd48700f1dfea5ea088cfaf013af55a5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dcef34c19361007447a8e53d49d9f8b94dc7c444e9d573f78def1a595af7c2b0f52e0e37dedc5bf6d5792219f466648f43a6b8d26f53b03fdb4162a053740a789c26d37936768329a9d759a32754;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c35a8315d6649ec3d67ebad807a4c6b80613ccc2a3bcb9f26661dba35ef76624a578e94c96c8e5a069614127fbaecef420860ca2914d1852358e33fbb097c06a949cf3b85d2bb89d51db4a3cbff7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e1250c578f08d5e665efa59f68c9f16d5c6dbf4af2473006d23af266ff701f0c850bdaf147dbbbc4794f708b42ba4cf72d9fa5066311f4f97d3cbd9799d8e8f4c27fa86b44dc90fa1961fe89fca2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h25de70670ac438560bb2e1912f5a69bdabd15d51ad9d700ebb7109ecfbfbdcbf2f3ec7125abfea8c0a74dd18c82e544bf8785c8c580c75e9519c7203eddcca3091d260a15f14b18bae2c74088214;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6521c00b39e39b8333cb3476d56997ddb70596591995586158a0f3c3bcd4a5297b6e77c819828c744144637978bb63cd7d8e0931bb1601cff755c5d6f120fe1a3fb1c04fc38251b0514672e3b696;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1be871467bc56e0032340f456ee886c999dc39befb023c9c317764c2213e14102eec0c68e3793e0174e507ce398f769bca8222e0422e01806db43ca6b6f74929fe2449767e5bae3db306e98fd83b4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc22d5e05517362c52066ef64f63e39bae043263f6c05c379a335c80a4f483513129dcbd761173f4a07a915832228f31a7c53a2bc9a5818cb8833e75731cd6ee98f7ad7432fe45ecde3e380ced1ec;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12ace9d70ffb3114c6d4d4c04f6302cb23dd14fde0879583bfd0486612e14afae5ba71e34ff3c9981f901889da0053a9beaf99a2e19bec1e8949eec38024e5c39d29f3a9ebecc54808316e8fc6967;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1356c597a607fbb49ce231f11cbe2b5bdb6d66b1bc1ee3aab632d3d6c1edbf9af854bb221370f5e3abaf0e21ae3285f358f9f16919c60a5dfa069571f8a808a958a14eba93ac7c0ee5c2a231ca02e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9e6b9be135897bdb5d22282aafa7f6f8968e5c58c5d69c91c658504d9aa8915217d9c4cffc0c4ad2a1513e8b9872e90bca60b8534f2f1a18f799d787c36906697fc8968c67f0bdda79ea10340be;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19bb296601979a7795a61684c3cd7ce9f2f1cf96fa40a6ca34398decde5e7fd69ca8ee9e3ad7acd58297d9eb2c873d327f8ed275da0d7e4c0a10e28c5a66f120bd0a5e84ce3ddf859ea5b7243c89f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h508ee0c89866f75d284ba6c8a1631514ec1d4581daef7ab57e9164474b82e4052c95d325e5194968e669c3d07a4d1b45f4a47713d4d291815cd4f70e5d666d0d0ae10ed95096fb7e31ae7b82aead;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a040d59d70e3c8fd7a4ec90c763210a17a03579a55f1747d6e34e41a89400c6eb99f60461dd321651514c6f09ea5b3b77adc5584be99a994864f76a60017b5db7473cb1d587374b68d7791447a3a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1427d28ab11fcbce811e87b911afe00cd228af4f8d1d0e731704db81df377607a3b82ee097370366ba9dacc09be68d9c7cc25244fb34781e9293d25f060124ba96bf63a99becd063bf36507b393ca;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h25a6ea39711567ddecf9545f2d93742fc6d50c7a244c7ac382e02c9a94f6ada35f174be2dc62ee026cc2d24566d6da3dc6268052ce8028e9202391dd70a247dfd0130d762943c2bc323f5b7925f9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a52aec2a8897abff1efb6ca257c82427c2db78859569338235c822741a1a0f551f3907ffa425a5798fa773f46ec9e44f2ef505e8e5579ab8cca07391882d0588e7430492143bfddb5fe0422ca5ed;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd9b29dec65c449c9e0ca828ce413fa60e2918d235a9054f7b30abe8d8db3510de376a2a97350ad0885444d77062cbb30148146e468f4152a8bab458dfa29701a128dfc552e7000841c3131a04f74;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h43fa51a944226471b62ed8c5302799c12209f6c197ed0787c08ab61c583e5cca8be562f34af1963caca0e8f64fc5fa59b3aac84d15d4405bac626f323611d3846f9ceca94540fe08de78c9271a8c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e4f674ec4c41b3a208b62fdbcdc501e90879194de14e68c55d39ef1169fed75a07cacc8892f05a3431916369aaadf3f5b819c4f58ca232ccad90080e6d014966aa8e0b0777cb6a5b74a0bfe5e701;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h170febe0b5a80cff11248928a54e53f1f1362024c6db699a7ceb01aa6d2e39927365d9e8f3be2cae627e9e7e6b65f7663bc830d615fe74b979b8de828ca52dea7743b597db99b740de0b40a4b7ba9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd7e7794162aa6f55732bfe9a9666f19f87da0c8ebc8d12afa9fbf89bd98311b8625a4b575ac15b9f4daf24db231aca902a6c4f1c9768ab748fd834f92897b3abcb2c1ed2da5e2379198b05dd90ec;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1be923b08dd281927f08601658b22a25eaccbb24e89639c002608807c3e863d6169804fd4b92279f758a59550610e27cec6ef2a0d562e8d0ef81f307f520e8b38b2b9f12918d27684dd8e32d7abc7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3ab17b4033d725caade4cfb79ba1b4c62074d03b5103a2275edc0e33d64e28a2a60c3e62bc3c09457fc4cceac44294e1641a17740f6e6ef2afd6b82994b1bddc27990e52905c4af31bdeda4f507d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heb5833476b3a289cbd6f24b0900806eceeec9cfa4906f14e637d75cbe2596af4bb3a23ac0954db2518d6a7987c9e2ae087984d00713e25c2cbd59b04ef184aa92e7cc3e914500e74026b71e3b2a6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h113572c33b8ff721733cf27029e5043cbbc8dffe32cadb33899bdcfc3e92c32b7895d64fb9a3706359518ff0bee2b8f5bc1b747fab5de82e9113d8cea8be7e8919fa9b37f482ee0204d660fea1c7a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5ee86acdcec5895d2f99c205bb9b961ffa4b79ba88fc82cb5e747e419a1ed482eefec0e7699e98c3470ad24b20168d69cded51e680cae155b329991e126b50edd3cf3a9d3c3e0b30e410c8d07bd4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e8c8a0b5b10bfd39aefbef29a960bb8c93601a503763cc47354c58d9bfacb1b2136190fde9145e273ca2cc70320ae97dea06d8029a732ee58aaedd555673716b8ab5e72dac7e28c4c41c2b73e39b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hec5c1cdb111ca20c8dcce69e4cbbfa7282b5f12db47672f2e552fe7d2107e906038868984b123cfdd22110e092fda3cac820f7353d9f95c4c1b79f8745248b2e4c1dd6b361e911466f084ce60c02;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h107fa76c94fcc7439cecf7498c01a85d7d423dda5280dbf3ed8008c55baa7900e0ddcbb5730cdd597d34504a20925aef6a375241db0f042efeb17813eae2e93cc23ed8c1ea2316ebbb75067808dc1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h727a2c46b5e58e3ed6f46df4c02335a54bedb067a0a7070c73d95774b4e1bf7d63d3c0fc23d0b853d75ca08049c3fee92ce0f8817eec379d855f2cf95705510316c44d09781fe1870e24141412c4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b7326caffe13f3222522ad2a4f33d5c734c22510a5eb5861157efa309d10c1d3db8cf1635482a6dbab1aa736af572e671c8abd767b84cbaf60710c77bc1f5775ed664d8d843603b0e58135b4294;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5686f19c4c7258ffe478237a2155a24b81bb72fbc45c39fbe3ff6a317dd23d3c8e8ea21e4970859631d627cfedc7b9d408e785b718372cac5819112a1db3245f2c1cb77b24b9d2e05cb06510673c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hed5144905d2f8170a97988bd9240a0af750c3d5248e80835e4df706bbdc93ac7dc18642d8cee254112356e077681807c0aa0812cef3107922a4d80a853cd587d4333a4331764a13dab792eab5117;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e0c7ba02593c9b2f1b01ea17e404bf638a01be36c4e5a0bc226d31b6db40e011750761d785ad30153fbd0e41a87525cdec09e8fde8b5a3ea4189a40706158c9024853161f15dcec2b3a91624367e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h83eac528b3bc9ac3aaff5237ddb55caedd29f8642eee60f22b911a1738c1f32c377ec44c2696ddd1fa4e6690e89fc75f7c5f585f4aac2f52e6e40e66a83c33d4e90a61c6d22e5d055cab327a90ca;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha86dd9e1b6bb1cd6349fe9d9c760994910a7d744030b512fc16062d7d0cb56182c8a3a74e6889908f05dd5b9e002ecf2eb994e53d30572dfd0bfa8e10677a75ba2e31dde1feff0088c6c124a442a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haf62c231ba5b5a28daefe624f90e17d9679b2625157a4d2f9c31a302b4bcbd432edd4195a861e0d11fe83a89123eba1383d856e75e304a3612ab26b0561d99be8f1a01a5e85993f9ea9fa4fa0117;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10e777aa12bab0328eba51ea639a36761e5c4990f007a9d9ada19fd4d1d691a7b1d8f74d931b9640c5c058a8f65037480c05ad17e0fe0a8c1d6e51a9644ac46c0aecc019f2e7a6212aae7283b2436;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h78927494bacfaaea782f331981730bc874d9ee74f3575edb323469fdff23857da652fab84f008876a955398d26b3d44466bf73812ab046420e6aa2c137d8b3e26c793b4fa62058b183e206a42068;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hff7ebdcf049cfb507b9a5a41fb2b84be44de4b8c6983453d93734386a3eab617608e35937fc4c6fa66c00c677776ecb48581020ed802c0a71128984ba6a0f09ad67d7db5da4745d6b9e8e5f60e78;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heab85edd1710aba14649c2eae0de9079f952242ce67208ab5e22fb02759b916887a6ca4453a7b2ff834abddd79516e27cfb5d07f1174a84281337640eaffd094a3e2f547d0234d6df1c109fc958a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb04002193886ba34ff1606c69a3fe1f9343ae3424512bcdd04613b9f3e525219bc870147a7cf690acb73a7febd398469a4e3f500745589c2e92acee672b4036fef30d22502ba43abbf96e7a49b38;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h641cd23cfa8699cd2f92ce42d29efc53439d5fe5fd7321cd41fc3fff0a053c09c8c7bad41871c35ada49369b0c5a64a027b0a9cefd2868bf719713ac3d4bef29d45352f724f8ed8ac1ba84eaeb7d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1451763e958a451b42b1db1b7b5855beb6f4a67287e393e96aa4757662b98d7c709507cb347323a384809db452bc2a48168d2f725cfd396ad42d5f0db5b4233d347a9f4ae394dc053de2ef00c099f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h122b002cf958d177c471ef3ee07499e2e3d09ea5302005322fa2a62ba114cfe8b9d5d03fc4157efe07cce596c9f43867ed159ea44ed3bfd90d2059e3f11564b6edb55871d7d731876c81257c7c8e8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12049d5463652f561d190775e67d04cabe0de69b836b931a253f702ae5a1a09e1fd4a322213dd528f27ae0c2fe91d90eb32a704b72e4ed8dc78fef5677fcb367f5db37e529a2462599de8c62384c4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8e120b260c108589de82cf283da706b732e5534eedf56ae05c0784737377461206e1d7a678bafda9e7e45aaf9ac2f74492f75001473c1eb70d519527729bc7ede704a426b3bb319bc544bfcca78d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9192ca17a633d10a2d6b23bab56d8a07dac2d930801b4444424989c9d24c02498a84375e5615d9dd3773535f080b3a5eb67eefd9080eca5de7693cf2c5a38d182373cc627330b472a8ea52aee84b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hff01451eebb8e23acffc72e27d585c824e3f140ce6d0215ec0be1dd1feb4a28714c7b5ba26941ce22d574f1743559a2cbdf447fd415e8398110316db77dabc4e7f6b6d206533ffb87a666a1b2a07;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12b7d80b6c1c42964334e4e791184bbe09bd553484f93b78dd6a6e5f9725e3ec5fa46f34020c3b22d44809716b21d6e004423658a8617407a6697103d3389ae0a9acfb6ce864be83ec957a1cb869b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb2ff898f601b107b52d1c67594093e855c1b540b5713b3d5fdd035f0da9e27e421b01e64f215ce2760d25fffa6d69e2e07e740d4030cdf279159f21aba59fe6a71201513ec32d0d231fd5fcdc99c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h124e7aabb4fad2e4196de933fd1b3ce1781176de5aff696e6713d32d597342e16045d0680abf4112cab3f85a3e3f3313cf153a3b0dbaca55f596a4a7ad5e9bb2758b31725f85767592c3dd7eafcb5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h61fd93b2807d6219e6a1fb183c9918b1c130eb3ef3914b3f687186ddff12e1ac2a1c7efd386f6104bc46c90e0e793438fa0339f563ccc2e11ba938a2ab88cf155b6f27cf34d1b95288bcadfebae4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1229d87647307d8f18d3fbc51c965fabb823274ed40016f0b0f7a37af9f789421d493d70f13edd222f3ba88e44238e0eae46222f3fcf7f6175f2d6da7106854657452662d59aaf562455f20fbd35b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8caa5e7cd2c4fb3f2ceba6d448c6e1a6a8c5a0c978c38e285017a0a8c148b9d06628dd4fac16b6e3aa770d2a16bd871d792328c341ad5f4b4714dcc0158fe58e9b7002fdb1d02b0825260b306c4b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h411b784844ab3895ceeb8cd69a7a3e3bde93e25b918ca508a489e2b73ace765da66716a8b3c02b69dca4b6a54fa1af7a862e1d8e508bffde479518737b190167346b5ff821a84fd283df84d6776f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9553ee5d4784612cc84ebf84e49ce298480c34fb132af5cac0549f7e549b7c693d5f2d1a95f5c174d2186648a712c73d91b4589e6d4b72944d065f0560daeacacddde971ce46e28505dc6228c4ee;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h40b977d9f92c5bea311d909e5c92c93782d6ff0b7f6c6ec3d63e0c10060a47d68f3b24cc1cdd05b73d290f55f64d59d752d65f4c00687370aafc0c83d6410eb9eff0ef130c4f3249d34c3859d55e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha690a85b37d4eafb973b2b966dd34a831cc05294ef47de3c65a5c2d17b91015ebc5154148666d2ef9b8fca8d31d640ea49cc9aaa3d87765f6c3a43036af757c396171f2857a26b31649492b9bb2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16ea53297da9c1bbc33524d7468519646748dccc7649115dd21dc7660063ca75abb4bb74e14967026202d0fa8387d2b660a7b3ec0a091faa07f4ba3cfd8b070abef4534635de113d1f73fb622a5bc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1baecc4e0a768025a88afa4e0c71e33bb7686a091fa278fe6a8fb4804665ccfedfd03de5b5934398e62a1265f4f0ce0a01d1ff13642aecf4c294a50f65ddd689ab6e6a8e1d472cce749f037302cdb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b230ebf0b0f64672177d7abc8717a970574d79ef8017a68f62710185d97d64d9ab08950e993fcde79034c8da737391dc5a3850a45d44664d9e874f967901f860b2d4747be0bf7fb22e5c9e0d4733;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a679959c265c25141cf5fcf8fd525b7bcb7dd30bb16965364e4cfbd8db0eeb1dc689eacac5801f9255168ed7d0edb290b0ed5172e7fcbc8d14436b3da359885fc2e7bd99a00374e5d1796bd46bb6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17e6f77738173f83bb1b8178e18928413c50dcd2e4d8354842e925cdadb1179736a7592cc46b59cd939c2e60e43895dcf3cdc2132630ac55bc3230525a0b2a4aa9ec150c93dec58ff1f1615c2e9b3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heb4b5753467e60ac99f14b0631db382e7b8cd4214eed3766dcfbf76dc36bbe6c18575ae1d5c9e8ad177c4a5bfa1b34533ce296778fa9ced4e4e339b3a4a8d7a17a5c2a022c6d5d58b02da2bf4c4c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13a9743f433dc833bd65a9d876d778faeef0a744d600710781d84561dea567cb76ea96bd17afee72a4530bfd8a76c0585e8166a288b0f6ce702bead0633dd3b4b3017d3ca3b38123899cf1a74495d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd758d8627db45105b25e2a02152d316cbbae93bdf561362e59914c61aa34feed31c661559537703e70ca9838629fecf3800372822fca41da11b90fb886070e7fb448a49c56f9cd684e76f7fc8009;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h96a0627989f815a66a4015ab21ed66dcdb93d7a630cdbc40b884d2d45fc76bb12cb7c8b4596dfed1368d2dc37aff6269ae573ad2a73e147d7a56da4aa4cfe2eaf9682021f079b64edf4af0d5593d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h97c1bd3b73e750e078f0800335b61d66f0d3f172641f9bc2d8d5557538dbc028747c3d945649b3292cb446dd8dc05e1ae53e7fe278fbf094b4249b044bf243e9e73958124b30227be47538d3f2cc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e4acc509a0006c163c1204d5bcbd9f2629567747cd95c8357fd14db062b0ea6557890a0382bb8eceffc639a18d923ee184c2f77b5cf09e566d2ba702cd02592ad27ff906a589d8244fc9fdcf9be7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13f295e9ea68991e47f6418b17b5aa1173311c7ecc605a7c8314c9042a0f488b955c25a4c031a6f56a5294e1468ee30f54bf17578e00d23f559d74daf790a2dfcb0a4844b23c53e71eea981401834;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16076f5bc9a9abcfd5585ae1d29418bdcffd4cfa4ae3714cb38364face936f0a58e591a129fa4eda293c2c12917a07da9878f3faccce7c4eb278f9ee8492fab4b74c4c5152ca51267c7fdc12b7d1c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbc2bfd4b7e3ed393c7126f7b75eedd6fd28dd578c6678a35c896e8569f4252f561cd6d7b9768edf5f8df20eadd25babdea9a633980b0a55f51f9c327d25906f4f822d6d1c10248f779c5c3052ad;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9194430c6b9c342eede803011a4e3fe2882483ca8f466ea49dbb24d0402747b3057dbe3bf12d96a3b338b35159ea03ac1b7d29a89a169bbeffa63e757bd2d4294d6d7f02b7a60e7c90fb19910079;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf5e7624b21e3e245af0d578be1ed80ee4a395e1ab6ece879138f4bc6e7afbee3331856133422c698c25f2f9afc93d63fe1950f31c28697de4c6e3b91d605a201c7f02037ffdcf4dbcb80dad924ea;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cb3ac21eec75bc6f068bd64d5bfc1b03a9e3c70a8348b4508191b544e74ce644f7125d11b0ffdf7a1126c54e8fa3b73876c25a9b427e843240880be95f75c2a1d0e4831f2713c1fe563da536dd90;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb2eed3eede2d8c4714cf07e45ace0e823128f0ce215002cdda4e2aba2f8ce1e434e8636ea6d1d5745f786d496fd274a33f9999deb8fc9715c79c2d8820b40031b0f1a0a4b33fea14f0945c32e138;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15afcde10686a1023640afe02f64c73e7a59172fca16f138037e5fc24184fa4e8163eed63c3a2f8e2dea8cd57a3ffb5d5f9dd7b94ede4bbae7b007d8e2eaaac8d58db0057128cc7274c560ec4a61a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h118716084a290ce5e98243d1c6237257af0d78855cce1d7aac7b96c6cb232e6d999b2f17bad4af406db003200eacfd5189e51b7c6e0fe70f3d991866e3758d5a3678779c4d0a82258e2a73daa4701;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdb19de87aae88f7cf94fd2d71e46e55b6d4f61238a3400dad63382bf66c1e6f279d9fe6505919e40f2edab6d28b262137b97aa31cf1108384104400d4fd884af3d954af406b0cc172a7bf350a6d4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6867c24d15e0a295ef1a9951b0865cbe8691d3371f7077419edb8a5845fec77e3c8c8b4bcd1a7a96b417a01fa15d8fdc68bd535bbe34f492d5f09b1536c8897e2a915987a1d409fcbd9b15aff040;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h87f5540a629052d29b4515a09a15b06e5e8acfa47bbe1c820453831c21f5923efa5f3ce55abf37304ec0da9c17d45170060a2c9de701a2db4052d724906448f45d0e5fae8057c1d436d99cb1b30f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3d90a60293f3dc6187f2ea00655c9517b122b3362f8f5a13b612c21aff31d8ef0097123be87d9ece2a628b29864093df210a0d02ec5db82e07e155c0f1954d1441180f347f576cf017b4e592be7f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19f02359efed0d8f0247e9f4b47d23925b2fbc45f7a26fa4a847b87257e67c68cdaed3a29747de686ef8df3126577621e0a94c7d75960cb8bb29ba426579092b3359e3d4e44c6b053a7b67ab0e4af;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fe72b3e3855215d2e330af10ec6597ea0eed5394137c4c7675a001385dc4ae83b48b4aff0c7a73a4f345cd4eeaf1c661b3be8e579c5ff064928b9b90fff0ab906f4766fcfc3c8bcc51c489b855e4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10f70b70e84d7744366bf6fb04c8500d74d3af467d914d30f463512d39067c2c22dcb47033bb3d54e0cd9de4cb377fa22d9e038ca204c28d1acf30b2fb784e881b95a15ada4f18fba6382dd6eae5d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cf4e78e0457383b003ec109d008db8bc2527ea5b508be4a90395aa2de6a63ac90791482b9a0f54458924bd9b47f2901430cae45745b0f08186287e53eaa71f75f9f6b8f390b4cbbc46610c2dd95a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7fa5eeab64d15d91d5b16940e48ee01694826a8666d832262022dddaca9a4ce5c3ab35f54e3737053f4cc7866d722b2fee12c193d8dc966cc73ceda6eb2690b7362b8decb55967bad3a1a6b394d7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14a0f2e3af6b0b63f5c15a47dd2a8625173c4ec0822b540e6454d3dd171eb978a5677ca05315085d8d477d9b435be45c0f71e0ba54ea167ba63273d7a1c8857f15f41f36f7d6db4e08a6258bcea04;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11e2b5e742cd2c188daee37caf4b50991dd9c0e3d11cdfe934f743285927c878080706d4f9be86c79b8a467cd202717cf0f98d2e4adee7bbac29d179a5a3333fa18ec0ccde224ce94c5ab4de25ab0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd7345f9f2fb1e4ac78b355681cf4694cfe875d60c07351ebad366788e54ecb557270cdf3223550a97f39e814e2f4e8f3f2351d1eb6f67cb253af807cfd0e8dd55acbaf048e2f32901ef10d713e4d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10480b2ae073ed7eef01be570475f55fd049b0d576a351e921b020d839fa6474586c8df28dcfbc854c6b1bfcf737b441503e4c2c32b09f1160d15d35a17691e5ab3301868f45f1c194914a3287561;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18a7bf06400bb46c691814d5f5fea06129376f4405ac6cb38627176d18200e7ac1f6be296280302130e29fde53b7b6668e2b2997565a18689271e96eb88cee74e27ddabb89a9aa6ae85c948c80875;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h164b427eba9cca4270447e1a590f65aca810a2a1985ff25681de0d81eeeea085b50d615f01cc00fd45e8b365e8467fe2c041b7fca04a213c40e21d69b3b7f9acee1e12b2a5e476183947ef63e0939;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h28c4937a63b8e7dfa44fc118bcd93c9de897fc5fd44927d5eee3ee7f4a65ba3c768561a5dcf0acdddb99c049a8fa90c42a6f46c4044a1fdc2b6488b6b2a4bda616b947c554f8da03b7dcc52a3887;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1caeb7f658535652c3a131a1884ae0042298f2174c12ac4caab2fddb398f424e4965c66eec4a34656971c92440909e7949e99ea68a7d869b99936a0ebab401cba2e82691b99af1619aa80fb006231;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h93784d8b09664c241c9cc5bda7624c76fe82b1bad30d6dfa00415fbd975ae01502df64bd376a2b2768b3d7d1e7493880da8f2600812351524cedb373652d67677b2f1f5da65d702ba9ab7086818d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb5b47617b556578141ad263dff8bc7fdaf7444bd81fce782edc45e487884d3ae587733c16774f97e2fca633326650079ba0bf1365d3143070725b595a923e3dd394af716ab67649bfaa182d96910;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hae44b17015de0402cf2cae636a96b614b89344823c7473f78f4b5e698f82f3c3ef28758e050d8c015fa571af793c2fce24f45089f72c83f3ed600caa03cee44d1a973faac53e0515d5550deefcd0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h165eeaae24b6f8c99e568a2408e93351bf6207c9ed80fa5ef7cc3ce88d11d8a301821978e64c5423cb8ac9206852ad442a60cb198dddb6536af65e40e890bfc8db90a670ec02c63be4bb9a495ca66;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h62b4a340759d89d023f6bb29e510a7bc27cdbbc94ba93b14f4ca3ab7f93656a0d934766c68580e730c2682de033e9ecab039ff6141cb9136fd679238aec6b71ce666d65872837da929d81bfa9bfd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a8223d382084b5ad45c7818418b4ba854521a636fb0ca9206ac159aedc6d97449a696ed6061abe63ef6dc28027c9991219330401825eabf6ebcf3e6b1be2fff19a6092f139e8a3a5ce8c15a7a6b8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15d1783cfe6fdc0ed34f2de8319dae3002e892954ee8c390b40310651c7849dace337b84dbc766ee4a0f0e37362017bb44dc18bbb17e43faf9fb9f46f674765fc79e22ad9699d984d85ccf324244f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12b9d730b9734fdbc49f9562d97973f117b1b12c6ef6122088e758424296a16b32a95b958f4fa21535bd9fc95fa5f437d525d8e00a90752ae1bc85cc21099b98c57c12024bcbe3a6ef497cdadc55c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17b2c128b4ae88aefd3a4a4d9ce105b9afe6c8a84b21a90b3beaa92d5b6d50eb94cdb80db149a913ef8877aa2b465697830d9a872aab2ccf38c9c6bdb320686bc24da5992300cf445e17f38a8f63b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha13a7c9ebe54e7805dfc8db4f4e9301ef285c69e483a56600ad4824d95d06a016d2e4cd9395225bae5cda0dd01687dfec4d7086c92ea28c160c0dc87c475c224e1f6ed8d9ca0bd5178167f5745ac;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f354f95d3359b424f8f9d7074de17e66fc53e32ef9046482b3e993b10d23c1364bc37d3bd4fff7857f61d78221ebe4785285dfb788d59389c1ceb04e4dabeb68a2f042993b7b04a52319d63841ee;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1058accfef467a22ae18ad146cc63499f4a0cca6ad38542d4b2aaa2775e96695e580c21f998106d53a3b6d0cd90ba5d39836c25e91790842809a4a54ebcb50614dbdcd05676d4ac67280e7fe462a1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7bc724771767c291c83a1b7367132aed13bafda6f6553cbba50cd5c71c9cb358a3a355531e9f15c43d38adb562af29aeba0e8374c753aa2f2cfe66eb1d1eb0cf7cdf4fa3ca4feb5e48c25326513d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h68f6f7e5795863ee35ee9d0f7ef69806c2445c8a65677c21299b2d86cc2c1eedc5b8df3d852797581bcd034e778d5f50b515bc9da352f77dc3d0cc7250932909cab2553bd0f906b2b028c621eea2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h114c46f577b1d3e7fe1139d017fb71f9accc6fc13a41019a1c017425350b680288f45ae565c96c77c395616698ac05c7ac4680fef9b60dd5e1a4d7c1f7e6a327847e5ddc586c2b726c6c96037aea3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4c5203ceb0a449b17920678f1c63f304db20d42bdee5b3f262f23f9604a76892b27e5bbd7ef77a791bd20dab223f16af73d440697de307d78067ba1d851793de27cdc40bff28ad32c7bd111af19c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15475af272926570831bf35af9d0ce16c00d7d36ee0a2f8576fea73bcdcb9aa0bec4b2878be848c4789172fd3ae2e46ddb5a70a0694e58c81c299183a62f05b8c9d0c3778d56ad93a57bd82e44ff6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h119d2ef903f019ab2f784a37698dcbf50fced3d3ba9a8a431a29a082396f7da4a202bc2f74dcd2383d87101740a828fd7e3c52c91e2baed4940ecd05f1c1a4cdb1f709ea4f984882fe80e4bb4a049;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h96a666907eb773076281d6005cd8dacd253bdf63367e71cf921ff2f384947ac4a0ef2fad16f05f6bcaa54ba3e89bc471a6dd97f54d76be0aeabea63a883d0c353ca914d11a0bb7925ae5e0755055;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10f546384832e47d4cc3045ebf8c88d791fa9cef2cdc970128fe5eb38534bbfc8dbd1ef4d3febf6121289f1ca82cba71cc6b912e28fd1733f68f9682271db4337dbb2b425f74c3a0d24cedd90eee2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc65363f479ea20e092be5b145a14ac43c65d4d1f9ae37d380b823473acc79227b7436a38f12d2d3fb4cfaed0e9cee6d4ae51cf1042c0713d7729d4641c2761f6d615ac2de589cb968e531f3d568b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bff703829760365aff1ef40bb8b8c51d72223a7455d74992082ce7c31e524866b0d849a1f9e7e5aadca05b6b26fab8a5fb9c1165c9c897739c41688ba5c8f6e0488cc74cf9b529f2f1197ff09328;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5297b26f2b6e9ec79b08b13077bb41eb0ddef560b0fb7059e0f09e509bc93c2b1aa721008abb28d755d528b799ade64c5294c55645974164b6b7a961af21ab7efcd77e6c8acec4cf91ef40480a68;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7764fae501314d4d30be07bf8a994281df8f318ee7e496604343f075ea5fe0796258dee55861ceab91f6eeff05fa9733efc91e3e49949fd983f8d0340fdd4a8e172fe2cc39d0167156083cde8abb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcbab99e8919828f2ff7639b72611e3b13da94eee837c83f59abf47f59a368c167fa4226497c1e68620807f00fe740ff353d343c9e93dc46638c22451dade32d5c49acb9c860e83e63e6993207a09;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd83844846b47350e8261974904ad061e09caabfcffe0de5a6773456abc5a94532c40f22f863313c85f9f4210edc9bb917aa57e31fe6e93a1439389bd79e1354df1a6c5a2df1e1a1f595108e4bea1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18ad8b033d94a740b281daa4e95f332e6a26ea8649920357efae733422cef3aac9af40d7db92d8ecfbf23cef0a2677b1b9b9c743cf6cdc9cde516e1e4d773929a2a6380a32c7367ea7ad2e8e3c2c2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11b5386d6f26c65bd28c1db03c27b500b5d059f2c6f4a171d9484da6858af31924c1134f536cad1dec498e93a73effd31100fc48a2e44781db598dd23f20023026702b2c81215c51708373f9b5fb6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h679f36b0aeec171ce9cdebda6aac4909ac144ced16b606fd1749e9faf827472a5bb5a14a120e155928fb79deb55868e9e04ebb884546cf89e4005067f8c41f03601172161172ba89126f1dc097b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcdc8563f3ba309076afe760d685fbc11a95b216e7aec429f6d849bc859905a3c1d44b2c8383080306be8466816f28466a3d46993134772addfcd93541e197c78e52d6b938e58ce208a27d1aadfeb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dee4ec7c579d864e2dd85f1e7617364ce1ff661734476392b27307ab08c3d627da99fe6ecf7afc7b9333dd26ee9b7da7961768cb769aacef19afa377f27b92d0cb3b1dd04460f97df3d47bdc11a4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6f56107ebf9f68f1c97cd83149f7d0f0e8e4bd3268940aeb3b00722f3066d955541d8f75835fcf8b8d3e6d5ba0db9e6e9f8b1387d6145b084a67d50e21d2037faa6045be57d555798838a78cf5d1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4aa93ed41d3939f47688ba633103640219257ffaa63c58a1d886309e8341ae90111db244add3667ab3767f36c5fe0eccda85b1f8c2082786f4cb36f137cbd1e2e82c1a8ef53b70d28db7e9bf015;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hee5eacce2e26b01b275f91e0ae74bc812f45af7d8e5a1023c33531a431a4053a9fd6fcc96b8c8204000e58037b6f5630f9c1f7d128844ed64cc441508c21e363e9f532e6e8c97fa384d1995b8bf9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h71eaf4521436c1e137b47718a18e9e98cb7b6cbd38b385c74e6513d668f3fbd92a2d6fff517012e73ef0b0404f73940b651f1b44537d0ecc31d2d87f40867a0b95165cd6f81750ccfccfcee32d23;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he0b121d96fe2bfaeb0d36acc0424f68f51918878485b946215554a5da23a5adb1288bfb7bc03fdb1e899652d813b6ea7a794ca1798dc360d275790faec379d42e39b4af7028544f860d9c81a670d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1120197bfcb80526481de93235c500628a03d4ce1ac042f9f7b4d3fbd060b8558df08cbb17dc053287f769bb50c6b1742f67a21f47e3796dea92137275000a911f19b1e81cd5f10d358de760a04ac;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f50b053a19a763a9bada118f3647f7166bd4c1c67c8ee8f29cde470c41b2ea52ce99670115a04dc485b5f3e18234171671344026dca28fd5c5de5779ccb42f6dd2be39a9e5f9793eea365c01bc8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1072e930c77e60054cb0b1027e406206fbd25d46575145d3a6cbd91b0a09ac833f5135b6722cad3409fe9bbfd738f800ca2ca86303bc43c93f09360cbd92331877fb0641788919d2f474a2519cf6a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e3efabf179b6650c6321fa35d4794ab7424a7b12e8874a4b0ad7c5be60a43812dc06f736ec4eab28353ac00f40d290e1bb549b50808e5200bd2a94a9f6845d70f1158761489e86a4ae94d5dabdc6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdfd325a3462048fa6b76c6977a0cb979124dd0eae9c89eeb0a9e95d340671b52155e899f10d185166d06f02e1dce8ed199e33ea34df74590bdee713db660b7aaf2bef25e64fca2e6e309e84737d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10d1349ccd94b3c2a4f69182b89cd82aa1cac66ec3bbb0175874b0fae0ec2e4046b2e504e80e53d4e9894d6d0736ad3b7e1843695ba326c68c37cd84673421937b7df75a789e1083245bc6c730e4a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3443274df97e44d774e18a639a4ff6c028af8280905a375808fdd3193e45087fc10528fab21d6966d85cd616c4a7a7f5dc6fdc10175b538a9373d27f4e5825db089d4570be440675edfeb65902b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ff7311169aff8763f0762ef460b9b4214e368c5c7d856d2a8c7539b7d85d5dc5985d69f6e1cbbce8d2b9c547ea0f8400bad03840a0596fff7e920c02636ec01978697ff749bd6e68bdf05f350e3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdf9597fd27a32854cf4f8b21e4d9a751bbb73ad7444f7e2dc5f8b83a65470b7b7a16ee45af21530e062da2f10dfb36307904f7bf68242254938808e0916be0495f18d59d7d68e2f4e75181c01818;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4693a72e291c8868f5c82b0104061769ea3fe83e654672b0250303763e7054a59e45cd02defc39945d10f38770ff51836b0f342e8f8d1be1f2726d93ec9cae5745557d45b11a510dbcab6b02452d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hac48ab45b10169901e79808c491be2b02a33d6365915cd4a6e4bec0e024f3af8051f1b83c5e93a446161a69cca98e6805ef60b2fc082f8e99f0eef6dd21eab0822e94f8617cb96b31edbc8e85c2d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15478dcd1e70ab7f675b0ef039d679ec6ba93f4ba01fb167a3b03e89f888cc4f219fec50eb500d053f567c984fdedd2b20e86074012ebc653d3d0d2c269509eaae29837acb2229898edcf29071583;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17786eba068e62b68279008c8e7340c4d15dbc7d77491e5d2b4282c4037c7654ee398a6d9c8353d7599c693ecc40ae1637d1e89c8c28bb99bccefaee8f7dd45125d903497b51e775efa17ea879957;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc04914fcf5b73d3baf5b9165b1090b4d413ee2ca69fb82ab2e0ff9c28c1467aa245a707d0ab2c05e20c21073ea9dde0287f28d0f9b27a8f6c85d555825f1954efe39c03d71b38bc578a6ef8c4a9d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h180e4344eba4456d1e1df18f1741315d277985087c51939059e90cc396a6652bb85a2032750f0ad1dcbbacbf8c5d71496476a31d4a81937a0bb44c0e5063fa797165c38fe63149772b4253528c82e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd8090e5f27aad0ab5fb0cb2814afb72b13547c18695347cc2d90ab23f4e87edd02b641db3e3814f96f93eb6d714fc3d820789cead891436beb366225ea6fb447eff4279c0f160444a2aa4c467de2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h183dbeb041b7a0f03551b3aee49db670729343366bb5691609d2e42725f8a3354975e13bf4f04be9e36016162236e4d4d2f52811422f3bc19ad528d217dfbb4d1062366c9e2d1aa26bfa54c2585ee;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2b2e3ca45d4949ddd5f1ddfe0eccc1cbdaac5e35fd29d49ae87cfc336bd69177118be9aa125ee2809870c4f4cb00dfccd780b00f141f22c00beb45f2884ca79a53ec011161334ad64bf224f041a8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19f406f8f8eadc49b60c2fd8a50c80dd3359cf370cf940c3fb0fae1e5f4567e79b49a1ebd21a9d33a1180916eed0a154facb2fef8b2dbf0dc7dba0635b62f3c180c01654ae8f52d837a248dec018a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1153b2c905473ebe895f2210dd69e4177f17baab3692428854b4368620d6117c505afae41b8515011da980b45c6389c87cd1a7a2387f017685d0baf2d57434453a4cb0d8bf27d2d05867c6bc90a3c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10ecceb8d1d3e88db3195baf7c62fb40a583533ef13259cff4d987597835a9ff7c44eefbc1e2347d20ca566a37548bb82a51cb584744e946d93c4b978e127629c4e108adb1af9499b3df4acdf1f7f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a748971e0f3b133290bd95aaf9876a927b0ca7433fe66c431ee018f16951771dc4dcde1b719a997692b0d253f1123caabbbea5a756b6a49f0121dace26f66cab5c2fe41ad9faf6d8f57792fd97a1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h88955670de8f576cc7368f3f59c89b39e7e31992ca737173852fcc06378506e104e563e5b8e2fc86ae028a262017f5bec3dd9d3d611fe9e5b7bb8e0c7ab112d661d1715dba14c0b3bbb67b8200ec;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h107ce0c5dc5731d98aa885871f910be600fb0e93aabf03d3cc849a774e47a1ce606ab86b7fc096a82f139c545205fe9f7e982488bf9d9717eadeafb03299734195aea2082cc1eb2a523adcd81c7b2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fa7b18f7c871b35151fcadb36d66b474d48671e1e55c750c133301707ee0ecd3034d0f7911d07460352c20c79bdaf68dcd315638a4528e76a41c313698c659c414fa3ed68a265ff56f69acd84c89;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dcaad01f80c6839520a9a45375b050a9b62a480745c9b685ac104219cd4083da6874022408200ce3a6d532aacfcb37bf2396bdf5960aac8d06c78aabc80c9b4f9141b38044a521994ffc704056b4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h24fe19a10343bd122bc3b900634b68b7394e7d42686430b51b687d7e7fa3c4d87bd0fac39e7ac501097cbce503bcba267f4f3b20114d183ca7efcd9066e0b30fcb9c57d0ef9dfc3558eaaf0fcbe1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h730113fdfc151f9583467b48f7c07d56a872ff7fdf685b6e24b3e22cfb85e05c1d41f9b8166739bf145d1469c5ea00e9abb9a21f1752e09dec1814099affe92218e40b29054ff048de6e5f734c5a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ba21c4b1d748bf3d2207710575557c00f7284f1f9e69d2077fa0eb1be5d95e6145f3df774c37ffc1a4dcf6ac187f67ace11471dcfeeb7449a5ed988baf7afd64143c3942c8f6f4f12c2e154f5e62;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13806c173dbf3f7b6857a66884b8a5b273518aa34bb50fe9bb98284277f7ceec00d49b104f6fe0871569627e9b1ba6616ee7510b5429b2e137dbe50f47a75808f2de2d0170180df6f1d5eabf9547c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haa3d4b29137e16c31871b7fd73c83200f644acb6a42b97c3a82bf7537d880c991fee726de4702cce9f8fc6e52c638e1989d09a097a5efa3f27eb792b057584674c5b5b1f672781cb9b87cff968cd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bd44c381d9729adc7a90b693912271eb2a61be31eac8fb3fb3c95660f75fd316a4e0592a7da52b081a1088fdf1172fda8dcc71e8269726fc5924a3c5c11f1b1e821265fcd4960ec78821af55b8c5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13877efb405dc11116b2390db472bb9017c68889c9a3e326ba2ef1a4e7c223daea94e2ec9f90ad06ab749247320260bf3c78925bb3eb8d44a85fe2c20247503d55000e65ff2c2c5987be39ccb2ace;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1de5107e2b835ad830bc7344c83e92ef1034fbb4bcdc495976c9e28f5823e704e96b9a9c76744028e2d56be9b4dd1c55df6a0df17a6110b21f9f0bce7f7dfd5d51e1eb7f3544a2418dec3d9d16ad1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb0ea282cb75b4a898a189505b2549753311e78a42171b3cd90f5b5b363b2c36d0007981feb3c8d60980bcc5388e79922ee889eb45376600861180ff8ed764f8d12b99d2dd2f2e034bd0007eb88f5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h133a6a4de64342e600621ae198762bce4d4cbc1e2a0b1dea950068d820a47a6731273430d0534893d2eee793d789f055705f0190d338bf71fd3abb1baa10ecce25ec152c059ceb5244a5266f16e2f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e39ad33d894a836c98062c1ad137cf1fcb68722bc49907c66ff8ca0613082e9d55df06ccd4cd7886933a7f034d6bd70ca7f2c08bd32f8cdffa9af5bcd002a79f59c4327ae6b92d0ac0bb18c5dec1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd564a5888e28e24b27e1db2863437a3675867bc53e5e28e9c362c87006d17cb9a7b89d15d14334af47815e69cdce834668351689bf75477bf9beb36880f4b8d7544dc7c9deefa6f9d2229da54c7a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h91d97efa905dd8ab589957edb4718940ac1de92c3d425e38fcf8a0c9048ac3905e0da458a6f046b1f1e4dcf444a92e57c0ab804b394f06d0d86f71f0b9662739df179c42e8a8b5e89d1cecb272a3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fe8f0eaaa080cd9e2a6ecef320936e6f0c2cf9e182bb44f7d560904d783227edad584ece8bf46a9826930d0d3ebb4069e54888887102ab31651d24842bb8850bc795da326f516ec712bf6d7af298;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h60bd4d9e7cb16cddeda3023c1fbc5eb0b5e610d8762c9d067d80d578fbf05102b9bbd1564c4340a2d176e84dc502691a4d2f8a4126d960e7a00b41be9ad1c4917f2a7c4ec1fff964f727867f6b0d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h195218f6f240c69aeac4f44e13232112f6fe504cfcc2c61bccd42a10f8278a7e3339ac487d0f206ecd70e36bd970d9887cf3954887b367a8f269ed330c4fe229195c479d0ba4d9b2fcf6c12683d88;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16b50e9c7565a5839eba2fd2e662d786c6cb728f80a6df64deadaee59b6eba584187488a9c708ef4dce17f7b6e482d051ab139d5e602b17638a592feebf35ccd486db0910d216d4f59ae850c1701f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13bc011c7821d6952487922ead33d951b5fd0941f6008bdf46c3ff462b5b9ce5d768e2549d4f08f463eecd2e06a2a0fd994e45c4f3635e382af432b8fbe6ac86b6e671f96c7904bacd8760c453cad;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h761cffac9033c113940da7bd5a3e44e02e5957398c882ca83447e02771334c5d2174a81f71a620beb6bc8041db0e08141f1c9d55373a38c0023ce465e9695440b54d4d9b102858aadb378f82f156;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc04579d27f7f27d98c1f5174e27ad5919ae68eb2048badc2cd867861db0ce65ad72fab131ea2299a0829e6128717841aefe4a40c73e0ad587f373db7f5dce5ecd279d0e1b4dae6550320167e5784;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h27de13ba16b99284d93762fcad1eabdf159dc6def06cfc64901bfd19f67c6334658f26506801d2f4bed2ca9bdf9fcf1d36475d4a3647be129917a8f4b38ef2de3b88156ec3dea78329345d7c5fc0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h194ff23c73865953dd09dea6e8d4523ff9c454eea680571384d9a633b5a4374c4d44270820c372ffb64e8e844e4c2f2faf88b2f5d23951c63a1db6349e3d3628c174ce318162dad7e2779066844af;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf8c6c70fcfbd708aa86c3c19bf33331a4ed34058ed0511d7da30a346e1b3aa788ffd6f9fa7dfeedbb4abf84d11b937cbc73fd309beabb0c128d4b29282c94a3a6da7e9a85811903c2094ba5fca5e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f6dae4714e0fe65fe2f1e93ec856506921c718f3a87825bd789c5ffe25c570177e98472d803fb4e837fc309e3455bd36a55896327628b924b0ae254030351313923a2f06250f3d21e64c8ba053a7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b17c01bd19cacf13bacd186addaab959e9523b49afee8f9fb311cade06878a324e69dc1b19d9ac35ff848759ca3d791f03813d033582e56f269c59a15a8233d4930ea6c4cb47b396d23fcdd1684f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e4fad8a2f6cc02351a281ee0a8499c7c69e927c4669a6725fbcd1e6d610546983264b821c10ae226d687d5135efadcd5d00f1eb546315a92fc0c8c6512bdad7b7c2b0aadbe91ca496fc4140602b6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b562ca0c8d1a3fb9b92cd33fb0af0d03087bee20ba6580b8cd45cd94f15ad9304fcc11f85524dc717b007bbcb6366d43d536ba9c5f54c8d01bbc07510d33e36b4f0be7b5b7f3282a67d94e4ff99a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16eb5f08586b3d608d0a2aa0f6c01a6dfb17c639e857e88dc56d7081389b0a23f5c14ca023490d046af19ac8ae65d21d2859d8c100616614f3baef10171800b55cd3fc8aa2cbf10a294d11bf61913;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h168493fb66def60aef410f032bf42ace18d7fff764ab20bc88d8e9fabf7529cecaacb1a4a4cf2befe3c4342103d3ee5a868cbdb4c713ccdb2004e6c45fe72ebf2a47f62df44c4424db4cdc02a8103;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h35f598f96a05f2e0daaedcc321b49af29dd389d859c52c87d395fed2023e67d8f48923f1271607b7a69486627ad4c62c65468b2ee5b2ce30cd05e0db0fa541c5e759ddf03a19d6c908fe52a32fc7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11d324f30c266d1137f2ebb4d3e703d34c1416f55833259d6f00e1dc7dbc693bc5ed07bb291255350767c6b285a1a9b8dbafcf3a293d330e9521858f7d2b36cf611c4a5bbcfac5043ffe7892efb93;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h30e97f3cc5607de1f8af3a85bfcf1f79c012f42609123b7494147ab0d700940e752e11b7dba36390ba5dd71c6039734c359e61b641df5c920955303f8250b6dd320895f1d399d6a53940b3d7434b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdaa30711b6d7319192c7914fe3af76f3361a4a733d9bad6159436acc2ca1a3cffb68c0e0cf88e1224f07bacf36fe0e1fd15298ef1751de622bc67b7d9abe0640dad74c1864283d5e385326ab589c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6c5c7cc586bd101f714b139b1f1ee0980876cdd95730261a8089f774c66e33b5ca001a4228755874778f2a4f0418540e9dfdac9c9fa40f4945eb6899eef2bb544ca72188c9a216bc8b1affae6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h847591761213fd35cb5f1e419cdc3859b07d2851009cbe40f2b054b6e3fdad49d6576319137d5a019146e433b5a0775eba3d10be4354191c241900e477f4337eb07ccaafe78afee6284ea4d284d0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h98f374057a83aedeeba459bb0629e55ec298fe89eea84a8346c465a285b6c3eb10a7dd2842ec7523a902a1c34162a7dd7a9fb7efaaa3976c6cf9a756b058240057371d2929c1856a41c1d625faec;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17666ec5642f8b8e5e04833d594d66c339b64f6afc459eff914797dc34f36b7bf61968137b2679c94860e65508177618c5ed2cc507d74f671d2d12fd91e723f07a1f7ac46f5b5b72b37b4877dfe57;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h188648700bd952db8dcefe5edec07f65e0538512edccf0ab67e465c6f9395eda3aa67979a45971d570f15be08873d489bab15004f65fa49a59cfa2ce68f6a94f6e157351e3571315fc966f5308ba7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1963b6eec0f84103fb5fe47f100cf16b1e5263e35d3a6dbc23c09cd870bb17f6b7e0333617b40b134e91fee20a9f4225268a1000eb9d28960812895e069acfaf5c4ecdc1bf2a80b129ccabc03f5a0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18b858c25ce5f6a3e0c91a9f67cedefa917e96e26ff29c02fac7c2c3f62c55cd8515ad7a2d132599a2cf1fdea2f6e5eac30f48898352ef1be8ca8bfe24a706ea9924d148e2d305b4cf78a3fa5bdc3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d24f12d0c24e6e57572c6b533d0b77f39063c970035f90a4f60988999a54d3b6d8adcf3d5af87dbb9535245d17799aa275028755bf22979820c7a9cf3d5f7fc473e9409d0b10356c84ceb20dae9e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1652c8dead3e86fac9f100171a09c01e83d0db29b3025b34e53a53d50c04081c70e8ad12b5a197287c99b194de62f182b8b6c80c7230899124024e8471255bcc907722f737add79bea0a39310ad48;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h276b9d4edbabe5fe931ce26d8ea19455e4dd3c3ee2ea506a944a4ced579d0bfc800d5e63571bf16d44d96df7621147870864a16a16369c1bce0b6ee8bb94c0de0845963a7f19837fa3943ad3ac18;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he7ab691d7d20315a8b58e22438247aa46672b7de8f1384f356128babdc04e1e0a5cdbebf2e0536a0c70a5af74e66d9778819be409b9d10ccd9c139ea855b9266ded73f6c9dcade951f6659b77899;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6923d24ca396daa5cc682bc0acfd42e2207713130e7b5e432362c98a6b22c8e85f5b48ee67e6e58a880c80abc0384e7815f8eba2c0ddef680587b739f15944ef64954166987f9d17d7b5179804d1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16373a7da303daa7f5f603e2ae538e5f8a50a404a14dc9a8f1fd56321af3b9dd909237689919d790ec8673af44db04944cc8dd8e08af4285bd03be0d965553365555fc2851382ec962762b971d38a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10f321c0fe1abc4e5f5e1720cf2949749fd748fa951073a4d28a9526863e92bb306dd219039b6c8f8d7c9a3b375460eb86911069143333004bf55bd33b9dfcfaf32d37af63203433764ccbc24cf37;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19e069a81baa8c6ab47e74f3cfa53c30c0cd7a4ae726ae17ee3d32b5cdab8bb42ad5c8bebf7ba56dfa36e81a0aecc2d89f9a882cdb2a09b42b5a3c5b8625a4babe0cd3d25c2dca8a7091771b95b19;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ea5f2c7cc69b675350f29c092dd91fa88737a9732e88de0216d5c876060d9a62380dafcccf787c2c427f0af1d5edf610eccff24e0f51553cf39a49d509bd7b004c3e24c10b5e69f33ea33703dbdc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h42e5e96ad060c45916e1b19a6e7375a20a755750eb8af4ddc69d466728464dbf311292b14869548f0865e65cb973a2df23267ecc45b5566834dc3f76924ea2e843d240b71aebc3d926d3d32ec2bf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3211109ef82d4286f4f190cb15281e921f97508d7bd039a149e52482c80736a2aca0b4124102cd0932dfc06ece8b68dc8f09ea2bf366f24d230d1a276a80b9a3dee842522b0deadd0d269d11e82e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h54110c3a11c7fc2231c046b5017b64d026e63fe37292a604a845a41aaf94ae38aafe65e9e44b5675ae85c1a8d1d1a51008de9eaf497056807ed73bc8a9710493dfaf0f91a60f7a83e61e4a201f3d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h80adc887d5e8a50bcc233a8a94f33db208790bef0646f34446649f069ae5265508c196b94a8fa77eeeeb2152786e83abccfab9bd3ea57e5ecf5c4404daede94f156fe5671f8cb0d757cfc46679df;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8d8f1f723951cf15721af6e2fedf76f3da37cba812de7fec41381fcad38c1db17ea954d03f79f6f29b36cbfc425170f843ef8ba1b92d8fb26dbe0076f690354f1d5a22c3528f043ed18b6bf58159;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb0a96ea610abc5d890bf421abe0ea6171d131da7aa2c5198fe95871d5332b609ba9cb2b3ce0beac1072321f03a633e8caf561592d31c9e8e0b72bbe18800f357fd0d4eef8b57b33f68421bb69f01;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h73055f23deb74d9ba73538315459523e4534ee4bd43643291af72a2ae35de6852c37326d8b459b74ef9185acec7bdd5d698672be6d4b34db701b6630d28bc13e8c34b296113c27cc764d68ce10e6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h197570a2c1542f616de9a21e9fa1c359b3793f13e460eb8a974623bf8dca2c8c0867ac83f71a9e71e49da87c35fc23f40927e4cd76e1a93dc39c3a8e16c267048daac919a24e1b18d9bff1d763692;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2306f7063fbe7b099bb24b17c8cd3a15facee6eeab48c77e865fe4a3a3b236a53c9d92b56e3ac67446cdabc86dd512d91edc95f91f981217a47e500b26f7090b4be588022fce68a257e8bd9c059c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17da89285eb5622e8793f8b8ae653b6637fbc75f5c911f6f22590040de94c747ad3e42e2651fad634826e1e2ffc3f0f5d1d51294dea67b1be13664c4798160719be51252ade98453516e936abe723;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c7d94cad20f20cd12f156ee715a87454d9e94b3b25c6c7ddf803ec25d6e5f653fd3eccc25b1e92e554019be21e3d4d29472797c2ce9c2d07c80eb052dcae601a23378b3ec85617917919527614e3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17f31abe9f3d62ca6dc8452c8849fdf5343e4ddac04ebd617f7c9292dd49c744389ef98d9d96676865639881fb668ce00c6fd7dc2339fac6c1f4f74315bacf4b228fe441dbb4c2744eaf3c22115f7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h146e4488bc242a0b1492f5dc24aab5847eacce6ad7593ddff145a2e233b0271ea467a86fa8e685d2d5175249f70715077f94e4984856582dedf37b34a29751e345ef0bd168f1ff17574f85bab4080;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1172bd0dd1599d650df353f813264e6b039f2829690974fd29032fea16521a530ddecbab78adccd379a089585640bf7c9d880f5890105c4d00e3b59889142e6519c9b471dce537ced4e084f56e2d5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h180e5a7c23a9ab091e9151cb76b85dfce973cc5ca0e7b0523746a399d74eeebd6ec2ce94fdee1d28f95771c9210cad2507bd64d6a8334351479f9079f5888b711fcfeddb885965efe8b513f086e2e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aa49eafa1b9fe80df2c492df3a6f0b42889afdbb94916c62338374e0ab2b683f43bb6bded43ea4cc8dade083b5d2934088ec739c3c9e0afd1dcdf5e82f3d6ebe362a61c6f6b7285e4bef10a099b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd933131232ff2de7d62b0d5209fc92b36f6c9d55214a36dce21c83decd8f8158db81df64f5096fc88d1d160a60ae0e3d354bd6dd4fba70c23070042b4de1ebc9d5998f6d4eb4fd00b958667b1a8d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f1fcb9bd5df7d10d0df0309ca68a3a3fcc1532d3ddc60f157108fbd0ae75e0e1b86c51b28c60f027bc1d505eba7e049bce26652adc2fa27ece289d40c6faa396f6984ef872a267e753e428c9d30c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e44143359d54a8bcdeed35c51c4dabb4abbe0b1c680cdf807b88e9a64269830d338b36f04698dbfeb58324706cdda6f20afbe7cd3f8579eff4b4119853c1d3e0614e403e50ef7e5fba26067fd3ab;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haf831aa9418c6c34c5becdf50ad2ebd1f0a1bd72658586c52804b434ed0f2f6436f19475ae18c1229637e5fa9e27b02573b89a91c012470292c3f5ab485d9d8dba12aa2c22a63d185a5aff542b94;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbce5d10eb6af95669c32aebbbd4a2902e9dce0b5e5b4f565f01136714156221f9e70251bd7e1c351a6ab5a7da14c6b6344977781ccae77c035fc7908105d3907e2c48ce96aeb17c55335b5ea735e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1da388af6274fd91659eced1d9c560fcf6290741d4b427ef773645a8c2bfff9eb00d810bbdbd0065e8f3fe700a29650cea1beb69d3e19b2cb54666425d79563e91ff965a276851c80f2755ddc78fe;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ced4d95def9053e4f1a6ef666ba8556f17da6d1b11552e0c69a46315bceb88ff60376890b7019e41c992009ce1c600ce3aab316b58654561075c36c973e6fd1a00180c941164865ca9d756ca28f8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h45a207e55a36354a929358a338becaf3b19601fc150beb2fe86d586122a6058cb8ac71b70764eda6bf718c9ec0e5cd4b5404f3385815d340652df71d7088c3a686dbd820558341bdedf13755af96;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h46935d35f89eb92eeb63f7a6895b044edfd55709b8cd00ecace94a19aa93071cf3af573ae42eedc7d06a1903cef5a5c8913d5997bad758b473b0c1290c00512ee1766ca291c532223de7a0f1a552;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ba8fbb8ab2c7cd2a482f9076dfd0cb0369e874f691117bbda071236e6dc28893e38f0997c1334b3287447f41c3ba008f1dae63ce3954492e75255f481ff3bfd76c8cb6ac5187a08e307e3b6940f7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3bd4d100ffdfdbec056e5c10df2fa9a97594ead00f32b6d4ec52ee0a1182007a6ab7ab4d3e7747d18ea8498e9e8733c37c6f10c5270506afe7e7c0b6270c005cd19f584db597cf4bd8ab372ea951;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h62ecf3c17caf703f72f87900b79c8e501d9ec73bc8d9c001c78b3bdf61012d75fd8280e23b7d3b89d364c389c054158d927b8ab4a80ceb82daf7df53b425d3cfa9d494c93daf4bee97caa8d4f08b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7c401dcd552a7fec3de14351b5e39574eb34b5a799d67effb2bd6789880b9152b7ff8680ce3c398b4771456153819e763b3a2be10995668c3ae8a3d324412eabe19ada31cc72415b332458fd832b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h40abb168b630f8a31441888351124f52beb192d1aa29920878665f91109018c9614dc951d0ad67e72542ffb64879488305c39586fb4baded6356c78bd0e4fff4386a806e9ee9454f3f09232a98b1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he1b5201b0716485bcaeb666fa3b731c887d512a2885a8f2ba940db52ea50974e4b85161b6465972f84bbc976a10cd5499d16db07aec1a474330bd55b5bffd369478072d69efa776a0e830d691b05;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18a7fdb2a638fa9774386757b7ac7d02a802d5367a33108a5fd572b6b1d17166faa84fba50ab17567e58b4abec8e5836dbb813090f6788c68b539d340eee7c335410c1c216b3a62d8a45933baf415;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fa25812b127876f854b292117c549329f8ba8ac8d71cffe800f7417f1786e097e529a54abc491e0fd1fe7f885503b33d40b556d771fe4337f0557ad42545cd1b3b8570858588f1665bbb8543c1e4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c7c6d16b46d1fee320c8b2c68edf11b7affd77f0d8ff53827b1f0f49e96eff44848dc903b8138805930d6e77dc483640fa97273405ddb8e86347a9150f3f466f6d252c16fb47d774765315636fb3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf5d73e5a9f8b7c039abdbc716ce4a99e1814e7c5a07d9aef460998ee6a12bc769541f18392517d4033f3838394ab57f36f82b1d5ce4a8cb55aa9d2b50b42a2dec2f27a1d7dae5da4f413557e27f5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8e1c9ef60cc92af71e22cbc1abc39015501b9b412b80c695bc9059329fcc2f1b50803e453c5aacfc2c6d8c7d59df95d9e31ac96a866f2c59baf0da34e7bd495980646c9b8948ec852ec6bd62d9c1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2643e74af0cf4414a3772ad85565aa2ac64207d087d64c4512614dda838b4d079835e7570ba5ca42479a2adbc6e4be0acea4780ed571ae1ec32eb8b337c920e7565e2061b87c51141bcb25d86da5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2112e8dbd589b6c76ad94ca91c3309a763ea02598f7a3ec0b0caa610c0830d7f6c97a52652e792f49edcd41561765853315525331140f5dfd3cd6d85a819a4a7393426cec0cad1f1da2ec0eec475;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h149ef5408414257ca1fd965acde226a67fd2303a40fd880f0f12476fdb450e1cb221b5a74450d66443c6b5e78ce385fbbd66fbbec6140a09a50e95c58c4acea8299afc45033647022301b39da2391;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcc3ec9f637eb81ae4df4f213b2d124decbfc247efc423b547a6080e9fe3f9153e7aa69744ae6c27f758007f4428819727fee4cc66c1b0b71ba348c35dc7e2e68a3ccf073cd56befd2fe90a45bc74;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h47f096c6d501094e24d8b85549ec13dff9c96c6eccdad929072e3a201c4191bcebde6b16f3ca00d20c08e2a508e8f1dfa434a1e1fe60b6896a267df2539ab57328ed3c76dc3bcf3c0ead0c05ed8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbcb6a49b496a0c5683fe4d00f130ad451dd9e5598fbc254b5dd54692afac5d79bfb60691969013f4e5887df40be7fbffadebd1a2c539b27f2e9b7b42154cb838917beb5bb68a250668a6e98664cd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8ffdd29c67c43b381929f614388ddb517ecb476be9f6272448b909fcaf8f254ff90b5ac3c06430dee39e5607fc7575d767c37f3913f83b296769ff58a9a48c8377be543091a57101869e80878ecb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h94c95c25ff6767efb4ae112ab4c240aaa3ba0cc01080d2f2d9ae14fc6f0f927d087af0b6c21d4d3d8dffa58fad5853ef97a46e4b33f7455018179a7adce8e1846ce654f86666695a604936b21468;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf9f07bde27b2a21bba334458437b8031bdc37653aa5987ed66a4b76c07ae24d47dc572c167d711d547e3d7976dacd7713a3a8633463fdde035c16f23cd8aff7f6401210242dd470228fbbd29008b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hec2b511ab3b3665ab3a8fb7c7d8c45d680746039211d9aa3fc4159b754d705d72d7d4f1290b9b9d5f233acd9a0c75f556f984378839d286c7f6ac18f2010d46fd7e822ea3e8426a0a940c19fe9a6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd7c49f79365abda6f788ac17e91572433fa79992cd09095a87af7a848377acbda26f926a27824d9d8902e91d003d1dcd27ac2b183f261c6968a881da8b7467ce6a7b98f375bf0f7e1d86b04f3fa0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdc192656808a857dc1e81a223077275ae309fc8c98e0a2f7df4513551bf19ca163db44a6e650fecba5a2bd57433c9649c6051e25b84daf8341537edba24cd3b32b83224ccdd6d25d727f59ed9c55;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd46e193772bfb95719ae62a2da78b543c9e870f520a56e87962cc6e2639fccf3a74cb417ffc6802c29a0edfa9799baf70fb224b1182e1f624b62020eb1d2c9f79f1787f72fabdd882ab86efc22cc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1db5e08744861bfeb9448c5938aaf580b150e928300dcf2e9c6cd01a1b8683e2c0408207b5584f9652d165f2a138367f69df0f653d49288f1c3d0dbdef67a9eda2c615d77e6057fb3604e1a95d295;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1978724309421ef26c7b8be940e6302b38980196a8dabc13ce9c3af73bb192843938514c54bf5bffb8be7e1b6ccc58674f664e3b03f1453672f1b20e35f986e57b328059c2629cb325f793a432a66;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd6d8158096e779b44fb87aa0693475dab2474b9443c240a59f063dc9f863290c4219692dd7c79ae267dc92dd252c1bb1fbb5b42b16c6467af86ced307acaf9eac652faa322a3bec3f5330c69cbdb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7556392e404cf537db1730b085c4577dba13c9e7d01bb389d8be71ab89ac3f2bfc410e4cb6e9a89ea9ea54b80bd4b05a18dc9cd2f3864012f60c9846953ab656d95b85e615bf9fc5565871aa9c45;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e6e2b17346215e2ccfd556e0ed3cca59a50e0d8a57bb7d005cac60cec91ed3f77099c98fbc623f2c353d21083c1e16003e2749479558c83518e46f03c11e1dbeb857a53854446f5627f60c581df1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc31275aa5ba62a35fdbcdb57c9ff76184f63941bbe8965be27de1bf9a5d4948bfaacd9df0992004ca0a84b0aaf359edd51205bca26a8b3014e76e223fbb023390e84df8939d186e92702ab2f5fda;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb7af4637224948d5a9f4f903bf167691fba9207973941d182c54a23430cdb090be81475a8dfebf8b25c0f919e13b1c175303f44e4b2d1ea653c73bd8d64836a75e6311ff533d8bbe45dd49d79648;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h110dd39d78fbfd21b8518abb22d793d060bacf7bf5dcdca820b32f93ab55849d4594d6456b6be1e96f029817ac03bace285dd86250f6c95d7e34075ef10653b71fd00dc508fdcd90541bb1339c91e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f0cbf9845f3d0030f75f8509d5adc7a9fa2baf14e406c928970bd77386b923bef34f8870d9469d68975c594896309b55ce44afbfe8bb3213a29ae21e89ffb4657ccc0fba06471e2e2a7a1ca350c3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13ef05f38a7470d9d6c5eecae7b1577d5799b45962e42e2ee5bbd2fc699d6daf51a9f9aa7db2ddcd6792cc981cc67278eb7fcdb8fd62bc1c6e3e350c4cb70c661c82e0dba8ef37e162756cede315;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcb1965c3a3151810626500df2a68abb9ad07437ed2dd80e5bfb00c37a8c002b241aaa09923c388334c2f3a842f6b5a53f319a7de89f9773e04fef291a51db151a1a27978ce00e3cb067da643d5b7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf864fbc9b5bbc0d08df5c51fada9651b5dabb34882ff842c79a5505ddcfe374b20f19219a1a5ef3b65e1473eefa914b4830a22ac905a02210f042e635e7cbe5fbe91e489a201fa714bacf0da4fbb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17344203eb5986522326ab0aeba09704bb9c5095ebaf8d87df4fb707e839d0bc7e62449707db3b571baa163b7c096139af0ae475bfc73ab9573d417d0aa52911d7edc3bde102fd1b7f76a5641b891;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd487bba53cc289f092a4a1e8dcb9efbd0c42f917b4e1112d9ba621e42d39b5d087d24ec89f6cd366302ba856e421bf53414145209f83e809c11e1f56b3a6c17831d65e87bf09067255805f6364d5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h197d9a444f21b4879b8f325a17474cbb10d4657a27dcce094bb1c8e58f089e19d35f79901d57f2b1f73e3f1d255a10a1f52fc86c3ec133d984ee0ce42aa0c0d974fb2d632bead6139e88378723288;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcb3e43766855ec8279634f30fc79572f357266604161eba9fc99041c09622c0cb6a9fc0c5f3e83d2f4da495c35c8a29287f6be5f1727217cc170c26054b8f7164e3d7e2423031440493697163cbd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h91c826ce2f648ab0a78bf3877079a828aa737c4235cfcdd2e61734fb110e801b515f6cde4a85b57580ed894020bac99ef81311176e4e0232a138ac8a3d657559e33c0fbcf3076321b715ba3d434b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8b54fd7e90c80a8d9d5c8f12e3b08e4c9d91e9143a2cb04b0bda2e41be5ae50cb1be88af253153d6284d49aff1d48e2d4ba611e6f365d8ed0fc0547461c664db8262c863d343235027159848e019;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d85f45714fd08b8d9b3825c2b87179ad8e2762f9279cef71705968e705139c414109a78a9201fc24e2f387c827c6000142d83f2c0905a0c1b9b6555d54eb836cb61a330d2d36fff7f5fc150ae761;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he907b0e4cc738fdeda8a80bec8548d5ebf3c955e4027550ced68435afb2482a5b0d9d4f77b5cf6662160bcb7acbbe03f837ef82ee1a4e3c0467e200516001b2c17a4ea3d11d39a705446c687adbe;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14db84c86b94594f4c5a16d63cb824574b3701b9522b2318c2b30b2c31d225763277c75a49e68cc474bd774e30a834ef0ea909b3edef30ac9df2761da9be319fdbc47ebe4ba7deff7de65528b7aa0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd7dae87a1a4390e98bf29b171262ae6a31939affbb0114aca49d3731a68bb38aa9d355742e40f1b989702153034a2545723499e7c674b5a06f81ec8b81deb636661d4746474cb1e7abdb80823659;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbb9f6221e170b13c956238f6130e9cf95ad41cefb8a1f7314b3c95de89f5653f2588ca059d3e23779f3a7b2cb18e7f679ae5c95d7821c7531c657062c071cfbbc969936c6a087b9eb8a885d14aa8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h49e234f2b7996acd72821e8f57cd6cd3f5c22ad3e5f44f586d72c5eca08cc2cbc66c2ec4d3ca3649d2ce07c27e61242284e6eeda412b3bfcfb9df27ae96a91f7b63fa733679926ea40642f0abbb9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb13de837bf41ccafe80dd031d456dcecaa5dcbd407887828941325b5b2dd706a541eec074389725fb08a1d8067799ed7f613a8dc19713331650f74996f979c0c48a5277fa4bc48557747e9c171a3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h124f761268b82eea884210b614629ae4a1d6f8fd12245480ffa0a07b0f798506029b1f521e82ee3cd82d3ec1eda9c537811da0ccfb7a8f063a3e2bec9b8a1931dfab7c3e48a90ad8a9faa8bc375b1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h125a71a07bb57c4002f25bd17d4a64de7a7675e17b8fa578992805f211ff9a0f5fc4fcfb53bd4bb5ae0a0d4659a31b9e895c56f8fc71db30438d98ca30502066343ac06ddfa9ce9eade0e95284a67;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hce8417283bbad36b1a2b7a14b6488b7cbe53b1f13546cbd3acbbba5ffffa5312646abf2774ce3cc782c8e89358efb5dc2570a2d92cf35a2d592a7ee14853efdc7858eb22b415bc236807f6571b28;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f5060568eda5990b799a440adec2ca06433156021e47cedef7ce9f057d9865b58178f43962e722ce1dcb417095e3fa8d3841f0b17e5f1274bb8d911bac5c7e552215dc1f5ab8ca6b441fb22a2085;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ab2fee1f56edb21c4034d13164948ec50dcf95aac987fd224c2e602f72b8e5df59af3fd8fb7bd0a2feb339e3277e1ed3e21aa58f96c82b7f5bc1c83215a698ab39834e0defedc52e5d8722b0e671;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb3141c54684f9c898960408e273673e18ec9a67434bc055012f28cb71c264a6e130146992a331f2591cfd96aaa40d333ded7e2d75d98f3d5335651e43da91a89cfba3c273760eefabf4d4c66589c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h259c68ab7b2c0d96d984a65049d321f59a755099c9e3d4cbd9a782e49e4e696cf729e160f951ce343814a263625cb04b6f630756575174fc7ede87061cc13df8039efd4a550e8304b68d1d5473f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17e04cdb539c5229164335946899d432afbbe857d031022539600360da0240c55a14aa8b47a042d02b122c630d12a5001fc1759cbbcf9fc3d4dd2454694cad2eadbfda0e410b44e5872ab7445122b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1db66104f0c58995089be643561358330a4b24cb4fccd09575061d88553573807ead4f4a89a9660227d907ac3c8cec6249757f2fa36227868b03698232db1d498e8ac0caee8ed8205b49708dbde12;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14a9297afe1cbd94b9bac804f6f4a9a5d53c18faecf1839c13d6a587395c67c6968aa3332683583ce121727485f0658ad829e45026a985b83054026e6ce6e3305420f8421d6cc96e4481fce37c1ae;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1302a290c29105b8b10b9fe8337524c2227264a3ed409a96a1a877ad5f160b89848834bc8c72925a88aaafc7b613acffbfb02cfcbafed21e9f3263cdeb1574666d25bb185ba4b4833b3bd37201cf2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17c39eda4994fd53db52b6ac9d86135964d4f1d45397278b9313a03481d4dc6f5696fce285b6a5974dd6abbe661849e76c3585ad3358ffef54c017c0c0fef3561b69f1c9a80bccacfcc1c33794a2d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12f0f4839414f17cc19738a48af50d5e188f8c23044ff2797dd2dbb827750768982067d228db8174b8184f0a0f5c9db290dc7f3e679f441dab671039dc553de3b695ef4d2501344e1b9f55987d170;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cc3054c1e6d86c0f7036da709116c544ed2d9074fabc277f3fac594db8243321cedfb3f74bbcf80650ca43dd063db3dd5fd10ab69d6320add54b034f684b7ae7e231e89878db5f0aacf6f62cf651;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e5b67a760a73c6b67ded7301d775f40d53ea113d29f67690e63afaaab747d5117db1a3fae71a2e6d8e08794d6f5961f8c00d7b208426dfb161a68c4e0acb6ca1e5c547251d5a18b06a23ce643555;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e86eb811426745346ee96604017016fdf3c3aa6ac1966d072f0273b39d0bedce1a87f6ddee6acb85773451b5bbd07eb99501870d8f445d064f302951b70a20a49a6f9368d6c476efa01b28b27df4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8b397b265f932c127e7a563b867de70a45b5477798024bd8edfd962bc9d7a69ac4e682a573cee4f0cd092644372f66f948e579c0e8f6c445db5ec58ed036a61cdf5ca50a4ef777e27015ce792511;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3c571e8db38e92c04475e6e3dd3d9612bf4d3cde483e54db7b0495ca7db759fbb6aa585a6a06172bd2db2dd5ee182bbd13b08c24af94ea45d85ef9b222ee7806c3f38bf64a97c61b466e6e0cfadc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18627073cc385972b50516425fca97d3b029483bb7cf1474a25738fa9c164ad7cd7845c0172bad0b77ae2554541182f1aa3160c21251f300a5a700d380ed56d3dccfd7deb453a26c78605c9023856;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1512e540c54eeec4d770bd54fcb422474bf3731fdcbd576752dc68a9b8b39aa291fa171f5811a71e720ca9bfe842311006e57314032e101e09761f5039e467cf58913859920126a47f84ed06474f2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fc7f4759d2b220466a226fb4c255c75bec5c4c2ff70f7c1f74c1f8541d31a86479583ec42765ac4835b84122943edb3bcdb7cceacf3700b47d1fd8ec3d6e42fdb936eada913a97407b1f37d68af2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h119649506da2a980a55e2ea829ce234ca0764b423d37d37fa6af40b67639331b9331a33d662a1ccabae47e604107f2c24f683e8c0426d1fba42d7ac7591e8d5e5419820c2a5f7369f292c6f788217;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ab2895af2f5d2d9bb68a7063eea7822f1f128967b1d699ff1aefc53d180e5c457f1fe75f1b5ff08b7e75e4ea8397c09c067f701d30f802f072d7fc99aff08fb2900055a0782bab8838d08fab0eb6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18fbd3ba01d23d2c480d61727339a8d926ac8c7852c52a9245642c75d41beab59286cc30514a7e691a0c2a36ff8582e20eef22a85bb6c9ce9a0454cd7d6ff867571844e9603ccb53a85cb50259e63;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16794b9d6be964dd196623e525488ba705459c19e4d64f5b347c466dfd918a532bba669192b28a1466c91bb951bcce7a693fe1d62f6694024f2ac25515975a56ec8e0e3638a897a57d65110e49fa8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e939e8bc3519b6c4d9f6ae4ef845d690657f48181953aba6ce8bdc8f399a3ed4e794d18b6cb8a527b8d4a4a68ecd86e7f26350d62addfc7571575f9af1c714fffe97b71afb981a64b16a220109b0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a2d7d7190d0eb707d6a5cb9423623b45ca7f576c4870967079a0e96b458a7139fee2037a5591f3a8d4a0695c365b2b82d7746abf12fadb5f1b3842f9b395bcde07385d06dc89a17a40750af04cae;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h339c0c6a2c2b53f8ae8cf33f7437bbbc129e73751678534b74343628534bac4834baf230491541b71ed6ae50f5f0e521f76dac007ecaa20218ffb01221920d06c78d2e4122bdaaacc206c95ca298;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12c3d18244a43affe22bb0ac83826624a0ededd4edb5b50b3af919cd490e085eb206a1dc556ca5e4a8432666c5ee9cdeeefb7b3ea2005355e21da2af73ceed889ec79ecedf2b3b3f80147d33b06d0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8554aefa5379ca22193bb19ead4ed8262e75730095c9b86c546d1004d03ea2b6c02b0578d4f76b5d7e49c1b2234c4d232c87e21e2f925ec44a477988b449db68f603017f95234f3e9306e845cbf6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h44ef5d59e209496ded495900e6ce7488e32277525fb555825271a8f569ff7652c5073a8cd36b9bae765cded16d8b3b6f6e70b4ab7b629fae7895e6c18ee0a632a311a8d7a3af64f13d7ec7aa47c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he0719a2d4c4a7b9d086c921377577a0a0fac03ea38044904201c98f15152723a3453c65fe0f7b684702e7e9e426265db79a5d0fe373a498e9c78cf7ce92f15e723891ab91809c20a0e4490a9e7da;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1253ccc81ba70c0883a992754f6e2ff63458c955326cf972e3a26c2621db7c85a1ebd60957601cb7b6fd52ecc99e3bac3b9feedc1e26ec12ab94478c61199f60fc0de3e87b64106711d3f821c69a8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ce26a6dd3b5c526a4afc7ccfbcf477b00b428ccb76509fe53bf845f32f64992a1605997386edb7addb150fe7b489e0285ea9e3a033da9ef108757b6bc467f1cb9020c7bf742031c2487db7e6b042;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbb9b065e2dc371c7767b6ba4d008b785c97a309e029b67286a1bf0f14aff71b862594bfbb9f8f4de4bd3b9caf55fedb86692674d0d50c6161d428bab46323e7bc0595d750a0ceaeec2171c0d8378;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd02f8c971ba9912330492a98b9da53cc1648370eda660e556158efbfb9092b8bc9b6ce416569d622f6e91b386f68c74a61b991979798191c78a8c9f7f86a594dd0a7074bb6abb4db1a6f9c04076e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbd473a75665eb39f5429880ea27ccdcb6100cd9b9650645c7e09d177699c373f8b11f46021ddb22068a66e7fa9a6ccbe707fdf6c30fc0ba2be4ea97d54ced80b3a0fbab5012b5bc5de173d395dea;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b560319834104be101e2b836d5cee16a50f3e69f4e87cb8a13cd816819b7c90181cfa8bf129a5041d69084c48462049402efd168e7bec5c8aac3541f07a9bc26b9bc234e71138f8a668578912908;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10e4dcc1bee6b1b155a1cebff203689f391194818dc32937134c132ad56e9ca9653036a2a69f33e4a3b7cc4405337d83db4a60a0e2b31bf31fcf54a661e0076a505fdc8870c8e788b21a95d3eb1ab;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha77dff3caa6a2c161bfb71639a87798cea2ae52a49a88d296a51a4d2dbf3563464ba2a53eb5d651222cf6557a1acc9fdc65d92225c058c0ea72a0352116e6c8c35c0be4a0277b253c51d2637f8ad;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h132abcd95971e5ca5ccf72d2b91351411e25651bebb9168137668a6b84e1c22307ca88d1fa58ed8ca1e9fac50ac1cfda88229698ddad40686c678feef790ef6c061e510f053403048b992d93cf370;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h606dd78c777982e8fb5672fd00ea3ebc8ad7826ff47ec166bc37a008894bd0f6af5e45cc43d9ca3bdde25d86586811ff0e1d38ebd501e6a555edc683bdb6c9cb5d2d7764d2cfa377f84775ff533c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a200fa293d3820dba6ac99f1758a52ab739e325fecfa75791affcf3c7ac6669d0ead891adc2c6d8a98ed45eafe723a81149194720f31fd74427a917f950d8a28817c655b9e9ace0ebb2b4fc3f6c1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18518fe111dcf08278724e4b311bc75276826b39590c27d95c7de37ce51920b7cd839d8aecb042067922150bae3425e6b6a2eae29372a02caf9c0342ea99236b2cc609fee4b84651f56b45318b104;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd6b35f326b2c89aa6cdbbc08a855513c6aff087210175769f76a8875987cb2e29466fdc523eb70547e6a5e8e45c2fc36a7c89d6eb21ecd25e9e639a7feeab83a07a709653c89bf6d6431ef460662;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7df60d40b047ee49ef1acab61e5b8b4b448cc82d1aa0f7ed7ac776fbda4cd90b4425c02a5e59727dfce961bca8bb84ed1eaaa8a59d6fad20b9c5547ef0e6d73c5a429cc4806ea4e53f3b53c81e21;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bb16196588370a9bc64042f1184fd62cfdb6b204eece40dcf7b4c65cd780dc15d626668223f5b257da76da4c69dc680548d363e8d579fdb1e83e5501559a4a87e004fca42f714969338c7d484d5e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hebb7778c4a3700ee1961a67a254b35822f76dea59727c1c33860e8b9f9b2cfee7a164676f5049d6ba6dd9762bb63b68a472ec0a6a1ae6b33267bbe5e634520370b6237b6ce53f4eb1d2b995dd794;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5ac1ba75018e28210f70533d40c591faa056aec97d71d1cd9fc1abd90546527975791645d27b3878f921d09ff2d5ee71c25135bdc23d0bf827b0ff140ae7d80ed448e4f7f1f7d8693d0e7a518609;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12b883c8449efd16d9539d989ed246fde651b7d9db6aad279b036ba2b4734a72b9bf6943a1cd2576f86a59bdcf6dd9e093ca7f0feff574602c4171b498f09de3f6a6ca6329db5c1052431e2b77661;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc684632dc28697f05bebf8de5dbe84c93bf8e8221b0c3c6bd307d2c0bd3166ab74324b23322b4a531cc45804d04db68e9dedd6938b32156ed28929be488f46cca9edb4f01ff4e15000d3a51b1976;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h85b6cc2b25b7b0a03105152888a0a03bec4d9bde888b1942c282d8b5f2c95bc904d9b2e3e58cd6a5b9a1663bfffc9062960a327e6439046e412b3729da04728b3249a3e87c2f7bdc73bd7b50853c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha6d077355907b7aa2a1e28158c539279693e7e6f44b4d38836fd934857c6a009744632d1dfb9dc9bd91cb1199ced04641be42d465eb0867d87f736983b7c977d48f49253743e77078d3011f74521;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h58692ef2d9628ed02e2e3627a70bb2c69bcaa386b8839a66efe477986d456d9c33dac75890190e82dbf6975f71e59897d36f947f394fec09a744e95bd08d3f4a941efe6063b1ae3b003c5c75f02;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8d7d607e77a5bd5c48b4324fbbe12d1d5db58c7be46f02ec5b6fb296c95cd212ec13950e3102770e0afafc4f4d0da279b6a9aed6302edce7df6d0d7f44d318e518487d0c1d84924e113398521f92;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3c06f88c8f8311e502b5de1c8bb9c34698a0a12be76a45122abd77d3190ef755919ba37b8ab2e19bc4b94cfd1eea1f4ec0cf57a2c3bef17c967f0868c4e9a1aa646e72ceabb9da156d2bba4f44f1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h92ca4beef9ced8f9bbc59023b90be56089be4a58435d0397824f39edd6495c85ae690dca7baca6026e74970e7695643d23aff9684825b526acebb67351a9e6b292e06144623eb40337b0bb7e6aad;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1133d0bd8e6950a676397872259ed65db5f9eed73f37d1fcd3713b8d139946af4415d0291b091eb81addde0712e59bda56fe26839996970a7c8caa04c02ea820b897d43526dd3c62c9958df50f3ef;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9d34f0915785ccb844e11362537bf580e192480f55394fe0e9dc80f95291ae05166a5ee0797811e8a54a7fbb46979aaa9e57ad241ccb3914abfb34c2107556b72ea412d53972a4e007a1f51db37d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19776b3c98e2caf5731aef898cec52585fd0e576ac422c1a6d774c77197b33adf0fe94d2bdf393c6eb6ae9f693531503b0c321d87ad3b91c64f0207a0b604a964ddaf9b5ad3d88dbd878dc9f27de9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc71c51e326ed967c8211f282bc4101eb22ee9f9c4d5003a35eda4aca49051f0e1ec96b4012c1b27df8966abb023708ffd22b9807433175041cf655cc4f93df6b9285a7a001857f16e0b2dbf065e5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbceb242589af10feb68eb00c73582741577ce90a0c9701225ac27395ad96a82ef234a8033f16932f446459feac1943cfdfca8f5cadb1fd0d57f5b30c9e471d7dc60960b7f389b6f23c2bb20919c1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10adff4f19c6b84138261e2d2c6f134b7915c7ef37218e0ac6888477b6e06b676c5ce3913e0e79730253fc21b3d6edb42d0e8cd2cee68ff9e8e34d18d9506b79a7ff64b0db0f55fb1d81312d39d4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h181db2093b944fe19da11ca88e0453d12f3f3fa8509e8c6223f42ffb2f66e01a7f682056f033da4beec605ce2c9414662b5d69f89456d3f7c74a0301b526c9edbb05668bc0b1693ab5321fe8b63b4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h951118fadb915ebc4af19fad62fa09f0d6e13430bf1c32af0bf3a86f4499c9e21703cb61b7ad60023d66877168bf117ef9e78f8557d47be124ec38b959e5e82f28f7024b481c6f5c0440ba0d07a3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a706f5ccc01117bccade66bd6bb8db3e130fa73b935bbaf189fb08647603fb1edae70f291d4386b807a415714b6cf97571897035e6c3ea618d5fe5863fa6de18bb2bb2d99abd4f86537cce3e05d0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1978885d5eb405c1a4ff8de5109c99941e79692cf20b9e0a534f758c956f320c5e70df3747d50c9f0f6ec7cc2cf4c7a1addb2b6893b4dc8de2b80124105302b5645fca5f2b375501035047c433b45;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h191cde0a2af2ba82dbe7068328cefdfbd4ec9e19d28d8d463578f942ac970e555716095d6e164029467c60d0aa3a3e7e66b1905c647d50cab18db29b7b060688b0edb052b41283320a1d1e0ea3b70;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c75a82f86acb781b509c260dce61c175dae1db80bcf3734b1d7cc6c7516a9c744a2c1d27c5b4fc0c80e54992100f688ac49cd402a1fe5dab56784c5128ac7b57d2868589a13c0a1f156ca32dff3b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h96324eb00f7a96c8b94fd6dde393dca3036c33337c13bb9559c29a159d88ab9afddf60e2e4d4aac1f110560fd07a5ed2c982fe0516e88979bdb0a70dc198c79f0fe84235ef6d030b0cd8993fbfa5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hacf8664d9ffb395ad7cf281f295bfe9d9a421d504c06ab2e13c6c1259527dd5339b7d4747e3ac61b5b2e4909eaa932f03ab16d1e5715b03d120633fad3d447f6552c21013a5eb7101ca111a5fd09;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha18bf3dd3a476c192c17eda463b93212c585f194c128d4fb7a5bdac08925f604df53e3de6d39f3c28e35303b436dd0fe9e4843a753dfaf92759e545162e983cb38c28e43df1980b8c3e4e604af7e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h137d1640af141aaf086d08c9e5f8f29d7cc94ff2dd99d2510145cd339a1e470c365575d3009f1ccb820ddf860e43518f9e161153e99dd33646a5e2296572f031f1b6630228905fd55cae9a95886bd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he3ddad9d86996d68d4264fa5700ea999be244f7aa2764d3ee45bfa2c349aa8f1393fed33b3a0a797d29aefd7ad12f354d8253c10b16074a1a80ddf3abbc6687cc86cfa754500d71a5a8f4226883c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d0e3682bbffacab9541464e066f57e08e5cf48feae0db7f27e50d6a0ca5342fba7cfefdf4b12b235135a2287d87f682a3c784bc707c33c228de8ed76749e7c6beec41ef0716372204af786681608;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h168e0da6b900a67b0989d437ebb76ecae5ba7ef3cc8d9cdb5268acbe537ab6be375f9a0cc930c805cdf116742b8673e28fb13e80f77dac356281c50ec6c26a75a7cb636711c8cbb207a4ee55be5b0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h100dfab4f78de28c43165e34068b58ed74d3490db20a5c8023990c05317455c18c50cfad3825ad2ded015348471311cbc898a1410485c8ad4119b5fd51c933f40d0760c4283431275301cafb032d3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc7781a40078232c2b1fa255db7591d8a2383458cf6c2db46fd437d7bd544d4ac131c2fc57fce3ca59624a00d13c25e501e8e7f7a5f1b9971bc24f775bf428c1e001d1e353ae0ae4f6c13f579a6cd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17cfeb21eb910dbf864c04acdd86bf151276f4137a6f998f44a7c98576b8b1ddb623e5954f20103f35fd8c293f37006adf1f768d9fdadfa45a84ddf0f3edeb819b6ffa15458ab655a2178a087dcf3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha87029bf3027ddbc1827d7f0fc31f1166a1331b4f86d80215a5f993dfa5d5489ad3a1b40e7e5d8b39a8013e2c47e65d498f2614bf2bfdd924ba1757f4366464a3777dd54b295cd3ab802991c9531;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3cfb660b76ce7bb6b348ed5badea2f1a0dbab7dd05b56580ff6a83943b8e5fd8ef139bad9d2ebb3ca2cf89939fe719f52b4fda1a4dfb63c28d97bf8e4ac6730a9ba38256f2d153eb9b5d15f4fb14;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h59bafb6dbe3ece087910c7469f39ba1e11075e53fd3b9e9b2a99cb506e8229350ee70459b4e21a888b482a29d83c4939eb210cd97e5c84409c4793c9a046c785cc591bf25095fd4f0e4aca6d2911;
        #1
        $finish();
    end
endmodule
