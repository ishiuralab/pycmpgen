module testbench();
    reg [7:0] src0;
    reg [7:0] src1;
    reg [7:0] src2;
    reg [7:0] src3;
    reg [7:0] src4;
    reg [7:0] src5;
    reg [7:0] src6;
    reg [7:0] src7;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [10:0] srcsum;
    wire [10:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hffffffffffffffff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc8fccaeb6dc573ed;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hab78369544e2eaf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h408625756aa038f8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4ff5ff7874e8886f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2f9a3e369cdd0967;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha9a8187662c58cbb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf92519b47e104b2d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hacbb121bebb6c3cc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h76a60490497dec1c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9d3674987d35fb6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb910b4451e40ab27;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he20784200b266191;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h35a1bec7c8e053f6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h66b6c9e66cd6a8d2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he4290109c4871aeb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hab53c87f6142105;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he83f21feb6e8c0da;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c88c7b390c2458b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h827c13fd0c142595;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd044ca8ade4c6c83;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h40b9d8cb4d912352;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5ab66e261df46f2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h61d320a8ef39bc9c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h731ab3496477a194;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4ab67ec444596536;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbd7e30d5671ddee0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he51f5f5421065b8f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8964cc29db24d73a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2bb3956d4f86bcba;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7bde5fa5fd480c1a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb8986c2962d9fb9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f318eaa4a370e91;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hed1686aaaa356192;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he28fc7e27e6fe9f6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc39095e7b825be46;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1e0df645a8734b4d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h47d740bbc27a065;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7d19878d02cac84e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h45e70682b8d53edc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2c50e3511e778f93;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdbfd12e7cb832149;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h41acdc100d3b9284;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha34155fb39d4f875;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf04d1f53b76b2578;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5f018410b9d229b4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf3e84bf181eb58bc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h290a8c3e51f3d285;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hab3e0166611f1e8e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h91dd78702ed65771;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h886ecd5cb37fb307;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc28994193c32de0e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc0343c648606c239;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h606ece4372455787;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h17f6a94081df899f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h942d166566779311;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdcbcab25dd8177fb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c75594cc2f7c1e7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h46682a4b263dd7ca;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbb6cdab6c60f65e6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h25f6468fddcff297;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2d6720965698fae2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb35c54a052b3c852;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6000519ac5691718;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h34aa51807941c541;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdbd73d311d45299e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha245875630d53334;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h48ee03d9dee10294;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h57b9c72d33b96d90;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h31847e5c7ddbae33;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5054cf054e954dd6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h454a2ac99bce372d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae16f5e292fd294a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4bc361d8f9dbc9ad;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h46c97bf8399da436;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcc446a579a53361f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hce169d6fff921e97;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9454d2595490ec7b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h246acb720c63cd06;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4d4f78707b7773da;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h82f576cb6f55e218;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h54b0880f141ed804;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a10373602b45adf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h346c60220bbd7e91;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h189119c42a5b6f48;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf06d766ed9979ba4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h552e464de0cc8368;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h218a280dabbc28d9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6bd7ac1115964e1c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2e991545db0ac7f9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd22bcbf19c5ad102;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e5bfa1f2cc65cb2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haad11a5825e44d18;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1701660200e25327;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb8a58dbdeff690f5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he7558217f78fe065;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb8eaa09e901b83a1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he590823b5d6afc81;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heda2cb8cd4b81421;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h789ea41d9862d18e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf5c240e8efa3a207;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he305c2f6e82c7d84;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbea2efff7281659c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd6de96b01d98c978;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd2814c63b0b55b77;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4cfbe5a99ed1a31f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2c59f9d29f0b1bd7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h22f93cc21affbc9f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1a8177dffdac3d75;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha7b793fe3791e844;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heeb57daa8ace0581;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9689c3ac5fcda0ee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h687a405b7b62f2f8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9df23b49393826dc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h87a1c69e7bd0b1dc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1964242aaaece1c0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h97fb74459131d836;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h709b5b35f9bbd4d9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hba2dfd8a3c928d41;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf60e867c735a9da5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h96221b9137f9e57;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfa83d4aa9d9cc0a0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5aa27e64d04063aa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8763bbc4df394d42;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha948870330ebcb20;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a49921cf7268bad;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfc2a8c3ef1da65d7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9e5950d4ea091032;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h54336113060d1df8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h69ec1b9dcf42220;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha03f605b84f99d87;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc1006c101b065875;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h55c32b7934756c76;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h840b043709fbdc59;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha2e0df3490750687;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h76ac2d775d98177f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h35d2b36f502a0935;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h41847b7e1474ec5f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4248bd6851a770da;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h412c436429209e54;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h742ab4b290ee0734;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf2a0f88b17deb72e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he99f7800e53112ce;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2f06c97da4c5605c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf821c7fef9fed30;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf5dff2e6be0932c0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h35a850382a1e395a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hecfc1efb667e609c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfe1277e304fab801;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b08373ee5b63a0b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h793c56ee75be522e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6968260e66678f92;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdaa1a4d98b70dd4f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ec451e9a8c6bde5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd63ac9b8f4e37292;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1934319675c170b0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hca679c893a99ad04;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4d14496ac5351af7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9d4b3f6d264550d7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h91943435f4336337;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4dd847ec0e2c2114;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec7c17e31136a2d8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h505a3d3e443363b6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8046335af75a5b7a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h31b0444a088470eb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f7af7e9b4167b46;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d921e4ebcd3408f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h57aec11dbd955317;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4ac9c7c6494c2392;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h963ea8c5002f29af;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h21ee7932c84f9762;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h48ce49127e5c2909;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfb6e511cf71830f2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d55d0c6fa84189d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h950213d6d9a66293;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha6d21985014e2491;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h24bba77daf136c1a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h645ba467157b18f8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1851dfb0b15528bf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6fe9ef2ad7a8992a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1e7d5d2293b24cb2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h10055eca40f5b2cd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf4bfc8a906c04ca1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd58a71afb13ad57b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf51f85e5297271cc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8842e8ffc717bd11;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha9ac0475a2e77434;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb0b6753a22b1db5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd7572f4265a56fba;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he19b68328fb32bc9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9c08fc8f16049a93;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1713b0f086ebe150;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd16ba91eead34ab7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd28e19a1ee361200;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha0c02fd8186b481d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha60b5fec7237d0cb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b338eef9975a038;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h153ea9f6f854b738;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3cc4e62297ed76c1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ba57c99baa324e8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha644acf1eb82cf5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8ef046d3cf70a443;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h99c0f7ca0464ccb4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h65b4173ea0972cc9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf735d68ec1d9d47e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b98deb73cc52f0e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb236826c6b7661a4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef95849f9e494523;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3c3c44f82812e77d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h45c77df9101b412e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h53bbf98a0a016915;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72f2a10aa5744822;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he7a1acd2090ef2f8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h94a8ed8a443bf1e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5c9576b6bbf38446;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h165d0f377ca7e1ab;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5d13852ddbd08c95;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72c36d0a4fdefaa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd8fc61158768342d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc5ff4f36da4beed7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3a68f8f73d06283;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h29161da1c3089c94;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h22367ebe4c1811c5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h242970acedd8cff0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h896705e109eb7548;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcc243c3b56021bdd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h43ac22f885102449;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf68f3c7669263b0f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9fc81964edd840fe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h713e07011169d6e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h33f43871befe3c3b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h38cfa3d36e3383e2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc8cca1d37c158a9a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2a48e7699a8c732e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h45b89c057d2ae61a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h558d828b30cfcd1a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1aa7b376c69bfe2d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5db6baf28105e8e9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c3acb579a941485;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he373e3ffeebb9454;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4d1ff2c348f2197;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h92920d868b5abb32;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h568a70bf2da2438b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd42e2f7f20fcd456;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h16767c07e01d6a97;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6fb6159c6df23ab6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7588a1bf2ed36e25;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h785122729d3c8798;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h20a51fe488c62b2c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha92c6920dd9db7fa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he9626b5cefeecf13;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h80901fbf0a553eba;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h942bcb35527054d2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h743bb77d11d05c3d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha3ff4a3dd460c608;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h49db29ffe56bc956;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc81b0d1fce383fa3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h285da1aea28bb5fe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e4f2b2f19a16a31;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hece6d9c379ec919d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he7ea8317b862af4f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h93a921d0b62da565;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h84c63b2409816b88;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha526c6f86bf4b383;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf9995ed840d99f7b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3107d05d299bb75d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b498a290b1646d9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h253cb64e479a636a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he486d4ab869cb3dd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9982d90b11446d4e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h302eb6cd53b58ca9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he80563698f025861;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h69c4cc31c7524f3c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde9cf6e42a52de1c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbc615e2dc902bd88;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb9639f908d925aee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9066fd7288d26628;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h843eb48b25c4338;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7db733a760d58bce;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4ba65a72d0c488a4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h568d56941f99db9b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2a9fb56bece17f75;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7c6292f94a392449;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h69dc2f095b849790;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha58671dd3f2bbd3f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5d3998e0c6723e25;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4ea9f9b036e3d0d9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc1994fcc058e1fef;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d2095f5d0a4b48e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hffd72e511477665;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf609fe098e7167f7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3787cd50435df524;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd6b18255787d969a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h720205752ffad471;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1f39e220a17401e9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he8fd4108fddfaa19;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he6214fb911c3606b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb1ed27e5fdfefda3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc94b6ad099da947d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3570f6c464da6cb5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4223c8c08942336a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf7e66d5b12dcb7c2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb1cc6a370a7ded5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc098eaacca152e17;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9011a17327cb437;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b43a256918f4273;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcae491fb0bc977c6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h68e32672a9ecee87;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4acd9b5a7d9f86ea;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf4cbe854f561214;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h14d7a87fda405564;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h78ded006b025a783;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc44c4cbaa681db53;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h46f2a8c3fdee0aaf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h92025472e4857d41;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4b4d9d10340a41c4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3148060a9213a8a1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4406686157dad451;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h28f145b702f41a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf53028aeae37bd3c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h127636656da082d0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9bbf8d806d9c07c7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h525546fb94eaad0b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha1687a13d65df05;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd7437cb1d269803b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h101e5d09089adceb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb7663b2fa54c8e0d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h59d4b713a6f20246;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha54d5668672c4559;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2fb2eb1ef37222a0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3357793e67521ac;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbfe2c23782af8b0d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72983f71f2b53c23;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h841906882a7b38f4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6d153824c0739ed3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf16e23a832fc8463;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd1a39d463394c9ae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h26a26d0eb9142dff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heff6c395b87a90e5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf0ee94b79214ab1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2d70a82fde3a708b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc343caaa774afb62;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha5f5647ec5cf95e9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc65be389a0ca6f5b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h21d3c05b59444671;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h96bb89ae7e5dede2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9766c5b3f7ec5146;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha3cb040c2f655e51;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h58d6e3ebf40889b9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d452373acc42094;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h50860e771c238ae3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1194431b964fd0cf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h71fc1d83a27f35bd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha4434137f4781270;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h32202f78d52c65e8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4031f6bb44590935;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb31f9724f1c4713;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h99d89b74b08b1673;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7a19c03d9b9c5c18;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4504426f03a4a6fb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1613c3ce12a288fc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h66908c13f5dd7abf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9c84415f0d4b957c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha6ac332daaba4c60;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he540be6f792ea059;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h51e9f77dd6595d00;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5fe2961cad97dce5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3ed64de98fe2997f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb959202f22d8caa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h945dcfc3f2f06e0b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haad074b20db4ef26;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2ee441e9f46cfcbb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h481ef0917629485a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a8ba19ef7524a7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfc92c81de1582f16;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h624b2aafc05bf938;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5d9904df7f97921e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h44c48464f0719fa6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d02934502891964;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf93caf30d519b2d8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2fa80728b79488;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3dd9602c65409b11;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he737b9aafa1704d8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde640394162e0ec3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbe4be8e3a90367a4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc4fd134961105ca;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h440a5472d7b2c330;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb9100c2190a6f25;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6020f457219135a6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec33b3f1361d8608;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha57206f681a65103;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec53fc38bd2b6b5c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf348c66cb2019e96;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d83da51a6166bfa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h728c808d5d41fa48;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b7023e43fb637bf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h50676549898a604e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hca1dbdf0be669ead;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h590b90f0e5611770;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3c3b4dd0e65c885e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h700a09a04fa67f94;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6117fbc5364aaf0a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha922d55f91f5b7f8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb496f47e997a40a9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3b0f5134d979b276;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h46a02ec9ae6ef3f5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6df22394239a0f91;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heaa37c176a6df247;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h49f0f14902357d3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha619475586ffc3bc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h83a7f7c964d02480;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1beb26a858121417;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8aea2416ae05da0b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc12a605e4c3e36d0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7150a8ecdc861d9c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc7df2cb94775579d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h799ea1f758198f1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4e3dfcc969f6e1bd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3082b81109daa521;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcdeda1de12f8236e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7debfffbc0abb17;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5c514e32b92339dd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heacdc51556ad801;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4ec080c2910caa28;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha138ce1abefc94ae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb850d1ff5b5f12b5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72a66deeba3206fa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h419a7202f5a74f4e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd7257975f3a53e76;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3b70e9f9ec07c2da;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc8ed2d4126889e4b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2ae04a2d19e41878;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3ee0c722ead701fb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd615b4e76153597b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb45e7c80526c0ee0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd1cbcae3642aee7e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcf5ea9ed34e2bd5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc08bff48380275fd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9e8845abedaad65;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h774190694f4929f4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdbbb77f1f92432fa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd4f01051f5244b33;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3a64ebbc32b6a178;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5f580fe6b0f603c6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc573b2e888c51ef0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb6bba47071819af;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d0267118434b4aa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf908b44b96444bb5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7e48ace4b0773f03;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h169708831cc60ba0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcab9108dc9371abe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9bacca430f20a960;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc998d18f827eb73;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9171444af84f3f38;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8420a856810c5bf9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ba41162cf29b034;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha5b641bfcbf64fb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5661a9e7e075bd87;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd09a9bb06c72bf5d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h61be121676351dc2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb1b178e85b22dc52;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd2805a1dad9487ae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f074f4ab964544;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb12bf4fd6084719e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4d6cfb9ec261533a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h658def8f78391184;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h84d1ceb9a3d3424b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b861ee60f82365b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h321a132c09251e4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h918be081057ad1d4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h57119801720ea025;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2797be72151f5d61;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h505ab6e5f552ac23;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h93dc993bd2584852;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5263ea90cdfd7781;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b1269cdef0955bf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haa32394423645a43;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hac950d8922890137;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h166a1f5571a8d34f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6ca30dd763f5f7e5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcc3ce83806cb078f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h39746c3e99464bf4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6d6ebad2d7bab126;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h48625bbb24c30bd3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c0896e964734432;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae176767bee208dd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6b192548b676328a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h83653f9ab2a5ac73;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7aab06ff67ee164a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd6a4355eb3f806c3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he672ef582f67c1a1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6163b8e546460a91;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h678c9b67146a5aa7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc8966bc6a3dc0930;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd895987cf260cb65;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h454e6f3ced8a512f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hecba276a62c364c0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h15bc0f581d30354a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h68d7ae4afd8a0cd7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h28d1b913dd4b6d64;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h93d84792b61a6291;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6f20b66c44ff49ec;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc3193eb9ca105a61;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6342812aecb71621;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heee5163652eafb41;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h92da92ac84fb0dd4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h675221a635edef5c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4920aab334cf69ec;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h81f612cd616bc530;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha058856ff26bafb0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbc884984afc9a356;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfb5376897cf5c195;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haf7bb9b062207442;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'habb8278df88d2659;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h451fa76a628b5d93;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he29827b86f6f5bbf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6e23f8ba48f80acf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc1e5b05fb54049d1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4b241f97b4c3cbeb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hff9b407c5e6ec4ed;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef769fad8e0b3b5c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfdbbfa0befd48425;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb1210c75c7c1675e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee84d2259949e636;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e5035b88576b2a5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb02f4b170df147b6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb2e92d013551f9b9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h68fe89f419bfdded;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h808f9f2717ec9cc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hce6c0062a8467d62;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h63e460798fcebc56;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha7698fdd5c1863e4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf523e50881e6306b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haea65e9881e4e422;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5fa62764b3706a2b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h951e90a0d06cb626;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb3f2817b9e83f7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hce12f64c80c77ea5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf92b098a50fbb9c8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h51e48ad77a5b5d65;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h60cc16fcfffe181a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcdda797b9670ae23;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he27a05fe0a9b7fd2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef65d8ed01f9483b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc066b72841a045d5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h317d852eeb685153;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6c84bb294d22dd0a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h805d7e26ad085a2e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5092021d9c2e5d51;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf23ac5dcfa0465e4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd1968646faf2e290;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7a6fbddab9d5309e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7dffb92a11cabfd4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h95c6e626b3f77d57;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbf3acf06d3bf9e58;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h20f6400ba4c2f8d9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb4032f42e86e9fe0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3169c61bc796ab9b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6b0ade99f2bef9ea;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h549ce0ba8e877d48;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h48634267ea62dfb8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4eb0e70ef3de252e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he75352d64bde184a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha6c75935928ecb90;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb3d076e7117a238;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e41ba4878f6d19c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2e2ada9b0962b510;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h15e2015d6b94f4d1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h59e80ac0ab41e7bf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5b8cc71f627568ef;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h44983121a4e83111;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h46b8eb45aff7113;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h803754d78d4d4dcb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5100daa5f24cec00;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hac71ac8231b95d1f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h442716c31defe213;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a11c74aec9c2ca7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he8454dae4d955b8d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2df8ab01369feafc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h66c3cd76f021c54f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee8b6c23792a5211;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haabb783dea1a9ab;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2bf5da2a21ee25b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha78a14119be015fa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6b20d4ff1855cd06;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hccf7c408b176a2d3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h156751e7c3fb6134;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7d0c72284f22e909;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f2061a3f6dfb36c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1bbf30d13e26a89f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbe2a52921d4dfbd6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hff5623bb91475b65;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4f3aa681dcb82f3f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2c0614c0eb782798;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d566c5471c5f58;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2cd4439fcd68f22b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3e94fc8241e3470;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2a7373756ad7eeae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d1a6c3cdd62efe7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h17f6ce9bb001907a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2769bf798513346b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hff0ffb4f9c12734f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h68bce5fc949138a3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he39f87d84c437c03;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb4b5461a43ddc4d9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd97f39fb2d6c710f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd18071a892cc3e2c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc0c425f0d7dc236a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb9e1dce73a16611a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he0caf2b7dc3336f4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf6e0d76772c5c9c4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h910929bfd104e8c6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha5bf803c83919057;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h50e3732e59ffc92e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5ea6a10c6878ff83;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h187a05ea14907876;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he4ffbe13cdbc293;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h294602990fec7dbd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf44502edcdad215;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h10ebd17b09ff3a0d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6103c15c1ebfc88d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbb1c01364edb6e61;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf3ccba03e2c5c14c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h46b0cfb6c968f7a0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7d434446fc882e1b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc978542244c2e5d6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf31c8232f82cb736;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h47e947f021bb26cd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h732cc92c251d9cfd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc0e90d81bfd47064;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcefa8e1eaf67c77b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h416f6d99b3e871f4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h14d68435edd28b6a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h858cb0d33186853d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h58068d16968512df;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3dac7d800787d70d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbdcc71c37ffb4a78;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hffed476a8bb6091f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f63c7d7c0b39063;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf6b13ca1bc676426;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2950d6e8d585a5a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he691aa239a2fe1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf0d7c6dc53c1f042;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1e760caadc8e5ef0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcbdff64bf6e864d1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb6f8704fb0b8de2e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h589a45723ad4f352;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1bc192a60ac7a417;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1510476c6cedc416;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1e52450506ef8492;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5c6d3c43ce3f688e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5c045511b451116b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5171b37a7249e80f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7dc908a9571ad81d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1da90fd44f894143;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha2d08e26b6c07754;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7dd7ca3cc870274c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h902c193b5fea3239;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9394b7417f5774e0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h977aa16257b57245;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h70b9ca40ecab0eec;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h840137e4310285e5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha6f36f72e3d10d36;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h80887765035dfe78;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7e3d1b781c883de9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd72990928ab61258;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfa0daba93b3c58a1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h51a80298051213da;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e9696c5a3564d01;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8323a7d8d9554271;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h43929f522128099b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb4c2319e34fdc37b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4411d6a90913ae93;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcb979cbecec67579;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3e2edfd64b9fea94;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc0de11ce5ead8537;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h87e6f136dc4189b7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb6ec53f292d30ba9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha1911079b6a39df;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee160de3cb2aed2c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h401131205aafbdc5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hadad99a16c5f25f7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha16f7a47813c6fe3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee2128a38dc8a294;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf59fe67765c95949;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haaaeac33a685dcb8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h895cf69646d29a06;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7987e96ae86cfdef;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc336ea97b85fa6c0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb675380fd45283fc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb94fd119e83263d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf7d84cd35065ca1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf428f51b2006ddf3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h90cadebc0376033e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6e7430a709c5f8b8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7bdb80853971f7f1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc0e43df2ec852811;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h822a0b9f4949072b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h914e0043eb9f5347;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h29139e8f423032c9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h33cbcd4384b3da21;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4fe5077fa1e925c3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a7a086762247193;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc3beef1ef1fff48e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h853ae30b64b05ee2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1d43f8e14fc6c8d9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2256f69afa0efb74;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h37fee7fae7818f7b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h99774c530f39af8b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee3e933fbf188b94;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5f906bd0f341eb5c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbcd1e813c250f7a5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h617366ab74ab242b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he29600ada3a3354;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2cdcabd7a8455311;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcf67eb9d04d48d75;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf1e9af24c70ff083;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4ca05afca5c1c653;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc61530627f865ca5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha4f0a365d3a4f1d6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h75a81dedba5d8481;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7d44429744dbaf53;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcae8bbdcdb5ffb65;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf5cad46368def6ef;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha741666865e2d266;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdfcf4fc215737f2a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbc906c47bbe9f7f7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h722a1f92a916adc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h223b6573b0363cc8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h752e41634d53eb93;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h144450a0e041f113;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8811f867576f74d4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf8f8f98d82580b1e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha5ac863d6b0a38ee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3b9b120c08813695;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb67c08972abf494;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h13582906297eccbe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h64b9ed328a914863;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4bd873f3de8c3d03;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he6121dca3722e31f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h847a1d0196584147;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3498ba2aaa50ecbe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcc48a6e65a2e46c9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2ac4dd25ddeae3ad;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec05f390a121ca54;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h351a1362f5d3c215;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b9217559a2a396b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd27f02f0accd6292;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha48613a5c688fb22;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2005e69d7e586f00;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h87cfa6b5b22346fb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h59f02f47f141d539;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd10e25ec24b865f8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h19da28c282879269;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha72a1baee7f92799;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h790e61ae4c64b2ce;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdfddb416b3ab1eab;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h37bae053b09a026a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcdbeb314c3ff51fd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h16b4fee55291fb46;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b0f4425f57ff3e6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h63f20ff386b2d94d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4e39ebaebe30b917;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3aec28b1c7904768;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h47bc43b024d47de7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbcad63e329e2735f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7472a21c1e3bb4d7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5b1db1a0f879b00a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hebc297bea4ba3fbf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc829af028ed6550f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1a9119ec938f6de4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4c4c18bfd55544c5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2068bc5606969ccb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he8dbff53c37ffc79;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd0af7c224ac3c0d0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he345b3c8ed8cfb6b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h195e33b60fc99e99;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd514717e3a139248;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae42035c6cfc6989;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf017de2d29583442;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd5a8e9814160f7f1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha90a09b926993709;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h40ab44f3f534d025;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb6c1c0ffd58d7e7d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha80c2ee85b969491;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h18b662e5822f6938;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h21680aa4602ac025;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2728ccae42b34589;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7d4f0abf48e64d81;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7a3bfbceae9704b7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb1f38bbc004379b5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hac3287ef5db4ee2b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5f6fc40f9bc42081;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he716028ded8de0b2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h646bbe04e32fa68d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd03ac2b3c1e02a9d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h41c22e5ac4ec462c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6e9a6a8c6e00e09;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcb13b4b860a3f5ea;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b9c15ab04ba1538;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h96c307325d3294c5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h40cdb2715473a8cc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha85202387d5c19d3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e809557e136710f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d0c9fc2eaaf297;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdffe764b47c6312b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec9b20bbd20dc76f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfdcbda14a72a5c4e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc14a920fddc9d813;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he14a8d774ce1bedf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3b7fb302c52060f8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha96b0ceda862bd64;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha497af0badf895d1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3260a8bbd04b3ae3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc0709730660c74bb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haae2e3f50087b9c9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb11efceada847eb4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h80c564df8bd1a325;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9bdd417505761f65;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b77cdc6e64c5c7d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he179d786b3bf2aa6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae486661eb3ead8b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb3ae7b5e747ae583;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc526ceef040f7f17;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbfb7a38cfaaa00ff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae146895605768b5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc740e6769f3556d1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haa94057380a00245;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1e8760d5cf063ad1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'had6f50acce50ca3d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc757d634c3a1bc3f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h860d19e828a3cb0c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbc3606337c0ddad9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6a6f46fd8860ca92;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h29acd7d87f323480;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2dfe5027c1df2ad9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f651f836dbae8bc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9584a553b67dfd13;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h83ca077da18be9cd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd1912dd9da69f12b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5fe6f24baf39c52d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd900be2bf6ccf159;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcfea6977ddd54167;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdaf5bc39043a692f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc0ac65d64349c060;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h17e84e1f7fb91ddb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8dc702d3c969fc6c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h69083ba9744e8bbd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h983a42c1741c2aa6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha2f05edec207e5af;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf134bdda4faf50f9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h74a886bdebd36887;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h210bbffa85ce09fc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4b09be713afa1a6d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h40626b4341c8d2fc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h76862a59b9e9a211;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hca51434f8ffb4979;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb78b209568d139fd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb0143ca6a1a68c3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h53184d192938144c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4b67ce43b5f5f69c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2501c2b9615345c9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcc5c6fc2c3060cb4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd476c6fa239bf20f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbe869f0b9fb7c2cc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h166e2a73c07acb1e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfe7b6eb3dbd8e8aa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8eddbde82e53bd54;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1d5763a60c767c46;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h39ff1626af3ca404;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b56b5fef5207fd9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h105aa2834a19542a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3ce7485274e424bc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h351b9a61d018e61a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3227a0b406a03507;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h533d0dfce6cfd63;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h276f1f8dfbd1e8d9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbce34fc1e3f7da1f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb34900969ba725fb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdec7083e78384547;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b2916553a2129b6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9c6bad344262939a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6f0c75e640cbfdb2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6e450c9c83b56f0a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd0d3357c90ad83c0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6dfdb3a9c47bf3cf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h569e6fe272b9da70;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h12141093848be084;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he08900bbb25fd9e5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc1670f9eacfa8746;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3b905c711eaaee6c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h10a3da4175279c10;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hca9a8b32c91dcc53;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5405b9f718a0881d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha108043b03265356;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9bb3d8e66686526d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcce2e47ff4fccaa3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hadd65adf19b7fb55;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heac19ae8432617ae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6318b0cdab42c52;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h560079a8ba36d68b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9fd8dc4d4c833304;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc4d2b3989c1ecefd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8b4ba62ef1eb756d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd9cdbc9e07954583;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8cd1d5dce4d95b14;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h64196375cde2efae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6268bb046e259f28;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6efe120979e5cfe8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h84e8c93f0c424d26;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h96e40e6ec162c4ff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h69aa430ce96ed180;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb42b665654973cf9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb5189354a40dc7f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hca0007cf9600255b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf1d249afab2e99e1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h19d056aca4228105;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6d4cfcdcb24336bb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h65e1560788392e40;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5d35a2444f0adf8f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2241bc013cb455eb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h458d457478d31510;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc93e41e50d765d66;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8cedd09d78347294;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h241e28434461cc35;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3ac400cc265e637a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcd5ffd5d1ac3d31;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4e7c7380bbe7445c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc5623733a1e4b22;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfcb5ff9929fe0375;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h85583129874cba0d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h916dc2abad6fb1e1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h589354ec2b2145b3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h683ad05f9328f785;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h99361d87e5a3880;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1f0f982f7894a83;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'had92d1afe8ed7876;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he1e80f83940eb1da;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha35dfc43d877339d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hce24d61208202c1a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5f2f738fba8bc04d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb4c926bf912e79b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h672c0192965cfdb5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc521492925f53b3b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h53ef55a93ce26be2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc925e3ad8cab5a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h27f1a7323cd47d5c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h67b0804e4d537715;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7c19d899f89373e6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfc1ae1a1fa24057a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc9f32ac3a6e4f5ee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h57fa0145a4396f43;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he6e02f771121aed6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7c8a7eb9f13494b5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h891728811bb5a367;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h158765b6472ebaec;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1a61674fa4f88853;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h18ab3a61326f306c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hed099a8f2c168517;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1f5287b35c4236cb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcfac45f63478607;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8cdc7fdd1dbbe236;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he480817cc2827357;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5b2bdd3080c2e98;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4060f89c7b35689;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h22e2d9f74fa17ac7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5f680f543494585f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f17420a7c962e2a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf6ae85dd63b9975f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf964f9122b5a0767;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'habfb0d925c6c572a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfef1934ba28a3d10;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h26c2d03e65bc2df5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha9c19813e19a8e3d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h83d213440a9cd1dc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he3da60da0f88bac1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b8506354a9a8501;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha174c40b6f09aa6a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcbf6cb680d73f438;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb47a0fbb919617c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf4866528afebe27d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd64862d9a4926d58;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4ea49b39c3eda1e4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5e58d4de8f2dd278;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3521a5a0a2c26cb8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h95a4f1f88f6ae134;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4d4573dccc3b1e7c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdfd651ff9ef9f278;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h33d8b4fd67035205;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he69b7569705dcd3b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h668354b70babd476;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h55c8886180d588f7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7d70809675560cd1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h442dfd3de270ffc0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc16eb01b80d45dbd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha798e78896360767;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h78702153e4e18;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb3b52a723810c897;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1405979c9443731e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc772496bf1a33633;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha6eda68d65af939;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbe5ea72562f69610;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f91d1c0ea776765;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he0bbdf52913d087e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1fbca792880b0ab4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha1811922bb3ea03b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha52ddd74e953db3c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd615045a2f3aebde;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6231799a55479af8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hba7856b554958ff0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h542949cabe1d0199;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h450f23a775883ccf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcaadf135ff774640;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3363072b7a27e5da;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h108f084586ec822f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf2fb93e238a0c06c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9df5d277959d711;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf36d636cb1823e5b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd1935cf0430ac535;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4da9394ef239964c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8eeadfedf0453286;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdaa36cd02c4df78b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc50560d3724b8f58;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdbbb8c18591afa64;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h32a5e0e3ab095fec;
        #1
        $finish();
    end
endmodule
