module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [18:0] src20;
    reg [17:0] src21;
    reg [16:0] src22;
    reg [15:0] src23;
    reg [14:0] src24;
    reg [13:0] src25;
    reg [12:0] src26;
    reg [11:0] src27;
    reg [10:0] src28;
    reg [9:0] src29;
    reg [8:0] src30;
    reg [7:0] src31;
    reg [6:0] src32;
    reg [5:0] src33;
    reg [4:0] src34;
    reg [3:0] src35;
    reg [2:0] src36;
    reg [1:0] src37;
    reg [0:0] src38;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [39:0] srcsum;
    wire [39:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3])<<35) + ((src36[0] + src36[1] + src36[2])<<36) + ((src37[0] + src37[1])<<37) + ((src38[0])<<38);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h305ff8d56c58ea95e8731d217f4a47758c0786bed6ac1895f3e6bd2620e0e61e8d1546ecd770601a5640a6a98af752252f1e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf2215fe9d7c9daee611944d24567d3cf02de61a5f35ff58d2f42f542ca6d92009cc2693b5130f1c3bcda44ed518d09ded3f0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha95c75b9f849589705a44d3c2c0ae72f338dfebb16a629a9a3cac8ec4e95144fb32eccaf6cb500cf5a72c3dd23d5d2f039a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h95b36f777d293e7df44e6a035eab95fea7807fb68c46346079d689b2c2b32f98acbcb64c8c4ab76ccebc322d66b8df1f255e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hca08eb622de5dd03d1458e7edb2feae844ba25305f125fa572f5db057fc3adfec601109094d1d2b8dc432e2928c40ee307de;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h728a48ebe09e24a01a1cc22e028488878e52ccfb9a97fad908e758c8e7201f4de567cd1cd3424e22d843652f50e19b8f2fa9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h539bd6edea0dc522fc0b27f7166a6cdbc5b258507bd15722b4ae44050270fd881cd1c06e37229179c530fe2b6b2bb4ed9988;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hde9fa0ac7c1eb177a3dac11f2a4347aed8e3cc5d52f8ee715279cc4cedda57761c3ede8aa505cc0b7effcda3d0e000eff447;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha47707d1a2597d1ae643c47ef30c9f22db073395b8ea58f767aeff146d64c908bdfe03f1b6458e8bf44b39426f1c3ce7331b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he347a34a8c8e1dac4caa570b4d5674473b63bf8c12db0c35d42fa0c15f75b5d963ddd35036b5f2afc74d6155a7186a96caa3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he4c2ab24bc4bd748d6b6c347dfc0cfc673b27e681de210a9333c6e4eebd8b2dc2b9a2f518df34b54f9f1e80a5b8c0b58c8e8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc47fc7811fb4b8c256890aa9ed3837f8f687cec2b6ed10613c420f194ac0fabcceaca24b4a506bf71f71292ebb6636d12bf3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h87f269d0d94b11869698d1ec3df0f1de9142b4165bdd96d8510021503d92b89748b90bf5fe8152aebf4525aff659d96402a1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h86e89ec170fb34587691812cf83b4d9b545478928a9ab86f143e6f0a5afcaba17cb02a275a6ef32544ad176f3c5f5c0b83be;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf50b0c7fc408e4f35cacc3122723cebdbd554009fe2f9e1714822e6faf26bed04a695d80f8d183cf05f461d5c756b54d78a3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5f23bb0e63a36b3f14f8107c8a204451b8f765710b818d57745c20e2da1993b6d3ce3e554127b5f16d3f54d0396bc91e3e71;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfaf10c4b907e243853e391dea2da6d5a3db0a0a60815c4b75d3dfcbe0b7f2cc0053a7a4d6c314568ef0dbc9a48058e25c80e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfba37f2d4701e8d453affd6f1ed0dbf5676fa584b9063498ecab66046b7d85b64b445e6ff8fa996de207f880f9e56f8bbf5a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd7a2117c36e6f581271765c3ba210fb443295e14bc4d4d17eff83dbdccd51cc4ae03b813d57450b54f8e6dec86a9eb9095f0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6dd6828058ab0acbda1b64ccaef3879f0ab677e846797605f92f883ce5ff7fb6a0dbef252a6bc448d9adb56b67ec6647172;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h58c9ac7406b66a6d6a2d286639accb328f317c817dd7a04db5675f1d894acbbce50a2baafd012049de1c701f1737a0f88c37;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf849091f13b8026d2523534b927db4f32c434e01677eab9c260ca371e894604e5da7689a2ad64fe55cc0ee35645d78c103fe;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h55dbcb4bce0ebdf3de6952b7b3e86c276a38832b1b763d2400abb38ad594d5a1c6054fea8377ca4950db95c233ccd2a4bcda;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h70fc455fbde558fa5e46bace1e6aed830bc446667ea5e525e3f94530dbdc80e374e75f2e159bcc95768a8348f6e114139385;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcb958eb1f8c8cea1a440024a9eb9c854c83d7cc65f6021e73917059e4a3209e44439804304bec4d942940a8c4ef655783586;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4dce887735c6939bcadf2d9a50ca1ce77262328a7f031865d9b91f9b0c7c3a28a1bd2bc2781d3811ac6abd7e94af0577ae7d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hccaa0f3d33f8984a8125d58fbbc5059be1dc4736557ce4f0407b98188e876427616b894265dc0e53b5606cc4f78f68b33bc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4d6ac3e17eea9d3fbffe51fac40a62e709e95cb08e55f9ec9a9fafd4fe45faa17604e941619b11e12db96f5ae07533a16fb6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf048fd9e4dccb15c49bc6284a0807e105ace1a922920d9aaf42cba9886dfaa21649cdc29c7784dba1f9324c4b076149f189b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ce5dc14b57d46cef3a04e538a6eaf0b2e1c1d848f5d1d7de553f1d7894a20f93de285dee138293893a3342c815482ebfe22;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hef6c76556516539ede01a6bfffa9dbc09a22e7f456646c02b7c8dd081676741f4612d1ae799c7a8c605d356e372a7a11a0c0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hee0c1c0055ac9e4ee27ef8db5b4c16216bcd462447dec5da00cd7eb3b9b02f1186767b2103adb4026ba26b4a17807e13a6a3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc1f031c7920985d2c105cf05372f08fa66ab7146f5b6ae44a7b4175c4817f190c4db16cefc51147307b801afe1789d7c9ff4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he80179c0c72f9750e31a2d964882864087d45044a236424d25bd7c4f1565dea0855fd644f49b6452984e9a9244bcd733d81b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hac95d4f6f753f220a8db783bbca35a423c79a076958539b812c87c758382fa6bed0c5da30321034a70989fae39b837a8265b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb5b8966daaaa9191e1208416f1f8ed94711277a8d4f2312b7a17d9f0e04dbeb9b1f3c486200b5d1d838c4793782676ce9420;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd1eafe570f4aa03c0e56ffb22a566736576bb119d863dfa7177949ff561536c53b7ac500f5a799f17f85b03aeae1f52dfa05;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbd4aa2ec482e1e70a9b782bfbe9b33b8a4dbf74faff12b5665ba9088c6c4d9dfbbe475dce9dd7d048e92a5a48264ed92b76d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5576002aabe2bc16a12118295bf230d9bbc57d45836ebc0dc06bbb8bcc2ab8562f835bcfc6dcd38545215cd32ec6f16aee0e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc486ff91d31b87fa825be18a7b4d4532ee3ff2c09323dd4a03f1798c5ee3069da2d4e40b074d4e5ab324ee7f362f423917c4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h117ba7b9cfb1fe646777bade5f1e6b8ddc53012fd1064ec166a1e0b70393008c13c33bef871a247a3c2643449074774a141b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h11406e3fd29a2052c908d1f3fd99d1c692152432a042bf85a9a12e45c065dae5e5b1c592454d14d7a803bc7e7a183a5beaa9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h308dd49455174824a4a27506da8b34225efed36ca7bb8fc2f047c1e5041d443f3ab143ab0c6747b9714f2a3e97700732d386;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcfca09f24b1639aad5c8e236c8d82bec016fb1cf6f422a109e09d410f84bad2de70d700a8fd4de7d04e3c50e8408786c2d9b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdbeb5b14a0356c97ea91f28da9be6abd6add3fa9e5b9e36d32db3b7e769f7c5277df92301accea925bef91815a9ed7262ecc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4976863d5d75a1cdeb80a787791c4f638fae0b8445ac6392021786545432faab290be93dc7b64b3d174ef0acf9229a50ee9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h48ab5ed4a62ba990d458ca88135d95b98a25f045e0b6bf3d7c83b6d8593d229532a470aa0ac3f51d359a1ab8e132fbbef453;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha103990842ab050e5ec0779c58131284f4b2f55ad2534b576c3ae8417956a69fa7a1b5ed0317c3d65cc1acd156d7a8fb1ec7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbb7fb309e05f3aff78f3cb01f253d8a1894489d3d2bb5cc342cc9888bb06223d860a7f9cde19064fad5accba9a4826714e4b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7d31d2ec015a0ca5da4516f9aacb24b9e0ced2c1afda0da696c6e368899571b4896455a674e188f5adce97a0e9240cfb618b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hea27e3eca7cb4258e3eb2c6f9fba8c05edfd02513bd037d44eff5105baaa004ae1ddf6a8635b4008e4c2691c55328046b737;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5ff3d5e947a719ea951227368d5ef439ebc22416c755182b5ed26386aa8c4eb3ba5adfdc6cc4df9927944572409208aec5f2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3ed5343cead70d84e7279418831097d388987be5c88f5cd78fe213ed969d990a27ed1fd619affa83fa5a7abdae2228c0938c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h79044330917f98a7b51c73bf1db32e510f688a6b84fa49b6be9c70f888935c27d032012df455569253b3148675cfb4f1db15;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1d9a683378d0ef685914e4a613ea40da22ecd31d7d6ca7d9d87442cef823da55da91e1180eb0b23fa3026998b7d2c0fb18a8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h327e6977153313835f7af2bd13aee369af6712a92bae26b985db251f4d55edfc899823d8fd2ce71f8bc1f4fa13b53d31b260;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcb62d53a4b6824146da5cf67399c6dccde914e4eaeee4b1781236631132c3c12403032ffde250c3312a7d02123368a779352;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h16eda8ae8d7c1c5b7d27215bacb40496d075e663b8639dfa40cde72d289afcb4cb333c68dab4bcf9b17d444fb948a1c91f94;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9292d29f1879f62bd6126157ca7f8063dad57925ca7e398e9913ee9d6994471bc955ec3cec698ad25bb84c946f35eaeb2ec2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb2ac89d463ed60219d73060d9292e528e3fd324a9e0878654948baf7bee9c0ec31975ede34b182f8fbf027fcfcafb01f1a48;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h835e5174d83e1131c4955e5d0b68e604de7fe81dbca554c2213caba6db2bea336184b7d1d7c65264a7155ee880931fcef21b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b89ce438670fc6776ac7009edad60fe1f1e17992d729e76f49cfdec728c957e27d54a7963eac8c9f4468fcbf127fdb030ee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8fc4549ecbafe8a8d0e5231a6783b2a8b8415239361063b3d8534ac1862ed4e6c6cc36528c993b166904a7a6992c08ede17d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7836d8c3507484b78813b8939aab47f20d70fe7c731c871b943c01a1db0a67978b666e89ddd5d5d3830795f494720b29d73a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd98ac1409c941a9237220b00e89d7c92481fb59f87c88d8b0c97cf566bfa97f338d431df88eb8ad935c1d85971e6053705db;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h486c385ff3de58b5d093272d5400d0197e7ee20f93a274694b1e4216ac7be862b335a7bb429ea929ec614dc50b70788e2d3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d97d35bafeb8c7820a48b6eee0dcd873031c1ced2dddc4cf2270e595aa7addb7d60f330bba7521b25e32570310f7417ed79;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d47b67d8108a9388ee8172bd7fd94f3c413c7c2f8635588ccc274dbf8499abed3a2b3cbb3c8d179b36fbe71d84b7d239bd4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a294c6f24f5992ab1fadfd0b9aa8e950f5250477b1e8324edc77bf720c654b75d219a9263bf4605aba3a85551b3576824ac;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he30743d3e8f40e5a3a4b98f4df6e71c980e87fe70167aade90d2d61fd4c97bdaa51baf2bde7c21758dff68c1f0b8faf209d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3e709ec7f6ed62d9f599cdb88083be11c74f5078d6148012239f0923f8f8dcb08f99e9856a6efc91001ab758d204937bd86c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc85d13d9a359383465e80469b587638be68c53032f4ebf30e9058c1a5e86bc57de6cc0b1a17169e749b0c45859907777a1ce;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7f26080ab09bb85b8116b449e79d98b6a641dd71c9762a431d09324b046936c8579e2737fd3857fcf7647dc05c360957e946;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he0c31af021011952df95eeb800eb516af9288d171a00277c2912e010af07e822d87ab5dc50bf7749b6511607e8e8d1303fef;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h34b55443099ba14d4aae21739c3622bd439db544068b48dab729922e8ca1c5663d0ad12acdcecc069472360d5f4cef18c122;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb4e43c48b4673f6d96473434bb71e82d1e5f301653540703f4e40d93ec6ae51747c3a0b7740c5e80d1c7f2a7af5648165d25;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4e018bf228a3435297986ad1e7af7b4ba0cde3776fdb741aa4cf2a849e1b256179e603abc2a9d3b64dc431967cf78d089d82;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf29741ca0e299b66d04cb7cab6367e598ffeb17c01f60b084afc1fee3892d60cb4424113e790439b3a41d714a9bccf4f8b87;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec9a30eb84251dcf3e6835976711ed950be82aa5464cac21bad3ec85a830460291968d76507ebbaf3743c29b4f3521f91e90;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2e853deb6f729c3d4d1fba361d21bef04609ce1243e0db63e99865bce09cdc3d11753d89f5e86fa263d0ed06913ca6a1a147;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b6fccb6b6ba0a16d0e1fc050fc8df4267635c2b1612f7d8c4d9e80222a75da3965c127a48a5c810072cef040e30fd8011a0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a4955145e8ea22287e92ab1cef4ab7956b17848833cd0d9f311389fccf6f4618cc3b444f03f6ec04217d144bf76fa11d341;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h633cd2c6ab81d4e772dacb7c955436ef969482b72d82de1700dd854d22982b3da5e6fb9a0d6bceecfcdd49a177b9723c4851;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2973a4bb43801ba7a70a6d90ee4d07300bebf4d50aec3e44d59fed64bb914633aadbc92f0a6c53dcbfd8d8226affcd088c64;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha50f0dbe47637c790c7cae36dcb9c7b181d6b9d45548fc466495c488ed3287fe244d50225d84536257d23ffb613cce6c4f3c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h419a793b671d70e8147dca29345fb15d26d73b1667396eb36c9ee34e0583d9deb9b07f44843254a6074306cb0ba70a403bd6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8df92c22572434f41f096e55524da6fbe22c7ef2c18a5891deee7e7273b470143839c7b58d65a621190401d110d3ec504317;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd7247afc345786413307768358d487887a742ab35b9d20c64f0cecd12cf91eee6cfcca0ae653c157fec94dceb1cc3f093590;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h582c483cad65868712be1f55e7e4dbb743ab181ea1e24413361ae4a544c8153eca0c9d3109f6119f1f7600a1666c64f22322;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc68f058b84a292fed2b053f9737beb497faa0f52fcf7484808f9750b3572fb724dbd085f96630403b548aa851cef3f29fc5e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haa902b37fd92f6ac1ada2529f98840fa1577cdec4996e70fe897d623357644ec400b6003f1016ffa5b4709dc08daaf93673c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hba88093578578ea40e463df4e2e80332fb346e18ab3ff5439d49e172c9d1aba4589e8ed5340b4b7edaae9acb5a21973cdab;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5bafe925c31a65bed7afe8676f63f433108155659c06f52edaba10d796c9354cccf144f3e962d6e05dd6b6c08ad37718ac5c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae380c5ab7416543407ed20ab7afe205c6f435408893808556c5597f930d393beb9f90c64b5d849b5712d9b89391e52775f2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h60778fd4311f5688edaa1588a27d37b9d0b6feac444dc9a39750f0b23d2ed527c98a9bbf0c2de25a212a4ec8ba91c1145475;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3478d2fc7808871c25d78c77845e46e96f324d88334e6a58ce3229f37439eb4248f1e5158043897bf4f89e3f952cc2f2c3cc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6de75a5eb2af5638f16747c7133b7ea0ec5829d42b5fa7d55f7bbd5d2acac759c159b212c3638f3f38d80c35f3bd6c69ca41;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb52ae1d1bbad7cb26e3645205aa079086340d612dce0ee041d1ad1e0a3912eb91e3b8f79796d05573dab7bae47f9a53cbf08;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hba99c256cc858114b12fc8833b93c0bfeb7c6c916580912b080d636ae8db3237b289e594e42596643dbcd81753436d2288ab;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h804c70161e4e683ca34b72566a54ab84ef5c1a175687aaa598eebc1576a3be87bd6f98cfc990178d3b4ab99303d9e991bb03;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfc5f7888f2f82332c089d01133c25691716ba22b18afe4e23773beb4bea0b60b4c7e4a7bb66d3e14e22939788ce4be1a0a4f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfeedecbdc9b40ff3bcb8b2cdfb78ac008087ab6a4e28c3233350f9db657de220d185256a41f430565aab4b809053ce664b4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h23c805d6a96f42cf51b554b9b963e25a20927a4925decf8adfa2c8643743dd99997ae54866d2c2151362cca45bfc4c205bfa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9d6911d37e4c97de900e79d26b374f33d91e12c60f1dab73bb8c3ef63f548b8d73f3f3d381793c9e2afa78bb88cd0d9adb56;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1bf3b7cca5e1d0c0d3e3581616599a0cd4689f58a2f2bb61552139c96ea4b3af613818a31b1c9b1511ad72c7cc42ee8c8526;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc9587bf7ab01232dc2ec3c658d17485421258593bd1a50c4d0c939b150c85fd3fe740285c63b3b4a0b269a78c9e40053db04;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he196a5f1ac752c8129f3df8f6292a313f77c9cdc6ea24dfb9a78e611f02e266547d4182d38a78084c6694d9001366e39e4b4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb12a66196726e7501d9d5494a7705798338a3ac97269a4fe807b0e678a6de218a9d418ab345533c92cc3543741ef46aa1b2a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h78a38053d11444ea5a5a6c107a1b5c068461b2d66f8b198a970004832aa894805492473125404dd768f2ccac41a6d9922fab;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdf29cbb2d9a9264d4b69f4909daf52bacf98d1c46256f3689c8423d72059ab02e16cddad5b18d02568a4f0b5fec0e2a48cee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h24ec8fa3c98b452b188473e8d999ff54034aa975e90175850472fd562309be0eb40f41d3ef79a64de4413b3188830ebe8099;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h10eecd8ca3aff8c9f9b4a19fd3398525e3a150375380b79d3d018f1f401fb6513fd6ff15b8076c7e16fdda5db2603e5167e6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd9fc7bc6fe2834624309986186943b95aa6ad5e3f247b4a0410e4c6636d2026bade693f09b128a2d5dc7f8281fc2a95c8a40;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h642831838cb0094734e8f245dbdb55c417679c9c9a31194e1c7baf173a150ebccb9b4ffea58b0db59ecbe6b460ba18f48dfa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h64510fb0f0162c461de4fa7e991a735636156d22b95f1b499c61828e3abd19a014e66e2b1fa2b079cd9dd5e506fe9703227a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5516392b792b772a07da5e881e9e6a8e75329419d52a6bceb9efc3525a588f353206a69ffe83789aa13edcb9d3c5af664c06;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb3700a800df559fe9eb6c163dd7ee7e396cf35b43a77d72a72058f3f6a854e3dd5e654889159347f36d83dc366d28345667b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h85ce5fac3675cd51b0be34c6a122117d1504797ab522e01da9b3a672a119b1c2483d12aad024cff1c7ab50f62777adcb4013;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h68f69b09fe0166b5f8a47cee27dea25b4f74213a5825748a9ad6527346db97718efe1bb1c3682054772d5e1a2d51f3c92936;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ddb642f5e47ff4da6c4d111d9b24365acdefd966b23aa64cfb70ba5148b98932cbad513eb73cbab99b01f740cd7a33a7dfd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h61c2ac237f04b035448b06c915af9b41da034b54b83bac60baf0fd529b8b089edab7a46014ea842a2da9b472df1105465f64;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbba4dcb163c685b62d98eccbf09d2242ad3642db0686b0345dfd5d90976c4d616e0f0ae2970f5d6f192437a0a56b2755a9dd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9fc1edcb11f89808850e0cc1a97f0871c0f3bb3a196401903b029f64a9adf1be4de7ea3495e1efb8999431cef433fec1ff9b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h29b4a1a654e116dfe1a570c15088056bab28f4bd19ffe25de505cfdadee0ac0c671c43be6897e9c118e52e32c121112d1e80;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb09b2b9ccf25fb9414e6c81c2a5793f09a9485263b05daa25d76cf0f53a9d1cc70e059dd8d998313ca1bc4feb108b443c6d6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h675005c1d8a6309ceb0a484cc9ea6d740bfb96b1401bf5ee7e29c16fc6f6c16ba26b499f67f8867b53eea98fd1ca9b03a137;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha8f5cedb970ee86d5d2bce6eae2cc790161e21e32126e1f04a2222486294d1c605cc5eb8e625a40c1dc54d41df19f385c252;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8fc6e06295408ebcf0c8e48611df57e85695e2f54967f96d91b22603f5f31fffb16e433d27e091f89bd817e1a422adc13460;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbc292636cb63ef5e4183e04c8048ecf6342f4775600cbb1f1178c209be98f84498428574c85ba7e4263181406696f7dd80a6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hedc4101c22f416108c39187bee9abb6533ccb07126a01ad81a6d046ab9345455ba17ef52684388579e508089dda534240557;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1890a1e8137dbd4d01ef3645f53e8f7a07528fb38f9c9a305ce7c0318275cee712cc98b8c24f3ee2d57a7b070fdb3e8e22b3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ee2d0f005107e76fb51dd0d86b4980246d2ff27ccad806d8e676267c96c2aaedbc03819d7f54032c71223f99f6d2f243c74;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hac1dfef9b761cbcdd37a3da13d900825f1048ecf1fd37576426cff42e26f3dde0b6755a20fcbbad97f5bb58f588de9bd5292;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4d789911decfb435c98c6f2208f7db95182178b4211ee79e6d28bad22fda27d9e6f0da8dbbffe808be80c955e2172869135e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7b78447f57d5fa02e3680c2704ba4315139330109e91c2ba67fd5a78e98ba4eccab96af76ed4bbeb3d15d22af7bb5ce16ff1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9c49b400853fcb77b036159803415f7ef267b2ada51254f3db97a9a802bc0084579403a575c75604ff06b286857dc6a39d96;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7383c51b27e39305b4ba6d64fdef469dcb475d1be5aa64b3c0342cd97be0065ab0e5156d21da1c7a18cfd32a1c009f01000b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ba4747037f1ff5d88bd7444dafedcec82350753f1aa7f444cc4d1a6afb646962deabb21edf686b9525ee97c8722aa416ada;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he434b4cd959befe9c05a577fcde2ad868fdf92e3010045095c3c88b265f9319c83f52fcea563cc80a0d7f21e3098e3bb28e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h40dcd700405dfe7464374cb4783b58e1a04084f8aea91436e1fc491a9884757e74cb356be4491e9009a5c41638ae4c85ef52;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h51974104770cf4c7633ca194b86fd4460c9bef2188a9341a65450a37a074de512bc633af4a80882144f48e1c3723f5080a10;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf849f976988a93611dadeeba06efb55505dc1c9fbd6113ab63ff231d01a6482653be4f0b0b12b4cdc72f7a9cab544125eb7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb9f8a58ed65f991f2382ef43b737eeafd2efad9850e1c92d1c01c5c6d20f5020d8d1808226b95503fd056d7c81acd04f6cd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h760d34b0b98b61635d23b59bdd0d0594bae56b1066163db0d14185c4316495c9ae94a7e747715fc5e29e868a8bfe56fce359;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h80c6900d1a06bc56800381dbaf162ea0f50ba971b51b75dbcc35ce2c7a39bf9307313f68f482f6debd4d88d6fdf1fb274ce4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb72d6b78e1443a76a627fe6e7cb4aeb60338b2a5c7b8631753d0d7af27f39111ec9f76ade200a48ac98847d28d4ff6ca801a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8fc5b0b5e351a57f2584d46b2edeecfc80fd9e6a87ce5503283379a0939d4e8cb1129ad54fb94384d8216f2d78b2e0e96b29;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha0bb49ecd159891c86619e9e973932abc0b94b0b47acad712a8cbbe536f80b66a50e8cf633504f3e7b50fee34212210cd4b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8660b82c84da1508a8b03cb6eba2f649870e053f5d5f1d2e3475dc7327654eb71ea7c375f6c01fa41039a7da287812751b48;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3c227fdf89159cde825cca58e1e46b11279a8863bed5d7367e01e1f9a18eaf4d89b08a35001f5f5ad2bec5cb285f37d963c7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha58eb7512cf64e73d4fef7351eb109a3e2c954e0b700d452f5ab4769510b8cd348a62a1e3290fc18092442afd4237ef9eab3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d70b659e9563a4b374c2e35f852378d6d55a7a28bb0f49b716d6cf2e7437347d6638fd142c34d70aba3df8abe7388b9530a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he8e2e4bc464115e338f32b2064cd6fe11bda108693bdfdea9c7e7ade158652ed9abf8d104b24470ee1228533246447488c22;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he1ada4fd0108aba37c99952628bd468fcd8d82ab079f910fcf8432cfd7e0772d1d0a5182dfeb4f49d7dc791aaec77b43ec45;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a34bda450f19a23115e3b9d131320b9eb699873a168df4e6cf3eb47ec4e5d4d4718bf6d1286c7efb9f8c8142fa805ffa59e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ca98be8311fcfb96a1996c3cebcaa55a5865152466a3b584c2896525a71b47741bdff2f8d2782aa8f09d9a54972dc62ad4a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h69350210c16725323b142a0a757d5abf18ac26ab9903af3530afdcef2d97d6b3d6b806c9da1ffab9509adfc66512a329ad10;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h841b137fd9c4b2d387f53086d2acaf94f4014611cc2940315eb57e931d94df4f2a80d04ed76b7bac8821eabef94d06dbc104;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe7ce0d9f281f2fa187810773000357fab991a2ba16684794d92c04a16d96a581b14e16c40c90743498fce639d8f2fb9419d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h133161c1fdf2390627109597ec40834b13addf536dda634028d33ed2abd10c4175ffdaabcdfa5dd7a6db6e5afd3c2fa379ad;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2e7f046a114f004c476ff9511068be7dbc2086012bbb2fc95b87f178040075b58b7b5e099523bab5fec239a30c629454e0d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h18ac67dfb0225464547faba265be12b325a80191d015784dafa47b006b69f976b1a0acb578950bec682c7a7a296be6e13c79;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1cfa50d82ae61219161b6180be8fa2707047cfd7828a0426b878483f667b7f330a5e4e63bc755441c6042d87fcbd6939951;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h56ac3356307bd931a12252fd843b5de39bf306541818127482b1779298c3ea5dc6fbd37e2290119db5517b10a03648e10fbb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4c4de529902ed3d5f41fbd468e5a7ba3c13f23f55bae1fe1f359b5c5770c8895d2e221d01bc9ffe9c4f774971d2b95fbd045;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d9e7d857d1275072955dffd7cf06b9af1cbd6e1260cfb7b5b6f1facefb10ff3afafb4a40032a9e6320b9890733aaa55f6c7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae14c370ad5fbd9adac84dc956caaf6396a3138dcadb4e2408af121ca03dd86078b6390e00d23069ba8c9bd71897a6dd9533;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h101ab8bb041b604bcd6aaf6e3f66c8e06f44d9a726904405a4c77e61883cd1e7d8d07c1244665ec42a43953ca83b5bd6133b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h56b31035b6039f5284c53082fd5346e318c24e2372b2d7879e797c4c4bad5bf4c2580283b45dcfc16b33ad4a8ab61068bca0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h421b498742b0756542dde65f2afb60dea0ee65303b129729c7030f2b91cda61828beb3b07a153e15f67851466e52b42e8b46;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haebe0d8c3e19177b83d45424327be6f58c97b45f562252a244e3813e83d3a14354c52391e54cb205500597185bbbe9f222d9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h253428250348aad8b4bd4621aa2d8ad6a9b6bb749ef1e7a32cf5d5b24107b033f0b11f0fe26943a8d6456763715d16d7d690;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3a48765b6f5abcb0da63814908dfc0687b282129f069ad24128ca356d4e1fce4877e69d052e8b9756d8f0628e9933462cb7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d005299f06e6953571b7dccffae858a510d44c7bb596af50dd8ee3a2e7c1522d6279c428001af52e36cf6a72742536362ef;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h480964c12a235eb5c1894bfd570703416d64728ba6963153f621b6c61a91dcf11885ccc7e22760b310713c424ea75dd4a8e0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h98f7ce1c458cf4414268d052af1a3b8511adbaa3a7b886eb1c4c071d588b2a49c8134036a2ce70fec0a99a09647b7839a35d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4e1815db355410a12b1332131749747b839e0fad35fb66cee8485d446168df5776dbfb2f7cb0b7c2050e9f1e2daa3e6a5382;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h962f814502b1ca1b81db290c80f98ba0e4ea5ee0da5b407cdf512bc5ee3d1f0cec833be0963e0684028e36236b6782987bb4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb92d8c410990ddcda30015a67125ccf6270d387ff53036e16057574e79ed46a9b69d8b55998726559169ddf140829df7ff52;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6564c42adff7c73a9c07e4457f49d5c5372ddd164bb9dbe085bfbbbdbc8be1472310f2c7e81e0c4e5fb2e107420ccd4301c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5c9038c13df208e0efe9a12f1ee9acb171aac8d4fbf4f688f9bf4935b81f5a1446517fde21ae822f103ae60403d874cf3238;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hde734496e98ea0f5ab84cd43a65322e77559dcaa495d2f5baa2c9e36586db871894e759dc57bc57e05a41fa796be8f8fac0b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hef09ae771f152fa8b64e898f4555547ef894c2b6feab085a37bff41a5b64f177e3f03d84f12b926e52bef92ff1ee792d89e5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd56cf96093e6ec89deafb862b90afa4e1a17356f172e26e31975674fb0807611cef7c7219cf920a05021e4d94d70be9e6717;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf5e4ef8f6fd4a35b215468a0697e67e5c550833b6a3e88eada97a56fb1b97b5d89e98d2fab878dd73ef1704811718a4e2af4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hce48972ca9bfd8be6c58c8c56ea0117f90782ac32918c3e8cd89dc23e7381d66d882594059680048d7b0aa1dedb108d43547;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ac284cd652abcf0a8341434045b8c755306b8d3bcd2f590bcd468b95d1cad922f8614b16e6e4a00df03cb87ed9a04862a73;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h66b4daa8edeeba1d66ae623e883704e89405cfab5b040906803266fe94cc682294d5ef85781f0efc03d585be264edfb00820;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2bf1b85e3fabec6e7eb2cea41acc0a327332f3c28d8bb9f6bbd46e933cde22ead440780e4a685862a6456a0b499b303ea215;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h73059ba5957b2f050ec5b82acc4a56e6d97da7764aaf8191c797da92a38f2fd8537f1af102f0be6808e008b6a2b0859c9ee1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h33e7ceca3a781fc4dcab98a697deb5101ecaddee23b22f7dee29e2ac3ecedbee6fe6f18d5fe19454486656879122e5f16406;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h90fae9207cc80ddeebf9dcd86a9a6faaf90cec6372ff86b89a9971be6684959d2a60ad313bec9a0c9040d59480f3f829ad59;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1fa36b1edde7e0a60570480ecf4914cc1984010596e914a57a73e15e484168a31bf0a94592fb7e3dc64542bf32dfae8de89;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb6ee47ac236278eb2999b25d559ea01c752197716a7d6e2d79465e0d3a7aa0e3d9ff10315f372516071dc778535fe3717397;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h933e4ec27271573cc1c850eda4cf70ea2d8d789ad26b26033bb829a3ec15207fd8eb8a610c1eecb81577aca9e2ac1db7ccf1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5593706df56a9d8557aecf750ebb32221023e2e3212493175eb1f676d942967c4c22575350ca7a445afba56f8105dbcdb48b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb73028e665140de08392c25bb6467d48b5f68158d3e9e9a8209e6857545d1537e5b95de66d06041f32a51c30ffb52342e13e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfcc692162a10bfa7da9dc70738c28589be0655866b50f24a0ad64210aaf907aa817a08182692c6f0f9c3304b11a2bdfecc28;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdeb6cb7c6a6e77d7959086e24623602e58f6c798070fa468963ddb3fc21194f752646e5e1ad9416a9dbfa62e138d590d9a9e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h961c54e7ed63a3e685044e0cca8d74d8319edd8943e95af5cf98d551da425e2b73a44b142196e5f29420f66b9bc94d7cc52f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc7135427ce3c98816443586dc84ca5451cbef46f8d1ac7524eeadfd89165945f975012dbcdfaad1e2d9af5d2e39157290e31;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h51908b5732783038eae432cc55a6757aa36168ebac0556b893d1cc9eb6fe43cf53b1f3e58612701dc61b68fc62e19c3e2e99;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h24a35c26014cb71264a29ffc6442cb14d887384cbaebe355b178958a61eccec07a9e6e9ffbe9e33ec19a60cdb706faaa4fdb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc3f70241f35f89d505e15cf032e9c6b1e2bb258905b1307e44554300aa30a07f83ea5b05be09418d44cc05000420bf091164;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8a09b464429993dc229d04b20f8b4e4bc7d5adcdde15e352c82767f8b43e3d904bd7398633a9ef4905a2e3633681496160ae;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h31d1190f932843e2662b21a181a722b997b073a424ea4eff4e299abb34878817c8e6e4899a68efbfd2897446626598ffeeab;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h19c6f94312c4a4056c9df7ace70804302aa4d86fbaaf66939f5b933b1befc9bf15a7b9b8271df703691365b158f13fec935b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb46ad428fdf2eaefa4839d3804a8f49ad65b371dbb02417da82299f7902fa46a25876f93fd8e1eebd55dbf0578ea024380b2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h34f6a3c39b97e42bbc11621aa038d91f785117734d0567034798cea72f7314da749ad904efafeeb37361f89854ad3960964e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd6fcef474790b1eeeb265e07e734176a5687fb8b7204847ba9bb07644eb8e4babf701d2611d9b8bc89274106e3b50cca6a3c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf3ff6b24c112200c317775085d605e6d52958fc1269588213f53410657410df456074a60d14536c883999dbc99a2be7a2eb4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h64fdb37964ee6833f20c88366216f5c3755447ab73412ac53bcc05cbb505bfa63eaa8dc588c0a391a19fc256e25377e37af1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbffe476926abe6daea94538dad646af8be965b4c6e90a2e49f2f8636f52773f8197955333de58efa5425fec00a5c0b1c8557;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9b357ca8b0f411b5fe5ed4ac94304302af65b1b8effe7a0667c1289ff525d7cb18a57865ce06e6ebbb155035f4b52fe8da18;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ea138e1e895acc7a90826066de63191660e4eccee858e3f31fd5e3641f68dbba00dcfa4c064b7fb307cc6b88b0c0f820ecd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3bd6f6bdcec35aab043ba02873a3350cd562b96fd06a2639e055788aae6a7c69ffbf75a94a7d487f91555f1e5e47bfd4a5aa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc42a0fb5517ef22cd0642ad1621b0ea0e885aea7f3a4f954c3c5700be82561a08132766a84f0fea1a0a6d459014c0aee4f72;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha257ab58d6b37cab5764fcd11a66c4ef19fe20e4b8ec7ff92a34a1f3f2dfa1e3b6f700466244aaf864526ecbb790376ff11;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9fcdf4b9c7f183d346d590fb45cbb7ffddf529031fdfaa92ec21330e0155e38f24614e38644d0e2d9160c9e2a22893d84498;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8219f950b4634e320e87861cc19025bc2ef1fa96663394a8a507511d96937cf8b38b291b8bef932d9eede282ebe80fa8d00a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h49b3b43afbb9a2f47373f0d11b103e5d39cf4eec755547b6b691cf3d4cdeebdf34521b49d1423d89af31a1654d28e10d8080;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5aca3927c1127f7c742f79e4189e314ed20db9fd518e4ec62d91c0706e44b617dc35009f51a944f9c7d2a86230124373fa58;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcdb536f9966cff568327f29ca11f4d71aef6890410dd6a6c38698336b57a48848a0459c678c42a46dd738988639bdd6f91f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf9c51bcf3636d862e3c3fe2b380bcf00ab7d62d272b3051e261371619591c43ded5dc96888c1b5b7c7c409647b1a8b037654;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2815e666cbcb2ccf8dbede95795d6c1a7854486b8654cb6c5f741482367c262bf66d9a0fe0eb7a29e9afe33072ba4916a07a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7505fc61861bda046b1590d59d0c0edd2a632a0eb0bf8df9169029037c59ec35737e64b6f6cccae0b1a22193c6b33bf2c0ed;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1f7fb71b00fdc875a3428f62e70845dbf3a497914a6abd7725722271d1130072e165218b654a6c5c8caba7988b4bc74838;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1b57cb94c79979d4ef1aa946b5de2cbfd4184ff219d969384c9f6ef8345f0d1f32c1a4978aedb7536402229461143ad11333;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1d58ae177cea0c8a7e0f7c91be8df0723dd86c63c21005c330125de4abff44418f04fc149d5bd4c164c8ba37307a82660257;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4ce09db2daab17075402a9e108f2e92b9d79eea5566116745f357551b4c84e977fffd3383ed675182f153f2059ff864da7b1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2cff46861732b6f8db582b6d274b4856249b7f6b48f3eedddaa2737c7ecd404e1eea757e4793fb9a8140cc80345c7e6ccf78;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h163dc20a4821d26f1b22a257af54fd19b07be963017d57e42cc0558b9d72333976fbeb4f6d86a2061f808fa081091e5f6315;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd9f268406c58dfb2fccf2215fbc8f2281e49f574deb7812f21dbef70ea782139519a6458f30c4c962381e3d622e773df06f7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha286d182825a9b32b7ad5e266451253e06ee8b4e0262092c15af1167adbaa3f6a36959cfc85828c14a2511c99dcfacc6b28b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3cb4b83aa0c42a9850c387d93627d20e64aed41526fc1994029760b232ce1a98af354901f8015f536c7bc2b8f3a2041a59ea;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h289316be23f1a49f59ed7d2ac0351cf4f1fb6d177e033f9d7c301954559a76e93b19765294cd13984e6edbcdfbf554b711fe;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26cdf530f0ec0475058fc7f8635ee15de6caf9e23d354a7fe5a44aa6ca03da7fae5e256be95c7e4c47a95ff4c3407484c718;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9979b62ca3479a6e30e07833ee499ac3a43202e980398b13f8045ca4646d4dc6d756a64ab34c26a61cbf4cce1eb587650321;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h428daa397a4d106e22b6484c7ffb47b5de93ecff523c39a3f8e56689cb2c596f2a309fd08116be0d9113b2a1701f3f15dcfa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h37d78566ebabd603a24cc1bfbbf156d2461f877afb5c53fe033135fc3a85708116fbff56f17f5163787f0a235dab8bcdcd1b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1301c82b4b39e39fccba2682594407858cd2daad306fb72ffa8d968f29a40f0f3df3b8be9701db83b907ba534ef733e1834d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1da75a576d8d5373e02baa369cf3904620cb93bdd62ad870defc6e506dc96164c8b298f4588975c02f1255061bdd6e65d395;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a600abb3b94ac296b32a6d429c2ab6e6f8868788d7de7a837ce192c056ee5aa6c681fdcd380fc71a70536296c0761abc56b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h91cf1bd8f7ca2208b3571e6ee5e3c69958b291972c8a09443b2d9e4338ccc3ef2f36c6c6b02b274678c4c9c75a9a61d17af6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h22ddb08a36d65765006f88d35d4d16ba832ec05bbb228361b87df26d33fc59c8712ef0b8794cb1ed33c2d8363feedd47daad;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h34d2625080b8e517e5b392a3125c28cae35d62193b4df735e94d39555a444d1dfc80434010367c327dc97f6946bbd7b6f7d1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h51d1d0e206c3ae615f68a14b3ca9d6dca6c117451b1e7b34e28105832abf8417ccffd146790c8d6b15e9b7bb6e50fd3f5446;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4cf65d016ea744165ad8bb2e6157c116aa05d7f97a5a7ddd328cc58c0550d8e4b13cb0750cba38184d390dd4208892c9fdb1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h15aa1525e00d1d45632ac219a02b7f4b0732523ab512fdb90f8ff473c9e64c0927aad292ec59f27afe4d8a97225dd05e6b03;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h41be1259f7bc9eaec13f6878fb163329cd4f58e50901e3b2d822e4f9bb2f8f31af78e2e7eb6d45f2c3d3615a613cd119d3e9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8a3289ccd88f781e98124c9d6f3efd47d464fdf82a18cec39ee92ca620e0ab340ad51117db1932744f67d8904c1e82af936c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h96e2c947dbcfe6cbc7a6bba20ad57d62fb82f6fd3b74496ba5c25e51168fc5611faf4ebdc25a57ffb6c92454778629920100;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5028654c6ad0ed05dc590af4cbc7ba935c10817f6effb99480421dbfa5ae20935599e2230f54f5d1e9462921b7bb5f3a533f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h277bc914f98351231379122445cf72207cdfebeada6ac59d25ddb2391dc56310372e5cf593a9dbcaf46351b21116a37694a2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcff4df441cd2608853589fa464d0238680a7aee63d64ebf89ad1221fda26a4529f53d267068e7f3a52783cc0007ec2e09fab;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdec7d17f661047e3f5d957729e1ec10e3102c465acf45405e6233012b2a173ac9186a18464cd8889ca3c2cc64cd7f7c95709;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h626e63456aa3e16b673640445d680786e453e51e8b00483faf2ad65e73c42c3d93102e322f99a437bc020f363e045118da0e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9386d9181bea2a5b1fc5f99c7719f98f00c6a83ea4613ddb0fe50338bde8aaf3ae963a310e5d5af69063eb434c639d96e8aa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h90d52a477cafda23c668ba3a1a5beb4f730d0cc5f4d386e72d068aa76008da50764b05f525281815ec31d88540bcfc922f7c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h64fd2d298f95587a9335299978177be88d0d64745c55ac3e1bbae30cff8ab066d673777906e6aa47a43f1f214191f1233431;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h57e8469eed8ceef40372cb54817dcd3264de36e1964d03589b580097d412d195fd87aed9c91821d3168716052e0e10e5c6f0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he8c8b59eb164fe3bf349b066119f41922cbf2e0dff52d16616170b88318f08b6d0f562b6bdc2c6ce76555f8538dfaacfb051;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf20ca48b747f84767d949fe5e3aefe5ed6ffaf8f6bc4aa2e9376c0dc82e3d88614159c721aee177006fbe5f0523fb855f406;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h470bca2906b12575f1aa02dea2278e0fff54e041a8043b7e049593229469881b7eb4086d291d1ee0ad8f446c662808ef8315;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf90171ab7c8cb8b696d118bac42b64935255146b71a8e945e41df7d92bfc642622f29e7d8a81bd381c0e5afccb14514e0375;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf979377ebb4cc3aa32f577a68eedbd8921148d313f0393c9220f6e6da5426ffd2ecddb529611018c113d9ceb6ce130be5693;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2e4e73534b4a45a02dea5d594cd71215c0890dca9ba6ea03cdf38a5bf6c76e95a10515dc73fe3df79d3e76659531642de57b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7f440cd67be7ad2ee8a86b7e3ee8b8ea9f4c5aac4b3a905153cead9e5e68916e395d653188cf48238026ec4b7ee79dfc4bea;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdbf8d7454fc35526de1f5462f4bb4c5d24de3b229aea5a7174309de4752c1d01073a9f56e0ec6259ee49072bf9f9eed5df56;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5c10bff983ae8b7f2fcc55b60f240973fe00018b169249e6b0e0f0c507761bb9bc452ebf3266452863749e150a2633284a9a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h75d57ce66c75bd8d4841203ee606b2035c942be9b9873e3914b8f6614edd683008474479aeb3dbbf329a7b3a02374424e461;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4a9f1da2162d0c08ce641f76811526be083ab7794a22cdc1bc1ffb8524c73865300b341f8f32265aa527e0fc4fcadc380070;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h50b0eb2a81a9a987a84db7e6eadba2dbef0bd424f4d4e0338e89ff7eac4ebc975aa0478dd30d0e6486fc212cb97b334d2acf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h36a86e40583c46d4f7cce46e87a531ca674eca0a80fe4a9fec0f68be5179bf125a44db7b045f21014ce2d4553cb452cc7917;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a8a0a17fdec316065b7dc629834769e1184a7d19982f2069c4cddb409bd2eae86ffb0a7f5e5191024609fc0fbd9d968602a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he6136eafcedcdcacb888a0fc48d4d66abca312a3369eb3616c50c8b90f9d82f24c5dacc825b5df4a8c7d3ccf3a1e96a5fc6b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7acc99f1f3851c13a1f199467e349aa66a30d57ce703970185082998679603fbf0e96d60438c77dffca8d0af60f98663c896;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h81cd18a5c9d20a3b7991d2050a00035950ae5f3d79468e4c2e5eba0b887b0bdcead6af24565b7b72a1af02eb0642a8ba8bd0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc5e41ca9ffb6ddf56840378a259b4f56e5734ee0dc19ffb554a5570e3cb49ad7477b02a0eaae8df6871505af6d74718d6d1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4c0171f99834f8b2c6b82763fdc0090265879fe30bbef1de7b60845c845a7108f095cd8e31941d4724726e46b30fed0f217d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha4969e29149c3a5f34a3dcd1341452f09ec7802d8f26a2d261cc533144e48bbd2b881f62995042fce545b3e3a0a428280d80;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h530d71d832941e04242bbf70dfafbf3ecbe32cf41034890f2379e53dce052121ab46b193720db2e899718443cd0b27ec40dd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7de6137eb42a559e1746ddbc664e5cb8726a82c3c8d42a6178dfd7427c624355ad08d838df89e0de9210973a2de7220351d0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd506b976d84f2bcd1b0904630796453322c5dec6594e3579db5092ee9e0400d17ce2a626626daa01f0fdb37f9b4c57014dce;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf93c0671e7ddef414c5ca77c5ba89d158ad337dcb8cc45d339a60138362cedc925a7a8368fa8caf1feb230251dbf67f73a8c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha38833deab245f447e6dcb89495d266312dfd253a47e515bf155c40e333a2956e1dff1d80208765c80e875805e8b4a511800;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2bc205981a5e30b3884a0aba9ca41342ad24362a997be8c1a3cd542dfdff3c57d2ecc784d6c2fadc095c79a3acda49f02d1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4a19d00253779bf5581c443b4fc112a5fc386186d8191a5ef5ba1836d360c63da26c2e1bdac8ec7f9644e81342886e9dcb84;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a71547219e7afd4aa74eca4f6c070dc9d5ebf3b51e6a21bf35d2d54d32d003a5037f1ffe2f429555a329d54902d7fda3884;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcf1a7f0916534bc3b665c8d3d752eb969622c8c33657ce3fe609db58b0322a9a3a36ad3b4578a8c96c46bc0e8dfc2f382ab6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb47cc75eac8ae3cf3e4007abd52e5990b12698775475753b93176a95a4257ec94dc30095541df00a4242860543772697bc11;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdbf44561c739fc379dede11208c2ec8898930cea3b5ec8576d4406abe1dfee8f319f13563e3d00bb1ae3e93184a80fdaa783;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha8ea22e36c61d98227165dd8148b63fdc1bc71c851d18e92b40acf82c309f2c64389da788ebd5855df75639da6d397208d32;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd95e94f0283fdf7a7e737e888ec93807f559d1feab740a457aeea9eb128cea27aba7c8703c0a6a1794dedc758b71ec6a6456;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d465e6f1da912be5d08f444bee3ac9d0f022f18c782930e496329cf3950ece9e0759a32e290302c5a9eebd61705cddc897c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5dc9c48789bef4bf7a3f9fc415811e5e4b7212b4c4b717b3a5c6c046c88d0b6951aa207b966d9be96c3d6d447740d6c697de;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2cad6327936dd5a752f69bc547a5a7223865904172100f39cce5fdd3e8c7590ba5259a2bce544c117512b64dc6643ffb3a45;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9ed825e230142cbe79c911476532464dccd2f41f0430927e83c10a61b34277c29b0ad7147c5334e2a8334fdc160524d7ca79;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4354fcfc3168076cc7f062b30be9fb3feb277c0f3af95b852de5b84e7cc38932aef79e2388d7fc51d94da0ea2b6f630e1b34;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf3e3d296154f11b39fce1cb438b90c2e00cd41a9f0a60ee7664bc44c4769fc79ff17a522b8b936005b447bedef017cc787d6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he06b61368efb1c8f9b8a8353cf3ebbd4017a10dc989e4042c1197183a2aab4072aba0a06b3f8786914ac4621fab5ca44f0b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h61752409d276c4da3243f001b25ed7f8bc630d1f61024ff750c4c1a0384073d7175e7d1fb0f6b9a3e502b1b2b9125bcd9b0d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6170c7294fa0fbb5222000fc7626a6e220e313ef4d8a8d3422d0a6515bbc9030ef8e0c44c03b030d699826576e75dcf32d8d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h34989d047516f37a89e521e81429b99b32ba9df16bf953e7ccbfc0aa19ed1a71c4a3ac21ebbc057cca7d0cd70e5d5f3f37b8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe2fab00cc483bd64ca17e2bdc721131f9329eacb1b6b360feebfcfc5f489bf2e29c92e39c54de72dbd2a59a2ca1f009f1ec;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8361d34ba97b77e0fe8a86f3a31daa4b0fdca5b684cb370c611b474f134b100a4ee8eaa162e5cdd1d3224d8c805157c4f4a1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1fca20acd3446d15fd39bb55dd213d3dfeaa6fdce9b2b0356df755e65eb7cba1feaaed8f234b34d10db61d07cfc7be4080a1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hacf6108e48e3ef4e4ce2c33b88edf9a69393b2d3db2aa9f00010e5348de8ae1511d8652ece9ec0d1e0ac890d71f0eedc44bb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf0dc66d68a07061b1e987ece7def129dd335dfc296382d6ae2589403cbbbed7e1c82815be378a2f76bd7ef6631152ae72b9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7b15d90e1fbbb2554b3cad5406b716cebfc5ab95c35b58373ab22753c27afb6428e4498c9172420afc9fb81b7db1bb86a0c8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h629c90511020de60c1f977246bf3b6f997e7d524a0e45fa4a1e70e5442f405f2d80a2e8177b9f8fe8db8f00bfce3aedb86e3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec1d7b73c037349eab851d88275f5a329e7c89452ba5a81857d776ac489f5e83d40f6c318f56e8dd82ac68e2a8b2505de623;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc95dc72d7c8d0aa0d1a4f8758f4263c1570774ad35e04e2805502b301b5105f57ca6c676b77aeb6e575047e1ff24021f79e4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb155061873ab913863af2ea8c1a9ad60605abd46c2c9e39617edd35e6730e959f2f16d42a803677bec29e683a4d483f1ed69;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd7d16139ae78cabfff0307395eb949eab4197d4a705a19ef3e86ed73d95c80d5d8a97e5dd716d8dd6023fde5d8e5f3e4a1cb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h277980d856d552b68c2742b3c4767ef5dabd1ff1bde4733d0d6a7d52308fb10432dc6c2899521680c4e76df70035cf14dced;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h97bf84051cc48999f62e4ff2cf947a19a748f04f368094ee144fa86b55012a891772f14b4b1f15a94fb98063a6d955767a5e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd039bb546b1d71e7ae865a961211c530a75e160fd58be9b2aab707a2f7714df4da901d4780f3c20d33032428c997200e16f7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3ad06bb84e3ae38f30e379a926baee76a20427e6bdde3d68897951c9551e5c05c7673d7b5f2b1e5e3cc8c4c83d0c633fc4f6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha12f8530619c8ee2f804b9ee980ab62807c6a561c71ea81ef7e6ee32434ff53b0bfc1a2098b8f4eeeaca5d40d1d9fe1184a5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf489bc5fa7607aa46b6e932007ed3596f8d37c1861fb3f7c2e2825ad773fa93d8c34c709094b11b264552229139aa10c4fed;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h47708acf369d0a0c37a90a244748f68a99972d0032e5453cbd39eea9933faf453e6d53a5826fb898d3a1f67b9b6259cfe034;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfd0d98b9009381da86b412c63de62d85cc17b0783505baeaa2f0208e4de3cd2bde3d06152bf7b127e87a339b167ba67b313f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha31486dd0ac0237a42e83d0a2b42bba3ab0ac92aeedb667d49c0906b3dbc7b6edbbebae891f56d800a54e9d2ae27fae614a5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha0f381491e0fcbad92070c40d10c67c429e80312232f4c3468211c139d1fe637f711c5dfb568fed6a2860935a05d97d7a4c8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h40068413321249a9a7ff218324efd6a609108f332e7ccca6ba3b2b6300ba631184512fee7411a0086267dd8cc90de53bfe79;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h36c7f18ebeb67a58e244b50f7ec8e0a73dcbd9f624dbae4ce058800f0f8dc693d21cb65c9a2eaa929bb24ebedc558ca7867e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hab2f1092de0b2a885b91163320e8276d88892dab6c2e9f98f384e5a8a5b84c9a5986a691f258302dc9037d54f2502dc2e42e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h373822381dca81e94d63a40b4f1b5238cdd5f0cac3286142e480d7d2af51b9be20274c0fa4f7358a45b99d1051fd0fc5e263;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6c656182f62a5636194a7ea996b858b5e8b92ba025d5a52da45579affd4a83a076934c1ab5a79d052eddf499468c9ec04500;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h16dc39131d4df3f1749d4a222346e45f591410a079ba6c636da46c555bb88167ba20788d93d0bb61a7f12edd3470621b382f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h77227aa11fb52035097e310dad7d20817d07c30dd8d433a6617a2321b6004b5258155b8d0c87eafb4db2c398ace9c699d27;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7f976610bc28a949b474afb9e958fe7abbebff90ef00b4b8c749bd3ef4ca2eaa18b3b081cc35dd3e51a09ef1af2b5d697f5f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h25bf3ecbc8f9034505f17dbeb61c1f2e4ff27de91344e8d011668d7b596eba659c17fb9da200b9e32ba3f4e042fe7db734c7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h86017cf4aba4a4b57374eb87987d8d1fba798872cafdaec8895c6f60544f9be66cf1e20eab48dae6eab7ab044536f3c3d55b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb93ed22a4370ed1c10ef01680aba433b75b1d861f72186b662a9486612fe6323760c9464fa30d6a94259b0f1b83e9e3182fa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h98a1ea5ab2e387779671d60484fc8bfc8229ec75dfd6c21adbbd88280a294f74b27ed88e6217f57d9d87ee7c128b2bf9fc4f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d5b3f1995e80717f1d21a706c05f0acfa6fe064b1ad3539f5783b6240ce2114c24631c40cb1979d48f58d51a6836b57a326;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d85bb9c9dcfa50e50b3f008abe9940fe7b00cef86edff958e28baed23f0ec25bbbca96521ff30783e02c96cb84905b496ec;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h40bca8fec853d62c43f89ab5f2815f1b2ee6f784c7a69a710da5604437a636942f489940392bd2f4f26ab84e4e86cbdbacaa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbb7c3e19c2fdd4ed0a902aa2819e4028db7ed1687edf99cdb9013bbca7f4d2bf0e02f2a5dd951dd8409c57cb0b86f49fda43;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he991ea4a05e8f156136ce336501cd156fef77ed870be54abc97f1546f8c12fbe370186f688ece867da77ee4888e06db8da8e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9c998ca23ecf063e46560aa64745a7689bbc61983d1ffcbebd0c8bb455958bba2c83a3fb496cad43d521f99c4f7117e8969;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h409f5ad6d41da849456980d0265f1363cf4cf9151d3c2289df4009e3d2be22d602d1f7315cee8d15d1c7d20f881dd7704180;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd932565a6ed7e7cdde1a5bee58ba3db082aa9d36c21641933cb513736a03a261f2ebb4d12a9da0262483373a530fab399515;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he383defec6e978d79e2d66ec77957cc819aeac76007180469f2ec8fc3045e2783c1cea6941c9c128b5bf58aaf3c8fe684afc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2fc18421c94f7a6759870b0b0e4128e37e1c2a62dbd60ba42b24f2f7148c304ba18efc59b3e388653694c40390e0ec85f388;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h21208f7b0d533a0cf666fba114c6c39d0540de0d6ea2fe341c4bd929578f4095656e3b2f66c0cf93758875c150614de76ece;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hef75fcbe22693faab9a8e91d4e55b4ab11eb2130fef1c46fc45fd518aa6d7317a1649118fecd223c086ba33a28ac33393984;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc751ec009cd41c058310281a7ca364e281f54841f75a5562c3db497a0ff5829a4331a70685045d6e1b7c68657069b31ee26f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h83e479dc965138ec7afc9d7fc29e4eed8cec5e16a08b76f70e35b628f00b18e99d3fd1a4b102bd9e3fb48b399e99b796d05b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf3438ced5af752bdf6d7fd9d90b1da07f5df388d35fa3dd4d5de8aeb2b262a471c785b662a3ade559a5c3cf893e325b0c418;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h264efc05aa491381a1bd60dc922d6f89e6f70648d0ded12152c7a6d60352d98bd34a8121ca734102ba302f94331c480c6036;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h14483599fa460b937c9f49ee96d48da0a764b34a6321c5169270554095028879120b1f5425d0145e8299fb3b09250d1adfea;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7dcb7167c8fc0a551f58472fdffa29655861c989b311612be624d7e8961884c965dbda23d88fd2ee848f9ba67c843ae5407c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f762b23555e778369f707ef3e72e82ea745ac33d2deef761675c4b0fe06ce57b5458b3c4f733b931dbc20030dc9fae9c38e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5689dfab3694406afac89a719378edc7ce1a496042e41286e5ca42ad6fef0fb44f6b7265c178b2661f92e91560659167c20a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3bbe767b5bc2223acb90e08107204eec51edfda4e11b6a91c4176bb72af5fa47334100d6cbb9fb22fff4146c18ea6e9d431a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h30e3c4eb28567a42a44a3444832469f547033c53f622794de4cb1e1122573092b8d30e89ba3d64addbf03047772a152fe3cf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h49e64afb9e0e7ef3eb4ae1d8dacf9604befd08fb48e566b6970be2eee312c1e99f5bc6ff7274e28a7031237e7538edbe6056;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d636d8951fb1845028125ef2e6efb2f04989a1fc812b3f1b39d86685886c0125f2b9458f96769f18de864ff4946501b15fe;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heb7eca08903492c73c565e111a3e20005be7615e9d7c0124dd6f7b4fff2f0c5f06c5c9c63b983a8235b045ad385ce91514fa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcf9ef36f411e7a5710461f387df23506434088f6935f28022e75318e49ce9746365d5ac446886429cd041c955a11144b3e76;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h484ec3de81626680dcd0a729c9bf6133c21139e71ab951b880e7a3fe163fc7617e566c5339e73b55398c64476aa93d1cb3b3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2006d300bc8f0762bb8a612523dbfba819b5a3104ee60c0489bace4fea87e91e83cd75563ec637aa436fd9d3a564b32b4b88;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdafea5e912436e6c358c31a7e8db8ad6a7062efe03d422d4d96d83e324ab6487920a8407e9fc6a6b0a4a7f2a6300a3be8edf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd2ee61de6cffcfb0f96e50028c5e749b0f7bf82f994b653fc84e1d523a6e06d421432c5da463e0a8980a94102e6d7d7c7660;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h991e5ec47a0acd0b15858fbe93429dd08f72b767b01eeea1fa8eceabcaabedd93296f4b6267c4be42910a29f439be343b551;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2475937b57ff8605f9f57c98996f423089617e92a88d3484bab446840a09d7bc68e8ea1e3b7b849f0da6d8c9a1197fa701f1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h23ae15fc5db7e8c0b401e6c6b7f0b28a989fc6cd2625c011a79d5dba286c54418c52227aceefbc7dfef95c06e32b697807c3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h82fb2c214fb743594f433a2a8c31d7808fc3cfef7e8f670dd372ddd9da9829d83f29e5c28c82961811fa325cbcff2e701c30;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7bf007f654e6c4d8ce5a7cb6353622c5f7239019f613809d18d345dc8bdf4287a9c303faa495240c69f0eac4417ca64a017b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4369514e661e7deba3571ff2160ea5e92c3118bd28b146d3da2ca531dbcdf130079cd3e74e21a6afc1fc75fda9e4f8da266c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8c9c3dc0445c98c9effb3ce539d34114b96096a3a73c528440341bbb38cc8c5d9fdf247ef530c87c0f3cf1809d9bb36311d4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha628749fff493e2f7c9422a52dbceb2dd231d95924a6e8d843f6dcdede5b2bbab037f04daf4e6714cd356228bf7ea48be27c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h905f4c7a921aaf341b8d18f66555d777c84f4d4e6b5c358452caa9be8d38854f6d1a66667c0524a4d42ea6c5fbc59d6a33b9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h929f7a50cb47f571b8ee2d68c2da72b9bb60fe23cd0763817964e45dea66e5f52772e2d65a2d0aaf5cba622dfcd09b911358;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h299f0e678a0bedc0d310eea61afb7b31894260572a08d9ed248990ebad243e2e6ca82b71832ee3e600089569e8221cca60fd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h18e65db30acd819c70ec4464932d6abc4bc283d78e6897edebb1c3c556ef038717351a110cbd4e19341647d4644646b5e594;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h61cc94f269699b6eb85cf8be52c313bac2c1832fc83c0d594852422ad1ccff1b13fb2837b122b6127e5ed97109adef4ba982;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd8e5a1371570d0ab5d54e716794e7cf69d0dea2d684f82b5acba404b785fe7becc5c8b1f9165015a9169ce18ff47f33fc4e9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf5adfd8840b4dfdcb24f5c27e333591cf5d3a0d096a9afefc149de9d0900d47788eaca5bc50ecc40618de57b4fb5d8080e6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hda22613b48c78c6a102fa4e006b00134eedf5273593ce0b9119b2f4022c47759b61ae6210e55a1332c07bde2de1fd44f9b67;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heceaa8c5ff7bf0037b6c9a146c3ec41643ccaacb151c8d1c5652c793d5bb4454ce9f264047c06d3296f6730d1406974d0b0a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heb50d11e81e6786fc98bf62a7e571b04ab46be61cef1528dae444e6e347f784e625a235b5b6bdce58880958a6dbf5d167eec;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb144ad54883875f9e359b9d8cc32397ac14db375f48ece69c93f76507beaf5ad4cae0ed1b56d853d9ef342a20c1d9c7cca9a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6c3107aafca22d90612e6dc0dfa0a1c580aa5d645aeb249e1bd8d2728f856551e1de75fe73686563fd01839a73beb3b5c09e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4a9424a3ba1aa2a129e7a0785c87579e0eb28552f50d51e30ee087fa9e273f3a9dee1b139224657b2cdc5c96bb42054cde76;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9127b42d1b06d1d7e2623793d97be947b4cd2bcb24652cb646c1521961b342d3c7c0cfced1ccfebc5ce0141b9d065c1ada71;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h22026ac571ff6851e7ef8c08d95be55db089bb755cda7ba823f7cf8263ae25522fe306d723b202c8ce2f78d4aca1e70d0f0f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h301870c146b34939ff05bc2250081d33f5bc5492a79199f45ae3fde66af0c77057c1c0cbe62a5b20b1c22e22f5da7c9c7bee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he541f82542284adbb9562405be4b1cc027f2bd573a430b89df4d769a07d2aeb6a0e686437c426f55ffc3d43d9125a4d71a89;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b875d43aacfed6b2e94b5978a276d8d2782c8353c5b47f11f9f09f2f43a649d9fddf1e0ddc0ad6431069ea277ab978ac9ab;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc10ab32c79cf17f90db4d1d3e6021451a165195867c9d2fb95db2fcfc06541bb61eb7ea085be6369489237d604211a9a65e8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3c945624e5982fc1079451d908115ec72fcea47598034aae87b64f0885b5e9bb57fc131a399e182a27d431e8acde0529b859;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h48b8ed6c9d36774d9f448192ccd0b83d9b40541913dd82c553e15983c96db3ab134790b0f3b22f1d906bfdaab5cda73adc4a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ef081b649c4180f45f3f8b18ebf6e90880bbb12425c692a23f2515ff863d1daaceaf60d188a58ed7a5c47b7fa7f8278ce79;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h505ec0ec74c3763794a5d44cfd9e4c1190049e6ee0deee6df6ed479c9fd5101d6834b26e95e327a6fb0f674690735a5aad7c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7ebe5f639f8191859d9e4fa9a5c8c57daad0942c6fda147fd7b83789eb8ca5cfaa330470711ae96959b5be5496c9c26edd13;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h92c3a78ad0b48698a28b989a59eb0a5092fb7d994929b1f6ad0eb37c555b6c49b891009f84843ee02c9dde8b04b95ab7afdc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdcaecb29bf06e96a670f836bfffa912442ee3fd5fbcf15d99d331658eeee551accf3e0eb23f4d0e7c1ce785849303fcd91d6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h65a258d398f20a63677a745b61fbc44f083466e816c0715df76051761582c8e18029d33674bb1ebeb5112b063611ffd8599e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf6f4d4e554e1a5664df6ee41903f8ee154557924c5e862fde7c87fb2694ac26ebf5c8c741f5ba14e9bf83800fd982bd5294;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he6a8b58883d23bb57ad4431a2d0e4a53de7c1e2311a4f2495b1ff50665850a9a0286a1909f1608b553cad5001612ab57d6f9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc76d397709a771efac2a5327ab041e53a0b46776366d9bd9e235b1102ca954b1d3696383cc59912db5b9190f9c9b38c7a098;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd3098a5662dd8b6f3be883b4f5a53339ba015718e36a32ec0b1fbb35b40ed927b5ab77d88fb7967614839ca7e6775efe9714;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1045f4affaf46f6bbde42878d05ce1cde5894aaed377f31940611fc9f144fa7c2332d97de24d28574b64bb1cc90cbff1f601;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2dae4bd5d321d120d602bfc24a985876f796374ee843eeeebc38ed7ac8bb1710d8273769669647abaad2e47c7ae7ad5c7c04;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hffbaefcf8b0e3dc41564e99e0ecb5a6306aba1d2476d9bdc5b06f6843db0e6bfb52ce5fb92bcdff0c72dbf4a6f9cc31932f6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he740244b205da552908c1b4f2e68a52bef42395d33155ae71bd52ba71a836106b13deff0bc9d16a6a468768ed147da74d7c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb06a6f2d9d37e1de036674ca9e1a56f084ee902ccb9fa6fec4949033b3410642a2533dc5a3b3e29d6d1342083a5b206d3363;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc74658ceb56fb627b8b067068a9d792aa4e810505faca4528b5449678277a83567bc436b3380016a25d9a6a3f897bb2a1883;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7006b6658afbd4a1b8040dbe8c8a19a419efec756bcc7e3a9747caac11ef9e1e8ba4cef62477aa104b93bddb76b02b1b05a3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hed1b2239be647d370affcdb0d994661ca3bcd6b7d4120f079928860ac78e6eb7bc8138f3b75bcd9f334738f9e0ee47b1953c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc4fe90b0e3ee28b673a4ca0ac7a88d1062df3d666582484de7724a39dd64279b08f2a8b52d47c40dc4336fd7a30d7523513;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc0760b89d41a884c48f2d6211b79cf45d7383444915e3ecec08c969fa3843290e31659633059ea10ebd540ac1e97d7d33e20;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd9a286ca00c488d8823061c55226dde6520802095fb010b205444e15cd41e2688a3d535cdc652a822fa4dac6528dab1d621e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd3e545fa01320f7ca175c99f605d01ee9323db4a9fd459a71d2d3db4496e3c2d2275fa2d0c9735ae2adb31c86a6b11ba316f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7889b10f2a89ad32b08f336177a1761400ee1ce072d090b19a4460774bac2bb758d4c2db03c40053d54f6ac21b97f9346022;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d23ebec722224cdc086b9b1936c2bd3041ac4f065cb970d89169c347ed5d31fb8ec103c6c05f5019c1045ee6f6b1cecf352;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h30277bd1bfe0548900916e5cb6d912aa8653e8561f87d553adf0e54ae098295233e606e9164f21278710712996760793a82d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc08e6af3c4329c2b65101bf720ca9cf5262bb2b0422a01ae5d920d58abd454df4caee2b903a54680b1a5a187c4e03d188f82;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf89b0463eba07412464ae4117dfcdbf68d3224a8960d9aa3edd664ffc92d086a36baa3bd4dd8e54caf639ea1bb340be66b70;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3b743dd6cf559dfe30880f26d51c9e4f4350311641593c5b2c051bc5a910cf2bac9cccbad24f6fa9d83c4725d980325d5a72;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he72e50305b448c68f208294f845be573ce088e0d26c657c5de40be391b60055e10de3e37e896c49467788f22a6d69af0c7f8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h416259a1b2809154610e76243fbdd8a38dd8c296faed0a90da24f4261af94cfea89833d19baff2602ef670778c7bfde20cfb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfeb9f9ea8d7be7584a80bb77aabf118efedc0af832773d7e55a7001ff961c9fab22cd28bcc4fc101d94571475108f8a7dd18;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hed24408699991438e4b1cc93c5da0da1f613bcbbdb044915b52928d27f34a81c64ff69618959175d374a102edba2cfd73b50;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc79a45cfefb2782364e51428c3c65475d6f6134d44013cb8d32e40a3511491f571a4bf2965100742f6594763ce5132be9859;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc24fea95c1da7eea40891f00a21acdb34efdf47fe6598938b4371d1fe0cde116803939566330f459fbe23ea300aee62b2a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf4305a4d76141bb1828f47df9749c27ad93ee15e58057cd3e8b8379a94e58365150241bbe4e176892fd12fa32bfe79040ea1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h81a1c96d6856aa50d67e9ad7e50216d52eed478626bf2c99cc06efd0120a180915d14621ff8380ff29206e5e33d38e016cb9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfaed97366f56fb5222c5b687dcfdcad641f2720398162e4bff1517ef3f90bfde9c524ad683c9b656a461abb13f23f6da743e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ad889c562c313a1f0acec1588d522208325846fc436960a7d4c75b4e905d739b9b65d9f90d8735973bb73a663520a85ed9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbea3d4185be598fd822eca95aab7b17e16c569263386d1bbbe3c589d3453e1b2680b05fc60d21bed71c57fcb375044104526;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha882fd950e9e468ce2c5d4f66258361b8355bd6067abad0514805bb82ad61c6344fc9ffb673190f3ea4b898648180ef2e0ce;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf5ab778d8b64439439a017a4f7a74c7dc743a6bd669f5adfbcb9e719fc95e1a8ceb5b8675cbe32e44b7237ba9ef3f409346;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h23d121b40a1b3d5b8f849f9c6ef2c286cd623d02489c518764c1b0dabe6173b2ffac1025c01c9f5b0a611384c729be26ada0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h711f59c970d21f3d1e1b3afba55bb51415782cc1dc4cf1e7e56ba2a737dce77cc26483df7cd1a2a39e2cf3246151e6fe0789;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcf3cfa56977dadf1b84f83912748f6cd79e69d4d1292cae2328814e122a05154e9a3bf0683291432122199151a80ab28a891;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h87a38b8fb2d0cf1fa264894f741b409bbd4a0f51cbb98718d0d2a0d6312b9ef7b37cb5e4e1537a0ce22e719a925b9809b2d2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hce805d98d740abeeef2acf5916d9587f8fe321fa76f3079a9499ba429142abbaa4a3f63e6a7499a80a624047f112d4732194;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2106f4aa8644cfc65aa6a4657d570dd52aa9a6394a3cce26dbf0f5084dc774997cac10425fedadc73014ab36f46339f6b67c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb59134cf8ba6043b5236091017a5ddb7685e8376b423ce06200d8461327a32df9bf70a8bcfd6dfb770d840cd8e129cff12bf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc9dc33214caa9c38658f311510005da374aedaba9dda90dadc4e37bd92ef0c36b39292bd76bf27327e77647dd603bebf282f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdb521219be51c8dc10a185fb2f88dc5347b10a60fbd676d30ac2619ee6743d9f98518e3ab6fa8929aa2d6d698f3cde9e8213;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdd848eba4b2fa8707cbd8f1d971df7ce73ec06376ba7744c19dbb904af17d40f4fa83ff37c961329f7b3153a8b11e66fa01c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h627a7faa0f047e424e42bee890f8764ab61668d05272a1a64b70f9fee088765558db635bb6f945c9c6ac0587c206329fffc0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h29a3ec77233828aa76572b1deb369e96c24287ec28b7622a18fa468b2d3a26a044a05580f93dc873af7cd2bc84985efa1fff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4cb9bb0847162fbb336bafb7e3acafe649ce53520bd63af8f89072497ecf9f606909c5ee1bbcec82352080f37bdb12892063;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfc4cfe583d718b1c1d6e7050cec64f54cf48fcae1fdfc4400fafc6458cb07b695c76b2d302236ad49fd7a6fe568a96509486;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcf0430ed3deae4e17cc3fe79caa147afe1920624b2562bec8e602d84f7a76cf16a5615c5698121678f29bb6e61a0461900af;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6b5b9d0b1f9c586becbeb4fb7ee72c5d35a0b8ad3e0b69b147b4d18d35e9d59305bad6c1b2ea1044d8a310808b5534037d53;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha7d9f94553d22f4a1f88bb70e30de4599b6fe898b9d19deec5ee44ff35eed4782aac66fc7d44d23f03e63c15a6ac1fd12558;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h656e4239fa24e05451ed063429b31f3097214d83c8895dca5dc178137f3ab7d3a72abd03e5290d04846d4372fdaeb70b9fb8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9cd5e1ac726d810946828e8bdd6c3de1cf8dc9956058b8e21435db0259fe731edbd0f83c9e2ee81720c3dd1ec29b85aff983;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4084bb64dcb295a9352f8beb47260351986edd860a99eb37446d4630c8654a6408fa7c864871b2c3e80342edaf12675de5eb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdef91fbe417cb840ebd0b97cb7d216d96bb05345c70a253041bf14196f77d9f11c981745e62aa42e9758f5c7309238e963f7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9e3001ec7484f253242e64193eed180cb34f2ebf269765cd25766540c1c92291348a33b41c3f5f31c75b4575ee3979565bb2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd4db6785e14c3127eada9c23b762946a9664805047c9b1a08034bfecf89b8081530fe013a82323656fd3e571cbb6d3ac1a92;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h87743cc328f2e6b7903c2ab2a24f965d33e33ead8db921307fda31d650429e8670e5d38ce3cd640fcab309db33101eeca817;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3b72b33ddd0a03cd040cca58ffac9be5f204b4537d2d57a4096916a58fd319d557d5eef41b11ac639fdc7ace4abd83911fcb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h74098fc95de864d0f2c9e2ba84a32f84002db0dd0d7561f1fbd6edc3da86f69f3c155a754059dc1ae5a6ee2aa9125c27bb11;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h628abb92a97453f5679e99874951456aa9e9f111465ca21a851513e25509649cc3537b75c0629170b751ca0893d7cb58c417;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb2275ed2afc2b563a48cb22deb6769d6f74032a19c7cf7acb03deb5041dd4b1fe51419181f094a981edeefe4f195d1e1936e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hee808cd53cbdfffb7bf964052bb39ca7a62955cee74c1182dc33454067f6a762d50d6f7fb3a51c4ef98a30a3a4c5cc9b66e2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f22d11ff6bcc09056e6f02979de6844ffd191516f0675616636ad7b6991717ebad47bda220af7c43c1511823cff1c22d817;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a47a99a25f646aae6f38f9429c5fd7f1b2e8096927845eda8fd3333ee8e2c3b2369ad56fc03aeea18b3ad42455e73a374a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hce1c5f4844576b55ba8171ab6584f237ebda4898c61069ccf38986771311b5516e300cf50beea04adb0a69f4bbb212dcce0f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc505abf2ed72d30aec35230b11fc0f5fc1887a5dc3002225fd2d538e5bece753ebe12d7cd54a63009a786873038432eefb61;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfdbf821cecb55ebf51d37208a5e94c02f7322fd0be319c4ca79eb58f87154448203b5bd09b72f12e78f437488a4ed59d5a32;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd6136f73c89d2ab83b81eb4c1074382aad7ac216f3665be6bb0efa287a898246bd064e35398a892eb4c5310ccadf3b5c4f09;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd5c9a388f1503c656bf3c9f2ed1622a99a1ee7dc49ab1efb2b0d986df4c0dc54677e564464ea445e7c940f27c8385d206b43;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he371d3635299290c0527f6f3005bac9202254fcbb9f647744ed2267091a3ea29d8ee6df7c943cdf3a09e64b6226dad79c317;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h50b5e40509769e82d3e700455c5fa865bb196fdec238e3e9fd8735c97e2ed722bcaced0fc0c44145d85333e56a9e0fe0c5ee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hef4abb2d7017a118c4b70a4e5a0fd24f903e4414de66302a6d2e5a9f27fc335bb426d20e14b2f85591fb31b500f0e1854eeb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdb0f9878db27ef04423cbed9516f19477ab43cd3690b9e193a009e1d376c1a94a83f00f485cff18898f8d69ce86688d7dc3a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec83702eee2d5f5a059a25c34a30b063b5e53ec0cdc3d398425d12d19dcfa11f73524ff48cbdc85e8b69f50e5ad6c054dae7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9979479f781897113098242648af077338f60d6cf56e7a8ba8885c4792c9665ec3e31dcb25838813f6295fba55153c040023;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3fd060ca9c7b2978ffe2c95cfea29ebda891e844950a5d8f88dd04b939029b4302c2990e68df496a604608a56f65c3c74fec;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9e77802fb6767a3280c1211ead3af8defeac2f39eaac629cf56bb6e8c25c8d4c8cd1b496b70c1d32f7d2649a36f278d46510;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7934055001957ad1ccfcac92e3630922df0f1ff4c3124fa7b935330868324b58f041c5c6bb1cc1fc6aaaf5bb6c0ae37ebd26;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h34f1cd3f6846a51271002ea941125d918a79ce3719ed705c09aeb421a7dc4b7e268913f2b69d38efee93e610b8ef9498376f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h38021f8135007be95cb9e63109035c3caf197f50a6fd1f1cee0450f3a126474f34ef7d2bf4abef6b9f3d7ecb44e704c68b01;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h37039dff5be18e1edc3842fa01750360003b65aaece4ed3c581bc12cea869d1653645bd9aaa1d1608f9f8ce055c298ed1f69;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h28a97777bc5e9a98144f2f70d8e538a3b96c191c14c6de59e4e899db25af72c8e3bc8dbd151fdedf4bcd1ec3191d5c6b8a83;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a7efdd3fbd60f565fce8c4667927b4a949979e7932116d697ff21f1e37b72ffe392f1f675ffe0a3822b69c6961afbb2012c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd50a777373012101891ca1f0cdbfda70c6b370a5c929918ea48998031dd78017812581c7c11edff57e2c72e94bcaf369ba75;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8cff3a72c2e52d4b6d4a1665025308a090d194806d846ab488e6ffc346aa34be066daba2b5e0d05e0bfefb9fffa94dc1f7ff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h69c36eac4ccbb41ce594fd673450e0c11508f41d08ed3c8c9d0b32823b041279a520bfad4a18f60e2eec548fde1b3b1aed56;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3bb66fe53a461097dc3fbcf22692161d3fc21e40d674c574e07b321b406c8816b2db5595baefd746f9d8864159120c5a4a88;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hef6efa3fbb9b9f4e1ad67cd11bd4d125e9ff17d90762d0a53dced3671ad30b6babb12c2bf98e071951df4663499ec35aecfa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9c7a93a8e4eae015dce238a06c37f9e9f32c710b074887261b4c00491ddbe832cd93294482d2bab81f6957739a1d11ff4a91;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7d6179e3f3e17ada52b54932146bac5e3119e4da11b975651712087241cbe65bbef612aa2586146da3d1b5e5ddf3c35513a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdbc2856bdead799120a44694ce1ae94e32676fe85d3b9190b05cf9d606d0a5311dd96deea20cd3bb56b8f58731552b7d7b9b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcf7615786cda91e4d2090d1908f0f90596b45e46dfe5683e2c669e9ee7ae489b600df5f3d280d51a567984551bb2a3de7d30;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1497d2cb14d3a0278b6edb02735d9028798db9abadf53c1022a037b316a3e7d7bb10be52b7d56240c31021493a0c53ffa422;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hba9f846c096bb3399e89331c9fb68bb3c63d4fc1f4126757375336b0f2e9e9e726b9dc39433b325dc72afc54c51a6e186d36;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h635de1dcf3fa91072d7f950f2ed7ee8beb3878f06b064281600f7dddaaffff6fbf33d5f8f6e6d2268b43ca10a0321601a36d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h70868f73038d93d59972ebe86f89f7fe4643f299ac89dcc00594b0c4a8c91f460c3a5267fb493cc82880b13374d6b2f5021e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h23ab098b82276311cdcc8c46bb5fe18cad7272cebb303ebdd54d81fb4f6fe401874984e77b76e5325ad95146852ea42bf3b4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3ed653a0d273bbb4ddedc3c43d719ae1efc22d9fa061bcd1c0af166cd7aa37337e818951f4270805ce0832cfa1f520779735;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf16ce2eeda16b7d1867bd480dc1d1fc73a9b6eb86a370da140809512c4b88eab8f91b99f0ec1f44c7ceb88e2728f8da0e7d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he41872612efb1f0519cd27d22afde74d48ded401e30c2f90ae463f8bc8a7c7eaab9da3451d4ff90fecebd3ab6eb771097d71;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd29f1e77967f855f61273ae7fbb26cf67005fb2fbf26fc9da80255925ae730f6834639d992d704cb0c1180256742f4286f6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2dddbcb7b944c80ac283d3ebbb655cf1b78637e760f1663c4f56267d36e71cd8b3806a4328484a85de3701001b79158c64bc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b7ae9bfdf8dfaaae5d2128eb419ea7790bc30fa632e78706f734f4b7cebe68154411d21a3b32db7d4a743e1d67ee32b27a0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h148a1579848770f1be814490117b3a0894adada8dfc65561127c89cf6f3b65af4f1c3a3e404a6846e6e6d50413170d45b8ee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h80b01b52dc5f7133a1dd1fcf53c1d45dad3671ff77762adc1e04be3940dd323d9955ae9cc084d3379c569783a9e1ff2984f8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h79bdf2a78db36082a78531529de3aff700b8c7816cf193c2894120f4ff1da6e3a8367ad91fa69dddc2d32be6d0820563933a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h72d01eef47a57a296158e5d3474514b9bb1babd5fead8ff0ecc2ac09bc97a084d34b37d7c55a378173e182acebe597024b4b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h91adc38c722fd5cc9edb6cab1210eb3b2e490a4ca845d663deee4cbb079f985503da8faf38ad30a61311c9e5401a3117fda;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ee9eccb51145c3602e78e526d9eea288c514e270d2422026523657467e2d70fabf4c87fcdff3f054cab5fcb4c9562ad0ac;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc99835b0e16aa45fea82e0d5deeeed8bb20ed37685a53a654cec08b829648dda69d71b3b53bbe17753d839e2b030aadf5624;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h24e1b36d13e8b653591dab671f6d73f8a77232c0d39a40f060266db0b505e30d3c32caf2a094b18baed7ac5e257f7e712018;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9394f3bdc7fb4518df3ef7efad59727cb6ba0cdc4f257bdc07ac6e84dd3731048f77afe48ff7fc7ca54d67f5dc5580476a43;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1500fcb3c7d06d55259863ce5c4ebdbb46ab5659388b321c92d428fe6ab4ab2b67c4fae3fa15bfc476c8be4aeeb69515e3cf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf724a7197138427a3791118ef9e55900eaf053538403de3cba406ed4e0ca6f7b119a1e42bac770b6015a2b7a8ce4abbc1a7a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcf733d43e891a9f3a16d257fb42ef2c06d0a4857823d30814a378b61760fec78de20f3e155484e5d7b36b3bb390dd07784e3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h402cfe00e30c25aeadc3f70b4251b138c15742d23df8c2c97d4c3a5bcb07495459e7b55f6fcb4d32cdaf23eb9df73ccda311;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hed9ead37145e0da7314c5235bb56069c930a4533741380a765c855a194f13cbc8ef4a61e1ea1a2a3f3b733e3ce8184473d77;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hce10060f27e4ad2458c0996230f2ebfad9879cd5a4adeb783726db88b9751356f1695de7a39e4fafb335ddf4d43596717190;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7be9c420f4605ba94791a8dd391a814cfe493adeee2771a31d705f09998da123490ee7074de600ae154e85619956ad52094a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h74a6419fcf6cc0b5c14c93098a30b95e30313371f5c371b8c6765c148d5d8811a29b02d26fbfb01aa16ffc9f68b5a4da4269;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d8f5e0b94d746cf26cb4685156f9415317dc749d25c8eb86bd8e325358e5f7cecfaccefb356072e80f025dfce983e35e5a7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hafc1fb3b6bd028275f6fb5ec17263920e6c89874afaf74cd0e6aa132c999251f7a3bee5f2e4d7e227b008581e1d4c08f6de5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h520da7174b4364213e564c45281ca1c4e45a5f3257f340ed6ef7f02984e6671b5889d6121c38ce4d5086c7e8f52faeb77c4a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he4f58ef1738f1bc86fd7fc53513da60c2d1dd32f0e6ef92d3e89dcde91632459f483f5221c5400c8d93e2a58d4395a8a6fcf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ae479eb7011e6fa6a3c990a8d3ed31342a6230cb595faea48463a83d4425b5486c343bfd452344a21f66b6a1b5b7d016272;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h12dd7418b4547763d6f7a78957ce776fc012b2515d624a127433c241591fd029fbd68a9e5916b70a46fc63a97623df848cb0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7d3c863a6a034726e8a706d5ee75a165367a3270cffaa191e0c349139bded92bb60d6444cfa175c35b84ff072bb4f7c2c99d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h54381beddd2e580da59ee4c01e9ceae8840dbe7a567e4bfea85fbc39a6796c10fc650521c7948a1bf9e55a8ebba43a2decbb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha8d6ad03c33da0a03a621061a5a0b70dc49d98519e1045694a9112a669d921d70f66a88c24c25e3ddada85d2f94dbeca4e75;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h124308696bd034a0e259dd02e141bad19a6ed87ec700d249a39cd2a8ce2919d663f9f067aa2671720953a3faa75427c36eca;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h79d1559a52cb581fb80a733d5f1835dd17704bde8981a01dd123cb89bc2e5d3284123e85a95b1e8e26a0a7b46614673a508a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d67440ba8781fc18cbedf36f00c3c60b278f78586cefa6ef6430f409eb8a335921253a186c65bb4b4aa25ea715a0e1e1fc8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h54682f487c798892d633b399ff605667def62d6bf9547e99a7ec8635c793623e7786b68e1eacb5a6ac91f2af6d71c3597561;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9e2a94c02d688590d2a9f519b3340ecaa90a0434ece617fe9a64dbb2a93b43922a23ff68a93edffa2d56d6df97721f9b8978;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h254ea07bd38b74a849d47ef98a27eaf7467233b2de3087a9da820cd8231e1b40337b235fbbab41e74cc411c0eebe33084943;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h47689d90c9fb998cb79363abddb3839a82f1da288d710e3c63f863a0362102ac2998eccd7865ef9ccdc1b1fd18180b91e09e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he647897581291a945f0f67a71e84b78d83dd94587a48ee6f77e99da7ea9d1f1e506b4ab3cdf8692504dc82cd4b9f3f1f9597;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4d4302ae7bfc84d96b5da96cfd06ddd0fffd9e6c0203473571f363eb2b01a2f39440dc964c761d4b2f716855ddb4e4b052e7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1fcfa3c3b1668aee7b451f851319380c6f9aadbc01dadae699581324cf7fa5aa7c7972aa7a7f2981713067773648ed9cbf5d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfdfaa368229cc888ad1f22e9673343fc5f1b68efd151e61adbc7e7bdefb8b1680dcded3063a1c259e65d7a402a9842a3e01e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2577956e936e4655b3fe82ea43b4cc0123f08c197602e74a624b9048e5ad353ff3f0a5d83b9861ccd09b5f9b1be598e71655;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2df6fe177c2621ff3db256b340a50ee4b15a9ca74b6fa6e415415dad8ae4fee0d92756e42046231eaff7e31da79a9bfb6125;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9e1a5d57e3b0666f4d930e2ba20344432b0391c658836fedce3d1515da24def7c7c676a0a39099331cded8f0888fe732da4e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he13d340214cc0ce4c5050107b024dcea3c3be467593ed962293252d5b321d677eba252baa4eee322533ca6d192760be0c837;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he350ed8d554072a88c11b9c3abd8737ce7e90336e8d69ea0ed28ec7e11cf7797160ceb5faf09f015808289b954b3df5e2e4f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc0705c66fcf664ff69ae55581cb9bb3234c8a837919fffaf240d45a4e16b3fdb72d478f5fa98ba0107713a87109d78f497f0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h82dfaaebf48b3fa77462e80e1cad56aa7eb86c50dbc78d83f4d3eb0ff44d1203b7bdb2376d0995eb49d43913d4d16f53e7fd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9fe41a6f546969db51c713eab1ea6ff5b575c79b3908999f232f3b531c4e43cd0e446bbb79a613c579f2fa42c628fe38f68b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbd6222ece55d4d08a510a51fdba20586cfe4060dbe8bd568126ec85e658f8ef0c0ffea13751858bdb5a9d08fae1b1e768fe6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6965607f7bdeaecf8c1c95af2299dc4fb0c6524f2d9bec894f7cd7dd8dc80079fd36e97f6db49d5f633db2cc7b69f26321c5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h569f8f5a2e39ab68489f2177fa9462c5b3c65833a9ccec5ee89fc643688d953af24f23d6911b525e75fb16c0a52786df6222;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbc6bfe5825881ebec8bcf9cc85cb2194fd98beed7a94093ad5ce69df613247c64ddc922d2345a0ed6f6dcb23639cda7eb071;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc6827395d82ebae9156c7d20688919ee4f3b3d89cca4e0dd634f2e38d114f72d7a84f2c648c631e9d7c9d4d462a9eadbac68;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd929d2488a2dd081d0e66776371e6ee19c1ff23720d88e15644b9c630e1541822280672fe3a46e8a130413fe54231177ceb8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h79aec6c03369b11b55a27e01fea1b75b5c11fbdb352d24a5754e76a346b907fcf40be97ef622c48b48f70add9f57f941d5fb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd394bde5e46b2bb567e3d924fa4ab17c0b5ecdeb8153672b6b7b7dedc23fded381837ce8807b7644487d685484e18951d080;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hba6b19a060b28ec8630687199b13b44a930e3afcee6603f2fe20d5812d5ef9ff93c5440eb83df7ed5cc0b96f9085c3f1146a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h60b17d6361296be5d073cf11198cb06b7b22ef398ab51bf37c2f2bf49f4a30dd935ce8d7aa21f0c7a92a8edb939cb9b4c003;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8bb9200c3beea552729d63b595c7fe5ac7d5b60f181c70bd1d73bc54a198dd98367fed468bcce55d63ebb3a4fbc3a9c1c3bb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8e6eec38681e76a7dece2fd730d837ca5f2cf3509079ac9d5a180bdc928b7bf0045a7597e4d602afc77fb76c0d911cfb43f4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4aae2f1cee324820c4651047825b2f3cb34944be654fab3877c525fa7fac54d61f5ff3c7c5d52749fb0308749e7883400b26;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf2d48e2efb7b98c152eb0c9dc739e889f24e0ee1b2bd8b56da0413461e126268d776f70840bd215f4282f6001b63d04cb7b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2c117f6a845c0f7d259c6354c06441ccef5130b4d74a88f255ec446d9070c5a514cf81101eb10f7a5186ec2c3339884d8f8a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h95ec26f0e83e8d8aa2936473ac767bf1bd3bc982fccb0c53f2eb813b24fd09cb6fb6a7113e75907ffa3f5965368a51ed7d8a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h35b4e254b13b6afdc15fb15c6c9ca3d6ec807bc4c11eb1e4e36d68d96ebdb80b1d46066a4b4200b1fcd8220fa6bf25fc1d97;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h10f5e97469aa76f91d5624e622e3adec22f570c35526714611d171d4d539a8607cffc126fbac6a14763940a9138a7dd3dd16;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd22c2f1de2c6d83d016de076f7cdddc8fd4af6cc8619095b3c2dbeef3b36cbcbdb7342721eeb44f8bd236104f6b04c0ff1e1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4c7d819bc8eedd3375211ed072e87b1ef97bca493e0d7058993e11a799d5a27badb9771951990a40c79a2a64ba20f8aa739d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha96ce9ac11f8917ca128d9878b4f3dd66275a6a539f8068e15a42e807c59dbc814556cb786c6ddecf04e9253eb6624ef7fb4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h531f466a636adab9ff073dc1c03d660876dabd02bccf56d2084a257fa96ebc659faa451ffbd2c0cc9e55ffbf4ab6e7c9b97b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7326dd2f64b75d10ef79644ae73b99b9338f9912249aaadbfeb0e2ff1454fe40428e85ff1f1853e67c6bc3ab54ed25b6c349;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcc110c67c6e594805bce3dbd42e76cd1c258818be99787d0e577d2060fa417aedbade55b81609bb855a5516bcd9ada7c4a51;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb36c9dee65810f89c7844bc693893f1c531fd4f979519a9e627461cf118ae6ba26715efca2300540c8bcfb0467182603f348;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1f34f75e0757d176af00a60c20ce2a4ab5abfeeb7793f7f7776e19e634896cdf081546edbc3beac1855fc8c728f821d19533;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h516aaf117149e0858e9755cf1b663c449f619a8eb560538c59e1389ab93997c4b6cfe88492d2a0b146e9a5a81f0349c4b661;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc62939b2f5de04cef3a5cb666d746ee0eea097bf15efc625606982be8f7021b4bd03bf1bf6616efbe1507369305230f1c4d8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h92a5c2ca6737a5b59fbe85db5469f0c0bedaf171dd8cdc4bd684be63fdec9ed6906428a515f82cf3fd445777f3bbd21dfdd2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9e54b8fbdbac03dc3f74a77aa935896c890cc2de0bdf911baa723cc466c357fb5bfe5bfd9b847f5177e025654779f3572cf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hff2ba4566f57c8e722e7a96639b6b0e4c0d00ca96979f24914b73873a2838a5f70e8d0570985ddb53cd780b662a66e589577;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h660c4112b63d9afdd7aae98a6ac15682172f8172a36101a719d4ec3d04a4d01962d327bd192acb907e3453340c7b77ad37d9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h73210d1278c233e7b5ba093e557afe02e10fe876c1d9dd5e79ffa5298375ce3478ad6a00ccd4736ba002941cf85762f16c9e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he5cc033a8d9409ac3fd2ccdc64d53eaa1195735ef55ffe0a8d2a87be0446981b214d8e4db75c869c691c3dd3a9236c0be7d4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1f908500de2f56f8936a21feaf5a0edddaee4e1e2b504d5007e1cde5847786cf254ffec64a52cf773ae26602104fb95b412c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4e9656cdf1a6a48b86b1d639bbded086153a9e36a1e9166254701f063271540aaff5576a7f1d88864e3cbc0fd3998982bfa5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha94d087728606aa1eaf93a4bdd98709c50ff0e045308ff9e695e5dc2ca6a05f6b0aa52f9752912bf455c79cec9dcb75926ac;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc9ad12c78d699ae4d4b0252c0da266fa91000f2f29e392c8f18026d8cc9143567b89e820ccf5645f5c06b0554ad3bcf6302a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha062f3ddd13d054505693bee1366a3c1ed4985759971f5d879165b9c23e3dafef04d5cd8b037c6135e844d3a9518fa7cb1b6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1dbbde880c91aea680dcc4b1af5d7e0174220e2a76108e69b9087027b22d11c1135c6301c522e74f56aeea280c5a06e20fde;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h36cff8064f4d0a43a8ec6c8abdd05a31060e813d6ebe3d6c6eb1fb55ae7801935011d41da4255085e18c776197b51d76e36c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a289d87b1d8ff64d58b98444831787916e29f0e4a9d3d4f9a7a2232743dd240b228ced35babf2889fd73740c7d7033cd3e4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha649cac858e1343b913cebcc019cb6bef6903e51987edd5add96cfa4a3d6ebc6970e836b1772e448740e8a1105749ecc15bf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h58dbdf92e6d72f639be47590abb67b5dd1494ad87265d3f0bb9a54c883700a66be113f6df2b5c2aa7a1bdc8908a43239d9f3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7578160c9ef05981ff6766cedb37c5e33ace8e133e86a2bc3b4725e80c9a4942b0d7948cd3de26a24a68e535e58c883953f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfd4aa83d3cd9341e0ecc4d60fa98d5ac8c402385a7fa936519e224d49cd1126e4c0e203458b9ab2243f6ceaf36600f8cbe36;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h83ab059f6812a930097b6df8be75940b0f3a1e709ad86c72effb9ce9a92a3d296bf2c3f7fcd0d10e6969944d01933eff329c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfd8c7eb24fe7c021dba7690d07291b482f75a5ade1cc81056f9242deedf94aa1cf877e874e083e93e57264c6e916cabb61bd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h80a2ba8133caabce03a42383ba000a3617abaaf31d93fdd80c0df464f2d6089bfddf9d3cf63c4639c4c6d3b3e1ee00be0854;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he069452c3f6b052c61bdd631ee0d655d099d7ab41b7ff14f1f905cadae845faa7a2ff500025bdd0496780c17b1c88e7bc19;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha0367f0f9bcaeca56eaf5946faaf6c9a134781c2b5d2e0dd8cd2419a61156c8a673805cde1d2bb70744a952a49f34c7fd4b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h752eba2ceec6a542ec97eaede447c2450d236710a73346beddf3f627198587e7a0acb32361ac315faac85d42bf04150a6495;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3429d812d47aedaf26302aa03f94fa990629a6cdd81198cc0eb90b171bbfea532ea9754e53cd25c8dbb48519475e69c7959;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e1460df82fb299a32f470489088222e8a63837db7e88bc76816ba0677689138a88d04c5048cef4b5f87e942bd4458147dab;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h67cec17986512136655618fd867c6ed04be653e205f00416c3dc694b26feee73f35851e0d0092087f6e8930c3a0d3a3438a7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h12b9ec243c2aec89fa365b203db32de4c4a00604befa750cb1de317f8df25b944cfbe12c12ba5aa51f29c06f9fd1898dc214;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h589caab38085984e515f4f6108ceca90265204639a11df2d7b8dbe56dddfda9847b206aafb923e4ccac1bf550ec6d8515d60;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4f273b781a7fefcdab989a4c3dcb62030b2fb1a1d1669993ee3d4d009b72f20a0404351b43e8046e8bd80e9b22e1ac581d5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfc60f2534294327b5e8b2a2db4e5525b58ca41550d86a423a55c82aa1bca0c33de322e3bd60071d26655b20bb0541e5e6a29;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1835d2f2ca3e61f1bbc60caaab7109b444b610f66af1f899eff60209022e400221ef2e8b8de767ec5847d499c983d3a770e7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h48d28f8493ebc32619344efc1d62ffb6ce030c6d50f2baec536e436e133d4a20104ef31c28daeaf1a5fe0cc756bd02f98da9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h57a09cd7f9999281e773e21c323dd07b679f5eff18b107b1cbb536a161244f2aaf7353712a07625131e4841b2598c8708cda;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h90c34db87acb6cdce755e8c86e77b715f716ec2a813290386ddd23704641c1207850380664ed4d9a0ca94e2b9f375d483262;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h573aabd252b30d5aea30c7976d1c65f5671ca27f131da89609d62dfb49dcea3393bf19efe29585408f9eb79a3906c08015d7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h55e583af5e56a3e70b98e2d1efc870d4491b95436d326a6fa9ce7b8c834501b6ede0d38d060188a191ab4ad4602efd9a78c5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h564b06c2140dbcd19b344a10ad4a1e0c32ba5e6a9abdf14039ca93be7a641f0b989b1169f8fc8673b7ecbf4d84dd035b486f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d08936d3cb4510627f930a2eee7c0a38318c598e324fdbab1689df258cbf4f7e5a470752a19079662e63fce1461baa4e54d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha72e487a42fd05cfc5a9ba233a7d320a275da013ffdec3f92547f42cf9b0f87daab75819ae2bc460d375b3941128e6d631c1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2cff84a87b308bc4967e9bd91aa625e9d49b19b200bb4b764a7f4181d4582bdb858d5497d1986e05b3b992eb04e1a3585ea3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb604130e9e229a1da35ed7e82a7238322c638b7468e2ba78ba66fb4eae923a91f21f023a7a0956325e7c36ed5b5750e85778;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heddbd0240d6dd1bb230a567d4b08abb9da8089e743d07614c507ccaf20b2f7746414e83231e9319e80f0724792d3ebf75b5e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3ee0bd9fff098b501adb9e1a20ef2b79e0236361260ed7ab0cc224e43f3b47549ad932013ea608903625635896d22ebaf31f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h74fbb9dd7ae852d601272025324a0fb1cdf3fd809dd1ccb51f0cbef1de9b4a350107839ab14eae1f6a7c152b7fcf167a1931;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he477f5757396c10d62b621b59d95a320bdc49f82d1fd2b497ab13e91dbb0833b715472d4b883b92219a0ac52bed1aac93303;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec77273e4329d9b9466f4dc81f38171649c4a8cb6529defc252595342cc3171b4551b14cfbde6fdc1bb31f1a073bd9f41605;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9dff16afd93924f80371d6c1d641f0bbb9cb9cd303b4e5d2dbdbe7a615b3a92185dfec1c84980a37ed1d1a766ddf1a33284e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'head1937783aa4b345ff1085a3a218cd42805824a9639ec9a919f1e0abc282c2ad36150f4e114b98bd89073985047ef2452f7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2384c07592d67acb37bdbf9ed819ac27e908ca486273d2692c5c80b16d7b6c87890929b620775a138eedfd325a3dc46ef62c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfa1d033d1ece81e36b54bdbf5c28b0028298b9e2eacc0e1e0d4c55e1f396557861a62ce27a104d280c96eb4dba2caf1f8300;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ba9259f4f476790ac486585f85ad2e998c2616f2f99748bf948def50317216a6381d9b56b3b524c5557c409c68b1e9728c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcd08b0b741abdc2893cad6eecdab3b644dcb54212b3139f6a5119aecd9e18994159ccc510222eeab10cb56cd146c730b7182;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h717c1dd92cf422190b371d9b2c470a8a55b45d9abc087a33cdf9bc351b32080b64be8dfaead557a6629b4c7c1accc8448436;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'headc9ec99150a180a88e3a5f674917d2e128161d9d1869b557aee1b6804f9ae9825ba306c724d3cd2d05fea1256c6c19f440;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f9b156c432e9acbf939d4ff25c99719127b1b1dcbcc06fc40085de37eb3dcbedd8eccc8badcc3931bcf97c8108c23d0eff1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8fa6696f233a51ecb547924f7211331822d73f8402a8f256b3d54ffd474c61e98bfc900d6cfecf0b68bd44395a5f9d1ea3f7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6b0f9032be9e94fae49fee57deb40a5edd2994f790e0e51c70f76f81966f8f75f437e99f201a27045cc76017a1c55483db5a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a59a989bb480a21a9b9d51a33a29592ca0fdb28d202f9463a1cc7eab3a7b7fb06d2018895ee0b385feeb7a949f78d1c5c09;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha056f63783085753342f3ccb232e1b573da07c3b3b71ae5d7e9cc32743d8a4cd9e60539ad769e15f8e6dcbd081f923d65562;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h654e5df676c02ef8fc534746b07bde01cd5d47e10bf0fa69cfed2c3f36a5cd376e46ea9540c4e1c081307c4d5c6abc77b64b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h49547b553a5093064c3ff87476dca58aaff75c2ca84c3a46a7ada6288ed39f821af47d69e676513b093f191c23f419d3c0ba;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8dc3818697ff764c42d643b097d4b29853802f351dd372bb087c2fad6e853eaf91abce1071222d03672a25e276db93b5546b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h602e942429a2313e1347c9b831a8918585f6879be326f0ca68f2f3e9399a683d22a26fb489db2ed66bdf38b658e3f3330c28;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1c8f7d9ab8a73282ac6ac8e42ae2dccd2e220e5f21a8eff1d20ccc266edb4a3a69e02108f4088b7ac2fb214d7a4df3d473cb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd50a7782940852fe65c60cce44454e8fb33452ac0f681e328994f5a311611dd1771aa03b25d0c5b1e859cd034d071b245773;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1ba8c8925ff6fbe7ea8503ae90572ed419187ee2ad20ced0215d15a96c0faaa1c6b4a0849d84c51524eef68c7b28515248c6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha8115b3c69c97e82334ef123c89c35c3677de0b5216391c291bbbd2acb574444e43d93397453869ddd45d9c2a0a32afc248;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9461e9da7cfeb6f4ad86b8b71b04bfe65aeeef823ce1ac0d7b42ecd7e247b83c3b7d5b9ae2bd56ffbbd553f741739e6cfed8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3fab779836eb4829b5153d1a895e817443138f42706318e7d1e727ede061190a0751e1fab84babf69b1f8c0f4159109a5d3e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h781006397fb16af7f013032ece90b591f7918efc6b40508406702b2fa7dbf70400778ddfe6e567ed1a4d43b018e495ce923e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb23bc12d3431de38c6bb1ff17bb0290341ed458810eb176eaafbf5e49eda8921b8e3c69d8b34f65026b323139727e5d067f9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h25b37ea6f2c4ae8ce2bc4133feae9123fb1c14de313358adcff0ec7ff0c3640140213de40f8f2b7475bfc354405ccc36ebd1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2400b504b6f41960755bb2bbf17310ece312076797ecdd242cbe0abd7e882402bf46001450195896461e42587873681dd04f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h62207c501eba147b93c801ae2c8ac9b3b6944ed20ce2c34986eadbd6b29dbaf6d417487c00a61378b07b6d09d25d281d3b94;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8b59998b5e92003fdde58a3724b96e2faa84e6493a5a480711fdeec74bc2af3bf40e83ddfeebac32ec0eb43678ee771144b5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7f8864c23db1626173be7c8c099a8ca8ff4c15839318d0940cc727d860b5bc17c97dcc3dc4649e8822dd83e3753c296dc2d6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbd68acd3f642cfcc153edd31665831b62bc6281cde3e6bf0f9f59bc4711fa4fd1a4927b22b85aa0a4dc833a2d04aba39b3e1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2602634523775dc42a4468ce57d8c8d148892fb0458121b8c9106a21a594042b19d4c43f289667459709b18edf9a7a7c0e07;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc6b6396dae63d99428e800e2db9d79956c96362377b01deeda6ad00022b26f14275b6104bdf95d09103bb5ac8f27b893d77;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd78e328fcd15fb0847ebdaccfbdd8c2ba1b8f0cc22b138870f83203ec0816bf57c11af0f91e1edde6b2eb10400d50fd85256;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc598a300c2b8cc60eae941d5d72cc29419f5d470cd013b8f1106b7fa8eb20c3396aa1b9c1704cd0a12ff214e02ac64c78ffa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hee3173822f1cbdacd769318a540cbd0a9fc6714a9f0813894a2acf30184a07809d35586563aaba9fc0ad613c5415e677a823;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd6a88ad4f5de3364377451e3da05beb2cca0cf1b56d8ee2041a90e1450ea91cfab4bb43698b5a469c870916568f1ae855378;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hacd09cc8a4f02e24a7e7f4a5f65d803a866173dc4107bcc1efe8c26df8dd0fde7fd892a39d81512ec3d9ad8f602c45aba4d3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ade7cfdf79995e242f1cb56f27011325eb07b57a107693c3174542be04e0c4defa7884943609c92b3c32fca9b29a7aa3847;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26de38d96a5c929d30c6ecbee856be8a700db5d7a55263c10059fd1ac62703aca78c18411e2ce47d58ceead26acbfb1be640;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd387ada05532f3e3ad1a875daf10d833f113dc54451f85ce60084a376edec0cae0a33ca62855f730adbd361d0cc604b33850;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9edc25e8414e9a3c1aeb8d584d0ea6d1920664cc3207e978bdc79cb11fc9e4ea632873963f2a81bdf7ff1c505639bd25acb2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h541bd6325182051691507592e1f2f5ea2c270cdd7018c85b15aac7aac8a9ed8c41696881f3ec7223e5375547caebe9a47b65;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h57cf60e85b3341027f2fdabbb638d37f817cb38fb000fe6e1b73f325d08df0e63451b50f45a8374d1ff4235ba3ecbf6f0e91;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hacec51dbc75be92c139bb4bcfa901c9fa3a2716a3b610aa11de5574b402ae166cc2aa52da2f2794f3cf2057a19e2a892aa1c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb9bd9fa61ab68905e5c870bb9b7104e647fcb1f34b8453b26eb6df53bc87230f362d75a6b7c63040832393b050002ae582a5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c2b9e60e76ed0334b616429c1fd3f7e185f72525b011444950b24c77df95247713afa7fbb9f50335122f44a5d0e8e3ed30a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h89f652cb2c1bd8f70385486e03b93c0c3d3fc5924468a71ac8ffaaaeda963f53a0b3141711d7bc7d69f301b9b6c9641a7799;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha99446c208ac532eab527b4d4a54d2a2f08804bd55d99e6dbbf0405cce380404ec3585fd5eaa0627e243842dbd9f6007f7b4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc71c7a23c5293e7ee53f4ae660eb48ebb2addedfdbb96ab445569054db5f5c8f2cdeb0e9790814dab60ae9d39a5add59a811;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h19ab65cb1cf570dd0f6aa8693d3d98c904f49695d12af30227e789795e2f2834cd44241ab5fe57ddabfa9bfb1b17e22f92f0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf397907921f9398d86739edad92837d391c94222d7bc6373c872c824846de69dd950bb092137f74b2b4ad70b079e3b360fd3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he7e1b0e1ec9218f84176fe75634be3caf7d927414a79d62f26a6074bcd02bd3ec62591844c7e47bc8df8d4690fc2d99b73e5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9e0ad2df05fb03ff48819076d687247206f0b747d5a8017fddc77866c3725de867f126e4905b9cdad5126fa87681d16b9f2c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfc38ba570ffc3f4b137d77d3e9bd8ccc91a1cfca6099074ccef68545c6381df82fdfdbc3da74cfc674567344604b21753e97;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h359f67052ac72017e5dcb9846b043dc97a0440b782b181ad6e826a2030e38e2ae72e30e0ffd453f4e6b4a6d7a509ea510fcc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e6419312084b7888bb4e030e82add9f5b5b44d4eee296ea22f6278d914512f158dbc7c74b520009dd59198fae4a595c9eb9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h19a83e3cc1ca79a84a919f4420e4dbb989d0742693f3f0ee12834f61e88da7f00228193290a7d229baab02cef451607f63e7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf05d8349f6d94b0497fd157d47cd77514a9231d9b81000897143f3015b237bf0702b9b1e8897aec4f0ba47c3057e0e7cfe7a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h23afb0ad6faef2bde9b4a0ef5c11feca3baa0e07500608de6830763b6178e0a2f06169f4efb5a6c4ebc1c247ed97dc7ff408;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h98c7c4a165c3bf4034c9fdb62eb14804078620a4e541fc34bb474c737e2f8922d31941beabd80a6607e3fe379c6988176db1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2a7ed21fd4615a3a7518f38e15780cdb35627572aec2b709aaa73e2559038e9a520219d50006b70bf00c4bf9ac0f1175248d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h11df063c42f230ea6fc4527dd9eb8213dd978d407ebd8b337eb5d9ea9d84313549d963b1d4382465b65a2e19b9d1024e1827;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hed2cab93f7c272cd71b5ad21cb1538fbbe9626f41e2aa60b26dd1ba379a64c40d5b596a40aee9c6fd6aacc059c7769bb5c95;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1151065173cfbb520d9ad4ec051d9e8415db04f0e5a0439d153f60fa66e9c795bc8f1136ac0838d7e7634b1f2d48a6625fab;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h93e652a445dbbf7d2a0360cecd0f69eb691f38a127ba44180dbdcdd9e20541c07f8114189b64bc4cd476ba2e7b04c2102021;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5c01f2ca9522b3bc4a032076c7aab1ea323df16ad1aa7c778aee37505c378676f83a63babaf90f9b9dba6b41f6eccf704a45;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha2a469775a32852158cec3086f41d374a0a5586f557f780886213af806d1d54926ac4716ed5729cd3e7ea78f777aa1263a18;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5943b164506c04d847d805cdf34d7e98c24ecb5fece247113a3e141cb33868305113b5171bcd4e72acef3a844be674b08246;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ba37e90661a858997e2a636f0c1f9baf1d1bd3576b3eb1b9b5e4140fcce7d6b5178bc7c97c85471419faa021f28f31ff797;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0ba48d7bdb2872b99ca75c7e7fc7768ec62a1fbdae76944305e3b385e46647387f578d799417b48f25cf469f2a81db897e7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8b6ac87ca9821f39293587234e984f52cfb10b4c57ef2f1bdc8e3d5c9dfb20789b504311cc57b05a883956d2fa25c4332b6e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hed80685dab04a5a9c134e230bacc42a402fca06a38b62c3cccb1ec3e45bf46f7d8a45dae5bc9227592201ddb1172006fbdb1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3066f44bafb50d5cef3f9594b228e6869742dfa929cd46e57483a2aa14eb1caff02e31feb24f4096b0320dd0e23c1f9b0482;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e17871e02cfd32ac9b08822f958889574e651697ff611031ed5b3888e3d42ddb5aab7795382f93bc8e1377bbab3b91dffc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f848a18bd6ad4dc6b96255f544ac2acd6d1b02fb6ca53d2f4779a1e0c69313cfe03299f5213798445e7dc9b9f2a1e6d3194;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf68a148e1427962e03f438965e82aa04af2e05cf3eec73bc4ef812b760ff430e18fedadc590a55d141185b5e697a84caa1db;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf3b25e682e2e5c44f1306da3b63b28c5043fb3dbe2d87240973b2a6130866bc59bb13955e768a0ee3f2a34e98cc5ba0ffa60;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2043abf18d95246aa0649e980da891ab42d6fd66d3a7efecb5e560c06bfd87c67ce9a29ead63cc881e53ae7ee7e0b737669b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h95d21e5f463047c00dea7768f6e8a00ed580881388afe808c426742d10a10771b65a9468727a54f2cd65df9ff7d998d123b1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8c09d7c3dffaeca5ca9208c47a3a21a51f4ee9ed515d590dc10735478865e8551e66c4fd952fbf3ad748d9ed78993fa032f5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha83b2da22fc80747e4b2d8b8ac16503bd1b25d1d9681d60605c8467b1d8990e02df20a2c185fadf9f8792eb3e971800215d6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h269f052d28c3e243fb41e2538e8a6bd1dac721515b913df633fd4bfaae22e0ccea99f751a290378aa7195823e6e4529698d8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdd95a7475a9e94e900ae6ed8abcd70412eb378118e18cb83f50209f0d1f4271a4677cfe70f44e59547366fb470e34e4d4ee5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26476fd496de20dcfe350e72c74add712e73aba8a18f2398b130fb0fe8c46fb8027ccd1860a9a0884fc3c37d0d46505e1525;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h19583c13a5c2853084926f1f9e516cce3591de141b341d90ad6d3340fee04ada4b214e51ac4df5d6f5a6fddb703b45b2b61f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h55a4f2a3a631315dadc9e200fef6d547209eb736999d9d26cce7e20be7fb5858e8cf3b78fbbe3d21c287b3c3c1ffb3a02d0e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h91986e0014ab01ec7c65d09a1ab2eea56731aa8c90c25eb2eac39726302020693a2929f64ea053d8f0af98fd50a6b855aeae;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9fe64d4bdde10a457901d911db9396d3e694fd562ddc88828cb4c51ef84dc2b10e3c457454a45364984ed574788718db50d5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h201bc0ca906fd543bbf61a63defc241cd0044c1a96dca4a2e2d38080fff6c9c361aa91061dca7edd03afd9d61d53b68292aa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9e7a654e872515c2851560eb96965ae1cb110a74bc71ef6f17129d1b9a410618d34a0982e4d137775464d14bb34ea6032c8c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h781980a7bfba9286ff176cdbacf5d3de5616ce25500fba28424129a229764bb675809c1d52fbb9a2444f7e2b9c2c2fc99bed;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'had23dcc603a5ff51f352e129a54e3e918c69d4e9748b44f5b1f103d1d8cb82243417ebc4fcc755fb90f7c15b4cf1f525fba;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1433865f9b88ded39760d93d503ec6f89f3be4fd5d265117b36d08238dc3f3a3cb119901fab9424acc2ae94ce4b4b323df66;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h28f45ce220ef677a1ccec058ddee248de58200ee7419da324d9f32dfc00828e20b73d6bb9b319d9bc93b320b8a5a6e0dc4f8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he7278f03a46322feba8face36ab092fb309d138a55280d945f0fd7d0a42fecf1ef84c8d20b6d0c349bc7f8ce3f933cb437e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h40ec2dbcd874965c694724874653ff149e822d0ddf988c7a57ac7cfaf8e7d7f9056124bb8365ccfd56152b3a9ffaa40d4b05;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hafe347625046792ee358f72c8fff93e955735df2905dd8b3d779ffc691bca6e4815cf47585e5a821416d20fa482b860ab130;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h379d4d90c47dcc84af147db184e92fff488ba535847d06dc1afb69cd046f90c23f13736e9e78e2a1d45e5468aaaae5d20fb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h60e18f0a53aa4251fe023e2ce3b7a3bd484f17016994c65f3c4708a7975f54dbefea05062348281ab47372dc9cd86ec3c098;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6b2206adca4c4b2c292d66a92bf6076dc623eaa250562c8fb2010584cddfc068a8aae2b68fcd8f6061854d80819c4fbfc375;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd961f0afb36242f54e3a398415d61c764746f4a81e51338537b7877ebff6909f6572bde78b459b71f34ed61851649022b404;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he75441f082e8d74f7b5ea00f1a66231cceed79111c74d60a5fde522dbd1059a8bbc7efd16da83ec3db605c9842e6695c710c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8e17c820c57dae55efced591dfce5ea67945dab66f40b00363eda9e7e1b7a50db31e5001b2f67a45882bbab3031a423f95ac;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf3de97e6708c1386646392346bbf0a310d14aa252e443f2f527711e8485a5e4ccd4c9cf0d53d48d3ce5859983cc8d91343d1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a96b9182d3938b1e571d66bae88b7c81a0f12706f04a9e00412e196f96eb43e985b220ecefcf303f4a4a6c93fd3f16e65fd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8c36cf2a302bc21704d6b3754fa35f7e100ac84639ec7be7fe9bd1720cc92c89f448a55c9b1bb0eed934499ccda694318f8f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h59aec485a40af1f205e9fa8a8cb802f0c103a24824a11eb92ffb38bd60fb61200529d224fa79a42dfa3f8b3c836c1e46175a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h11d0e0135fc45f0109ffce5ce3b890d7e842f2de5640a7783da7074e9c54bdd2b6544a52065c44f5932936caad2cd4a24054;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h892e64edfb6bd192ca79cc6343e90188a04f4d0a1eec0f2f253bffb403d6c3ee5388e97abb6c5d4a8d0c4f43a7d6e0b2a6e4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4f961b9902615168f4c8652b7810c22a7fc3119cb84e925050cf18428f8628a18cbb394c30aff4c3744adea36e80e90cfb63;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3418ff493ee281956c0d7e27e2257fefd2d9fc7bd958e804ec1a6a2b4f90b596b436434c9eec5670c5a76fad9a7fc67f3124;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb35d711de4507e4ccb5553379ede2197e0c260b3f17cdf7975c9de0648f1d73aab584615a38c8ea8a411e4e39a3af9f8ab71;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7f53c0122f5a6b9ca556cb1dfb5c8c590a483ffc2910785d88a6471b7a3ba127c557335015e2d86f55fd72cef853889627db;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h10551d8eeaa3c6c19c61b504e67ffe97f1b514f67c68ea87231dfd5efefe5a66aaa58823447a9e36c387dfcde09235e73526;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb76883e8c82fea934271605706491f74fc8e2acd06200f9098f40fe70f446669dfadd69482be00b4fa0926cf641a9108312;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf5e85985fc0b036033a99a9ab9c7db641c407ec99fac5658b13beedbaa5f62d94f77ae673eae20b6db53e4a35bdc00856802;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbc00f4fdaf74c35e04009f756ebcc132a479ed08e5f2dd93d97ed1d88b84523d093f65c62bf965d880ea48d69e3fdb99476;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he478a441b149d118788fa00e788eff207f5d61bdf565f9ee13746bce2f1a6a989964fdf4a56b0627b9c4eb4249567ff62e2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf3bb4ee6d444701a5b3644a491e29551e1b269e9bd12b43b8ee8400cec0a2499ed937038591237bd04441ecf038f52e363cb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha45d8bfbdc2dc49174465875ea0ce641be27419c3b44324194116c01d314ffe2c1068c2a8f07a74408f717bac24366545017;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h77f173a77fd770f24870dc6be00ea4188284a2a46c66897f3e82437faa44806b2ae8a442b5108f905c12512ed3b05583fbaa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3273e3c4341200e47b5a63ce7bf89763cdf352808752924b9bb2351cd6bf9efcfd71f495dadb3dcf92fbc92a5d4855ae081a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h217b4933dc16aec2322d61ae2554bdb29fc88ebfbe4ff6a4904e879977ce3ff951c871b9ba780fc23d76c6646bb04e86d080;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3402c4135f9a5a4c0b0fb2e0129d1125e56967de188aaa535cc7cd13710eb7060e7dd2a58cb9480c6c9ba8b80b9f69bb716;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h24e022bd905e6d9a68572d5f9985a0156e4e6e1e4956a863b176c8c0da1f4b566f98867d7645a988a369a4a44951e1730747;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4e71b429a431fe97b090ace4a0b26c49b8505feca2b714e9436b4872d1f350ad34a552f1e89ada8a18dd1b32486037894498;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hda9e2794579bb0a0ec39217b88daf4c0d92a1a05fb1f9feb8ee5db6fb990056d5f03bcfc49b345c5ba5e231dea930636c992;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf188bfae02a798b0d929305a15f4d900e43e09ab8f4195fe7d23cbbb630a6d6e46649dc160b22c3ae3f644e97bab456b91b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h561cac70de23807ca8e04c24f0139abc5a3f5f3978672e67f1f288960df4543a3ce72cb04d4ae8cabf52a7c3b11611631228;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9863e92551018e81cee86828d9f2ea784c38aa6e75f080b090142632e6a9e526c90904fa4c4d7ce230bd2cfaae1f4be64676;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9287d7720cc368c9c373f90c74aeaf1a89e539d6c7f86bfc54ca5e03ceeb5c54a8e85d20aa44deb7f00e9d374727213ad836;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4d0029de9086ba8aa3960a2920fcfe141c5dfa0cb24d9c95a97205c03f7ffa4973bc44833dc39c33a9580cc25f8452136c9c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h36c3a8124be336bffaaf9bc600095711a24bc232f95243075765db83e3e9dd78eeb1f9564a9cd2bbdc13cfc6f3a11bfc267d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae7ed191a4e671534efa58a02cac471aef30749e61388825e5eedd8f7316bad3e14e560ffdfad512b7f74a188e5bffd19e68;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb19b41890a4a9e97002306e78111de54889551c91d98c8d1f675b513a4d8619fb108d653020917f7a2a827d5eb92769ba3df;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfc44f3c0242115044e3deb4521bc7946e7d17d955f339937b6e37d8ef66f4fa2160ef8fd465043a768bb3c7cc3bff3df600e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h227138ce059dccb85d174c9a2fe44fd7c9ab147f4b549048835a0984c11084ad9acdbca4ed65d42267d3580bedef983b9d88;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he5b517f830706bb7d4543ed4abae593e35807394d64788574972967fa05a057a25c71dbe5342b81093d08647403bc372d231;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a8a9e4aa3d03a8ade991980628e8adf7f6fb9b5ebc2bcc9d2fffdecb26b12821c6d668c896be9ffbeb24e5076fe2563a6e7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc17aa81900f004371515ebb3657349ae552dc4c99741cd2ed2a4d1a355b31450b2f0759db0ad9f274e5be056edfe6ad27b17;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1692591874f06df5cf55aaeb7b319165d527662bc46d5e1ebcdc0a2bd7cf51d059291b8732e623bc17906162f2227e68882f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf4aa745661baa8a90ac966ac44e289849a903c6a0ef95d362befd3d0a7776b3c9b2245af3d6bc928db034fe6293cbb1f0deb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h53bbb41c7efca0a94aeebb063ddc7be946c2f142ba29c5d2d815540bcd29b2c1a34dc4dc010df25ba3d12179e1786f706d86;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h35afb1383318c10e14cf7dcd7c5e67cc28fbaa1b333331bab200af6f3bbacd72fdd793aa14993eb2f0cb6c447e1d539b6b3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d2ece1274214468c0aaf005d54808d45f331a4e9b316c9ff08d9d9d6b96d8b2aa160423a516cb0bbb83c0f2f53682f47a93;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h62a5520676cbce850ebb0b591f41a15867f49ee8fa16274145ef407f2366e3fb672b295c033822096f71b0faa70199a276b1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26a9774a1cff4f09624c31e3ee630b667d2184484450b37daf8947e437896de53cf8d0c1871719cfde21a14fb8cf5d290e9d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4c708ab3719a93586a299a3d0d344efdc8b8de88f4f4a64b0e9cabadbd78c268c3e1356375f0ea302b13ad012e7dc682a8ee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h63db5c4ce6b2afcc8cfab269491450288e1cf739a31046da846a78c7e39d0dc4c2d3b75e5b64da5ab19663e8020e3e8c0259;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h66458d7a4e9460cb10fb0b87c73e7936e67b28b107caa12399d98314abccd13dd5f2e1c8cc059d14d8c5a4dcb872e9d1c85a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6725fe863826aea8389795b44f7759ce53ca08b1d7482f93d5bfd8dca72bd8a4b8b0f4cc16c890ac62f8284b64a072c3f15d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1b97771a0a84393381638eed1179a1f81cf95b3c389b24113dd3fe959eb591fa5ded4b7bb2af9c91ae2f4abb2ddff3b5cf71;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h19064130c0a86fae66d08771f0498102a8fc0b6c7e946ffda0c64423f1a3ef3f542ef2d0a9c03f7eb02d2b37d55b52e4442e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f2574fb85e31b9a6f6363e53ad83eecbdcc72d0d57d88fcba62defdfba2f9677332e6b47a0af59f150bad595360f7e517af;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hda86e9e92982eb91659992ba15afa512d1a40cebaa9fabfa9636aa4bd38b9e4d5b3ecf5e6d2417a198dc4927dfcb11e72275;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h94cc752a445ca94b9bebec5707d3920657bf8784e03e929405dc0dfcea1884ac8d51031808d28fc44ec740e0bf3ba01e61d3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he1d91af8eb9f8a48609b0f93c86fcfe6472446e789c7fde0f78583cf6383c494b3a1bfaf628b1b31075de82ce0d6bf9d7754;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d9251decd2c4dba07c8fc0a94233a68c7a5354192e1a964371f2630fdfb9901869f369a8e271f34144a57ea443b08513bd1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8743dc4c6fdb768d15d425f1aea881f5525277ac86a2ca9ea7c18765019f12db9b45fe6577105efc85d60e5ffa745091e8b3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf36412364a21f568e3e8dc1b24933fbf8dbb08ba341cd664c15dd5cc61b58485776644db8ed7624543b4811eb3bc8fe6aa92;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h95e64713838e3a14eb15a42be4a15e2600a37657178007f5c452c3660476a1c709edeee45b001a129006df0e58d7df58c584;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h48fee3f6d224340bbcae7d6bd811eb9ad86dba9d41a222ca83a70732f993442385d3352d05be52c5217a460cc29602d297b6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3fc18436fbe93b652d4652ec0710f16d12dfac643c827c3e163ea5d41028258efe8d15ca4ee3fe5584d18224977f2ebe398d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf4d675cd36aba837239da7bc2237502830b9b0c541af70fa454ed0bb8559a28cee1ecb9228b6e073cda88ee0938f4e316dce;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h18ee828e447c611483a874da014f52c6186b996697642e14be3b2d2158050ffcfb3cef1404809c453dad1d321bd04c3764b2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha4eb39076b9b4cb9f9d5e967cffbe6dcb975177e64cb9cc1ee00de73fb76daeb08400e1ee302d2ece069fa8e9064245c1a9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5348879e5e748ed45ea5af154f1f1936a69e098b1c13207d9e508335c5c30d46237c5bb285643b9d777a295f148e57dc89b9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h935f1d869cf0041e1a5cbb3ba4ac57c1177b5a6263aef426c8dfc4412a05f3b1f78753809674e409e84ccc459d867813fa1f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b18c00690b47cb6d9c0fd8c8d2076ddec188d0d81027ff2831ea2ba1a5f1e72e46f4abf36c12f8baf2da2376933a95ea673;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4767e6eedfd4c054317b73a70e3c27e14a834a37a80e32fa8b18642cab33544a67517bf15bf8304f4a7bcda2ae31bbd0e402;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he07d32a5fb7b0aa0e9fa0bdd43998c24f755e4a67541a176c7860aec8ed8b9563f5c77b4dba9273002b26d37440ef6951735;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hef46f6020d9ae908e8a69212a3dad8d2395d068489010f6089767ac7329ed2119874a9de2f494939a9c4b78bd00e8c039dfa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a43ab6f8c762378ef74ea45c5241cee22ff1c47b397062786a7decdf725466bbfdfb91d588c5bde8d7ab3f2381c516f8d36;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he990fcb09806029661557bcd346584a8409516a45d34d01b58015af4dafe3c18e2584b29b4382b3bfbdd5d0f218a38b86514;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc09eb39a1de2b3a75c29e6fe0bf51e223e17bf86a5fe55e3b651d8807e6e21811523fa44de7c98afaa9d5a5b4cb3bf5d1f55;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe604166bf798e2f31bc7814665018006e0393c80ec6cb7dfa12dd6ea6d9aa893ada6f5fe213471c3bc52ed68cf5057d341f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd28e4d146d896c444e8031558223cb6d7040561b0163251a8877b3f527942086f701b9eeb07a26655dc951e5253d43333eb5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h51e6019f34aa02db1b0b6de2bafdd1ce94339939781ac7a8121905bebe7a4cdb8df445500c367c59503b7b3c40448d7618f4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2508dd4297612cc469d47d9e098c752a49d54b277992931dba70539bfa833c1cf487f5e8673a9540fb7f053b367982ea2372;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d7c0252492e2e18bef7a3b46e5228f75dbfe0e2d63370cd39a915ee0787a7dc95f8875455f6bac4c7b4be1a7c4670b15343;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h74eef6d4ff74758601cc3150d65e55b9280228c038a35196b511c1c3f804f0c773e1afab4bd706e556f3c371644dbf62a7dc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a3cd8743eff3c49e7ad35833f7303f521c28d583d0394a388385f38a1223dace5c4d683e346849c3808d6c802de12f5da61;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he9b8509c43095082f99ac7b4b194a30f1421c87c1a09db4c88c43a0eb2ec0778183478769e8149e25d8f9a7942a9895bdf7b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcd0057c32976a433c6e991218f66501a49c219f3add0b5dd5a22b14bad1d7dbe53b1b483ef210ec37ff5a61c081be990f2cf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hee73b6d45486834f018cd6e44dbb397ebb5d9b5f8e15009c5e4b7f3a823f1995ea927d7c9b16d7f6403b3a73d5c7bea493f5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcbfaf83ce06b3a44acb1853edfa65a3c257bad8b9517f3bd6e2073dc2432a0bbe6d69f0864352308dd7a3c51ae83277d10a5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h11783cd716da8dd18d54231fdfff55566014d7f31d51d2984843584f44247db8c466f1d54cabce7174a310041b800d3040ae;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8de950be7a64e0a2bf26fd7381ad3ae66ca822cefbd287e82efc3f721d34b833291be7e30894a47ac65fa548ad053a193cf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha912c8a8780ab23fd26ae0fd005ab0969b51ef999cb0d1ffceefacfe74110dd42089dd369c3ecb19db40124e192553345459;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha2f10a57ec8bd8e3e832702e2a252a7c625c24b820dbcf6feb012f155035d404d9de2769c6e7acd6b8517ef3ae0c8a79e942;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5c8eac6b8a93f81d6c8f925b056f8bd527aa1ccd0f31e856d3702b66039e7084bb7c8da523f888763596b7d7cb4b647d0fd1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h254e9dbc7f85bb8e45bde531c5d8ca35aff992d79daba4512691167846399b74626d00fdbc1553a6dde8f60331a5f7324785;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcc019c58b164e9bc8bf78f8d95f84a979f9cbc46816546787fdb98685bd1e51c052a54cb77534f59a5c206e72972dd596781;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha593797479f89725a1c6bbfce176837e694d82e55c53e63b283ce49c2773e0cff99a3857fa0feb8793d39123883ebf5344fd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec44a5e2f7fd66f2cfc1baee66e9f782c2c013c14be51171d831f6faffe169f03b11b3459907064c73f0fa6cc3bd9a8bd094;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7535e631b5d7bc90555a3dd2f92e123131e61f2f963bcb081299d126d98bdf8f15e9b598eb77ba7bb10e092ebbb1d21daaaa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h40ed23788927f5addfd25ee86346e81b73d931aecd1ffbdd66198e90de0ffe77bc4a50020c2ad0b0e2cdc67b381b1e1cfd93;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9ce607ccdf5aafdd1b82a3a8c6db236decc73f81ec97a9dc1061c0c8c054e63fed5b09cbf6d0afc44bee8acc51efe6c3ea89;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a33005765a7da490ce2627cd37f7d4c50ccbbdb9a12cc7907a9eb0a2b90ca165a3f4a006431b07312c222f30052aec1ce9a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h826fa6548846f82a5bca6da83d2fb555e9e26363a6511dc8a49b2b66ca21f506520911e6b340bd4ad15e992a851f3755d8e0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h28da0567f73115cadf709069af928faeccb096c15a5db3e3b1d71b179041b4f1a03a2b7a51835f8f5ba607d5bb40a743de7d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb0c805f27d3827fbdf4b2f6d0c18d5479bd13be3fb6f8f6820e3289ce35fa0520f7d4bd6cad4e949080384e0c6601bf2cc69;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf347f26be5d96456180051f06217cd15a4d9c7ace04ae114590b73d4279fb8c5c59debc1e1b2037c93cbcf3f7c9e9c5e293c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h268129f4fbce24f2e0611b176514ccd4ac8a03dd5690c2e9a331ea3e5d672894fc2ef063aa90d3f6d44ebb51ea05bfd951d9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcd13535ceb0fd8f24cd57d189e835c01ba62f40d21615d6e8bd369f85fde467a7b21904d280f319aa099df12df8b5338cf2b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h46dc1da6c605fe04c3f1504d67e9472aa5dedc1f5cc082c2ad2240be77cf399266f48492c0280785b63ab353b0deb129d8ec;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf92f08151bf30ae6d950af61ba5dd33fc2df555c62cb944af787f681c2a0fedd6e08a45d087e25ddcb03047428dc912779e4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h61df6663380de42a8d91bfda13b83ddcec1894b943e2c2de436835a2d1960270cd4749463cc97db90d9ad074d10bc54ea96b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc2253d54d81590024c8fbf7a8cd6bb2ab52dcf116132bb6481c9305395156ecaf9848e0880b1bd91eee71285dcc938d21abb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0001df61eaaa10959bd764488a42d5039603c6dc864a63b621462f6847abf0afcb1ae0076cbdeac053433539edffe6269d6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0d018f50e452d5affa639e2eebc9a98ea9ee66719971097cf3cca3e32c0de9875958a8e545d477002156249ba356fb2081b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfea8c19cb9b11a7704a3992a5b754fcf8079e310a2446e63d9ce0b5f7b34979ef71f59454bd7b19f8a7cd7706b8633cd4581;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a586f245f6156bc80c09a6ff9eb54d2dcb1663f99af106e1528fc0167e7732adfd2c4d9d8571b599951fa1498963c144c11;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha3e745d8af62d3557b2bce8544af8c1375debdb725805da021b20a7b319d901c4d4c6c530c14e8af4677c6b708872c76e80f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5afda0b2ea63fc530b56d3a39577fa717d4189b2f5f39efe36ebece6832b7850cccf34055b139a9440ca908c923029bba678;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h45aad1429efc08ef768f5eeeaf969698a057895172f5faeb0f19ff7f267d58205dbe69a3e92d7589fd7bfb3cfde87e42369;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hce629e0dd61f8ff3f09ec86964b83038b881612add036cad84519c84fdcc818667c20fd6dfe26b1b4e8a2248e960b5163107;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h22a23d8877721864f321d84984da5a539d84db5e5e849e168327f0ea3bbf33ab54067335ed5698e6ca9e0b092a96abb8f4db;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha353784d381eab3f9b0b4feede3ab2ddab95063b344b6864c7bbd90dc600516e4a122264f3e14ea1436974af485525e5d27a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h754ce68f5767d3b92fe36987bafb0fcea2963115767910a770e1b07a080d8d70c8784733a45e6fbe2af73ed0b0bc26f9ec32;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he1f1719ae4522d3b9c951988c1c332cf76f226c9d94e8d5d5506f1f5020299161b69d8723e0183078f2f126082dd3ef42cda;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb48297dc537d23b550a7b13982ddeb2af3ac7f329d2e5c998f31edf94feac1acae1f17c0054b61bb5871e1c8809583c20f6e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h42664fef56514d02f34cfd985e45ca732d0c51761db951e2a9959c100ebf511677ceb780fe0411dad2aa7dc5c023760e09a2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha7774b210ff02557af27f5814f425544955133e71feb62b66feed399736c07e20d91ac4a938417b7c25656800c473ef13810;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb1ed0c6ef0060c7e8b911428fa0519b5e30b8766a6d43d746c4af1d28cf1a0494eb3c3f4d7e2c484925249660862e5b9a92e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ca3687b7c6fb2629a823da9644a7197af2d8af18d2e52bc2d94b94431724641f4286c7a42d6c7d8d22a47031c34b59f6c3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7bae5f42886bb1ce8bb1c46386d279f99b1c88f0c5d135a9139ead72a57292f417647abcb9f5af898c5cac8210e8422d852b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdde356e75954ea4cd0e57cb325d7fecfd8aeaf97d0a0f9f8726f20e8be59b4edb72582fa9c44f6680a8e2e205f44e3adf732;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hebc46c3d4d5610f5911e6619088a8b2145681f9ab46cca8c7a0e31b3a0c593f01fc4be142e6eb15167c2bb2636700948af2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb8de3f43f8fa18b12875e11bfa24feb17d2b7eea1c6b919e469cb37eb37db647e80698ee75ae74d20316ee65fc1545a61a31;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h265dc75ed924743c7a43b07d440b260470fd471d4cfce0dfeda78327e128474d0e48e1a4762029538e7c8774899f3e81d555;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h285dc00fc986765a910c407052fc353d5f606f3c82f10949ca36b427dd63149ffed8b1ff89ea5612b65ab87c34f3fa3b10b7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h49bae9d39f13bc036314878ea3523465062623b09c09852617b3ce2329982de28cc0b3388b3d0523b615ce698173fff6afbe;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcad9fa8a5eb53c5d346b902d51944e81a14c35d277631c6e216cb33243b84622e2248c845ee1c7bbf3fef1e95e8ca0b3bc90;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfd21b6b72995ac60d7607e49b3aeb17e5231e87359b7ac8d512e01f56cb4b931c7c11c4e8b4f1ff1ab0d2e5874e2ad4b0be2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1cfcc807fd0716f723f98acb88f9db391cb3f7927a089a2d1d3c553be0c7f18c45adb7ebf7733a4425bf12965f3904603853;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h78cefa0e41bf7426433ff59f393676cb701be05dd1f255543885be07a08e741532fac3ab6904071afba8b1e5553c5f0b2d55;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb928e1d16517da1885bc6a1220d689d875ef200067703140b2322e4dbea903ffd8dd401c54c7c88adbdb6aa2875b58990dc8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcc1d1e22a1a2cb700aa03ccb130df9f446531a732106fbaafade5eb045bfb81b8c1ad531076fb4f88ed0d27e68b7a64042e5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heeb434835d91ddef9898f0f1b32acef41508633c7e8eb44fa1e129a3fc7f5950b807271c676e9f057c5a5d52e281c8478b73;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h67b894816a177d11b92bae1e0f8d73d8b1f6ebe52dc046134cf2bb4a4a080950d8219215c8bf25623f1f59e40006605493eb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h338dced9ce2b1e54bb6e926d17d20ac1f8d3ec1e255b69b2dd72b6d32413592c549043344e54f83fa3ced5470a14917616;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4e7972529f1cc78360588a337fbd9d068eb262d012ee9a9e12e8f98ea7aa9a425bfcfa6288cef2f9d29e6e166fa5a89f276c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he24a3272f38d0a7c5a2b64c0ef22ecb1f40aa3defc8ddfce04b6c1b664e9f48280addba3feaa23bf5dd74426992e2c26c561;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha873b1e3b395626c21c348803f4c782c654ad03c1b0585bb62bfcee33c7ee05fe61375ad4ce6381c60476767604aebb33101;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4eced6aef1849257f1728666b760b6cb12367def7154865b829a52c93ef3f828852cc46d9b1e7a2f7839fd953718a51e180b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4159a8a1cfdfe39645a5d2d3c5f63ddd7aad915231bdf0bf150b2feeb9c556b1858b54742608410d8e43d1291b5aa3bf18e2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h775f7cdba8ab551df6460e885393d4ba5b693bc696b847ee5f298812d6722298b826203dd1968b1cf42707032d2aa5467519;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3c61ace2ee3152ac42805f060ed2c50f0daf68f47290546e7619d0f4627275e9624e8e5033a692f3547930f551fcc779a7f4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b580864e49573a1fe1aea89eda368ed4983d9d290fae7acdef648ca9f06fa2f49386beea66aecdd9469db50865426cd25ac;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a04890eeec353385d863483c56928d1b14f22a9923a17935766f82616de387e750597dc2bfd1f7bf52c20a4af5239e51992;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd23bf43a9a8743b7ff8a6d1cd7f4995bd609efff57077bdc571edc15ff87926e02313f9b732ba52927a47a9165f9b9367de9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haffa09e1ea25cd2e4d17621712bd352df316a160fc843547f8d8409dec7da29cfb60e440494c49fb1974f979b230f4726ff4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hff5e5244d7f1e38606c48e7237889bd3ff8828ba8e35804bc72068ced86fc165bbe16b738b70f2e4ad727a641f7d7df2ab8b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb8586afd6b4b9d6a2bbe34635260c89b27c12e2efd0f029637f048499abd98df615db333faadb99891e608da76f40704ae2b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha0d8921b9430422f0c7a9236795af7e3386b7e42e979212b94b4e4324fbf052a7528a6c40f06c18823cf4ac25f60c5484253;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h77fe7593c48071848f7ed414130dcf557135d866a3ccfc3eb1f3eea5184e037387a7d1520522d3df65278e8fe1d249efbb24;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb66c43c50577c27a0c4e67f42ff02f82a2ee1864633e63c5cf0fcf6dc7adb0425eb48cb21239fb3fb03b939953b924da67be;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9d508f274562a91ab27f62be0f155375401ed436007c6c5ad72c8ed8779c15cf824c7409dc42023c58b4f09cba6d4d618d25;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0dbe0edfdb1e7d8b4c73455e4ca6057b5100e1461c700ea480c9de658fc9e0de20e92969fb3249132e45fb3e4731e15b561;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4606fcee0799c22b6a0ac6995efd7109559d6277af74b36243d6f7c2bf6c4b742b23f28fc13c0a3001575d196ad54aabfdd2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h162e700a0e450a7019cc876385a05882e8c6214b549def5f00ac6e78d1fae64c7d9c037f791964b0b2bdab584a4280a3aaab;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h386540095b8c87766a2de960bbbc2b6eb2fcec8f4ff3503c66c2c81fdf0905bf3271a781eec11703473d4c5943fae4e4aa8c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he7e5d3d52262d8d8e3d63dd12e91194c2dee9501b3ec4f34a3d13287604ce9d0168523ceb623c56be4ced0838ccf96f8a0ae;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf02c1f0d407392f3e76634734e9ee158319ba96922890867d1bb2484d0f1cd409b5cea49c6e75ee0bed88748bfbd338e213e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6b57230b2daf998fb09c84198c7e5d860d7c06d507c3e03721ae16f2a3b942709e8dabae4aa7bec9a674f189c373103e719e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e1cb7fb84bc2d0f5baf47c48f719ad1e98785844aaeb83eec73d196ab38f8ff11d24d2d51a3b04fb3343b563fa903018b0e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h62b84104e41d0309a70d1cd1fa86c5908311569e3406b904a3a9b964594e4bf2ec03c91ef940ada8dd7b029d49da60630380;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h73d1c31b8a999a5811b08cbbf035faa64f83097fe23e960daa29712f83880ce05f2cf9a6514f0990967f05f982bb5862d011;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf42a67fe63ba845156434fe3d9ccb24588d9bcb53f2cc36e92898e6e8b96a4995dd06b171890c89f8a925890fb2e1c8844c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h521ecc3618f9c3af2e3284f8ca7a95165263299228d243cfedcaa79586df5da13c1e8312fcb35c71c057ebc6b77cd0941ba3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h874c97d3633468f2a762204a61f350fb2b0d92454969f84ffbc87be4bd2e65f71c8ad58f7e6fd659091fe4e5149e5ecc73da;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h22a9febba1474728171fe3cb154353e8bd5d8e108c818b4f0519eb48604e71b61448963c09f6d3e40bafb7742f82d78727dc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h47fe63e77bf39ecb97493ed59704f4860ce18291294a9497192db916a7c779e9ddbf534c91ad78412870167df77c76cebbb3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h614e0a7a9dc70bece1a7083079d918ffb27ba4da0e1b27ed33022b7e832e5b82cf20555176d243839bc4ac5e979694100ec6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd3352d8d7f5d7521ddc2231e386a40efdcc801dc3d39bd586c900ef1c04108ec6ffc9db3723a81e2f00f4aa7bc54d65a7469;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h92c7cfd745cfa9ed1c3f66ad5bbbc7523edf9521d815c7d1c7a2ba683bbd14bda1c1a60a7755bb182107714309a446ede426;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9bf29db38b709302f3fce210f049cb9bd84778e7a2e394edae290b967d81cdf46b9bae3b36ef1617aabe49b0214566f8c6fc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7564c0856f0191b512dade12d85e576acca235cb8f6123c3da7c6b549e196f60ed2439a984c4ebdf977dbd5d9173cfbfba87;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6b1653c7d9d20cf58a7e18ecd6946e0d74fa17f75e23ce008381b468943dcf59d30fff359fc5208f46ae2473281cf16813cd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h39f3fa3c7517ec9c854541bc3b3fad65a5c468b85861e9d4edadd9286f0e7f66b504080f664f97e4b20b2c6b3436dc8100b4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h582bcbff1bdaa9b5058dfb6b3bcbf682bfab2148a79cc5e091fc9b78b66d90e27f92e05ae68f9b35c9c15c93243fdda1a6ef;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdf96250c02948e5ec9c607ca525b04e834626735e2723a11a16bdd8de302f68c0c6fd25cfe3be19589dd92f17bf580e89e64;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h87f847c1eeb2f7ec2b7a5da75bc9ecdbf516738ee73b0ee4b98c3e648af35eaad8f9ac470bf00ba19fcfc808519954661921;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h11d2a389bf0d15983d3e71eef2bd50815c69c23aa869ff3442f2c3ee1a20e83b55f9676c0d2142099cf8ea1f1ef92427b6b0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h843cfadc7f8ad2d2541d2388da8461b92e5d4498a448c9999cda648ca343a466d26133769fb18beb0c092d5910d948fb0528;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h418359ec778d9bec25df7c5710845041a7d0aa394139c3f6d8a022dc9b4f6bb016a95c232b744b43eee1136a841b5334f96e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7df41dcb07eabf98ee20c1be877da4efe5e0e3c878cb2c5d4fe07329325c92bbd363952162bdcccdafa13e4e13f0464edaba;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h211da348f67e50a685665606efc7130886ea5e913423a8e49a7e30bad23af9f9b0b641ec7c3147afa2b22f11cfa83f975814;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdd06fc467a95a05d1c93569f4919908c8c3f42f99296cf4efac4bf69e4a2cfc326239bb2fa3117d02ae7db02325c52f98f0f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1579bb27cc5b5614b94ef458809e18a22e2d866a3bc042fee1ccd8010f74f48ff7120cb26b2b7e80d85d7d91aed7b2fb9385;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc3da6910fa916b19ab09ff29f86205ddd4fa8c20f3ca290b5e7d0b875af11ae8382aa990bd00595c84b6c24bf2358eb00fc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfafd848bbafcc0ba6c6f6556bb2d37b966675a10d5bd04cf6b8f47557687ae3d84e0dbbafdfe4ed95ce1e2e88ebbd2761b50;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ba98c3fb250132731ef48be26d2c2feed692ced902f985a6d4f53363bf233a089148a86993b7a2e190ffdf5c35b73442a34;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf728b2955ebd5dd715e96680b3302bc85c2e748b693131cb7e522d16983a86922b6c1939006569ec0ea215b90e10825a571d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf3190c6c21013f020c6d6d23c760f53a86adb76850006c4d255d32488b85a78108770177f94823dab5edf5978d2ddfc96b86;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h796fc182e24cc605b097985c9f98f05186edc268208a501272ae86c479e9e206f43b79d6b399b1ea8740f448854ef1d57687;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha894862979be7b69abeabd2e98a68c5ae9556b278e5fd6f2c6b30ab11ec8a8964b692554ce51f1ab8b4258a9aeab9735e89f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8aff5ac8fb74d6831a048935ae98b5db158543089fa89e38adc0c1ae6f9d3502c579f0a590c4b330629c8178c317885d21a0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h89972443bde9af98efd6c435186fc061a37dac48153a66c6eafab190ab9ceb9309d1388e124cf3c83dac17175935b2ae3904;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc7a06be4ccd4a5690b09fbd9d72de0c5ca20919f9b950e328729bb35d203bf582f591123a1722a05557088c89c2b11e7b769;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h41f9828fcdc10decc26699970d4162209db1845e106c4aca985353c9c30fe76e50542f23f907184022ec532e61158d81e408;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc769cb634de467d9c1e6f80e898dc0df5ec64945274af46773353ac5f9e1526e74b3497a40f283315300dfb76aa3ecf40e16;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h25a839991e582e9b63bba20a45cc7232e2ed141de0bd9886e281fd51f819687d39a85277284212e1ee6d60c7ac2680a2d24d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h482452fcc7678c5786b7ca05c9c993e314998c110e372d79d230bf844600d376df6fc2de748a409ca2a7049069579eb2d422;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5839b96d08909ffc9fa53716ce98960efb46df11727c1cf3342ad76e3dc512f1f1d55f2d711fa105e234fd1404fbdd206c73;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h549e8b425770ba5342e13fb7672afc0b6e5bced122503ebd004444a8d277f7b7bafe01e822f045288d5fbc593235ca5244af;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h37290a616e5b5756a48b40468657314080a71bfac2557c51f30d867cc4982bbd586a9af22b352e91a1d44e2f53dd8fb957b2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbe7b02936d9570da5f7b08341c7540a5cc07f73607931b2ca9863d1c191fd5c138359e0ae8d23fec88fe0e4036f56cebd715;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3ed28b703cc53136f06c0fd7542f1b293c8779c8b646dfcc1964b3d3a6b0d146f1cbb26be6c291349db8802e19c6cdb6851f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha24c08ce25e47bd6452524ffde93dc8cd5ee2a99efd5af422da8b77501922de3bab278408fb5675474a39529324732398582;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h13a56c6dd6d602d582ad09325bf36b476057ea133219854446af8851cce8558cce01899d8bd747895570bb5cf179b449a781;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h38f082b0d33d23596603e0702577076d4ad9e8964b26c95c18c4d549b22858cdeb12741ec799ad36932a4393255edfaf3cbd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d104b7f41eba9b1afb99fd76d706c86af80fb0cc56f79da78d39ee2e60de650443c269fab171fad55a5fc562c7ec5ab0193;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcdf3f6a86a1b5d247fe3bb28b3d8548bebd80cf2120f166cb4352494b9c696ee9e42dbb3b3edd57b81b8e664da43956644;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4bd3387b49616602e878cad740b4e251b8f5ea57dc61598c05d3c1911e96461cf1e6537f5b11687dae3cd9307066b0a58ff4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3ddfbb766fc96e6b569c22fa700ab9957c65b26537eabf93ac4ac345575fe895db9d7e3214596cf114b5a7571e96a55d7f24;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h313a2bff9073c62385896b414379e3411537b2a4359a0f5752fb7228516bbd2973de81a672844b8be8f2623771c3e998884d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf4674dfac0982b3751659b31671e64d8f2e305ea1d0251cda9ff2c73bad71f69d4bf89d984d9655da73968ccd3a85f69d36;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a7f82b37a8f9a75bb5c54ba345b06ec48d376dc5ee3a12f812d20480fccd78248813f60ad3784753b5bd2d813fce184c44d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haacc48d770f3c906434f9468fc29ffe861d1e6e9fecfa17c3e777c0ce630222130da589b3f0c99543d0c4eadc6e281ab407a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd3c178a82c8d40c6bbf04695dd0de6f7f9a39337b67b0aae5b68f06473b9912cc1021ebcfca3942402703329dd6b0a5b2a8a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h563f78d2117f2dbd9658307153894c5bb6767db5ebeb9600f7976508f0ade1febb522f3c097fbec371dd031d9caf4854e3d2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7566121a2b6a01ac8c18cfb2e9129df6a9b5cb1e701833f01c6382ac92d9dbf2043cb7c15e332c2bae41b5bdd58b9819efb6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbb3cd61c91254acc1b48dd98d607f7b36d148b06b1025f7a1da52cd3a9ea37aa319215ad29e6d4832bdd70438c9be2e48b02;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc9ff0910d64c395195badf7ece726d97974945f8e2e896b92cd525f6a9340f4b0cd85cff9684e79fc55be4ceff02a60ccbd6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6c99adbc1776ee5e3b8acea70e08694fa27627c168df5c50d526c9e161e71efc33bdd398096f762c4b45f9f67129c3fdb567;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha0ec9522218166a42be2038db1ffc877805d0633c71f07dc68564aaa75e4f4409020096a4dce473bb6e376f8154977da654e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h892e632675cc16134a65805e1ce2f14cdf3bbe36f63161b6bd524b6cffd3e43592ac4ba87e7ff566721a07a3d38e374884d9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b1f970f5ee91e34ba3d1922629596b4709af7a9b11bacf25b1c09056372b1267922647979d10a34c53966e212aed26983ac;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7eda2072e561642970d2311faf4a981bf9d86674d2a347a594bf93da997f81159327c51f598855536049a6829cfac0d30dd4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h96273a514f2a5b19c38e58c9d5c33d4a52a5f433d469889d399b0440073878c2a23d179b7ac24e39fd6b9fb4cce42c1040e9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h515b9bafbdfa6568cd8be2a3259ead9be54bf60883b8c6ab9e7f6fd0b25aca20f00269577a4b88bbae2763e7b3936f1550e4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h48f50f98c9109a429419394d1d2898d2459a54294d3de07a93a9cbf3b106b6490288cbddb6549bbfa3dc5e7c2873ae15ce9a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha0bb236f8e044033e048103c4a44823b52fb09a833867067e4f111339b6d2bb9f7957e8e2e2103a76a2ade954f9c2bd9576b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd3ef96cfd57a81e5f725945a91becf0a3484b5b832e13c9852d5396866e00bd5665ce3c9a22d8628ed6ce4e0c2ed575892ed;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h87481eeb6121e4d018a03c5e99cbf82458192d2a3bb14dba5a8cc674f8c855758348ae466bf2a858ffb65e3f354edc187d20;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc76273545c772f025226c06ff90db82613125dc57a2b163ffc4fd5bd71532864af34229483aa89bc902d3f1e87454efbf022;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd37fdd4ef7f21c1db04932171bcd8eee962a5a72cde0a739419489430665933314fc1810d0908f24b743c11daef416fd1ee9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb0e9c060e162ba62c306128262afccc0901cf57953d1da518d0a4bdfb242500c8bd0d100f5fd53a1633e4be6a61cf76ec96a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h50ce486f671f8970a6aba2007cf5c1c08104611b3284cb561c6b962af318aeefcdf285ea3ff0582b90f7ecba632abfaf3cec;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc400e927c5fcff3b43b73452a5b6b25e988a2fbce977c3f8e310d9f1d98e930c6192d0ff2e092096135997b580506c4ddb01;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h63a4f5774dff5eca1fb0ceb548af2414e95e4a3208e06fddb12fb98cab94ae9ea7bac86590c6a48cd4c5910a8d03d3ea41ad;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf097a4c0b740a9184dffff18b710037002386f7f95d0286cc487d77f8a7a6b1ce0c90ae7b36de2999b1f3715f31196a8402c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h994f3220a756df1dce37fd392b5538ea463a20718d0f1e16d857c8a4c2f20cf7ac57c3aaa5b30b8f4e352153f0c28e86f195;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h399c46adda50fb93191e35d468919a1ac7b1c37c5f0f7eb8097ebaa4dee283fd969af9444f9ce39ef73cb10d46f66bd6796;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8fe6dfc9c089258e16538b529a6ec264925f88cf444a6e3771c6be2c2c4f642b6a1044e501bebb36190e21770e884ee44528;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfccbcea7dde98d7b9f7151f17f6d0a7072e90ba6aaec8f8a8b694d6dc9f30ca6f8f42307bbf99c475e3e9deafda510277f5f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h22c22da46962eb2a932c156b30d0080e63b7833847331b9dc21c14e8826661e7895660f7b126b2c2e3ba271917bc6e2e194c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1ce8cb90c4ebd328d62106c5d997099aaf7f2cfc00537a985f5e75e73162644d95fcd95bd29e3f56e9cb053b87c2dcbea95d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h481de9bbcc5215d8df5efd18ceb09cc4b934fe3a800ab0d4c2fa26f9d4a0c3bc7d7b0ec1b421df313a2a6dadb74f441471;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdb1c7c9e50bef8acae21048bd1c872bd8a807ce2fbb30a117b496d8afbb85c5f5528799bc7aad7247f943eaffdc4047c23bb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h927d25c56df0ce532386e262364c11a0e9a909b8e828f90178c4c2676720e2fa3a582f9eb9c99bbab59caa6d10e843591b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h87553c915c8012da7119fc625190b9572209af39a01517290c549a59c825d420a2c75b25e83367ee4b6855373a3ade0e60f2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb28b200b91bc4a9afe9ec59024ea326212c457354b4ee593e53339f6d71bdde6a51b03f7ff00ceb55cd877d26975f5ca3697;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8e2922b46e2f522d2617d78d36580c87e70e2b636f647c2ba9b5f9cdd957bfaee946c962bb1a157b8889185bef0f38438fd5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb1c007c672350c66bd5c1059ae3553d94bc4862d54650356dbb60e2033a4fa325aa85b939632ada22deea26e3ea28a2aca3e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb5ed599827171e361b87c7e35b69141daf66cf968537fbb8afd9f528665e1ad85886bf0695a8ddaca6ffe08843e3f4bea416;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h869b5609ad228602b349525754ac619ec08808164d4c2354beade5775bd32587c95d556f20ca4f822553459e7abaa662f546;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfea1718a9af1812591cb4b039def7eeb8bf00c77d7b20896071918c49c2fd5e19ae70a67c4226ac0f795c2510ed3045f4e40;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcc85e6c07efa5bbd77d58327d66dae05c163b79c3e9495ff41f3cb08582e2ce5893347aa6f21efadd997bedb5269e7a55729;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h338191f358d6b46f2f225eb7d19edfcf5396f1d81aaa4c2228a4d97098ee91507edf8c8281717dc18194f8d50bf177b98f48;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8dfa4167e5cad14730c6b43dfa1fd785640a45732ee46862fb977d1c5c03a1114d3ab7dbd6fe7478c593a74425b0e75ebdad;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6878ec5e31d42a67ae5592ca35c2d105cd8af1c8a0e08fc7f2515a894c459052e05bdb9436dc443b3f7b3a476b3769a4b6ca;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcc88169eadde139f4efefc285a579351d968454920eb50ddaa2aeda6d46575c6382b5187447b7b3158d8866ddadbff930109;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha21223b74a00d2fdb032060d0578196a1a6aced21de34cb53012e456a42a5025fd1280cb6c9c7b5520286487ba5d13c5a11f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he81adfe23d17889667148b9d9ae3a0828f0e266e1db76ef2a1273d04a7a98fa699d56796072f613381ec754397df32500dd2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc64ca1d30f1ce5676843c5b74e63727aec078a33649011a2275fa05f685f5fd2d7885feac732e49260492efd33546293bd4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h83e52b82e413fa02025277a214da0201b45f0ca160f18ddf6ff2b5241af248239d19baa99a0ea277584a8219571a6bab5ec7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc597475910e7e76090dee9b8f2ff9eda3ff65237cd5cf3b744a9ff6dd1ea45cfb5623caa6fcd522c90c6529f2d8915b5a8c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h32cee62f3c724061adca99b84cd767fd3e114817f30d405cec3282373347363d515ea0db9166f84188c69f3d03d86c8ef8f8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf32bb784350848e318e3bee1bc1b165482348ae1461a55d49a151676032e053a376811c411f0442f8727f996719f6423584d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc663674663662ab2515c83ef8234d1b3ce4d60401d6ce65993f4626f6ab8229974e359a45a2985b711cb8cc833bd45862e0b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a875bc30965e34d92cd172231582637108a30e9c1dbf87c674c6dfad7652da2705ed496d1fa2bd27e587996756ed3f5446b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26796a932eafd071cbd243d8d7f61ed8ab2bf2f29c37661d4bd2177d3d7803b5a555ffa510af310be1a2305ad43cd60ed780;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha05e688ef64fdccfaec53aed9054064b028c651e414d11142a88826f0f88921b7b292d565303c93d903a5039b61b8fb6932e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h85cc2149e0b4cabd149784e6e5ff8756711fd4e8937124e6b76cf7645d76db09ff0a21caf4d19070b6f5409a78f1cb6a0fb8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbfd9d97b0499ccd32200852fb8a842b09fcd2c7e73830662e3b94fee96f2cd90c212d9c76967a14153a93e16506ba82ad45d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf18bc8b56d09165617c263714e34bd2455d2e52420ace4998beb1915064f553409bd0076f91ca5e37b6b31b96fe5340a6eba;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5918813ddf65ee867238331dd1643bddb33da02c510903b79b1ea1e28c34255564f895100a43a5004691d45d053526bf644b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2452642fc36cb794f0fe3d5f11b0393c94de62b9a75dc860f19df652fdf9b2beb22ae3dc9dc973f51a0350dd6bf3ab3f3640;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha1a4b9a1c6a5501e8ea44ddd06523aebda66699312efcab35a4804db247d4620cbf2df21e3d10d90c0c1a453d7460f19f85f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf87922d07a01e2d22d6481a2b9a336a5a3e9f8adee6619c14d3192d3f6fa3f6219f30ddaf459a1efe669ab389c9f1ecd7dc4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2e60cd1bd313c48d33a317a1bf047d493d51da74f65ffba097f2f353ae419815284664bc82632c2cb2f0de1b4f4a4703dcd9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h68fd90d491899586181572ec4004ca77cab5ed1545752d1c86c59a2075fe0d14e93528ccbcdd7c63b6166c96f69dd9af86f0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2465ff7557f07701247ba98c99d2d6b413d219d7fe74c45d9f85e62464d28cfe1f66f8ff20bc793fe5500d1e425bbf1a0a31;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4dc9be21885b1d03f084d044fcccb26a644dab8719713810545ac391917af643439fad0dab8b4efb0d297d55b984f5e9ec73;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hedf367b887752530fa3fcefbada6a8dfc2dbcd0e9896e26581a88471e8594921f2522042852a27556dd663a8f7ca088cb106;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d338d9475013cf1adb4741bb367395a33378320b82a79fa05894b10d16dabdd743a21c63f0ea76dab7923ea1b4604a1c9db;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha795f031cb0438e190f5ef49f040dcfeaef7fa214e6896dff1cb6d63e11c8b6e87ce06c4756f8f1bfa42002843f8f6c756f2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h41c845c23a307822418dfd2cda42a6fedf22c043da4b20cd391722488b1d5eb2efe1d0b74aab7fe0dfce23abfd10b16ea0b5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha4757bfa960f0a0f7f2aed681d9f99ef2098f60f81d31c30cbb0b762fc9c1578d0d0a1c888dc2a716760c6fa65c3b840bea9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c9ade3ec6de723a07e4e5df8dc4b243c429892f54c8737a5c048b2896d97f95bf7de12a87c6326500a75e4cd036b4fc2318;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1b5295a0f290b68dbceeb900f5c96b40cfe190c7a9df990d5dc498b86478f974d0f5976602060ad89a8e5a34ce96da36a157;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h624227b26bd78436b5965416fe201618fd876bb1d5b138555e9942c9429786d2ac9d0bccc4360ad1beda4c8dd8b9f56cd353;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb7465dfce5891394808aad17238920556db7142d460f3133de19ebe0be820ebd30f28805d7b9d86aa6160e712d10d28e1847;
        #1
        $finish();
    end
endmodule
