module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20);
    reg [485:0] src0;
    reg [485:0] src1;
    reg [485:0] src2;
    reg [485:0] src3;
    reg [485:0] src4;
    reg [485:0] src5;
    reg [485:0] src6;
    reg [485:0] src7;
    reg [485:0] src8;
    reg [485:0] src9;
    reg [485:0] src10;
    reg [485:0] src11;
    compressor2_1_486_12 compressor2_1_486_12(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20));
    initial begin
        src0 <= 486'h0;
        src1 <= 486'h0;
        src2 <= 486'h0;
        src3 <= 486'h0;
        src4 <= 486'h0;
        src5 <= 486'h0;
        src6 <= 486'h0;
        src7 <= 486'h0;
        src8 <= 486'h0;
        src9 <= 486'h0;
        src10 <= 486'h0;
        src11 <= 486'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
    end
endmodule
module compressor2_1_486_12(
    input [485:0]src0,
    input [485:0]src1,
    input [485:0]src2,
    input [485:0]src3,
    input [485:0]src4,
    input [485:0]src5,
    input [485:0]src6,
    input [485:0]src7,
    input [485:0]src8,
    input [485:0]src9,
    input [485:0]src10,
    input [485:0]src11,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20);

    wire [0:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [0:0] comp_out19;
    wire [1:0] comp_out20;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20)
    );
    rowadder2_1_21 rowadder2_1inst(
        .src0({comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({comp_out20[1], 1'h0, comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], 1'h0}),
        .dst0({dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [485:0] src0,
      input wire [485:0] src1,
      input wire [485:0] src2,
      input wire [485:0] src3,
      input wire [485:0] src4,
      input wire [485:0] src5,
      input wire [485:0] src6,
      input wire [485:0] src7,
      input wire [485:0] src8,
      input wire [485:0] src9,
      input wire [485:0] src10,
      input wire [485:0] src11,
      output wire [0:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [0:0] dst19,
      output wire [1:0] dst20);

   wire [485:0] stage0_0;
   wire [485:0] stage0_1;
   wire [485:0] stage0_2;
   wire [485:0] stage0_3;
   wire [485:0] stage0_4;
   wire [485:0] stage0_5;
   wire [485:0] stage0_6;
   wire [485:0] stage0_7;
   wire [485:0] stage0_8;
   wire [485:0] stage0_9;
   wire [485:0] stage0_10;
   wire [485:0] stage0_11;
   wire [85:0] stage1_0;
   wire [154:0] stage1_1;
   wire [197:0] stage1_2;
   wire [195:0] stage1_3;
   wire [240:0] stage1_4;
   wire [229:0] stage1_5;
   wire [169:0] stage1_6;
   wire [161:0] stage1_7;
   wire [238:0] stage1_8;
   wire [240:0] stage1_9;
   wire [179:0] stage1_10;
   wire [170:0] stage1_11;
   wire [156:0] stage1_12;
   wire [78:0] stage1_13;
   wire [30:0] stage2_0;
   wire [57:0] stage2_1;
   wire [53:0] stage2_2;
   wire [83:0] stage2_3;
   wire [88:0] stage2_4;
   wire [74:0] stage2_5;
   wire [97:0] stage2_6;
   wire [88:0] stage2_7;
   wire [70:0] stage2_8;
   wire [91:0] stage2_9;
   wire [98:0] stage2_10;
   wire [81:0] stage2_11;
   wire [111:0] stage2_12;
   wire [51:0] stage2_13;
   wire [26:0] stage2_14;
   wire [11:0] stage2_15;
   wire [13:0] stage3_0;
   wire [25:0] stage3_1;
   wire [16:0] stage3_2;
   wire [24:0] stage3_3;
   wire [33:0] stage3_4;
   wire [31:0] stage3_5;
   wire [44:0] stage3_6;
   wire [37:0] stage3_7;
   wire [30:0] stage3_8;
   wire [42:0] stage3_9;
   wire [37:0] stage3_10;
   wire [53:0] stage3_11;
   wire [46:0] stage3_12;
   wire [33:0] stage3_13;
   wire [25:0] stage3_14;
   wire [17:0] stage3_15;
   wire [4:0] stage3_16;
   wire [0:0] stage3_17;
   wire [8:0] stage4_0;
   wire [11:0] stage4_1;
   wire [6:0] stage4_2;
   wire [6:0] stage4_3;
   wire [12:0] stage4_4;
   wire [14:0] stage4_5;
   wire [15:0] stage4_6;
   wire [18:0] stage4_7;
   wire [12:0] stage4_8;
   wire [16:0] stage4_9;
   wire [18:0] stage4_10;
   wire [15:0] stage4_11;
   wire [17:0] stage4_12;
   wire [22:0] stage4_13;
   wire [16:0] stage4_14;
   wire [7:0] stage4_15;
   wire [11:0] stage4_16;
   wire [3:0] stage4_17;
   wire [6:0] stage5_0;
   wire [6:0] stage5_1;
   wire [4:0] stage5_2;
   wire [5:0] stage5_3;
   wire [3:0] stage5_4;
   wire [4:0] stage5_5;
   wire [6:0] stage5_6;
   wire [5:0] stage5_7;
   wire [11:0] stage5_8;
   wire [6:0] stage5_9;
   wire [7:0] stage5_10;
   wire [7:0] stage5_11;
   wire [6:0] stage5_12;
   wire [10:0] stage5_13;
   wire [7:0] stage5_14;
   wire [6:0] stage5_15;
   wire [3:0] stage5_16;
   wire [6:0] stage5_17;
   wire [1:0] stage5_18;
   wire [0:0] stage6_0;
   wire [6:0] stage6_1;
   wire [4:0] stage6_2;
   wire [6:0] stage6_3;
   wire [3:0] stage6_4;
   wire [0:0] stage6_5;
   wire [2:0] stage6_6;
   wire [2:0] stage6_7;
   wire [6:0] stage6_8;
   wire [2:0] stage6_9;
   wire [3:0] stage6_10;
   wire [3:0] stage6_11;
   wire [1:0] stage6_12;
   wire [5:0] stage6_13;
   wire [4:0] stage6_14;
   wire [1:0] stage6_15;
   wire [2:0] stage6_16;
   wire [3:0] stage6_17;
   wire [1:0] stage6_18;
   wire [0:0] stage6_19;
   wire [0:0] stage6_20;
   wire [0:0] stage7_0;
   wire [1:0] stage7_1;
   wire [1:0] stage7_2;
   wire [1:0] stage7_3;
   wire [1:0] stage7_4;
   wire [1:0] stage7_5;
   wire [1:0] stage7_6;
   wire [1:0] stage7_7;
   wire [1:0] stage7_8;
   wire [1:0] stage7_9;
   wire [1:0] stage7_10;
   wire [1:0] stage7_11;
   wire [1:0] stage7_12;
   wire [1:0] stage7_13;
   wire [1:0] stage7_14;
   wire [1:0] stage7_15;
   wire [1:0] stage7_16;
   wire [1:0] stage7_17;
   wire [1:0] stage7_18;
   wire [0:0] stage7_19;
   wire [1:0] stage7_20;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage7_0;
   assign dst1 = stage7_1;
   assign dst2 = stage7_2;
   assign dst3 = stage7_3;
   assign dst4 = stage7_4;
   assign dst5 = stage7_5;
   assign dst6 = stage7_6;
   assign dst7 = stage7_7;
   assign dst8 = stage7_8;
   assign dst9 = stage7_9;
   assign dst10 = stage7_10;
   assign dst11 = stage7_11;
   assign dst12 = stage7_12;
   assign dst13 = stage7_13;
   assign dst14 = stage7_14;
   assign dst15 = stage7_15;
   assign dst16 = stage7_16;
   assign dst17 = stage7_17;
   assign dst18 = stage7_18;
   assign dst19 = stage7_19;
   assign dst20 = stage7_20;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc2135_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage0_3[4], stage0_3[5]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc2135_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[3]},
      {stage0_3[6], stage0_3[7]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc2135_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24]},
      {stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[4]},
      {stage0_3[8], stage0_3[9]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc2135_5 gpc5 (
      {stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[5]},
      {stage0_3[10], stage0_3[11]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc2135_5 gpc6 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_2[6]},
      {stage0_3[12], stage0_3[13]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc2135_5 gpc7 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39]},
      {stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[7]},
      {stage0_3[14], stage0_3[15]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc2135_5 gpc8 (
      {stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_1[24], stage0_1[25], stage0_1[26]},
      {stage0_2[8]},
      {stage0_3[16], stage0_3[17]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc2135_5 gpc9 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49]},
      {stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_2[9]},
      {stage0_3[18], stage0_3[19]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc1163_5 gpc10 (
      {stage0_0[50], stage0_0[51], stage0_0[52]},
      {stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_2[10]},
      {stage0_3[20]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc1163_5 gpc11 (
      {stage0_0[53], stage0_0[54], stage0_0[55]},
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_2[11]},
      {stage0_3[21]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc1163_5 gpc12 (
      {stage0_0[56], stage0_0[57], stage0_0[58]},
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_2[12]},
      {stage0_3[22]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc1163_5 gpc13 (
      {stage0_0[59], stage0_0[60], stage0_0[61]},
      {stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_2[13]},
      {stage0_3[23]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc1163_5 gpc14 (
      {stage0_0[62], stage0_0[63], stage0_0[64]},
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59]},
      {stage0_2[14]},
      {stage0_3[24]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc1163_5 gpc15 (
      {stage0_0[65], stage0_0[66], stage0_0[67]},
      {stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65]},
      {stage0_2[15]},
      {stage0_3[25]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc1163_5 gpc16 (
      {stage0_0[68], stage0_0[69], stage0_0[70]},
      {stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71]},
      {stage0_2[16]},
      {stage0_3[26]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc207_4 gpc17 (
      {stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74], stage0_0[75], stage0_0[76], stage0_0[77]},
      {stage0_2[17], stage0_2[18]},
      {stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc606_5 gpc18 (
      {stage0_0[78], stage0_0[79], stage0_0[80], stage0_0[81], stage0_0[82], stage0_0[83]},
      {stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24]},
      {stage1_4[17],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc606_5 gpc19 (
      {stage0_0[84], stage0_0[85], stage0_0[86], stage0_0[87], stage0_0[88], stage0_0[89]},
      {stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30]},
      {stage1_4[18],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc606_5 gpc20 (
      {stage0_0[90], stage0_0[91], stage0_0[92], stage0_0[93], stage0_0[94], stage0_0[95]},
      {stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36]},
      {stage1_4[19],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc606_5 gpc21 (
      {stage0_0[96], stage0_0[97], stage0_0[98], stage0_0[99], stage0_0[100], stage0_0[101]},
      {stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42]},
      {stage1_4[20],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc606_5 gpc22 (
      {stage0_0[102], stage0_0[103], stage0_0[104], stage0_0[105], stage0_0[106], stage0_0[107]},
      {stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48]},
      {stage1_4[21],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc606_5 gpc23 (
      {stage0_0[108], stage0_0[109], stage0_0[110], stage0_0[111], stage0_0[112], stage0_0[113]},
      {stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54]},
      {stage1_4[22],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc606_5 gpc24 (
      {stage0_0[114], stage0_0[115], stage0_0[116], stage0_0[117], stage0_0[118], stage0_0[119]},
      {stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60]},
      {stage1_4[23],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc606_5 gpc25 (
      {stage0_0[120], stage0_0[121], stage0_0[122], stage0_0[123], stage0_0[124], stage0_0[125]},
      {stage0_2[61], stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66]},
      {stage1_4[24],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc606_5 gpc26 (
      {stage0_0[126], stage0_0[127], stage0_0[128], stage0_0[129], stage0_0[130], stage0_0[131]},
      {stage0_2[67], stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72]},
      {stage1_4[25],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc606_5 gpc27 (
      {stage0_0[132], stage0_0[133], stage0_0[134], stage0_0[135], stage0_0[136], stage0_0[137]},
      {stage0_2[73], stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78]},
      {stage1_4[26],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc606_5 gpc28 (
      {stage0_0[138], stage0_0[139], stage0_0[140], stage0_0[141], stage0_0[142], stage0_0[143]},
      {stage0_2[79], stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84]},
      {stage1_4[27],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc606_5 gpc29 (
      {stage0_0[144], stage0_0[145], stage0_0[146], stage0_0[147], stage0_0[148], stage0_0[149]},
      {stage0_2[85], stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90]},
      {stage1_4[28],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc606_5 gpc30 (
      {stage0_0[150], stage0_0[151], stage0_0[152], stage0_0[153], stage0_0[154], stage0_0[155]},
      {stage0_2[91], stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96]},
      {stage1_4[29],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc606_5 gpc31 (
      {stage0_0[156], stage0_0[157], stage0_0[158], stage0_0[159], stage0_0[160], stage0_0[161]},
      {stage0_2[97], stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102]},
      {stage1_4[30],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc606_5 gpc32 (
      {stage0_0[162], stage0_0[163], stage0_0[164], stage0_0[165], stage0_0[166], stage0_0[167]},
      {stage0_2[103], stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108]},
      {stage1_4[31],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc606_5 gpc33 (
      {stage0_0[168], stage0_0[169], stage0_0[170], stage0_0[171], stage0_0[172], stage0_0[173]},
      {stage0_2[109], stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114]},
      {stage1_4[32],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc606_5 gpc34 (
      {stage0_0[174], stage0_0[175], stage0_0[176], stage0_0[177], stage0_0[178], stage0_0[179]},
      {stage0_2[115], stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120]},
      {stage1_4[33],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc606_5 gpc35 (
      {stage0_0[180], stage0_0[181], stage0_0[182], stage0_0[183], stage0_0[184], stage0_0[185]},
      {stage0_2[121], stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126]},
      {stage1_4[34],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc606_5 gpc36 (
      {stage0_0[186], stage0_0[187], stage0_0[188], stage0_0[189], stage0_0[190], stage0_0[191]},
      {stage0_2[127], stage0_2[128], stage0_2[129], stage0_2[130], stage0_2[131], stage0_2[132]},
      {stage1_4[35],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc606_5 gpc37 (
      {stage0_0[192], stage0_0[193], stage0_0[194], stage0_0[195], stage0_0[196], stage0_0[197]},
      {stage0_2[133], stage0_2[134], stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138]},
      {stage1_4[36],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc606_5 gpc38 (
      {stage0_0[198], stage0_0[199], stage0_0[200], stage0_0[201], stage0_0[202], stage0_0[203]},
      {stage0_2[139], stage0_2[140], stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144]},
      {stage1_4[37],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc606_5 gpc39 (
      {stage0_0[204], stage0_0[205], stage0_0[206], stage0_0[207], stage0_0[208], stage0_0[209]},
      {stage0_2[145], stage0_2[146], stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150]},
      {stage1_4[38],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc606_5 gpc40 (
      {stage0_0[210], stage0_0[211], stage0_0[212], stage0_0[213], stage0_0[214], stage0_0[215]},
      {stage0_2[151], stage0_2[152], stage0_2[153], stage0_2[154], stage0_2[155], stage0_2[156]},
      {stage1_4[39],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc606_5 gpc41 (
      {stage0_0[216], stage0_0[217], stage0_0[218], stage0_0[219], stage0_0[220], stage0_0[221]},
      {stage0_2[157], stage0_2[158], stage0_2[159], stage0_2[160], stage0_2[161], stage0_2[162]},
      {stage1_4[40],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc606_5 gpc42 (
      {stage0_0[222], stage0_0[223], stage0_0[224], stage0_0[225], stage0_0[226], stage0_0[227]},
      {stage0_2[163], stage0_2[164], stage0_2[165], stage0_2[166], stage0_2[167], stage0_2[168]},
      {stage1_4[41],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc606_5 gpc43 (
      {stage0_0[228], stage0_0[229], stage0_0[230], stage0_0[231], stage0_0[232], stage0_0[233]},
      {stage0_2[169], stage0_2[170], stage0_2[171], stage0_2[172], stage0_2[173], stage0_2[174]},
      {stage1_4[42],stage1_3[43],stage1_2[43],stage1_1[43],stage1_0[43]}
   );
   gpc606_5 gpc44 (
      {stage0_0[234], stage0_0[235], stage0_0[236], stage0_0[237], stage0_0[238], stage0_0[239]},
      {stage0_2[175], stage0_2[176], stage0_2[177], stage0_2[178], stage0_2[179], stage0_2[180]},
      {stage1_4[43],stage1_3[44],stage1_2[44],stage1_1[44],stage1_0[44]}
   );
   gpc606_5 gpc45 (
      {stage0_0[240], stage0_0[241], stage0_0[242], stage0_0[243], stage0_0[244], stage0_0[245]},
      {stage0_2[181], stage0_2[182], stage0_2[183], stage0_2[184], stage0_2[185], stage0_2[186]},
      {stage1_4[44],stage1_3[45],stage1_2[45],stage1_1[45],stage1_0[45]}
   );
   gpc606_5 gpc46 (
      {stage0_0[246], stage0_0[247], stage0_0[248], stage0_0[249], stage0_0[250], stage0_0[251]},
      {stage0_2[187], stage0_2[188], stage0_2[189], stage0_2[190], stage0_2[191], stage0_2[192]},
      {stage1_4[45],stage1_3[46],stage1_2[46],stage1_1[46],stage1_0[46]}
   );
   gpc606_5 gpc47 (
      {stage0_0[252], stage0_0[253], stage0_0[254], stage0_0[255], stage0_0[256], stage0_0[257]},
      {stage0_2[193], stage0_2[194], stage0_2[195], stage0_2[196], stage0_2[197], stage0_2[198]},
      {stage1_4[46],stage1_3[47],stage1_2[47],stage1_1[47],stage1_0[47]}
   );
   gpc606_5 gpc48 (
      {stage0_0[258], stage0_0[259], stage0_0[260], stage0_0[261], stage0_0[262], stage0_0[263]},
      {stage0_2[199], stage0_2[200], stage0_2[201], stage0_2[202], stage0_2[203], stage0_2[204]},
      {stage1_4[47],stage1_3[48],stage1_2[48],stage1_1[48],stage1_0[48]}
   );
   gpc606_5 gpc49 (
      {stage0_0[264], stage0_0[265], stage0_0[266], stage0_0[267], stage0_0[268], stage0_0[269]},
      {stage0_2[205], stage0_2[206], stage0_2[207], stage0_2[208], stage0_2[209], stage0_2[210]},
      {stage1_4[48],stage1_3[49],stage1_2[49],stage1_1[49],stage1_0[49]}
   );
   gpc606_5 gpc50 (
      {stage0_0[270], stage0_0[271], stage0_0[272], stage0_0[273], stage0_0[274], stage0_0[275]},
      {stage0_2[211], stage0_2[212], stage0_2[213], stage0_2[214], stage0_2[215], stage0_2[216]},
      {stage1_4[49],stage1_3[50],stage1_2[50],stage1_1[50],stage1_0[50]}
   );
   gpc606_5 gpc51 (
      {stage0_0[276], stage0_0[277], stage0_0[278], stage0_0[279], stage0_0[280], stage0_0[281]},
      {stage0_2[217], stage0_2[218], stage0_2[219], stage0_2[220], stage0_2[221], stage0_2[222]},
      {stage1_4[50],stage1_3[51],stage1_2[51],stage1_1[51],stage1_0[51]}
   );
   gpc606_5 gpc52 (
      {stage0_0[282], stage0_0[283], stage0_0[284], stage0_0[285], stage0_0[286], stage0_0[287]},
      {stage0_2[223], stage0_2[224], stage0_2[225], stage0_2[226], stage0_2[227], stage0_2[228]},
      {stage1_4[51],stage1_3[52],stage1_2[52],stage1_1[52],stage1_0[52]}
   );
   gpc606_5 gpc53 (
      {stage0_0[288], stage0_0[289], stage0_0[290], stage0_0[291], stage0_0[292], stage0_0[293]},
      {stage0_2[229], stage0_2[230], stage0_2[231], stage0_2[232], stage0_2[233], stage0_2[234]},
      {stage1_4[52],stage1_3[53],stage1_2[53],stage1_1[53],stage1_0[53]}
   );
   gpc606_5 gpc54 (
      {stage0_0[294], stage0_0[295], stage0_0[296], stage0_0[297], stage0_0[298], stage0_0[299]},
      {stage0_2[235], stage0_2[236], stage0_2[237], stage0_2[238], stage0_2[239], stage0_2[240]},
      {stage1_4[53],stage1_3[54],stage1_2[54],stage1_1[54],stage1_0[54]}
   );
   gpc606_5 gpc55 (
      {stage0_0[300], stage0_0[301], stage0_0[302], stage0_0[303], stage0_0[304], stage0_0[305]},
      {stage0_2[241], stage0_2[242], stage0_2[243], stage0_2[244], stage0_2[245], stage0_2[246]},
      {stage1_4[54],stage1_3[55],stage1_2[55],stage1_1[55],stage1_0[55]}
   );
   gpc606_5 gpc56 (
      {stage0_0[306], stage0_0[307], stage0_0[308], stage0_0[309], stage0_0[310], stage0_0[311]},
      {stage0_2[247], stage0_2[248], stage0_2[249], stage0_2[250], stage0_2[251], stage0_2[252]},
      {stage1_4[55],stage1_3[56],stage1_2[56],stage1_1[56],stage1_0[56]}
   );
   gpc606_5 gpc57 (
      {stage0_0[312], stage0_0[313], stage0_0[314], stage0_0[315], stage0_0[316], stage0_0[317]},
      {stage0_2[253], stage0_2[254], stage0_2[255], stage0_2[256], stage0_2[257], stage0_2[258]},
      {stage1_4[56],stage1_3[57],stage1_2[57],stage1_1[57],stage1_0[57]}
   );
   gpc606_5 gpc58 (
      {stage0_0[318], stage0_0[319], stage0_0[320], stage0_0[321], stage0_0[322], stage0_0[323]},
      {stage0_2[259], stage0_2[260], stage0_2[261], stage0_2[262], stage0_2[263], stage0_2[264]},
      {stage1_4[57],stage1_3[58],stage1_2[58],stage1_1[58],stage1_0[58]}
   );
   gpc606_5 gpc59 (
      {stage0_0[324], stage0_0[325], stage0_0[326], stage0_0[327], stage0_0[328], stage0_0[329]},
      {stage0_2[265], stage0_2[266], stage0_2[267], stage0_2[268], stage0_2[269], stage0_2[270]},
      {stage1_4[58],stage1_3[59],stage1_2[59],stage1_1[59],stage1_0[59]}
   );
   gpc606_5 gpc60 (
      {stage0_0[330], stage0_0[331], stage0_0[332], stage0_0[333], stage0_0[334], stage0_0[335]},
      {stage0_2[271], stage0_2[272], stage0_2[273], stage0_2[274], stage0_2[275], stage0_2[276]},
      {stage1_4[59],stage1_3[60],stage1_2[60],stage1_1[60],stage1_0[60]}
   );
   gpc606_5 gpc61 (
      {stage0_0[336], stage0_0[337], stage0_0[338], stage0_0[339], stage0_0[340], stage0_0[341]},
      {stage0_2[277], stage0_2[278], stage0_2[279], stage0_2[280], stage0_2[281], stage0_2[282]},
      {stage1_4[60],stage1_3[61],stage1_2[61],stage1_1[61],stage1_0[61]}
   );
   gpc606_5 gpc62 (
      {stage0_0[342], stage0_0[343], stage0_0[344], stage0_0[345], stage0_0[346], stage0_0[347]},
      {stage0_2[283], stage0_2[284], stage0_2[285], stage0_2[286], stage0_2[287], stage0_2[288]},
      {stage1_4[61],stage1_3[62],stage1_2[62],stage1_1[62],stage1_0[62]}
   );
   gpc606_5 gpc63 (
      {stage0_0[348], stage0_0[349], stage0_0[350], stage0_0[351], stage0_0[352], stage0_0[353]},
      {stage0_2[289], stage0_2[290], stage0_2[291], stage0_2[292], stage0_2[293], stage0_2[294]},
      {stage1_4[62],stage1_3[63],stage1_2[63],stage1_1[63],stage1_0[63]}
   );
   gpc606_5 gpc64 (
      {stage0_0[354], stage0_0[355], stage0_0[356], stage0_0[357], stage0_0[358], stage0_0[359]},
      {stage0_2[295], stage0_2[296], stage0_2[297], stage0_2[298], stage0_2[299], stage0_2[300]},
      {stage1_4[63],stage1_3[64],stage1_2[64],stage1_1[64],stage1_0[64]}
   );
   gpc606_5 gpc65 (
      {stage0_0[360], stage0_0[361], stage0_0[362], stage0_0[363], stage0_0[364], stage0_0[365]},
      {stage0_2[301], stage0_2[302], stage0_2[303], stage0_2[304], stage0_2[305], stage0_2[306]},
      {stage1_4[64],stage1_3[65],stage1_2[65],stage1_1[65],stage1_0[65]}
   );
   gpc606_5 gpc66 (
      {stage0_0[366], stage0_0[367], stage0_0[368], stage0_0[369], stage0_0[370], stage0_0[371]},
      {stage0_2[307], stage0_2[308], stage0_2[309], stage0_2[310], stage0_2[311], stage0_2[312]},
      {stage1_4[65],stage1_3[66],stage1_2[66],stage1_1[66],stage1_0[66]}
   );
   gpc606_5 gpc67 (
      {stage0_0[372], stage0_0[373], stage0_0[374], stage0_0[375], stage0_0[376], stage0_0[377]},
      {stage0_2[313], stage0_2[314], stage0_2[315], stage0_2[316], stage0_2[317], stage0_2[318]},
      {stage1_4[66],stage1_3[67],stage1_2[67],stage1_1[67],stage1_0[67]}
   );
   gpc606_5 gpc68 (
      {stage0_0[378], stage0_0[379], stage0_0[380], stage0_0[381], stage0_0[382], stage0_0[383]},
      {stage0_2[319], stage0_2[320], stage0_2[321], stage0_2[322], stage0_2[323], stage0_2[324]},
      {stage1_4[67],stage1_3[68],stage1_2[68],stage1_1[68],stage1_0[68]}
   );
   gpc606_5 gpc69 (
      {stage0_0[384], stage0_0[385], stage0_0[386], stage0_0[387], stage0_0[388], stage0_0[389]},
      {stage0_2[325], stage0_2[326], stage0_2[327], stage0_2[328], stage0_2[329], stage0_2[330]},
      {stage1_4[68],stage1_3[69],stage1_2[69],stage1_1[69],stage1_0[69]}
   );
   gpc606_5 gpc70 (
      {stage0_0[390], stage0_0[391], stage0_0[392], stage0_0[393], stage0_0[394], stage0_0[395]},
      {stage0_2[331], stage0_2[332], stage0_2[333], stage0_2[334], stage0_2[335], stage0_2[336]},
      {stage1_4[69],stage1_3[70],stage1_2[70],stage1_1[70],stage1_0[70]}
   );
   gpc606_5 gpc71 (
      {stage0_0[396], stage0_0[397], stage0_0[398], stage0_0[399], stage0_0[400], stage0_0[401]},
      {stage0_2[337], stage0_2[338], stage0_2[339], stage0_2[340], stage0_2[341], stage0_2[342]},
      {stage1_4[70],stage1_3[71],stage1_2[71],stage1_1[71],stage1_0[71]}
   );
   gpc606_5 gpc72 (
      {stage0_0[402], stage0_0[403], stage0_0[404], stage0_0[405], stage0_0[406], stage0_0[407]},
      {stage0_2[343], stage0_2[344], stage0_2[345], stage0_2[346], stage0_2[347], stage0_2[348]},
      {stage1_4[71],stage1_3[72],stage1_2[72],stage1_1[72],stage1_0[72]}
   );
   gpc606_5 gpc73 (
      {stage0_0[408], stage0_0[409], stage0_0[410], stage0_0[411], stage0_0[412], stage0_0[413]},
      {stage0_2[349], stage0_2[350], stage0_2[351], stage0_2[352], stage0_2[353], stage0_2[354]},
      {stage1_4[72],stage1_3[73],stage1_2[73],stage1_1[73],stage1_0[73]}
   );
   gpc606_5 gpc74 (
      {stage0_0[414], stage0_0[415], stage0_0[416], stage0_0[417], stage0_0[418], stage0_0[419]},
      {stage0_2[355], stage0_2[356], stage0_2[357], stage0_2[358], stage0_2[359], stage0_2[360]},
      {stage1_4[73],stage1_3[74],stage1_2[74],stage1_1[74],stage1_0[74]}
   );
   gpc606_5 gpc75 (
      {stage0_0[420], stage0_0[421], stage0_0[422], stage0_0[423], stage0_0[424], stage0_0[425]},
      {stage0_2[361], stage0_2[362], stage0_2[363], stage0_2[364], stage0_2[365], stage0_2[366]},
      {stage1_4[74],stage1_3[75],stage1_2[75],stage1_1[75],stage1_0[75]}
   );
   gpc606_5 gpc76 (
      {stage0_0[426], stage0_0[427], stage0_0[428], stage0_0[429], stage0_0[430], stage0_0[431]},
      {stage0_2[367], stage0_2[368], stage0_2[369], stage0_2[370], stage0_2[371], stage0_2[372]},
      {stage1_4[75],stage1_3[76],stage1_2[76],stage1_1[76],stage1_0[76]}
   );
   gpc606_5 gpc77 (
      {stage0_0[432], stage0_0[433], stage0_0[434], stage0_0[435], stage0_0[436], stage0_0[437]},
      {stage0_2[373], stage0_2[374], stage0_2[375], stage0_2[376], stage0_2[377], stage0_2[378]},
      {stage1_4[76],stage1_3[77],stage1_2[77],stage1_1[77],stage1_0[77]}
   );
   gpc606_5 gpc78 (
      {stage0_0[438], stage0_0[439], stage0_0[440], stage0_0[441], stage0_0[442], stage0_0[443]},
      {stage0_2[379], stage0_2[380], stage0_2[381], stage0_2[382], stage0_2[383], stage0_2[384]},
      {stage1_4[77],stage1_3[78],stage1_2[78],stage1_1[78],stage1_0[78]}
   );
   gpc606_5 gpc79 (
      {stage0_0[444], stage0_0[445], stage0_0[446], stage0_0[447], stage0_0[448], stage0_0[449]},
      {stage0_2[385], stage0_2[386], stage0_2[387], stage0_2[388], stage0_2[389], stage0_2[390]},
      {stage1_4[78],stage1_3[79],stage1_2[79],stage1_1[79],stage1_0[79]}
   );
   gpc606_5 gpc80 (
      {stage0_0[450], stage0_0[451], stage0_0[452], stage0_0[453], stage0_0[454], stage0_0[455]},
      {stage0_2[391], stage0_2[392], stage0_2[393], stage0_2[394], stage0_2[395], stage0_2[396]},
      {stage1_4[79],stage1_3[80],stage1_2[80],stage1_1[80],stage1_0[80]}
   );
   gpc606_5 gpc81 (
      {stage0_0[456], stage0_0[457], stage0_0[458], stage0_0[459], stage0_0[460], stage0_0[461]},
      {stage0_2[397], stage0_2[398], stage0_2[399], stage0_2[400], stage0_2[401], stage0_2[402]},
      {stage1_4[80],stage1_3[81],stage1_2[81],stage1_1[81],stage1_0[81]}
   );
   gpc606_5 gpc82 (
      {stage0_0[462], stage0_0[463], stage0_0[464], stage0_0[465], stage0_0[466], stage0_0[467]},
      {stage0_2[403], stage0_2[404], stage0_2[405], stage0_2[406], stage0_2[407], stage0_2[408]},
      {stage1_4[81],stage1_3[82],stage1_2[82],stage1_1[82],stage1_0[82]}
   );
   gpc606_5 gpc83 (
      {stage0_0[468], stage0_0[469], stage0_0[470], stage0_0[471], stage0_0[472], stage0_0[473]},
      {stage0_2[409], stage0_2[410], stage0_2[411], stage0_2[412], stage0_2[413], stage0_2[414]},
      {stage1_4[82],stage1_3[83],stage1_2[83],stage1_1[83],stage1_0[83]}
   );
   gpc606_5 gpc84 (
      {stage0_0[474], stage0_0[475], stage0_0[476], stage0_0[477], stage0_0[478], stage0_0[479]},
      {stage0_2[415], stage0_2[416], stage0_2[417], stage0_2[418], stage0_2[419], stage0_2[420]},
      {stage1_4[83],stage1_3[84],stage1_2[84],stage1_1[84],stage1_0[84]}
   );
   gpc606_5 gpc85 (
      {stage0_0[480], stage0_0[481], stage0_0[482], stage0_0[483], stage0_0[484], stage0_0[485]},
      {stage0_2[421], stage0_2[422], stage0_2[423], stage0_2[424], stage0_2[425], stage0_2[426]},
      {stage1_4[84],stage1_3[85],stage1_2[85],stage1_1[85],stage1_0[85]}
   );
   gpc606_5 gpc86 (
      {stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77]},
      {stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32]},
      {stage1_5[0],stage1_4[85],stage1_3[86],stage1_2[86],stage1_1[86]}
   );
   gpc606_5 gpc87 (
      {stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83]},
      {stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38]},
      {stage1_5[1],stage1_4[86],stage1_3[87],stage1_2[87],stage1_1[87]}
   );
   gpc606_5 gpc88 (
      {stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89]},
      {stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44]},
      {stage1_5[2],stage1_4[87],stage1_3[88],stage1_2[88],stage1_1[88]}
   );
   gpc606_5 gpc89 (
      {stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95]},
      {stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50]},
      {stage1_5[3],stage1_4[88],stage1_3[89],stage1_2[89],stage1_1[89]}
   );
   gpc606_5 gpc90 (
      {stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101]},
      {stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56]},
      {stage1_5[4],stage1_4[89],stage1_3[90],stage1_2[90],stage1_1[90]}
   );
   gpc606_5 gpc91 (
      {stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107]},
      {stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62]},
      {stage1_5[5],stage1_4[90],stage1_3[91],stage1_2[91],stage1_1[91]}
   );
   gpc606_5 gpc92 (
      {stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113]},
      {stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68]},
      {stage1_5[6],stage1_4[91],stage1_3[92],stage1_2[92],stage1_1[92]}
   );
   gpc606_5 gpc93 (
      {stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119]},
      {stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74]},
      {stage1_5[7],stage1_4[92],stage1_3[93],stage1_2[93],stage1_1[93]}
   );
   gpc606_5 gpc94 (
      {stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125]},
      {stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80]},
      {stage1_5[8],stage1_4[93],stage1_3[94],stage1_2[94],stage1_1[94]}
   );
   gpc606_5 gpc95 (
      {stage0_1[126], stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131]},
      {stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86]},
      {stage1_5[9],stage1_4[94],stage1_3[95],stage1_2[95],stage1_1[95]}
   );
   gpc606_5 gpc96 (
      {stage0_1[132], stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137]},
      {stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92]},
      {stage1_5[10],stage1_4[95],stage1_3[96],stage1_2[96],stage1_1[96]}
   );
   gpc606_5 gpc97 (
      {stage0_1[138], stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143]},
      {stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98]},
      {stage1_5[11],stage1_4[96],stage1_3[97],stage1_2[97],stage1_1[97]}
   );
   gpc606_5 gpc98 (
      {stage0_1[144], stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149]},
      {stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104]},
      {stage1_5[12],stage1_4[97],stage1_3[98],stage1_2[98],stage1_1[98]}
   );
   gpc606_5 gpc99 (
      {stage0_1[150], stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155]},
      {stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110]},
      {stage1_5[13],stage1_4[98],stage1_3[99],stage1_2[99],stage1_1[99]}
   );
   gpc606_5 gpc100 (
      {stage0_1[156], stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161]},
      {stage0_3[111], stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116]},
      {stage1_5[14],stage1_4[99],stage1_3[100],stage1_2[100],stage1_1[100]}
   );
   gpc606_5 gpc101 (
      {stage0_1[162], stage0_1[163], stage0_1[164], stage0_1[165], stage0_1[166], stage0_1[167]},
      {stage0_3[117], stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121], stage0_3[122]},
      {stage1_5[15],stage1_4[100],stage1_3[101],stage1_2[101],stage1_1[101]}
   );
   gpc606_5 gpc102 (
      {stage0_1[168], stage0_1[169], stage0_1[170], stage0_1[171], stage0_1[172], stage0_1[173]},
      {stage0_3[123], stage0_3[124], stage0_3[125], stage0_3[126], stage0_3[127], stage0_3[128]},
      {stage1_5[16],stage1_4[101],stage1_3[102],stage1_2[102],stage1_1[102]}
   );
   gpc606_5 gpc103 (
      {stage0_1[174], stage0_1[175], stage0_1[176], stage0_1[177], stage0_1[178], stage0_1[179]},
      {stage0_3[129], stage0_3[130], stage0_3[131], stage0_3[132], stage0_3[133], stage0_3[134]},
      {stage1_5[17],stage1_4[102],stage1_3[103],stage1_2[103],stage1_1[103]}
   );
   gpc606_5 gpc104 (
      {stage0_1[180], stage0_1[181], stage0_1[182], stage0_1[183], stage0_1[184], stage0_1[185]},
      {stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138], stage0_3[139], stage0_3[140]},
      {stage1_5[18],stage1_4[103],stage1_3[104],stage1_2[104],stage1_1[104]}
   );
   gpc606_5 gpc105 (
      {stage0_1[186], stage0_1[187], stage0_1[188], stage0_1[189], stage0_1[190], stage0_1[191]},
      {stage0_3[141], stage0_3[142], stage0_3[143], stage0_3[144], stage0_3[145], stage0_3[146]},
      {stage1_5[19],stage1_4[104],stage1_3[105],stage1_2[105],stage1_1[105]}
   );
   gpc606_5 gpc106 (
      {stage0_1[192], stage0_1[193], stage0_1[194], stage0_1[195], stage0_1[196], stage0_1[197]},
      {stage0_3[147], stage0_3[148], stage0_3[149], stage0_3[150], stage0_3[151], stage0_3[152]},
      {stage1_5[20],stage1_4[105],stage1_3[106],stage1_2[106],stage1_1[106]}
   );
   gpc606_5 gpc107 (
      {stage0_1[198], stage0_1[199], stage0_1[200], stage0_1[201], stage0_1[202], stage0_1[203]},
      {stage0_3[153], stage0_3[154], stage0_3[155], stage0_3[156], stage0_3[157], stage0_3[158]},
      {stage1_5[21],stage1_4[106],stage1_3[107],stage1_2[107],stage1_1[107]}
   );
   gpc606_5 gpc108 (
      {stage0_1[204], stage0_1[205], stage0_1[206], stage0_1[207], stage0_1[208], stage0_1[209]},
      {stage0_3[159], stage0_3[160], stage0_3[161], stage0_3[162], stage0_3[163], stage0_3[164]},
      {stage1_5[22],stage1_4[107],stage1_3[108],stage1_2[108],stage1_1[108]}
   );
   gpc606_5 gpc109 (
      {stage0_1[210], stage0_1[211], stage0_1[212], stage0_1[213], stage0_1[214], stage0_1[215]},
      {stage0_3[165], stage0_3[166], stage0_3[167], stage0_3[168], stage0_3[169], stage0_3[170]},
      {stage1_5[23],stage1_4[108],stage1_3[109],stage1_2[109],stage1_1[109]}
   );
   gpc606_5 gpc110 (
      {stage0_1[216], stage0_1[217], stage0_1[218], stage0_1[219], stage0_1[220], stage0_1[221]},
      {stage0_3[171], stage0_3[172], stage0_3[173], stage0_3[174], stage0_3[175], stage0_3[176]},
      {stage1_5[24],stage1_4[109],stage1_3[110],stage1_2[110],stage1_1[110]}
   );
   gpc606_5 gpc111 (
      {stage0_1[222], stage0_1[223], stage0_1[224], stage0_1[225], stage0_1[226], stage0_1[227]},
      {stage0_3[177], stage0_3[178], stage0_3[179], stage0_3[180], stage0_3[181], stage0_3[182]},
      {stage1_5[25],stage1_4[110],stage1_3[111],stage1_2[111],stage1_1[111]}
   );
   gpc606_5 gpc112 (
      {stage0_1[228], stage0_1[229], stage0_1[230], stage0_1[231], stage0_1[232], stage0_1[233]},
      {stage0_3[183], stage0_3[184], stage0_3[185], stage0_3[186], stage0_3[187], stage0_3[188]},
      {stage1_5[26],stage1_4[111],stage1_3[112],stage1_2[112],stage1_1[112]}
   );
   gpc606_5 gpc113 (
      {stage0_1[234], stage0_1[235], stage0_1[236], stage0_1[237], stage0_1[238], stage0_1[239]},
      {stage0_3[189], stage0_3[190], stage0_3[191], stage0_3[192], stage0_3[193], stage0_3[194]},
      {stage1_5[27],stage1_4[112],stage1_3[113],stage1_2[113],stage1_1[113]}
   );
   gpc606_5 gpc114 (
      {stage0_1[240], stage0_1[241], stage0_1[242], stage0_1[243], stage0_1[244], stage0_1[245]},
      {stage0_3[195], stage0_3[196], stage0_3[197], stage0_3[198], stage0_3[199], stage0_3[200]},
      {stage1_5[28],stage1_4[113],stage1_3[114],stage1_2[114],stage1_1[114]}
   );
   gpc606_5 gpc115 (
      {stage0_1[246], stage0_1[247], stage0_1[248], stage0_1[249], stage0_1[250], stage0_1[251]},
      {stage0_3[201], stage0_3[202], stage0_3[203], stage0_3[204], stage0_3[205], stage0_3[206]},
      {stage1_5[29],stage1_4[114],stage1_3[115],stage1_2[115],stage1_1[115]}
   );
   gpc606_5 gpc116 (
      {stage0_1[252], stage0_1[253], stage0_1[254], stage0_1[255], stage0_1[256], stage0_1[257]},
      {stage0_3[207], stage0_3[208], stage0_3[209], stage0_3[210], stage0_3[211], stage0_3[212]},
      {stage1_5[30],stage1_4[115],stage1_3[116],stage1_2[116],stage1_1[116]}
   );
   gpc606_5 gpc117 (
      {stage0_1[258], stage0_1[259], stage0_1[260], stage0_1[261], stage0_1[262], stage0_1[263]},
      {stage0_3[213], stage0_3[214], stage0_3[215], stage0_3[216], stage0_3[217], stage0_3[218]},
      {stage1_5[31],stage1_4[116],stage1_3[117],stage1_2[117],stage1_1[117]}
   );
   gpc606_5 gpc118 (
      {stage0_1[264], stage0_1[265], stage0_1[266], stage0_1[267], stage0_1[268], stage0_1[269]},
      {stage0_3[219], stage0_3[220], stage0_3[221], stage0_3[222], stage0_3[223], stage0_3[224]},
      {stage1_5[32],stage1_4[117],stage1_3[118],stage1_2[118],stage1_1[118]}
   );
   gpc606_5 gpc119 (
      {stage0_1[270], stage0_1[271], stage0_1[272], stage0_1[273], stage0_1[274], stage0_1[275]},
      {stage0_3[225], stage0_3[226], stage0_3[227], stage0_3[228], stage0_3[229], stage0_3[230]},
      {stage1_5[33],stage1_4[118],stage1_3[119],stage1_2[119],stage1_1[119]}
   );
   gpc606_5 gpc120 (
      {stage0_1[276], stage0_1[277], stage0_1[278], stage0_1[279], stage0_1[280], stage0_1[281]},
      {stage0_3[231], stage0_3[232], stage0_3[233], stage0_3[234], stage0_3[235], stage0_3[236]},
      {stage1_5[34],stage1_4[119],stage1_3[120],stage1_2[120],stage1_1[120]}
   );
   gpc606_5 gpc121 (
      {stage0_1[282], stage0_1[283], stage0_1[284], stage0_1[285], stage0_1[286], stage0_1[287]},
      {stage0_3[237], stage0_3[238], stage0_3[239], stage0_3[240], stage0_3[241], stage0_3[242]},
      {stage1_5[35],stage1_4[120],stage1_3[121],stage1_2[121],stage1_1[121]}
   );
   gpc606_5 gpc122 (
      {stage0_1[288], stage0_1[289], stage0_1[290], stage0_1[291], stage0_1[292], stage0_1[293]},
      {stage0_3[243], stage0_3[244], stage0_3[245], stage0_3[246], stage0_3[247], stage0_3[248]},
      {stage1_5[36],stage1_4[121],stage1_3[122],stage1_2[122],stage1_1[122]}
   );
   gpc606_5 gpc123 (
      {stage0_1[294], stage0_1[295], stage0_1[296], stage0_1[297], stage0_1[298], stage0_1[299]},
      {stage0_3[249], stage0_3[250], stage0_3[251], stage0_3[252], stage0_3[253], stage0_3[254]},
      {stage1_5[37],stage1_4[122],stage1_3[123],stage1_2[123],stage1_1[123]}
   );
   gpc606_5 gpc124 (
      {stage0_1[300], stage0_1[301], stage0_1[302], stage0_1[303], stage0_1[304], stage0_1[305]},
      {stage0_3[255], stage0_3[256], stage0_3[257], stage0_3[258], stage0_3[259], stage0_3[260]},
      {stage1_5[38],stage1_4[123],stage1_3[124],stage1_2[124],stage1_1[124]}
   );
   gpc606_5 gpc125 (
      {stage0_1[306], stage0_1[307], stage0_1[308], stage0_1[309], stage0_1[310], stage0_1[311]},
      {stage0_3[261], stage0_3[262], stage0_3[263], stage0_3[264], stage0_3[265], stage0_3[266]},
      {stage1_5[39],stage1_4[124],stage1_3[125],stage1_2[125],stage1_1[125]}
   );
   gpc606_5 gpc126 (
      {stage0_1[312], stage0_1[313], stage0_1[314], stage0_1[315], stage0_1[316], stage0_1[317]},
      {stage0_3[267], stage0_3[268], stage0_3[269], stage0_3[270], stage0_3[271], stage0_3[272]},
      {stage1_5[40],stage1_4[125],stage1_3[126],stage1_2[126],stage1_1[126]}
   );
   gpc606_5 gpc127 (
      {stage0_1[318], stage0_1[319], stage0_1[320], stage0_1[321], stage0_1[322], stage0_1[323]},
      {stage0_3[273], stage0_3[274], stage0_3[275], stage0_3[276], stage0_3[277], stage0_3[278]},
      {stage1_5[41],stage1_4[126],stage1_3[127],stage1_2[127],stage1_1[127]}
   );
   gpc606_5 gpc128 (
      {stage0_1[324], stage0_1[325], stage0_1[326], stage0_1[327], stage0_1[328], stage0_1[329]},
      {stage0_3[279], stage0_3[280], stage0_3[281], stage0_3[282], stage0_3[283], stage0_3[284]},
      {stage1_5[42],stage1_4[127],stage1_3[128],stage1_2[128],stage1_1[128]}
   );
   gpc606_5 gpc129 (
      {stage0_1[330], stage0_1[331], stage0_1[332], stage0_1[333], stage0_1[334], stage0_1[335]},
      {stage0_3[285], stage0_3[286], stage0_3[287], stage0_3[288], stage0_3[289], stage0_3[290]},
      {stage1_5[43],stage1_4[128],stage1_3[129],stage1_2[129],stage1_1[129]}
   );
   gpc606_5 gpc130 (
      {stage0_1[336], stage0_1[337], stage0_1[338], stage0_1[339], stage0_1[340], stage0_1[341]},
      {stage0_3[291], stage0_3[292], stage0_3[293], stage0_3[294], stage0_3[295], stage0_3[296]},
      {stage1_5[44],stage1_4[129],stage1_3[130],stage1_2[130],stage1_1[130]}
   );
   gpc606_5 gpc131 (
      {stage0_1[342], stage0_1[343], stage0_1[344], stage0_1[345], stage0_1[346], stage0_1[347]},
      {stage0_3[297], stage0_3[298], stage0_3[299], stage0_3[300], stage0_3[301], stage0_3[302]},
      {stage1_5[45],stage1_4[130],stage1_3[131],stage1_2[131],stage1_1[131]}
   );
   gpc606_5 gpc132 (
      {stage0_1[348], stage0_1[349], stage0_1[350], stage0_1[351], stage0_1[352], stage0_1[353]},
      {stage0_3[303], stage0_3[304], stage0_3[305], stage0_3[306], stage0_3[307], stage0_3[308]},
      {stage1_5[46],stage1_4[131],stage1_3[132],stage1_2[132],stage1_1[132]}
   );
   gpc606_5 gpc133 (
      {stage0_1[354], stage0_1[355], stage0_1[356], stage0_1[357], stage0_1[358], stage0_1[359]},
      {stage0_3[309], stage0_3[310], stage0_3[311], stage0_3[312], stage0_3[313], stage0_3[314]},
      {stage1_5[47],stage1_4[132],stage1_3[133],stage1_2[133],stage1_1[133]}
   );
   gpc606_5 gpc134 (
      {stage0_1[360], stage0_1[361], stage0_1[362], stage0_1[363], stage0_1[364], stage0_1[365]},
      {stage0_3[315], stage0_3[316], stage0_3[317], stage0_3[318], stage0_3[319], stage0_3[320]},
      {stage1_5[48],stage1_4[133],stage1_3[134],stage1_2[134],stage1_1[134]}
   );
   gpc606_5 gpc135 (
      {stage0_1[366], stage0_1[367], stage0_1[368], stage0_1[369], stage0_1[370], stage0_1[371]},
      {stage0_3[321], stage0_3[322], stage0_3[323], stage0_3[324], stage0_3[325], stage0_3[326]},
      {stage1_5[49],stage1_4[134],stage1_3[135],stage1_2[135],stage1_1[135]}
   );
   gpc606_5 gpc136 (
      {stage0_1[372], stage0_1[373], stage0_1[374], stage0_1[375], stage0_1[376], stage0_1[377]},
      {stage0_3[327], stage0_3[328], stage0_3[329], stage0_3[330], stage0_3[331], stage0_3[332]},
      {stage1_5[50],stage1_4[135],stage1_3[136],stage1_2[136],stage1_1[136]}
   );
   gpc606_5 gpc137 (
      {stage0_1[378], stage0_1[379], stage0_1[380], stage0_1[381], stage0_1[382], stage0_1[383]},
      {stage0_3[333], stage0_3[334], stage0_3[335], stage0_3[336], stage0_3[337], stage0_3[338]},
      {stage1_5[51],stage1_4[136],stage1_3[137],stage1_2[137],stage1_1[137]}
   );
   gpc606_5 gpc138 (
      {stage0_1[384], stage0_1[385], stage0_1[386], stage0_1[387], stage0_1[388], stage0_1[389]},
      {stage0_3[339], stage0_3[340], stage0_3[341], stage0_3[342], stage0_3[343], stage0_3[344]},
      {stage1_5[52],stage1_4[137],stage1_3[138],stage1_2[138],stage1_1[138]}
   );
   gpc606_5 gpc139 (
      {stage0_1[390], stage0_1[391], stage0_1[392], stage0_1[393], stage0_1[394], stage0_1[395]},
      {stage0_3[345], stage0_3[346], stage0_3[347], stage0_3[348], stage0_3[349], stage0_3[350]},
      {stage1_5[53],stage1_4[138],stage1_3[139],stage1_2[139],stage1_1[139]}
   );
   gpc606_5 gpc140 (
      {stage0_1[396], stage0_1[397], stage0_1[398], stage0_1[399], stage0_1[400], stage0_1[401]},
      {stage0_3[351], stage0_3[352], stage0_3[353], stage0_3[354], stage0_3[355], stage0_3[356]},
      {stage1_5[54],stage1_4[139],stage1_3[140],stage1_2[140],stage1_1[140]}
   );
   gpc606_5 gpc141 (
      {stage0_1[402], stage0_1[403], stage0_1[404], stage0_1[405], stage0_1[406], stage0_1[407]},
      {stage0_3[357], stage0_3[358], stage0_3[359], stage0_3[360], stage0_3[361], stage0_3[362]},
      {stage1_5[55],stage1_4[140],stage1_3[141],stage1_2[141],stage1_1[141]}
   );
   gpc606_5 gpc142 (
      {stage0_1[408], stage0_1[409], stage0_1[410], stage0_1[411], stage0_1[412], stage0_1[413]},
      {stage0_3[363], stage0_3[364], stage0_3[365], stage0_3[366], stage0_3[367], stage0_3[368]},
      {stage1_5[56],stage1_4[141],stage1_3[142],stage1_2[142],stage1_1[142]}
   );
   gpc606_5 gpc143 (
      {stage0_1[414], stage0_1[415], stage0_1[416], stage0_1[417], stage0_1[418], stage0_1[419]},
      {stage0_3[369], stage0_3[370], stage0_3[371], stage0_3[372], stage0_3[373], stage0_3[374]},
      {stage1_5[57],stage1_4[142],stage1_3[143],stage1_2[143],stage1_1[143]}
   );
   gpc606_5 gpc144 (
      {stage0_1[420], stage0_1[421], stage0_1[422], stage0_1[423], stage0_1[424], stage0_1[425]},
      {stage0_3[375], stage0_3[376], stage0_3[377], stage0_3[378], stage0_3[379], stage0_3[380]},
      {stage1_5[58],stage1_4[143],stage1_3[144],stage1_2[144],stage1_1[144]}
   );
   gpc606_5 gpc145 (
      {stage0_1[426], stage0_1[427], stage0_1[428], stage0_1[429], stage0_1[430], stage0_1[431]},
      {stage0_3[381], stage0_3[382], stage0_3[383], stage0_3[384], stage0_3[385], stage0_3[386]},
      {stage1_5[59],stage1_4[144],stage1_3[145],stage1_2[145],stage1_1[145]}
   );
   gpc606_5 gpc146 (
      {stage0_1[432], stage0_1[433], stage0_1[434], stage0_1[435], stage0_1[436], stage0_1[437]},
      {stage0_3[387], stage0_3[388], stage0_3[389], stage0_3[390], stage0_3[391], stage0_3[392]},
      {stage1_5[60],stage1_4[145],stage1_3[146],stage1_2[146],stage1_1[146]}
   );
   gpc606_5 gpc147 (
      {stage0_1[438], stage0_1[439], stage0_1[440], stage0_1[441], stage0_1[442], stage0_1[443]},
      {stage0_3[393], stage0_3[394], stage0_3[395], stage0_3[396], stage0_3[397], stage0_3[398]},
      {stage1_5[61],stage1_4[146],stage1_3[147],stage1_2[147],stage1_1[147]}
   );
   gpc606_5 gpc148 (
      {stage0_1[444], stage0_1[445], stage0_1[446], stage0_1[447], stage0_1[448], stage0_1[449]},
      {stage0_3[399], stage0_3[400], stage0_3[401], stage0_3[402], stage0_3[403], stage0_3[404]},
      {stage1_5[62],stage1_4[147],stage1_3[148],stage1_2[148],stage1_1[148]}
   );
   gpc606_5 gpc149 (
      {stage0_1[450], stage0_1[451], stage0_1[452], stage0_1[453], stage0_1[454], stage0_1[455]},
      {stage0_3[405], stage0_3[406], stage0_3[407], stage0_3[408], stage0_3[409], stage0_3[410]},
      {stage1_5[63],stage1_4[148],stage1_3[149],stage1_2[149],stage1_1[149]}
   );
   gpc606_5 gpc150 (
      {stage0_1[456], stage0_1[457], stage0_1[458], stage0_1[459], stage0_1[460], stage0_1[461]},
      {stage0_3[411], stage0_3[412], stage0_3[413], stage0_3[414], stage0_3[415], stage0_3[416]},
      {stage1_5[64],stage1_4[149],stage1_3[150],stage1_2[150],stage1_1[150]}
   );
   gpc606_5 gpc151 (
      {stage0_1[462], stage0_1[463], stage0_1[464], stage0_1[465], stage0_1[466], stage0_1[467]},
      {stage0_3[417], stage0_3[418], stage0_3[419], stage0_3[420], stage0_3[421], stage0_3[422]},
      {stage1_5[65],stage1_4[150],stage1_3[151],stage1_2[151],stage1_1[151]}
   );
   gpc606_5 gpc152 (
      {stage0_1[468], stage0_1[469], stage0_1[470], stage0_1[471], stage0_1[472], stage0_1[473]},
      {stage0_3[423], stage0_3[424], stage0_3[425], stage0_3[426], stage0_3[427], stage0_3[428]},
      {stage1_5[66],stage1_4[151],stage1_3[152],stage1_2[152],stage1_1[152]}
   );
   gpc606_5 gpc153 (
      {stage0_1[474], stage0_1[475], stage0_1[476], stage0_1[477], stage0_1[478], stage0_1[479]},
      {stage0_3[429], stage0_3[430], stage0_3[431], stage0_3[432], stage0_3[433], stage0_3[434]},
      {stage1_5[67],stage1_4[152],stage1_3[153],stage1_2[153],stage1_1[153]}
   );
   gpc606_5 gpc154 (
      {stage0_1[480], stage0_1[481], stage0_1[482], stage0_1[483], stage0_1[484], stage0_1[485]},
      {stage0_3[435], stage0_3[436], stage0_3[437], stage0_3[438], stage0_3[439], stage0_3[440]},
      {stage1_5[68],stage1_4[153],stage1_3[154],stage1_2[154],stage1_1[154]}
   );
   gpc615_5 gpc155 (
      {stage0_2[427], stage0_2[428], stage0_2[429], stage0_2[430], stage0_2[431]},
      {stage0_3[441]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[69],stage1_4[154],stage1_3[155],stage1_2[155]}
   );
   gpc615_5 gpc156 (
      {stage0_2[432], stage0_2[433], stage0_2[434], stage0_2[435], stage0_2[436]},
      {stage0_3[442]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[70],stage1_4[155],stage1_3[156],stage1_2[156]}
   );
   gpc615_5 gpc157 (
      {stage0_2[437], stage0_2[438], stage0_2[439], stage0_2[440], stage0_2[441]},
      {stage0_3[443]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[71],stage1_4[156],stage1_3[157],stage1_2[157]}
   );
   gpc615_5 gpc158 (
      {stage0_2[442], stage0_2[443], stage0_2[444], stage0_2[445], stage0_2[446]},
      {stage0_3[444]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[72],stage1_4[157],stage1_3[158],stage1_2[158]}
   );
   gpc615_5 gpc159 (
      {stage0_3[445], stage0_3[446], stage0_3[447], stage0_3[448], stage0_3[449]},
      {stage0_4[24]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[4],stage1_5[73],stage1_4[158],stage1_3[159]}
   );
   gpc606_5 gpc160 (
      {stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[1],stage1_6[5],stage1_5[74],stage1_4[159]}
   );
   gpc606_5 gpc161 (
      {stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35], stage0_4[36]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[2],stage1_6[6],stage1_5[75],stage1_4[160]}
   );
   gpc606_5 gpc162 (
      {stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41], stage0_4[42]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[3],stage1_6[7],stage1_5[76],stage1_4[161]}
   );
   gpc606_5 gpc163 (
      {stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47], stage0_4[48]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[4],stage1_6[8],stage1_5[77],stage1_4[162]}
   );
   gpc606_5 gpc164 (
      {stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53], stage0_4[54]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[5],stage1_6[9],stage1_5[78],stage1_4[163]}
   );
   gpc606_5 gpc165 (
      {stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59], stage0_4[60]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[6],stage1_6[10],stage1_5[79],stage1_4[164]}
   );
   gpc606_5 gpc166 (
      {stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65], stage0_4[66]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[7],stage1_6[11],stage1_5[80],stage1_4[165]}
   );
   gpc606_5 gpc167 (
      {stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71], stage0_4[72]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[8],stage1_6[12],stage1_5[81],stage1_4[166]}
   );
   gpc606_5 gpc168 (
      {stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77], stage0_4[78]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[9],stage1_6[13],stage1_5[82],stage1_4[167]}
   );
   gpc606_5 gpc169 (
      {stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83], stage0_4[84]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[10],stage1_6[14],stage1_5[83],stage1_4[168]}
   );
   gpc606_5 gpc170 (
      {stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89], stage0_4[90]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[11],stage1_6[15],stage1_5[84],stage1_4[169]}
   );
   gpc606_5 gpc171 (
      {stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95], stage0_4[96]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[12],stage1_6[16],stage1_5[85],stage1_4[170]}
   );
   gpc606_5 gpc172 (
      {stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101], stage0_4[102]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[13],stage1_6[17],stage1_5[86],stage1_4[171]}
   );
   gpc606_5 gpc173 (
      {stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107], stage0_4[108]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[14],stage1_6[18],stage1_5[87],stage1_4[172]}
   );
   gpc606_5 gpc174 (
      {stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113], stage0_4[114]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[15],stage1_6[19],stage1_5[88],stage1_4[173]}
   );
   gpc606_5 gpc175 (
      {stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119], stage0_4[120]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[16],stage1_6[20],stage1_5[89],stage1_4[174]}
   );
   gpc606_5 gpc176 (
      {stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125], stage0_4[126]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[17],stage1_6[21],stage1_5[90],stage1_4[175]}
   );
   gpc606_5 gpc177 (
      {stage0_4[127], stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131], stage0_4[132]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[18],stage1_6[22],stage1_5[91],stage1_4[176]}
   );
   gpc606_5 gpc178 (
      {stage0_4[133], stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137], stage0_4[138]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[19],stage1_6[23],stage1_5[92],stage1_4[177]}
   );
   gpc606_5 gpc179 (
      {stage0_4[139], stage0_4[140], stage0_4[141], stage0_4[142], stage0_4[143], stage0_4[144]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[20],stage1_6[24],stage1_5[93],stage1_4[178]}
   );
   gpc606_5 gpc180 (
      {stage0_4[145], stage0_4[146], stage0_4[147], stage0_4[148], stage0_4[149], stage0_4[150]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[21],stage1_6[25],stage1_5[94],stage1_4[179]}
   );
   gpc606_5 gpc181 (
      {stage0_4[151], stage0_4[152], stage0_4[153], stage0_4[154], stage0_4[155], stage0_4[156]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[21],stage1_7[22],stage1_6[26],stage1_5[95],stage1_4[180]}
   );
   gpc606_5 gpc182 (
      {stage0_4[157], stage0_4[158], stage0_4[159], stage0_4[160], stage0_4[161], stage0_4[162]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[22],stage1_7[23],stage1_6[27],stage1_5[96],stage1_4[181]}
   );
   gpc606_5 gpc183 (
      {stage0_4[163], stage0_4[164], stage0_4[165], stage0_4[166], stage0_4[167], stage0_4[168]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[23],stage1_7[24],stage1_6[28],stage1_5[97],stage1_4[182]}
   );
   gpc606_5 gpc184 (
      {stage0_4[169], stage0_4[170], stage0_4[171], stage0_4[172], stage0_4[173], stage0_4[174]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[24],stage1_7[25],stage1_6[29],stage1_5[98],stage1_4[183]}
   );
   gpc606_5 gpc185 (
      {stage0_4[175], stage0_4[176], stage0_4[177], stage0_4[178], stage0_4[179], stage0_4[180]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[25],stage1_7[26],stage1_6[30],stage1_5[99],stage1_4[184]}
   );
   gpc606_5 gpc186 (
      {stage0_4[181], stage0_4[182], stage0_4[183], stage0_4[184], stage0_4[185], stage0_4[186]},
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage1_8[26],stage1_7[27],stage1_6[31],stage1_5[100],stage1_4[185]}
   );
   gpc606_5 gpc187 (
      {stage0_4[187], stage0_4[188], stage0_4[189], stage0_4[190], stage0_4[191], stage0_4[192]},
      {stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167]},
      {stage1_8[27],stage1_7[28],stage1_6[32],stage1_5[101],stage1_4[186]}
   );
   gpc606_5 gpc188 (
      {stage0_4[193], stage0_4[194], stage0_4[195], stage0_4[196], stage0_4[197], stage0_4[198]},
      {stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173]},
      {stage1_8[28],stage1_7[29],stage1_6[33],stage1_5[102],stage1_4[187]}
   );
   gpc606_5 gpc189 (
      {stage0_4[199], stage0_4[200], stage0_4[201], stage0_4[202], stage0_4[203], stage0_4[204]},
      {stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179]},
      {stage1_8[29],stage1_7[30],stage1_6[34],stage1_5[103],stage1_4[188]}
   );
   gpc606_5 gpc190 (
      {stage0_4[205], stage0_4[206], stage0_4[207], stage0_4[208], stage0_4[209], stage0_4[210]},
      {stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184], stage0_6[185]},
      {stage1_8[30],stage1_7[31],stage1_6[35],stage1_5[104],stage1_4[189]}
   );
   gpc606_5 gpc191 (
      {stage0_4[211], stage0_4[212], stage0_4[213], stage0_4[214], stage0_4[215], stage0_4[216]},
      {stage0_6[186], stage0_6[187], stage0_6[188], stage0_6[189], stage0_6[190], stage0_6[191]},
      {stage1_8[31],stage1_7[32],stage1_6[36],stage1_5[105],stage1_4[190]}
   );
   gpc606_5 gpc192 (
      {stage0_4[217], stage0_4[218], stage0_4[219], stage0_4[220], stage0_4[221], stage0_4[222]},
      {stage0_6[192], stage0_6[193], stage0_6[194], stage0_6[195], stage0_6[196], stage0_6[197]},
      {stage1_8[32],stage1_7[33],stage1_6[37],stage1_5[106],stage1_4[191]}
   );
   gpc606_5 gpc193 (
      {stage0_4[223], stage0_4[224], stage0_4[225], stage0_4[226], stage0_4[227], stage0_4[228]},
      {stage0_6[198], stage0_6[199], stage0_6[200], stage0_6[201], stage0_6[202], stage0_6[203]},
      {stage1_8[33],stage1_7[34],stage1_6[38],stage1_5[107],stage1_4[192]}
   );
   gpc606_5 gpc194 (
      {stage0_4[229], stage0_4[230], stage0_4[231], stage0_4[232], stage0_4[233], stage0_4[234]},
      {stage0_6[204], stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208], stage0_6[209]},
      {stage1_8[34],stage1_7[35],stage1_6[39],stage1_5[108],stage1_4[193]}
   );
   gpc606_5 gpc195 (
      {stage0_4[235], stage0_4[236], stage0_4[237], stage0_4[238], stage0_4[239], stage0_4[240]},
      {stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214], stage0_6[215]},
      {stage1_8[35],stage1_7[36],stage1_6[40],stage1_5[109],stage1_4[194]}
   );
   gpc606_5 gpc196 (
      {stage0_4[241], stage0_4[242], stage0_4[243], stage0_4[244], stage0_4[245], stage0_4[246]},
      {stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219], stage0_6[220], stage0_6[221]},
      {stage1_8[36],stage1_7[37],stage1_6[41],stage1_5[110],stage1_4[195]}
   );
   gpc606_5 gpc197 (
      {stage0_4[247], stage0_4[248], stage0_4[249], stage0_4[250], stage0_4[251], stage0_4[252]},
      {stage0_6[222], stage0_6[223], stage0_6[224], stage0_6[225], stage0_6[226], stage0_6[227]},
      {stage1_8[37],stage1_7[38],stage1_6[42],stage1_5[111],stage1_4[196]}
   );
   gpc606_5 gpc198 (
      {stage0_4[253], stage0_4[254], stage0_4[255], stage0_4[256], stage0_4[257], stage0_4[258]},
      {stage0_6[228], stage0_6[229], stage0_6[230], stage0_6[231], stage0_6[232], stage0_6[233]},
      {stage1_8[38],stage1_7[39],stage1_6[43],stage1_5[112],stage1_4[197]}
   );
   gpc606_5 gpc199 (
      {stage0_4[259], stage0_4[260], stage0_4[261], stage0_4[262], stage0_4[263], stage0_4[264]},
      {stage0_6[234], stage0_6[235], stage0_6[236], stage0_6[237], stage0_6[238], stage0_6[239]},
      {stage1_8[39],stage1_7[40],stage1_6[44],stage1_5[113],stage1_4[198]}
   );
   gpc606_5 gpc200 (
      {stage0_4[265], stage0_4[266], stage0_4[267], stage0_4[268], stage0_4[269], stage0_4[270]},
      {stage0_6[240], stage0_6[241], stage0_6[242], stage0_6[243], stage0_6[244], stage0_6[245]},
      {stage1_8[40],stage1_7[41],stage1_6[45],stage1_5[114],stage1_4[199]}
   );
   gpc606_5 gpc201 (
      {stage0_4[271], stage0_4[272], stage0_4[273], stage0_4[274], stage0_4[275], stage0_4[276]},
      {stage0_6[246], stage0_6[247], stage0_6[248], stage0_6[249], stage0_6[250], stage0_6[251]},
      {stage1_8[41],stage1_7[42],stage1_6[46],stage1_5[115],stage1_4[200]}
   );
   gpc606_5 gpc202 (
      {stage0_4[277], stage0_4[278], stage0_4[279], stage0_4[280], stage0_4[281], stage0_4[282]},
      {stage0_6[252], stage0_6[253], stage0_6[254], stage0_6[255], stage0_6[256], stage0_6[257]},
      {stage1_8[42],stage1_7[43],stage1_6[47],stage1_5[116],stage1_4[201]}
   );
   gpc606_5 gpc203 (
      {stage0_4[283], stage0_4[284], stage0_4[285], stage0_4[286], stage0_4[287], stage0_4[288]},
      {stage0_6[258], stage0_6[259], stage0_6[260], stage0_6[261], stage0_6[262], stage0_6[263]},
      {stage1_8[43],stage1_7[44],stage1_6[48],stage1_5[117],stage1_4[202]}
   );
   gpc606_5 gpc204 (
      {stage0_4[289], stage0_4[290], stage0_4[291], stage0_4[292], stage0_4[293], stage0_4[294]},
      {stage0_6[264], stage0_6[265], stage0_6[266], stage0_6[267], stage0_6[268], stage0_6[269]},
      {stage1_8[44],stage1_7[45],stage1_6[49],stage1_5[118],stage1_4[203]}
   );
   gpc606_5 gpc205 (
      {stage0_4[295], stage0_4[296], stage0_4[297], stage0_4[298], stage0_4[299], stage0_4[300]},
      {stage0_6[270], stage0_6[271], stage0_6[272], stage0_6[273], stage0_6[274], stage0_6[275]},
      {stage1_8[45],stage1_7[46],stage1_6[50],stage1_5[119],stage1_4[204]}
   );
   gpc606_5 gpc206 (
      {stage0_4[301], stage0_4[302], stage0_4[303], stage0_4[304], stage0_4[305], stage0_4[306]},
      {stage0_6[276], stage0_6[277], stage0_6[278], stage0_6[279], stage0_6[280], stage0_6[281]},
      {stage1_8[46],stage1_7[47],stage1_6[51],stage1_5[120],stage1_4[205]}
   );
   gpc606_5 gpc207 (
      {stage0_4[307], stage0_4[308], stage0_4[309], stage0_4[310], stage0_4[311], stage0_4[312]},
      {stage0_6[282], stage0_6[283], stage0_6[284], stage0_6[285], stage0_6[286], stage0_6[287]},
      {stage1_8[47],stage1_7[48],stage1_6[52],stage1_5[121],stage1_4[206]}
   );
   gpc606_5 gpc208 (
      {stage0_4[313], stage0_4[314], stage0_4[315], stage0_4[316], stage0_4[317], stage0_4[318]},
      {stage0_6[288], stage0_6[289], stage0_6[290], stage0_6[291], stage0_6[292], stage0_6[293]},
      {stage1_8[48],stage1_7[49],stage1_6[53],stage1_5[122],stage1_4[207]}
   );
   gpc606_5 gpc209 (
      {stage0_4[319], stage0_4[320], stage0_4[321], stage0_4[322], stage0_4[323], stage0_4[324]},
      {stage0_6[294], stage0_6[295], stage0_6[296], stage0_6[297], stage0_6[298], stage0_6[299]},
      {stage1_8[49],stage1_7[50],stage1_6[54],stage1_5[123],stage1_4[208]}
   );
   gpc606_5 gpc210 (
      {stage0_4[325], stage0_4[326], stage0_4[327], stage0_4[328], stage0_4[329], stage0_4[330]},
      {stage0_6[300], stage0_6[301], stage0_6[302], stage0_6[303], stage0_6[304], stage0_6[305]},
      {stage1_8[50],stage1_7[51],stage1_6[55],stage1_5[124],stage1_4[209]}
   );
   gpc606_5 gpc211 (
      {stage0_4[331], stage0_4[332], stage0_4[333], stage0_4[334], stage0_4[335], stage0_4[336]},
      {stage0_6[306], stage0_6[307], stage0_6[308], stage0_6[309], stage0_6[310], stage0_6[311]},
      {stage1_8[51],stage1_7[52],stage1_6[56],stage1_5[125],stage1_4[210]}
   );
   gpc606_5 gpc212 (
      {stage0_4[337], stage0_4[338], stage0_4[339], stage0_4[340], stage0_4[341], stage0_4[342]},
      {stage0_6[312], stage0_6[313], stage0_6[314], stage0_6[315], stage0_6[316], stage0_6[317]},
      {stage1_8[52],stage1_7[53],stage1_6[57],stage1_5[126],stage1_4[211]}
   );
   gpc606_5 gpc213 (
      {stage0_4[343], stage0_4[344], stage0_4[345], stage0_4[346], stage0_4[347], stage0_4[348]},
      {stage0_6[318], stage0_6[319], stage0_6[320], stage0_6[321], stage0_6[322], stage0_6[323]},
      {stage1_8[53],stage1_7[54],stage1_6[58],stage1_5[127],stage1_4[212]}
   );
   gpc606_5 gpc214 (
      {stage0_4[349], stage0_4[350], stage0_4[351], stage0_4[352], stage0_4[353], stage0_4[354]},
      {stage0_6[324], stage0_6[325], stage0_6[326], stage0_6[327], stage0_6[328], stage0_6[329]},
      {stage1_8[54],stage1_7[55],stage1_6[59],stage1_5[128],stage1_4[213]}
   );
   gpc606_5 gpc215 (
      {stage0_4[355], stage0_4[356], stage0_4[357], stage0_4[358], stage0_4[359], stage0_4[360]},
      {stage0_6[330], stage0_6[331], stage0_6[332], stage0_6[333], stage0_6[334], stage0_6[335]},
      {stage1_8[55],stage1_7[56],stage1_6[60],stage1_5[129],stage1_4[214]}
   );
   gpc606_5 gpc216 (
      {stage0_4[361], stage0_4[362], stage0_4[363], stage0_4[364], stage0_4[365], stage0_4[366]},
      {stage0_6[336], stage0_6[337], stage0_6[338], stage0_6[339], stage0_6[340], stage0_6[341]},
      {stage1_8[56],stage1_7[57],stage1_6[61],stage1_5[130],stage1_4[215]}
   );
   gpc606_5 gpc217 (
      {stage0_4[367], stage0_4[368], stage0_4[369], stage0_4[370], stage0_4[371], stage0_4[372]},
      {stage0_6[342], stage0_6[343], stage0_6[344], stage0_6[345], stage0_6[346], stage0_6[347]},
      {stage1_8[57],stage1_7[58],stage1_6[62],stage1_5[131],stage1_4[216]}
   );
   gpc606_5 gpc218 (
      {stage0_4[373], stage0_4[374], stage0_4[375], stage0_4[376], stage0_4[377], stage0_4[378]},
      {stage0_6[348], stage0_6[349], stage0_6[350], stage0_6[351], stage0_6[352], stage0_6[353]},
      {stage1_8[58],stage1_7[59],stage1_6[63],stage1_5[132],stage1_4[217]}
   );
   gpc606_5 gpc219 (
      {stage0_4[379], stage0_4[380], stage0_4[381], stage0_4[382], stage0_4[383], stage0_4[384]},
      {stage0_6[354], stage0_6[355], stage0_6[356], stage0_6[357], stage0_6[358], stage0_6[359]},
      {stage1_8[59],stage1_7[60],stage1_6[64],stage1_5[133],stage1_4[218]}
   );
   gpc606_5 gpc220 (
      {stage0_4[385], stage0_4[386], stage0_4[387], stage0_4[388], stage0_4[389], stage0_4[390]},
      {stage0_6[360], stage0_6[361], stage0_6[362], stage0_6[363], stage0_6[364], stage0_6[365]},
      {stage1_8[60],stage1_7[61],stage1_6[65],stage1_5[134],stage1_4[219]}
   );
   gpc606_5 gpc221 (
      {stage0_4[391], stage0_4[392], stage0_4[393], stage0_4[394], stage0_4[395], stage0_4[396]},
      {stage0_6[366], stage0_6[367], stage0_6[368], stage0_6[369], stage0_6[370], stage0_6[371]},
      {stage1_8[61],stage1_7[62],stage1_6[66],stage1_5[135],stage1_4[220]}
   );
   gpc606_5 gpc222 (
      {stage0_4[397], stage0_4[398], stage0_4[399], stage0_4[400], stage0_4[401], stage0_4[402]},
      {stage0_6[372], stage0_6[373], stage0_6[374], stage0_6[375], stage0_6[376], stage0_6[377]},
      {stage1_8[62],stage1_7[63],stage1_6[67],stage1_5[136],stage1_4[221]}
   );
   gpc606_5 gpc223 (
      {stage0_4[403], stage0_4[404], stage0_4[405], stage0_4[406], stage0_4[407], stage0_4[408]},
      {stage0_6[378], stage0_6[379], stage0_6[380], stage0_6[381], stage0_6[382], stage0_6[383]},
      {stage1_8[63],stage1_7[64],stage1_6[68],stage1_5[137],stage1_4[222]}
   );
   gpc606_5 gpc224 (
      {stage0_4[409], stage0_4[410], stage0_4[411], stage0_4[412], stage0_4[413], stage0_4[414]},
      {stage0_6[384], stage0_6[385], stage0_6[386], stage0_6[387], stage0_6[388], stage0_6[389]},
      {stage1_8[64],stage1_7[65],stage1_6[69],stage1_5[138],stage1_4[223]}
   );
   gpc606_5 gpc225 (
      {stage0_4[415], stage0_4[416], stage0_4[417], stage0_4[418], stage0_4[419], stage0_4[420]},
      {stage0_6[390], stage0_6[391], stage0_6[392], stage0_6[393], stage0_6[394], stage0_6[395]},
      {stage1_8[65],stage1_7[66],stage1_6[70],stage1_5[139],stage1_4[224]}
   );
   gpc606_5 gpc226 (
      {stage0_4[421], stage0_4[422], stage0_4[423], stage0_4[424], stage0_4[425], stage0_4[426]},
      {stage0_6[396], stage0_6[397], stage0_6[398], stage0_6[399], stage0_6[400], stage0_6[401]},
      {stage1_8[66],stage1_7[67],stage1_6[71],stage1_5[140],stage1_4[225]}
   );
   gpc606_5 gpc227 (
      {stage0_4[427], stage0_4[428], stage0_4[429], stage0_4[430], stage0_4[431], stage0_4[432]},
      {stage0_6[402], stage0_6[403], stage0_6[404], stage0_6[405], stage0_6[406], stage0_6[407]},
      {stage1_8[67],stage1_7[68],stage1_6[72],stage1_5[141],stage1_4[226]}
   );
   gpc606_5 gpc228 (
      {stage0_4[433], stage0_4[434], stage0_4[435], stage0_4[436], stage0_4[437], stage0_4[438]},
      {stage0_6[408], stage0_6[409], stage0_6[410], stage0_6[411], stage0_6[412], stage0_6[413]},
      {stage1_8[68],stage1_7[69],stage1_6[73],stage1_5[142],stage1_4[227]}
   );
   gpc606_5 gpc229 (
      {stage0_4[439], stage0_4[440], stage0_4[441], stage0_4[442], stage0_4[443], stage0_4[444]},
      {stage0_6[414], stage0_6[415], stage0_6[416], stage0_6[417], stage0_6[418], stage0_6[419]},
      {stage1_8[69],stage1_7[70],stage1_6[74],stage1_5[143],stage1_4[228]}
   );
   gpc606_5 gpc230 (
      {stage0_4[445], stage0_4[446], stage0_4[447], stage0_4[448], stage0_4[449], stage0_4[450]},
      {stage0_6[420], stage0_6[421], stage0_6[422], stage0_6[423], stage0_6[424], stage0_6[425]},
      {stage1_8[70],stage1_7[71],stage1_6[75],stage1_5[144],stage1_4[229]}
   );
   gpc615_5 gpc231 (
      {stage0_4[451], stage0_4[452], stage0_4[453], stage0_4[454], stage0_4[455]},
      {stage0_5[6]},
      {stage0_6[426], stage0_6[427], stage0_6[428], stage0_6[429], stage0_6[430], stage0_6[431]},
      {stage1_8[71],stage1_7[72],stage1_6[76],stage1_5[145],stage1_4[230]}
   );
   gpc615_5 gpc232 (
      {stage0_4[456], stage0_4[457], stage0_4[458], stage0_4[459], stage0_4[460]},
      {stage0_5[7]},
      {stage0_6[432], stage0_6[433], stage0_6[434], stage0_6[435], stage0_6[436], stage0_6[437]},
      {stage1_8[72],stage1_7[73],stage1_6[77],stage1_5[146],stage1_4[231]}
   );
   gpc615_5 gpc233 (
      {stage0_4[461], stage0_4[462], stage0_4[463], stage0_4[464], stage0_4[465]},
      {stage0_5[8]},
      {stage0_6[438], stage0_6[439], stage0_6[440], stage0_6[441], stage0_6[442], stage0_6[443]},
      {stage1_8[73],stage1_7[74],stage1_6[78],stage1_5[147],stage1_4[232]}
   );
   gpc615_5 gpc234 (
      {stage0_4[466], stage0_4[467], stage0_4[468], stage0_4[469], stage0_4[470]},
      {stage0_5[9]},
      {stage0_6[444], stage0_6[445], stage0_6[446], stage0_6[447], stage0_6[448], stage0_6[449]},
      {stage1_8[74],stage1_7[75],stage1_6[79],stage1_5[148],stage1_4[233]}
   );
   gpc615_5 gpc235 (
      {stage0_4[471], stage0_4[472], stage0_4[473], stage0_4[474], stage0_4[475]},
      {stage0_5[10]},
      {stage0_6[450], stage0_6[451], stage0_6[452], stage0_6[453], stage0_6[454], stage0_6[455]},
      {stage1_8[75],stage1_7[76],stage1_6[80],stage1_5[149],stage1_4[234]}
   );
   gpc615_5 gpc236 (
      {stage0_4[476], stage0_4[477], stage0_4[478], stage0_4[479], stage0_4[480]},
      {stage0_5[11]},
      {stage0_6[456], stage0_6[457], stage0_6[458], stage0_6[459], stage0_6[460], stage0_6[461]},
      {stage1_8[76],stage1_7[77],stage1_6[81],stage1_5[150],stage1_4[235]}
   );
   gpc606_5 gpc237 (
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[77],stage1_7[78],stage1_6[82],stage1_5[151]}
   );
   gpc606_5 gpc238 (
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[78],stage1_7[79],stage1_6[83],stage1_5[152]}
   );
   gpc606_5 gpc239 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[79],stage1_7[80],stage1_6[84],stage1_5[153]}
   );
   gpc606_5 gpc240 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[80],stage1_7[81],stage1_6[85],stage1_5[154]}
   );
   gpc606_5 gpc241 (
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[81],stage1_7[82],stage1_6[86],stage1_5[155]}
   );
   gpc606_5 gpc242 (
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[82],stage1_7[83],stage1_6[87],stage1_5[156]}
   );
   gpc606_5 gpc243 (
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[83],stage1_7[84],stage1_6[88],stage1_5[157]}
   );
   gpc606_5 gpc244 (
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[84],stage1_7[85],stage1_6[89],stage1_5[158]}
   );
   gpc606_5 gpc245 (
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[85],stage1_7[86],stage1_6[90],stage1_5[159]}
   );
   gpc606_5 gpc246 (
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[86],stage1_7[87],stage1_6[91],stage1_5[160]}
   );
   gpc606_5 gpc247 (
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[87],stage1_7[88],stage1_6[92],stage1_5[161]}
   );
   gpc606_5 gpc248 (
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[88],stage1_7[89],stage1_6[93],stage1_5[162]}
   );
   gpc606_5 gpc249 (
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[89],stage1_7[90],stage1_6[94],stage1_5[163]}
   );
   gpc606_5 gpc250 (
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[90],stage1_7[91],stage1_6[95],stage1_5[164]}
   );
   gpc606_5 gpc251 (
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[91],stage1_7[92],stage1_6[96],stage1_5[165]}
   );
   gpc606_5 gpc252 (
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[92],stage1_7[93],stage1_6[97],stage1_5[166]}
   );
   gpc606_5 gpc253 (
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[93],stage1_7[94],stage1_6[98],stage1_5[167]}
   );
   gpc606_5 gpc254 (
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[94],stage1_7[95],stage1_6[99],stage1_5[168]}
   );
   gpc606_5 gpc255 (
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[95],stage1_7[96],stage1_6[100],stage1_5[169]}
   );
   gpc606_5 gpc256 (
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[96],stage1_7[97],stage1_6[101],stage1_5[170]}
   );
   gpc606_5 gpc257 (
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[97],stage1_7[98],stage1_6[102],stage1_5[171]}
   );
   gpc606_5 gpc258 (
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[98],stage1_7[99],stage1_6[103],stage1_5[172]}
   );
   gpc606_5 gpc259 (
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[99],stage1_7[100],stage1_6[104],stage1_5[173]}
   );
   gpc606_5 gpc260 (
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[100],stage1_7[101],stage1_6[105],stage1_5[174]}
   );
   gpc606_5 gpc261 (
      {stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[101],stage1_7[102],stage1_6[106],stage1_5[175]}
   );
   gpc606_5 gpc262 (
      {stage0_5[162], stage0_5[163], stage0_5[164], stage0_5[165], stage0_5[166], stage0_5[167]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[102],stage1_7[103],stage1_6[107],stage1_5[176]}
   );
   gpc606_5 gpc263 (
      {stage0_5[168], stage0_5[169], stage0_5[170], stage0_5[171], stage0_5[172], stage0_5[173]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[103],stage1_7[104],stage1_6[108],stage1_5[177]}
   );
   gpc606_5 gpc264 (
      {stage0_5[174], stage0_5[175], stage0_5[176], stage0_5[177], stage0_5[178], stage0_5[179]},
      {stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167]},
      {stage1_9[27],stage1_8[104],stage1_7[105],stage1_6[109],stage1_5[178]}
   );
   gpc606_5 gpc265 (
      {stage0_5[180], stage0_5[181], stage0_5[182], stage0_5[183], stage0_5[184], stage0_5[185]},
      {stage0_7[168], stage0_7[169], stage0_7[170], stage0_7[171], stage0_7[172], stage0_7[173]},
      {stage1_9[28],stage1_8[105],stage1_7[106],stage1_6[110],stage1_5[179]}
   );
   gpc606_5 gpc266 (
      {stage0_5[186], stage0_5[187], stage0_5[188], stage0_5[189], stage0_5[190], stage0_5[191]},
      {stage0_7[174], stage0_7[175], stage0_7[176], stage0_7[177], stage0_7[178], stage0_7[179]},
      {stage1_9[29],stage1_8[106],stage1_7[107],stage1_6[111],stage1_5[180]}
   );
   gpc606_5 gpc267 (
      {stage0_5[192], stage0_5[193], stage0_5[194], stage0_5[195], stage0_5[196], stage0_5[197]},
      {stage0_7[180], stage0_7[181], stage0_7[182], stage0_7[183], stage0_7[184], stage0_7[185]},
      {stage1_9[30],stage1_8[107],stage1_7[108],stage1_6[112],stage1_5[181]}
   );
   gpc606_5 gpc268 (
      {stage0_5[198], stage0_5[199], stage0_5[200], stage0_5[201], stage0_5[202], stage0_5[203]},
      {stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189], stage0_7[190], stage0_7[191]},
      {stage1_9[31],stage1_8[108],stage1_7[109],stage1_6[113],stage1_5[182]}
   );
   gpc606_5 gpc269 (
      {stage0_5[204], stage0_5[205], stage0_5[206], stage0_5[207], stage0_5[208], stage0_5[209]},
      {stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195], stage0_7[196], stage0_7[197]},
      {stage1_9[32],stage1_8[109],stage1_7[110],stage1_6[114],stage1_5[183]}
   );
   gpc606_5 gpc270 (
      {stage0_5[210], stage0_5[211], stage0_5[212], stage0_5[213], stage0_5[214], stage0_5[215]},
      {stage0_7[198], stage0_7[199], stage0_7[200], stage0_7[201], stage0_7[202], stage0_7[203]},
      {stage1_9[33],stage1_8[110],stage1_7[111],stage1_6[115],stage1_5[184]}
   );
   gpc606_5 gpc271 (
      {stage0_5[216], stage0_5[217], stage0_5[218], stage0_5[219], stage0_5[220], stage0_5[221]},
      {stage0_7[204], stage0_7[205], stage0_7[206], stage0_7[207], stage0_7[208], stage0_7[209]},
      {stage1_9[34],stage1_8[111],stage1_7[112],stage1_6[116],stage1_5[185]}
   );
   gpc606_5 gpc272 (
      {stage0_5[222], stage0_5[223], stage0_5[224], stage0_5[225], stage0_5[226], stage0_5[227]},
      {stage0_7[210], stage0_7[211], stage0_7[212], stage0_7[213], stage0_7[214], stage0_7[215]},
      {stage1_9[35],stage1_8[112],stage1_7[113],stage1_6[117],stage1_5[186]}
   );
   gpc606_5 gpc273 (
      {stage0_5[228], stage0_5[229], stage0_5[230], stage0_5[231], stage0_5[232], stage0_5[233]},
      {stage0_7[216], stage0_7[217], stage0_7[218], stage0_7[219], stage0_7[220], stage0_7[221]},
      {stage1_9[36],stage1_8[113],stage1_7[114],stage1_6[118],stage1_5[187]}
   );
   gpc606_5 gpc274 (
      {stage0_5[234], stage0_5[235], stage0_5[236], stage0_5[237], stage0_5[238], stage0_5[239]},
      {stage0_7[222], stage0_7[223], stage0_7[224], stage0_7[225], stage0_7[226], stage0_7[227]},
      {stage1_9[37],stage1_8[114],stage1_7[115],stage1_6[119],stage1_5[188]}
   );
   gpc606_5 gpc275 (
      {stage0_5[240], stage0_5[241], stage0_5[242], stage0_5[243], stage0_5[244], stage0_5[245]},
      {stage0_7[228], stage0_7[229], stage0_7[230], stage0_7[231], stage0_7[232], stage0_7[233]},
      {stage1_9[38],stage1_8[115],stage1_7[116],stage1_6[120],stage1_5[189]}
   );
   gpc606_5 gpc276 (
      {stage0_5[246], stage0_5[247], stage0_5[248], stage0_5[249], stage0_5[250], stage0_5[251]},
      {stage0_7[234], stage0_7[235], stage0_7[236], stage0_7[237], stage0_7[238], stage0_7[239]},
      {stage1_9[39],stage1_8[116],stage1_7[117],stage1_6[121],stage1_5[190]}
   );
   gpc606_5 gpc277 (
      {stage0_5[252], stage0_5[253], stage0_5[254], stage0_5[255], stage0_5[256], stage0_5[257]},
      {stage0_7[240], stage0_7[241], stage0_7[242], stage0_7[243], stage0_7[244], stage0_7[245]},
      {stage1_9[40],stage1_8[117],stage1_7[118],stage1_6[122],stage1_5[191]}
   );
   gpc606_5 gpc278 (
      {stage0_5[258], stage0_5[259], stage0_5[260], stage0_5[261], stage0_5[262], stage0_5[263]},
      {stage0_7[246], stage0_7[247], stage0_7[248], stage0_7[249], stage0_7[250], stage0_7[251]},
      {stage1_9[41],stage1_8[118],stage1_7[119],stage1_6[123],stage1_5[192]}
   );
   gpc606_5 gpc279 (
      {stage0_5[264], stage0_5[265], stage0_5[266], stage0_5[267], stage0_5[268], stage0_5[269]},
      {stage0_7[252], stage0_7[253], stage0_7[254], stage0_7[255], stage0_7[256], stage0_7[257]},
      {stage1_9[42],stage1_8[119],stage1_7[120],stage1_6[124],stage1_5[193]}
   );
   gpc606_5 gpc280 (
      {stage0_5[270], stage0_5[271], stage0_5[272], stage0_5[273], stage0_5[274], stage0_5[275]},
      {stage0_7[258], stage0_7[259], stage0_7[260], stage0_7[261], stage0_7[262], stage0_7[263]},
      {stage1_9[43],stage1_8[120],stage1_7[121],stage1_6[125],stage1_5[194]}
   );
   gpc606_5 gpc281 (
      {stage0_5[276], stage0_5[277], stage0_5[278], stage0_5[279], stage0_5[280], stage0_5[281]},
      {stage0_7[264], stage0_7[265], stage0_7[266], stage0_7[267], stage0_7[268], stage0_7[269]},
      {stage1_9[44],stage1_8[121],stage1_7[122],stage1_6[126],stage1_5[195]}
   );
   gpc606_5 gpc282 (
      {stage0_5[282], stage0_5[283], stage0_5[284], stage0_5[285], stage0_5[286], stage0_5[287]},
      {stage0_7[270], stage0_7[271], stage0_7[272], stage0_7[273], stage0_7[274], stage0_7[275]},
      {stage1_9[45],stage1_8[122],stage1_7[123],stage1_6[127],stage1_5[196]}
   );
   gpc606_5 gpc283 (
      {stage0_5[288], stage0_5[289], stage0_5[290], stage0_5[291], stage0_5[292], stage0_5[293]},
      {stage0_7[276], stage0_7[277], stage0_7[278], stage0_7[279], stage0_7[280], stage0_7[281]},
      {stage1_9[46],stage1_8[123],stage1_7[124],stage1_6[128],stage1_5[197]}
   );
   gpc606_5 gpc284 (
      {stage0_5[294], stage0_5[295], stage0_5[296], stage0_5[297], stage0_5[298], stage0_5[299]},
      {stage0_7[282], stage0_7[283], stage0_7[284], stage0_7[285], stage0_7[286], stage0_7[287]},
      {stage1_9[47],stage1_8[124],stage1_7[125],stage1_6[129],stage1_5[198]}
   );
   gpc606_5 gpc285 (
      {stage0_5[300], stage0_5[301], stage0_5[302], stage0_5[303], stage0_5[304], stage0_5[305]},
      {stage0_7[288], stage0_7[289], stage0_7[290], stage0_7[291], stage0_7[292], stage0_7[293]},
      {stage1_9[48],stage1_8[125],stage1_7[126],stage1_6[130],stage1_5[199]}
   );
   gpc606_5 gpc286 (
      {stage0_5[306], stage0_5[307], stage0_5[308], stage0_5[309], stage0_5[310], stage0_5[311]},
      {stage0_7[294], stage0_7[295], stage0_7[296], stage0_7[297], stage0_7[298], stage0_7[299]},
      {stage1_9[49],stage1_8[126],stage1_7[127],stage1_6[131],stage1_5[200]}
   );
   gpc606_5 gpc287 (
      {stage0_5[312], stage0_5[313], stage0_5[314], stage0_5[315], stage0_5[316], stage0_5[317]},
      {stage0_7[300], stage0_7[301], stage0_7[302], stage0_7[303], stage0_7[304], stage0_7[305]},
      {stage1_9[50],stage1_8[127],stage1_7[128],stage1_6[132],stage1_5[201]}
   );
   gpc606_5 gpc288 (
      {stage0_5[318], stage0_5[319], stage0_5[320], stage0_5[321], stage0_5[322], stage0_5[323]},
      {stage0_7[306], stage0_7[307], stage0_7[308], stage0_7[309], stage0_7[310], stage0_7[311]},
      {stage1_9[51],stage1_8[128],stage1_7[129],stage1_6[133],stage1_5[202]}
   );
   gpc606_5 gpc289 (
      {stage0_5[324], stage0_5[325], stage0_5[326], stage0_5[327], stage0_5[328], stage0_5[329]},
      {stage0_7[312], stage0_7[313], stage0_7[314], stage0_7[315], stage0_7[316], stage0_7[317]},
      {stage1_9[52],stage1_8[129],stage1_7[130],stage1_6[134],stage1_5[203]}
   );
   gpc606_5 gpc290 (
      {stage0_5[330], stage0_5[331], stage0_5[332], stage0_5[333], stage0_5[334], stage0_5[335]},
      {stage0_7[318], stage0_7[319], stage0_7[320], stage0_7[321], stage0_7[322], stage0_7[323]},
      {stage1_9[53],stage1_8[130],stage1_7[131],stage1_6[135],stage1_5[204]}
   );
   gpc606_5 gpc291 (
      {stage0_5[336], stage0_5[337], stage0_5[338], stage0_5[339], stage0_5[340], stage0_5[341]},
      {stage0_7[324], stage0_7[325], stage0_7[326], stage0_7[327], stage0_7[328], stage0_7[329]},
      {stage1_9[54],stage1_8[131],stage1_7[132],stage1_6[136],stage1_5[205]}
   );
   gpc606_5 gpc292 (
      {stage0_5[342], stage0_5[343], stage0_5[344], stage0_5[345], stage0_5[346], stage0_5[347]},
      {stage0_7[330], stage0_7[331], stage0_7[332], stage0_7[333], stage0_7[334], stage0_7[335]},
      {stage1_9[55],stage1_8[132],stage1_7[133],stage1_6[137],stage1_5[206]}
   );
   gpc606_5 gpc293 (
      {stage0_5[348], stage0_5[349], stage0_5[350], stage0_5[351], stage0_5[352], stage0_5[353]},
      {stage0_7[336], stage0_7[337], stage0_7[338], stage0_7[339], stage0_7[340], stage0_7[341]},
      {stage1_9[56],stage1_8[133],stage1_7[134],stage1_6[138],stage1_5[207]}
   );
   gpc606_5 gpc294 (
      {stage0_5[354], stage0_5[355], stage0_5[356], stage0_5[357], stage0_5[358], stage0_5[359]},
      {stage0_7[342], stage0_7[343], stage0_7[344], stage0_7[345], stage0_7[346], stage0_7[347]},
      {stage1_9[57],stage1_8[134],stage1_7[135],stage1_6[139],stage1_5[208]}
   );
   gpc606_5 gpc295 (
      {stage0_5[360], stage0_5[361], stage0_5[362], stage0_5[363], stage0_5[364], stage0_5[365]},
      {stage0_7[348], stage0_7[349], stage0_7[350], stage0_7[351], stage0_7[352], stage0_7[353]},
      {stage1_9[58],stage1_8[135],stage1_7[136],stage1_6[140],stage1_5[209]}
   );
   gpc606_5 gpc296 (
      {stage0_5[366], stage0_5[367], stage0_5[368], stage0_5[369], stage0_5[370], stage0_5[371]},
      {stage0_7[354], stage0_7[355], stage0_7[356], stage0_7[357], stage0_7[358], stage0_7[359]},
      {stage1_9[59],stage1_8[136],stage1_7[137],stage1_6[141],stage1_5[210]}
   );
   gpc606_5 gpc297 (
      {stage0_5[372], stage0_5[373], stage0_5[374], stage0_5[375], stage0_5[376], stage0_5[377]},
      {stage0_7[360], stage0_7[361], stage0_7[362], stage0_7[363], stage0_7[364], stage0_7[365]},
      {stage1_9[60],stage1_8[137],stage1_7[138],stage1_6[142],stage1_5[211]}
   );
   gpc606_5 gpc298 (
      {stage0_5[378], stage0_5[379], stage0_5[380], stage0_5[381], stage0_5[382], stage0_5[383]},
      {stage0_7[366], stage0_7[367], stage0_7[368], stage0_7[369], stage0_7[370], stage0_7[371]},
      {stage1_9[61],stage1_8[138],stage1_7[139],stage1_6[143],stage1_5[212]}
   );
   gpc606_5 gpc299 (
      {stage0_5[384], stage0_5[385], stage0_5[386], stage0_5[387], stage0_5[388], stage0_5[389]},
      {stage0_7[372], stage0_7[373], stage0_7[374], stage0_7[375], stage0_7[376], stage0_7[377]},
      {stage1_9[62],stage1_8[139],stage1_7[140],stage1_6[144],stage1_5[213]}
   );
   gpc606_5 gpc300 (
      {stage0_5[390], stage0_5[391], stage0_5[392], stage0_5[393], stage0_5[394], stage0_5[395]},
      {stage0_7[378], stage0_7[379], stage0_7[380], stage0_7[381], stage0_7[382], stage0_7[383]},
      {stage1_9[63],stage1_8[140],stage1_7[141],stage1_6[145],stage1_5[214]}
   );
   gpc606_5 gpc301 (
      {stage0_5[396], stage0_5[397], stage0_5[398], stage0_5[399], stage0_5[400], stage0_5[401]},
      {stage0_7[384], stage0_7[385], stage0_7[386], stage0_7[387], stage0_7[388], stage0_7[389]},
      {stage1_9[64],stage1_8[141],stage1_7[142],stage1_6[146],stage1_5[215]}
   );
   gpc606_5 gpc302 (
      {stage0_5[402], stage0_5[403], stage0_5[404], stage0_5[405], stage0_5[406], stage0_5[407]},
      {stage0_7[390], stage0_7[391], stage0_7[392], stage0_7[393], stage0_7[394], stage0_7[395]},
      {stage1_9[65],stage1_8[142],stage1_7[143],stage1_6[147],stage1_5[216]}
   );
   gpc606_5 gpc303 (
      {stage0_5[408], stage0_5[409], stage0_5[410], stage0_5[411], stage0_5[412], stage0_5[413]},
      {stage0_7[396], stage0_7[397], stage0_7[398], stage0_7[399], stage0_7[400], stage0_7[401]},
      {stage1_9[66],stage1_8[143],stage1_7[144],stage1_6[148],stage1_5[217]}
   );
   gpc606_5 gpc304 (
      {stage0_5[414], stage0_5[415], stage0_5[416], stage0_5[417], stage0_5[418], stage0_5[419]},
      {stage0_7[402], stage0_7[403], stage0_7[404], stage0_7[405], stage0_7[406], stage0_7[407]},
      {stage1_9[67],stage1_8[144],stage1_7[145],stage1_6[149],stage1_5[218]}
   );
   gpc606_5 gpc305 (
      {stage0_5[420], stage0_5[421], stage0_5[422], stage0_5[423], stage0_5[424], stage0_5[425]},
      {stage0_7[408], stage0_7[409], stage0_7[410], stage0_7[411], stage0_7[412], stage0_7[413]},
      {stage1_9[68],stage1_8[145],stage1_7[146],stage1_6[150],stage1_5[219]}
   );
   gpc606_5 gpc306 (
      {stage0_5[426], stage0_5[427], stage0_5[428], stage0_5[429], stage0_5[430], stage0_5[431]},
      {stage0_7[414], stage0_7[415], stage0_7[416], stage0_7[417], stage0_7[418], stage0_7[419]},
      {stage1_9[69],stage1_8[146],stage1_7[147],stage1_6[151],stage1_5[220]}
   );
   gpc606_5 gpc307 (
      {stage0_5[432], stage0_5[433], stage0_5[434], stage0_5[435], stage0_5[436], stage0_5[437]},
      {stage0_7[420], stage0_7[421], stage0_7[422], stage0_7[423], stage0_7[424], stage0_7[425]},
      {stage1_9[70],stage1_8[147],stage1_7[148],stage1_6[152],stage1_5[221]}
   );
   gpc606_5 gpc308 (
      {stage0_5[438], stage0_5[439], stage0_5[440], stage0_5[441], stage0_5[442], stage0_5[443]},
      {stage0_7[426], stage0_7[427], stage0_7[428], stage0_7[429], stage0_7[430], stage0_7[431]},
      {stage1_9[71],stage1_8[148],stage1_7[149],stage1_6[153],stage1_5[222]}
   );
   gpc606_5 gpc309 (
      {stage0_5[444], stage0_5[445], stage0_5[446], stage0_5[447], stage0_5[448], stage0_5[449]},
      {stage0_7[432], stage0_7[433], stage0_7[434], stage0_7[435], stage0_7[436], stage0_7[437]},
      {stage1_9[72],stage1_8[149],stage1_7[150],stage1_6[154],stage1_5[223]}
   );
   gpc606_5 gpc310 (
      {stage0_5[450], stage0_5[451], stage0_5[452], stage0_5[453], stage0_5[454], stage0_5[455]},
      {stage0_7[438], stage0_7[439], stage0_7[440], stage0_7[441], stage0_7[442], stage0_7[443]},
      {stage1_9[73],stage1_8[150],stage1_7[151],stage1_6[155],stage1_5[224]}
   );
   gpc606_5 gpc311 (
      {stage0_5[456], stage0_5[457], stage0_5[458], stage0_5[459], stage0_5[460], stage0_5[461]},
      {stage0_7[444], stage0_7[445], stage0_7[446], stage0_7[447], stage0_7[448], stage0_7[449]},
      {stage1_9[74],stage1_8[151],stage1_7[152],stage1_6[156],stage1_5[225]}
   );
   gpc606_5 gpc312 (
      {stage0_5[462], stage0_5[463], stage0_5[464], stage0_5[465], stage0_5[466], stage0_5[467]},
      {stage0_7[450], stage0_7[451], stage0_7[452], stage0_7[453], stage0_7[454], stage0_7[455]},
      {stage1_9[75],stage1_8[152],stage1_7[153],stage1_6[157],stage1_5[226]}
   );
   gpc606_5 gpc313 (
      {stage0_5[468], stage0_5[469], stage0_5[470], stage0_5[471], stage0_5[472], stage0_5[473]},
      {stage0_7[456], stage0_7[457], stage0_7[458], stage0_7[459], stage0_7[460], stage0_7[461]},
      {stage1_9[76],stage1_8[153],stage1_7[154],stage1_6[158],stage1_5[227]}
   );
   gpc606_5 gpc314 (
      {stage0_5[474], stage0_5[475], stage0_5[476], stage0_5[477], stage0_5[478], stage0_5[479]},
      {stage0_7[462], stage0_7[463], stage0_7[464], stage0_7[465], stage0_7[466], stage0_7[467]},
      {stage1_9[77],stage1_8[154],stage1_7[155],stage1_6[159],stage1_5[228]}
   );
   gpc606_5 gpc315 (
      {stage0_5[480], stage0_5[481], stage0_5[482], stage0_5[483], stage0_5[484], stage0_5[485]},
      {stage0_7[468], stage0_7[469], stage0_7[470], stage0_7[471], stage0_7[472], stage0_7[473]},
      {stage1_9[78],stage1_8[155],stage1_7[156],stage1_6[160],stage1_5[229]}
   );
   gpc606_5 gpc316 (
      {stage0_6[462], stage0_6[463], stage0_6[464], stage0_6[465], stage0_6[466], stage0_6[467]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[79],stage1_8[156],stage1_7[157],stage1_6[161]}
   );
   gpc606_5 gpc317 (
      {stage0_6[468], stage0_6[469], stage0_6[470], stage0_6[471], stage0_6[472], stage0_6[473]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[80],stage1_8[157],stage1_7[158],stage1_6[162]}
   );
   gpc606_5 gpc318 (
      {stage0_6[474], stage0_6[475], stage0_6[476], stage0_6[477], stage0_6[478], stage0_6[479]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[81],stage1_8[158],stage1_7[159],stage1_6[163]}
   );
   gpc606_5 gpc319 (
      {stage0_7[474], stage0_7[475], stage0_7[476], stage0_7[477], stage0_7[478], stage0_7[479]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[3],stage1_9[82],stage1_8[159],stage1_7[160]}
   );
   gpc606_5 gpc320 (
      {stage0_7[480], stage0_7[481], stage0_7[482], stage0_7[483], stage0_7[484], stage0_7[485]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[4],stage1_9[83],stage1_8[160],stage1_7[161]}
   );
   gpc606_5 gpc321 (
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[2],stage1_10[5],stage1_9[84],stage1_8[161]}
   );
   gpc606_5 gpc322 (
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[3],stage1_10[6],stage1_9[85],stage1_8[162]}
   );
   gpc606_5 gpc323 (
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[4],stage1_10[7],stage1_9[86],stage1_8[163]}
   );
   gpc606_5 gpc324 (
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[5],stage1_10[8],stage1_9[87],stage1_8[164]}
   );
   gpc606_5 gpc325 (
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[6],stage1_10[9],stage1_9[88],stage1_8[165]}
   );
   gpc606_5 gpc326 (
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[7],stage1_10[10],stage1_9[89],stage1_8[166]}
   );
   gpc606_5 gpc327 (
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[8],stage1_10[11],stage1_9[90],stage1_8[167]}
   );
   gpc606_5 gpc328 (
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[9],stage1_10[12],stage1_9[91],stage1_8[168]}
   );
   gpc606_5 gpc329 (
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[10],stage1_10[13],stage1_9[92],stage1_8[169]}
   );
   gpc606_5 gpc330 (
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[11],stage1_10[14],stage1_9[93],stage1_8[170]}
   );
   gpc606_5 gpc331 (
      {stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[12],stage1_10[15],stage1_9[94],stage1_8[171]}
   );
   gpc606_5 gpc332 (
      {stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[13],stage1_10[16],stage1_9[95],stage1_8[172]}
   );
   gpc606_5 gpc333 (
      {stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[14],stage1_10[17],stage1_9[96],stage1_8[173]}
   );
   gpc606_5 gpc334 (
      {stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[15],stage1_10[18],stage1_9[97],stage1_8[174]}
   );
   gpc606_5 gpc335 (
      {stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[16],stage1_10[19],stage1_9[98],stage1_8[175]}
   );
   gpc606_5 gpc336 (
      {stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[17],stage1_10[20],stage1_9[99],stage1_8[176]}
   );
   gpc606_5 gpc337 (
      {stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[18],stage1_10[21],stage1_9[100],stage1_8[177]}
   );
   gpc606_5 gpc338 (
      {stage0_8[120], stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[19],stage1_10[22],stage1_9[101],stage1_8[178]}
   );
   gpc606_5 gpc339 (
      {stage0_8[126], stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[20],stage1_10[23],stage1_9[102],stage1_8[179]}
   );
   gpc606_5 gpc340 (
      {stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[21],stage1_10[24],stage1_9[103],stage1_8[180]}
   );
   gpc606_5 gpc341 (
      {stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[22],stage1_10[25],stage1_9[104],stage1_8[181]}
   );
   gpc606_5 gpc342 (
      {stage0_8[144], stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[23],stage1_10[26],stage1_9[105],stage1_8[182]}
   );
   gpc606_5 gpc343 (
      {stage0_8[150], stage0_8[151], stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[24],stage1_10[27],stage1_9[106],stage1_8[183]}
   );
   gpc606_5 gpc344 (
      {stage0_8[156], stage0_8[157], stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[25],stage1_10[28],stage1_9[107],stage1_8[184]}
   );
   gpc606_5 gpc345 (
      {stage0_8[162], stage0_8[163], stage0_8[164], stage0_8[165], stage0_8[166], stage0_8[167]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[26],stage1_10[29],stage1_9[108],stage1_8[185]}
   );
   gpc606_5 gpc346 (
      {stage0_8[168], stage0_8[169], stage0_8[170], stage0_8[171], stage0_8[172], stage0_8[173]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[27],stage1_10[30],stage1_9[109],stage1_8[186]}
   );
   gpc606_5 gpc347 (
      {stage0_8[174], stage0_8[175], stage0_8[176], stage0_8[177], stage0_8[178], stage0_8[179]},
      {stage0_10[156], stage0_10[157], stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161]},
      {stage1_12[26],stage1_11[28],stage1_10[31],stage1_9[110],stage1_8[187]}
   );
   gpc606_5 gpc348 (
      {stage0_8[180], stage0_8[181], stage0_8[182], stage0_8[183], stage0_8[184], stage0_8[185]},
      {stage0_10[162], stage0_10[163], stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167]},
      {stage1_12[27],stage1_11[29],stage1_10[32],stage1_9[111],stage1_8[188]}
   );
   gpc606_5 gpc349 (
      {stage0_8[186], stage0_8[187], stage0_8[188], stage0_8[189], stage0_8[190], stage0_8[191]},
      {stage0_10[168], stage0_10[169], stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173]},
      {stage1_12[28],stage1_11[30],stage1_10[33],stage1_9[112],stage1_8[189]}
   );
   gpc606_5 gpc350 (
      {stage0_8[192], stage0_8[193], stage0_8[194], stage0_8[195], stage0_8[196], stage0_8[197]},
      {stage0_10[174], stage0_10[175], stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179]},
      {stage1_12[29],stage1_11[31],stage1_10[34],stage1_9[113],stage1_8[190]}
   );
   gpc606_5 gpc351 (
      {stage0_8[198], stage0_8[199], stage0_8[200], stage0_8[201], stage0_8[202], stage0_8[203]},
      {stage0_10[180], stage0_10[181], stage0_10[182], stage0_10[183], stage0_10[184], stage0_10[185]},
      {stage1_12[30],stage1_11[32],stage1_10[35],stage1_9[114],stage1_8[191]}
   );
   gpc606_5 gpc352 (
      {stage0_8[204], stage0_8[205], stage0_8[206], stage0_8[207], stage0_8[208], stage0_8[209]},
      {stage0_10[186], stage0_10[187], stage0_10[188], stage0_10[189], stage0_10[190], stage0_10[191]},
      {stage1_12[31],stage1_11[33],stage1_10[36],stage1_9[115],stage1_8[192]}
   );
   gpc606_5 gpc353 (
      {stage0_8[210], stage0_8[211], stage0_8[212], stage0_8[213], stage0_8[214], stage0_8[215]},
      {stage0_10[192], stage0_10[193], stage0_10[194], stage0_10[195], stage0_10[196], stage0_10[197]},
      {stage1_12[32],stage1_11[34],stage1_10[37],stage1_9[116],stage1_8[193]}
   );
   gpc606_5 gpc354 (
      {stage0_8[216], stage0_8[217], stage0_8[218], stage0_8[219], stage0_8[220], stage0_8[221]},
      {stage0_10[198], stage0_10[199], stage0_10[200], stage0_10[201], stage0_10[202], stage0_10[203]},
      {stage1_12[33],stage1_11[35],stage1_10[38],stage1_9[117],stage1_8[194]}
   );
   gpc606_5 gpc355 (
      {stage0_8[222], stage0_8[223], stage0_8[224], stage0_8[225], stage0_8[226], stage0_8[227]},
      {stage0_10[204], stage0_10[205], stage0_10[206], stage0_10[207], stage0_10[208], stage0_10[209]},
      {stage1_12[34],stage1_11[36],stage1_10[39],stage1_9[118],stage1_8[195]}
   );
   gpc606_5 gpc356 (
      {stage0_8[228], stage0_8[229], stage0_8[230], stage0_8[231], stage0_8[232], stage0_8[233]},
      {stage0_10[210], stage0_10[211], stage0_10[212], stage0_10[213], stage0_10[214], stage0_10[215]},
      {stage1_12[35],stage1_11[37],stage1_10[40],stage1_9[119],stage1_8[196]}
   );
   gpc606_5 gpc357 (
      {stage0_8[234], stage0_8[235], stage0_8[236], stage0_8[237], stage0_8[238], stage0_8[239]},
      {stage0_10[216], stage0_10[217], stage0_10[218], stage0_10[219], stage0_10[220], stage0_10[221]},
      {stage1_12[36],stage1_11[38],stage1_10[41],stage1_9[120],stage1_8[197]}
   );
   gpc606_5 gpc358 (
      {stage0_8[240], stage0_8[241], stage0_8[242], stage0_8[243], stage0_8[244], stage0_8[245]},
      {stage0_10[222], stage0_10[223], stage0_10[224], stage0_10[225], stage0_10[226], stage0_10[227]},
      {stage1_12[37],stage1_11[39],stage1_10[42],stage1_9[121],stage1_8[198]}
   );
   gpc606_5 gpc359 (
      {stage0_8[246], stage0_8[247], stage0_8[248], stage0_8[249], stage0_8[250], stage0_8[251]},
      {stage0_10[228], stage0_10[229], stage0_10[230], stage0_10[231], stage0_10[232], stage0_10[233]},
      {stage1_12[38],stage1_11[40],stage1_10[43],stage1_9[122],stage1_8[199]}
   );
   gpc606_5 gpc360 (
      {stage0_8[252], stage0_8[253], stage0_8[254], stage0_8[255], stage0_8[256], stage0_8[257]},
      {stage0_10[234], stage0_10[235], stage0_10[236], stage0_10[237], stage0_10[238], stage0_10[239]},
      {stage1_12[39],stage1_11[41],stage1_10[44],stage1_9[123],stage1_8[200]}
   );
   gpc606_5 gpc361 (
      {stage0_8[258], stage0_8[259], stage0_8[260], stage0_8[261], stage0_8[262], stage0_8[263]},
      {stage0_10[240], stage0_10[241], stage0_10[242], stage0_10[243], stage0_10[244], stage0_10[245]},
      {stage1_12[40],stage1_11[42],stage1_10[45],stage1_9[124],stage1_8[201]}
   );
   gpc606_5 gpc362 (
      {stage0_8[264], stage0_8[265], stage0_8[266], stage0_8[267], stage0_8[268], stage0_8[269]},
      {stage0_10[246], stage0_10[247], stage0_10[248], stage0_10[249], stage0_10[250], stage0_10[251]},
      {stage1_12[41],stage1_11[43],stage1_10[46],stage1_9[125],stage1_8[202]}
   );
   gpc606_5 gpc363 (
      {stage0_8[270], stage0_8[271], stage0_8[272], stage0_8[273], stage0_8[274], stage0_8[275]},
      {stage0_10[252], stage0_10[253], stage0_10[254], stage0_10[255], stage0_10[256], stage0_10[257]},
      {stage1_12[42],stage1_11[44],stage1_10[47],stage1_9[126],stage1_8[203]}
   );
   gpc606_5 gpc364 (
      {stage0_8[276], stage0_8[277], stage0_8[278], stage0_8[279], stage0_8[280], stage0_8[281]},
      {stage0_10[258], stage0_10[259], stage0_10[260], stage0_10[261], stage0_10[262], stage0_10[263]},
      {stage1_12[43],stage1_11[45],stage1_10[48],stage1_9[127],stage1_8[204]}
   );
   gpc606_5 gpc365 (
      {stage0_8[282], stage0_8[283], stage0_8[284], stage0_8[285], stage0_8[286], stage0_8[287]},
      {stage0_10[264], stage0_10[265], stage0_10[266], stage0_10[267], stage0_10[268], stage0_10[269]},
      {stage1_12[44],stage1_11[46],stage1_10[49],stage1_9[128],stage1_8[205]}
   );
   gpc606_5 gpc366 (
      {stage0_8[288], stage0_8[289], stage0_8[290], stage0_8[291], stage0_8[292], stage0_8[293]},
      {stage0_10[270], stage0_10[271], stage0_10[272], stage0_10[273], stage0_10[274], stage0_10[275]},
      {stage1_12[45],stage1_11[47],stage1_10[50],stage1_9[129],stage1_8[206]}
   );
   gpc606_5 gpc367 (
      {stage0_8[294], stage0_8[295], stage0_8[296], stage0_8[297], stage0_8[298], stage0_8[299]},
      {stage0_10[276], stage0_10[277], stage0_10[278], stage0_10[279], stage0_10[280], stage0_10[281]},
      {stage1_12[46],stage1_11[48],stage1_10[51],stage1_9[130],stage1_8[207]}
   );
   gpc606_5 gpc368 (
      {stage0_8[300], stage0_8[301], stage0_8[302], stage0_8[303], stage0_8[304], stage0_8[305]},
      {stage0_10[282], stage0_10[283], stage0_10[284], stage0_10[285], stage0_10[286], stage0_10[287]},
      {stage1_12[47],stage1_11[49],stage1_10[52],stage1_9[131],stage1_8[208]}
   );
   gpc606_5 gpc369 (
      {stage0_8[306], stage0_8[307], stage0_8[308], stage0_8[309], stage0_8[310], stage0_8[311]},
      {stage0_10[288], stage0_10[289], stage0_10[290], stage0_10[291], stage0_10[292], stage0_10[293]},
      {stage1_12[48],stage1_11[50],stage1_10[53],stage1_9[132],stage1_8[209]}
   );
   gpc606_5 gpc370 (
      {stage0_8[312], stage0_8[313], stage0_8[314], stage0_8[315], stage0_8[316], stage0_8[317]},
      {stage0_10[294], stage0_10[295], stage0_10[296], stage0_10[297], stage0_10[298], stage0_10[299]},
      {stage1_12[49],stage1_11[51],stage1_10[54],stage1_9[133],stage1_8[210]}
   );
   gpc606_5 gpc371 (
      {stage0_8[318], stage0_8[319], stage0_8[320], stage0_8[321], stage0_8[322], stage0_8[323]},
      {stage0_10[300], stage0_10[301], stage0_10[302], stage0_10[303], stage0_10[304], stage0_10[305]},
      {stage1_12[50],stage1_11[52],stage1_10[55],stage1_9[134],stage1_8[211]}
   );
   gpc606_5 gpc372 (
      {stage0_8[324], stage0_8[325], stage0_8[326], stage0_8[327], stage0_8[328], stage0_8[329]},
      {stage0_10[306], stage0_10[307], stage0_10[308], stage0_10[309], stage0_10[310], stage0_10[311]},
      {stage1_12[51],stage1_11[53],stage1_10[56],stage1_9[135],stage1_8[212]}
   );
   gpc606_5 gpc373 (
      {stage0_8[330], stage0_8[331], stage0_8[332], stage0_8[333], stage0_8[334], stage0_8[335]},
      {stage0_10[312], stage0_10[313], stage0_10[314], stage0_10[315], stage0_10[316], stage0_10[317]},
      {stage1_12[52],stage1_11[54],stage1_10[57],stage1_9[136],stage1_8[213]}
   );
   gpc606_5 gpc374 (
      {stage0_8[336], stage0_8[337], stage0_8[338], stage0_8[339], stage0_8[340], stage0_8[341]},
      {stage0_10[318], stage0_10[319], stage0_10[320], stage0_10[321], stage0_10[322], stage0_10[323]},
      {stage1_12[53],stage1_11[55],stage1_10[58],stage1_9[137],stage1_8[214]}
   );
   gpc606_5 gpc375 (
      {stage0_8[342], stage0_8[343], stage0_8[344], stage0_8[345], stage0_8[346], stage0_8[347]},
      {stage0_10[324], stage0_10[325], stage0_10[326], stage0_10[327], stage0_10[328], stage0_10[329]},
      {stage1_12[54],stage1_11[56],stage1_10[59],stage1_9[138],stage1_8[215]}
   );
   gpc606_5 gpc376 (
      {stage0_8[348], stage0_8[349], stage0_8[350], stage0_8[351], stage0_8[352], stage0_8[353]},
      {stage0_10[330], stage0_10[331], stage0_10[332], stage0_10[333], stage0_10[334], stage0_10[335]},
      {stage1_12[55],stage1_11[57],stage1_10[60],stage1_9[139],stage1_8[216]}
   );
   gpc606_5 gpc377 (
      {stage0_8[354], stage0_8[355], stage0_8[356], stage0_8[357], stage0_8[358], stage0_8[359]},
      {stage0_10[336], stage0_10[337], stage0_10[338], stage0_10[339], stage0_10[340], stage0_10[341]},
      {stage1_12[56],stage1_11[58],stage1_10[61],stage1_9[140],stage1_8[217]}
   );
   gpc606_5 gpc378 (
      {stage0_8[360], stage0_8[361], stage0_8[362], stage0_8[363], stage0_8[364], stage0_8[365]},
      {stage0_10[342], stage0_10[343], stage0_10[344], stage0_10[345], stage0_10[346], stage0_10[347]},
      {stage1_12[57],stage1_11[59],stage1_10[62],stage1_9[141],stage1_8[218]}
   );
   gpc606_5 gpc379 (
      {stage0_8[366], stage0_8[367], stage0_8[368], stage0_8[369], stage0_8[370], stage0_8[371]},
      {stage0_10[348], stage0_10[349], stage0_10[350], stage0_10[351], stage0_10[352], stage0_10[353]},
      {stage1_12[58],stage1_11[60],stage1_10[63],stage1_9[142],stage1_8[219]}
   );
   gpc606_5 gpc380 (
      {stage0_8[372], stage0_8[373], stage0_8[374], stage0_8[375], stage0_8[376], stage0_8[377]},
      {stage0_10[354], stage0_10[355], stage0_10[356], stage0_10[357], stage0_10[358], stage0_10[359]},
      {stage1_12[59],stage1_11[61],stage1_10[64],stage1_9[143],stage1_8[220]}
   );
   gpc606_5 gpc381 (
      {stage0_8[378], stage0_8[379], stage0_8[380], stage0_8[381], stage0_8[382], stage0_8[383]},
      {stage0_10[360], stage0_10[361], stage0_10[362], stage0_10[363], stage0_10[364], stage0_10[365]},
      {stage1_12[60],stage1_11[62],stage1_10[65],stage1_9[144],stage1_8[221]}
   );
   gpc606_5 gpc382 (
      {stage0_8[384], stage0_8[385], stage0_8[386], stage0_8[387], stage0_8[388], stage0_8[389]},
      {stage0_10[366], stage0_10[367], stage0_10[368], stage0_10[369], stage0_10[370], stage0_10[371]},
      {stage1_12[61],stage1_11[63],stage1_10[66],stage1_9[145],stage1_8[222]}
   );
   gpc606_5 gpc383 (
      {stage0_8[390], stage0_8[391], stage0_8[392], stage0_8[393], stage0_8[394], stage0_8[395]},
      {stage0_10[372], stage0_10[373], stage0_10[374], stage0_10[375], stage0_10[376], stage0_10[377]},
      {stage1_12[62],stage1_11[64],stage1_10[67],stage1_9[146],stage1_8[223]}
   );
   gpc606_5 gpc384 (
      {stage0_8[396], stage0_8[397], stage0_8[398], stage0_8[399], stage0_8[400], stage0_8[401]},
      {stage0_10[378], stage0_10[379], stage0_10[380], stage0_10[381], stage0_10[382], stage0_10[383]},
      {stage1_12[63],stage1_11[65],stage1_10[68],stage1_9[147],stage1_8[224]}
   );
   gpc606_5 gpc385 (
      {stage0_8[402], stage0_8[403], stage0_8[404], stage0_8[405], stage0_8[406], stage0_8[407]},
      {stage0_10[384], stage0_10[385], stage0_10[386], stage0_10[387], stage0_10[388], stage0_10[389]},
      {stage1_12[64],stage1_11[66],stage1_10[69],stage1_9[148],stage1_8[225]}
   );
   gpc606_5 gpc386 (
      {stage0_8[408], stage0_8[409], stage0_8[410], stage0_8[411], stage0_8[412], stage0_8[413]},
      {stage0_10[390], stage0_10[391], stage0_10[392], stage0_10[393], stage0_10[394], stage0_10[395]},
      {stage1_12[65],stage1_11[67],stage1_10[70],stage1_9[149],stage1_8[226]}
   );
   gpc606_5 gpc387 (
      {stage0_8[414], stage0_8[415], stage0_8[416], stage0_8[417], stage0_8[418], stage0_8[419]},
      {stage0_10[396], stage0_10[397], stage0_10[398], stage0_10[399], stage0_10[400], stage0_10[401]},
      {stage1_12[66],stage1_11[68],stage1_10[71],stage1_9[150],stage1_8[227]}
   );
   gpc606_5 gpc388 (
      {stage0_8[420], stage0_8[421], stage0_8[422], stage0_8[423], stage0_8[424], stage0_8[425]},
      {stage0_10[402], stage0_10[403], stage0_10[404], stage0_10[405], stage0_10[406], stage0_10[407]},
      {stage1_12[67],stage1_11[69],stage1_10[72],stage1_9[151],stage1_8[228]}
   );
   gpc606_5 gpc389 (
      {stage0_8[426], stage0_8[427], stage0_8[428], stage0_8[429], stage0_8[430], stage0_8[431]},
      {stage0_10[408], stage0_10[409], stage0_10[410], stage0_10[411], stage0_10[412], stage0_10[413]},
      {stage1_12[68],stage1_11[70],stage1_10[73],stage1_9[152],stage1_8[229]}
   );
   gpc606_5 gpc390 (
      {stage0_8[432], stage0_8[433], stage0_8[434], stage0_8[435], stage0_8[436], stage0_8[437]},
      {stage0_10[414], stage0_10[415], stage0_10[416], stage0_10[417], stage0_10[418], stage0_10[419]},
      {stage1_12[69],stage1_11[71],stage1_10[74],stage1_9[153],stage1_8[230]}
   );
   gpc606_5 gpc391 (
      {stage0_8[438], stage0_8[439], stage0_8[440], stage0_8[441], stage0_8[442], stage0_8[443]},
      {stage0_10[420], stage0_10[421], stage0_10[422], stage0_10[423], stage0_10[424], stage0_10[425]},
      {stage1_12[70],stage1_11[72],stage1_10[75],stage1_9[154],stage1_8[231]}
   );
   gpc606_5 gpc392 (
      {stage0_8[444], stage0_8[445], stage0_8[446], stage0_8[447], stage0_8[448], stage0_8[449]},
      {stage0_10[426], stage0_10[427], stage0_10[428], stage0_10[429], stage0_10[430], stage0_10[431]},
      {stage1_12[71],stage1_11[73],stage1_10[76],stage1_9[155],stage1_8[232]}
   );
   gpc606_5 gpc393 (
      {stage0_8[450], stage0_8[451], stage0_8[452], stage0_8[453], stage0_8[454], stage0_8[455]},
      {stage0_10[432], stage0_10[433], stage0_10[434], stage0_10[435], stage0_10[436], stage0_10[437]},
      {stage1_12[72],stage1_11[74],stage1_10[77],stage1_9[156],stage1_8[233]}
   );
   gpc606_5 gpc394 (
      {stage0_8[456], stage0_8[457], stage0_8[458], stage0_8[459], stage0_8[460], stage0_8[461]},
      {stage0_10[438], stage0_10[439], stage0_10[440], stage0_10[441], stage0_10[442], stage0_10[443]},
      {stage1_12[73],stage1_11[75],stage1_10[78],stage1_9[157],stage1_8[234]}
   );
   gpc606_5 gpc395 (
      {stage0_8[462], stage0_8[463], stage0_8[464], stage0_8[465], stage0_8[466], stage0_8[467]},
      {stage0_10[444], stage0_10[445], stage0_10[446], stage0_10[447], stage0_10[448], stage0_10[449]},
      {stage1_12[74],stage1_11[76],stage1_10[79],stage1_9[158],stage1_8[235]}
   );
   gpc606_5 gpc396 (
      {stage0_8[468], stage0_8[469], stage0_8[470], stage0_8[471], stage0_8[472], stage0_8[473]},
      {stage0_10[450], stage0_10[451], stage0_10[452], stage0_10[453], stage0_10[454], stage0_10[455]},
      {stage1_12[75],stage1_11[77],stage1_10[80],stage1_9[159],stage1_8[236]}
   );
   gpc606_5 gpc397 (
      {stage0_8[474], stage0_8[475], stage0_8[476], stage0_8[477], stage0_8[478], stage0_8[479]},
      {stage0_10[456], stage0_10[457], stage0_10[458], stage0_10[459], stage0_10[460], stage0_10[461]},
      {stage1_12[76],stage1_11[78],stage1_10[81],stage1_9[160],stage1_8[237]}
   );
   gpc606_5 gpc398 (
      {stage0_8[480], stage0_8[481], stage0_8[482], stage0_8[483], stage0_8[484], stage0_8[485]},
      {stage0_10[462], stage0_10[463], stage0_10[464], stage0_10[465], stage0_10[466], stage0_10[467]},
      {stage1_12[77],stage1_11[79],stage1_10[82],stage1_9[161],stage1_8[238]}
   );
   gpc606_5 gpc399 (
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[78],stage1_11[80],stage1_10[83],stage1_9[162]}
   );
   gpc606_5 gpc400 (
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[79],stage1_11[81],stage1_10[84],stage1_9[163]}
   );
   gpc606_5 gpc401 (
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[80],stage1_11[82],stage1_10[85],stage1_9[164]}
   );
   gpc606_5 gpc402 (
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[81],stage1_11[83],stage1_10[86],stage1_9[165]}
   );
   gpc606_5 gpc403 (
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[82],stage1_11[84],stage1_10[87],stage1_9[166]}
   );
   gpc606_5 gpc404 (
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[83],stage1_11[85],stage1_10[88],stage1_9[167]}
   );
   gpc606_5 gpc405 (
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[84],stage1_11[86],stage1_10[89],stage1_9[168]}
   );
   gpc606_5 gpc406 (
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[85],stage1_11[87],stage1_10[90],stage1_9[169]}
   );
   gpc606_5 gpc407 (
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[86],stage1_11[88],stage1_10[91],stage1_9[170]}
   );
   gpc606_5 gpc408 (
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[87],stage1_11[89],stage1_10[92],stage1_9[171]}
   );
   gpc606_5 gpc409 (
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[88],stage1_11[90],stage1_10[93],stage1_9[172]}
   );
   gpc606_5 gpc410 (
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[89],stage1_11[91],stage1_10[94],stage1_9[173]}
   );
   gpc606_5 gpc411 (
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[90],stage1_11[92],stage1_10[95],stage1_9[174]}
   );
   gpc606_5 gpc412 (
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[91],stage1_11[93],stage1_10[96],stage1_9[175]}
   );
   gpc606_5 gpc413 (
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[92],stage1_11[94],stage1_10[97],stage1_9[176]}
   );
   gpc606_5 gpc414 (
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[93],stage1_11[95],stage1_10[98],stage1_9[177]}
   );
   gpc606_5 gpc415 (
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[94],stage1_11[96],stage1_10[99],stage1_9[178]}
   );
   gpc606_5 gpc416 (
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[95],stage1_11[97],stage1_10[100],stage1_9[179]}
   );
   gpc606_5 gpc417 (
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[96],stage1_11[98],stage1_10[101],stage1_9[180]}
   );
   gpc606_5 gpc418 (
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[97],stage1_11[99],stage1_10[102],stage1_9[181]}
   );
   gpc606_5 gpc419 (
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[98],stage1_11[100],stage1_10[103],stage1_9[182]}
   );
   gpc606_5 gpc420 (
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[99],stage1_11[101],stage1_10[104],stage1_9[183]}
   );
   gpc606_5 gpc421 (
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[100],stage1_11[102],stage1_10[105],stage1_9[184]}
   );
   gpc606_5 gpc422 (
      {stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage1_13[23],stage1_12[101],stage1_11[103],stage1_10[106],stage1_9[185]}
   );
   gpc606_5 gpc423 (
      {stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160], stage0_9[161]},
      {stage0_11[144], stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage1_13[24],stage1_12[102],stage1_11[104],stage1_10[107],stage1_9[186]}
   );
   gpc606_5 gpc424 (
      {stage0_9[162], stage0_9[163], stage0_9[164], stage0_9[165], stage0_9[166], stage0_9[167]},
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154], stage0_11[155]},
      {stage1_13[25],stage1_12[103],stage1_11[105],stage1_10[108],stage1_9[187]}
   );
   gpc606_5 gpc425 (
      {stage0_9[168], stage0_9[169], stage0_9[170], stage0_9[171], stage0_9[172], stage0_9[173]},
      {stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159], stage0_11[160], stage0_11[161]},
      {stage1_13[26],stage1_12[104],stage1_11[106],stage1_10[109],stage1_9[188]}
   );
   gpc606_5 gpc426 (
      {stage0_9[174], stage0_9[175], stage0_9[176], stage0_9[177], stage0_9[178], stage0_9[179]},
      {stage0_11[162], stage0_11[163], stage0_11[164], stage0_11[165], stage0_11[166], stage0_11[167]},
      {stage1_13[27],stage1_12[105],stage1_11[107],stage1_10[110],stage1_9[189]}
   );
   gpc606_5 gpc427 (
      {stage0_9[180], stage0_9[181], stage0_9[182], stage0_9[183], stage0_9[184], stage0_9[185]},
      {stage0_11[168], stage0_11[169], stage0_11[170], stage0_11[171], stage0_11[172], stage0_11[173]},
      {stage1_13[28],stage1_12[106],stage1_11[108],stage1_10[111],stage1_9[190]}
   );
   gpc606_5 gpc428 (
      {stage0_9[186], stage0_9[187], stage0_9[188], stage0_9[189], stage0_9[190], stage0_9[191]},
      {stage0_11[174], stage0_11[175], stage0_11[176], stage0_11[177], stage0_11[178], stage0_11[179]},
      {stage1_13[29],stage1_12[107],stage1_11[109],stage1_10[112],stage1_9[191]}
   );
   gpc606_5 gpc429 (
      {stage0_9[192], stage0_9[193], stage0_9[194], stage0_9[195], stage0_9[196], stage0_9[197]},
      {stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183], stage0_11[184], stage0_11[185]},
      {stage1_13[30],stage1_12[108],stage1_11[110],stage1_10[113],stage1_9[192]}
   );
   gpc606_5 gpc430 (
      {stage0_9[198], stage0_9[199], stage0_9[200], stage0_9[201], stage0_9[202], stage0_9[203]},
      {stage0_11[186], stage0_11[187], stage0_11[188], stage0_11[189], stage0_11[190], stage0_11[191]},
      {stage1_13[31],stage1_12[109],stage1_11[111],stage1_10[114],stage1_9[193]}
   );
   gpc606_5 gpc431 (
      {stage0_9[204], stage0_9[205], stage0_9[206], stage0_9[207], stage0_9[208], stage0_9[209]},
      {stage0_11[192], stage0_11[193], stage0_11[194], stage0_11[195], stage0_11[196], stage0_11[197]},
      {stage1_13[32],stage1_12[110],stage1_11[112],stage1_10[115],stage1_9[194]}
   );
   gpc606_5 gpc432 (
      {stage0_9[210], stage0_9[211], stage0_9[212], stage0_9[213], stage0_9[214], stage0_9[215]},
      {stage0_11[198], stage0_11[199], stage0_11[200], stage0_11[201], stage0_11[202], stage0_11[203]},
      {stage1_13[33],stage1_12[111],stage1_11[113],stage1_10[116],stage1_9[195]}
   );
   gpc606_5 gpc433 (
      {stage0_9[216], stage0_9[217], stage0_9[218], stage0_9[219], stage0_9[220], stage0_9[221]},
      {stage0_11[204], stage0_11[205], stage0_11[206], stage0_11[207], stage0_11[208], stage0_11[209]},
      {stage1_13[34],stage1_12[112],stage1_11[114],stage1_10[117],stage1_9[196]}
   );
   gpc606_5 gpc434 (
      {stage0_9[222], stage0_9[223], stage0_9[224], stage0_9[225], stage0_9[226], stage0_9[227]},
      {stage0_11[210], stage0_11[211], stage0_11[212], stage0_11[213], stage0_11[214], stage0_11[215]},
      {stage1_13[35],stage1_12[113],stage1_11[115],stage1_10[118],stage1_9[197]}
   );
   gpc606_5 gpc435 (
      {stage0_9[228], stage0_9[229], stage0_9[230], stage0_9[231], stage0_9[232], stage0_9[233]},
      {stage0_11[216], stage0_11[217], stage0_11[218], stage0_11[219], stage0_11[220], stage0_11[221]},
      {stage1_13[36],stage1_12[114],stage1_11[116],stage1_10[119],stage1_9[198]}
   );
   gpc606_5 gpc436 (
      {stage0_9[234], stage0_9[235], stage0_9[236], stage0_9[237], stage0_9[238], stage0_9[239]},
      {stage0_11[222], stage0_11[223], stage0_11[224], stage0_11[225], stage0_11[226], stage0_11[227]},
      {stage1_13[37],stage1_12[115],stage1_11[117],stage1_10[120],stage1_9[199]}
   );
   gpc606_5 gpc437 (
      {stage0_9[240], stage0_9[241], stage0_9[242], stage0_9[243], stage0_9[244], stage0_9[245]},
      {stage0_11[228], stage0_11[229], stage0_11[230], stage0_11[231], stage0_11[232], stage0_11[233]},
      {stage1_13[38],stage1_12[116],stage1_11[118],stage1_10[121],stage1_9[200]}
   );
   gpc606_5 gpc438 (
      {stage0_9[246], stage0_9[247], stage0_9[248], stage0_9[249], stage0_9[250], stage0_9[251]},
      {stage0_11[234], stage0_11[235], stage0_11[236], stage0_11[237], stage0_11[238], stage0_11[239]},
      {stage1_13[39],stage1_12[117],stage1_11[119],stage1_10[122],stage1_9[201]}
   );
   gpc606_5 gpc439 (
      {stage0_9[252], stage0_9[253], stage0_9[254], stage0_9[255], stage0_9[256], stage0_9[257]},
      {stage0_11[240], stage0_11[241], stage0_11[242], stage0_11[243], stage0_11[244], stage0_11[245]},
      {stage1_13[40],stage1_12[118],stage1_11[120],stage1_10[123],stage1_9[202]}
   );
   gpc606_5 gpc440 (
      {stage0_9[258], stage0_9[259], stage0_9[260], stage0_9[261], stage0_9[262], stage0_9[263]},
      {stage0_11[246], stage0_11[247], stage0_11[248], stage0_11[249], stage0_11[250], stage0_11[251]},
      {stage1_13[41],stage1_12[119],stage1_11[121],stage1_10[124],stage1_9[203]}
   );
   gpc606_5 gpc441 (
      {stage0_9[264], stage0_9[265], stage0_9[266], stage0_9[267], stage0_9[268], stage0_9[269]},
      {stage0_11[252], stage0_11[253], stage0_11[254], stage0_11[255], stage0_11[256], stage0_11[257]},
      {stage1_13[42],stage1_12[120],stage1_11[122],stage1_10[125],stage1_9[204]}
   );
   gpc606_5 gpc442 (
      {stage0_9[270], stage0_9[271], stage0_9[272], stage0_9[273], stage0_9[274], stage0_9[275]},
      {stage0_11[258], stage0_11[259], stage0_11[260], stage0_11[261], stage0_11[262], stage0_11[263]},
      {stage1_13[43],stage1_12[121],stage1_11[123],stage1_10[126],stage1_9[205]}
   );
   gpc606_5 gpc443 (
      {stage0_9[276], stage0_9[277], stage0_9[278], stage0_9[279], stage0_9[280], stage0_9[281]},
      {stage0_11[264], stage0_11[265], stage0_11[266], stage0_11[267], stage0_11[268], stage0_11[269]},
      {stage1_13[44],stage1_12[122],stage1_11[124],stage1_10[127],stage1_9[206]}
   );
   gpc606_5 gpc444 (
      {stage0_9[282], stage0_9[283], stage0_9[284], stage0_9[285], stage0_9[286], stage0_9[287]},
      {stage0_11[270], stage0_11[271], stage0_11[272], stage0_11[273], stage0_11[274], stage0_11[275]},
      {stage1_13[45],stage1_12[123],stage1_11[125],stage1_10[128],stage1_9[207]}
   );
   gpc606_5 gpc445 (
      {stage0_9[288], stage0_9[289], stage0_9[290], stage0_9[291], stage0_9[292], stage0_9[293]},
      {stage0_11[276], stage0_11[277], stage0_11[278], stage0_11[279], stage0_11[280], stage0_11[281]},
      {stage1_13[46],stage1_12[124],stage1_11[126],stage1_10[129],stage1_9[208]}
   );
   gpc606_5 gpc446 (
      {stage0_9[294], stage0_9[295], stage0_9[296], stage0_9[297], stage0_9[298], stage0_9[299]},
      {stage0_11[282], stage0_11[283], stage0_11[284], stage0_11[285], stage0_11[286], stage0_11[287]},
      {stage1_13[47],stage1_12[125],stage1_11[127],stage1_10[130],stage1_9[209]}
   );
   gpc606_5 gpc447 (
      {stage0_9[300], stage0_9[301], stage0_9[302], stage0_9[303], stage0_9[304], stage0_9[305]},
      {stage0_11[288], stage0_11[289], stage0_11[290], stage0_11[291], stage0_11[292], stage0_11[293]},
      {stage1_13[48],stage1_12[126],stage1_11[128],stage1_10[131],stage1_9[210]}
   );
   gpc606_5 gpc448 (
      {stage0_9[306], stage0_9[307], stage0_9[308], stage0_9[309], stage0_9[310], stage0_9[311]},
      {stage0_11[294], stage0_11[295], stage0_11[296], stage0_11[297], stage0_11[298], stage0_11[299]},
      {stage1_13[49],stage1_12[127],stage1_11[129],stage1_10[132],stage1_9[211]}
   );
   gpc606_5 gpc449 (
      {stage0_9[312], stage0_9[313], stage0_9[314], stage0_9[315], stage0_9[316], stage0_9[317]},
      {stage0_11[300], stage0_11[301], stage0_11[302], stage0_11[303], stage0_11[304], stage0_11[305]},
      {stage1_13[50],stage1_12[128],stage1_11[130],stage1_10[133],stage1_9[212]}
   );
   gpc606_5 gpc450 (
      {stage0_9[318], stage0_9[319], stage0_9[320], stage0_9[321], stage0_9[322], stage0_9[323]},
      {stage0_11[306], stage0_11[307], stage0_11[308], stage0_11[309], stage0_11[310], stage0_11[311]},
      {stage1_13[51],stage1_12[129],stage1_11[131],stage1_10[134],stage1_9[213]}
   );
   gpc606_5 gpc451 (
      {stage0_9[324], stage0_9[325], stage0_9[326], stage0_9[327], stage0_9[328], stage0_9[329]},
      {stage0_11[312], stage0_11[313], stage0_11[314], stage0_11[315], stage0_11[316], stage0_11[317]},
      {stage1_13[52],stage1_12[130],stage1_11[132],stage1_10[135],stage1_9[214]}
   );
   gpc606_5 gpc452 (
      {stage0_9[330], stage0_9[331], stage0_9[332], stage0_9[333], stage0_9[334], stage0_9[335]},
      {stage0_11[318], stage0_11[319], stage0_11[320], stage0_11[321], stage0_11[322], stage0_11[323]},
      {stage1_13[53],stage1_12[131],stage1_11[133],stage1_10[136],stage1_9[215]}
   );
   gpc606_5 gpc453 (
      {stage0_9[336], stage0_9[337], stage0_9[338], stage0_9[339], stage0_9[340], stage0_9[341]},
      {stage0_11[324], stage0_11[325], stage0_11[326], stage0_11[327], stage0_11[328], stage0_11[329]},
      {stage1_13[54],stage1_12[132],stage1_11[134],stage1_10[137],stage1_9[216]}
   );
   gpc606_5 gpc454 (
      {stage0_9[342], stage0_9[343], stage0_9[344], stage0_9[345], stage0_9[346], stage0_9[347]},
      {stage0_11[330], stage0_11[331], stage0_11[332], stage0_11[333], stage0_11[334], stage0_11[335]},
      {stage1_13[55],stage1_12[133],stage1_11[135],stage1_10[138],stage1_9[217]}
   );
   gpc606_5 gpc455 (
      {stage0_9[348], stage0_9[349], stage0_9[350], stage0_9[351], stage0_9[352], stage0_9[353]},
      {stage0_11[336], stage0_11[337], stage0_11[338], stage0_11[339], stage0_11[340], stage0_11[341]},
      {stage1_13[56],stage1_12[134],stage1_11[136],stage1_10[139],stage1_9[218]}
   );
   gpc606_5 gpc456 (
      {stage0_9[354], stage0_9[355], stage0_9[356], stage0_9[357], stage0_9[358], stage0_9[359]},
      {stage0_11[342], stage0_11[343], stage0_11[344], stage0_11[345], stage0_11[346], stage0_11[347]},
      {stage1_13[57],stage1_12[135],stage1_11[137],stage1_10[140],stage1_9[219]}
   );
   gpc606_5 gpc457 (
      {stage0_9[360], stage0_9[361], stage0_9[362], stage0_9[363], stage0_9[364], stage0_9[365]},
      {stage0_11[348], stage0_11[349], stage0_11[350], stage0_11[351], stage0_11[352], stage0_11[353]},
      {stage1_13[58],stage1_12[136],stage1_11[138],stage1_10[141],stage1_9[220]}
   );
   gpc606_5 gpc458 (
      {stage0_9[366], stage0_9[367], stage0_9[368], stage0_9[369], stage0_9[370], stage0_9[371]},
      {stage0_11[354], stage0_11[355], stage0_11[356], stage0_11[357], stage0_11[358], stage0_11[359]},
      {stage1_13[59],stage1_12[137],stage1_11[139],stage1_10[142],stage1_9[221]}
   );
   gpc606_5 gpc459 (
      {stage0_9[372], stage0_9[373], stage0_9[374], stage0_9[375], stage0_9[376], stage0_9[377]},
      {stage0_11[360], stage0_11[361], stage0_11[362], stage0_11[363], stage0_11[364], stage0_11[365]},
      {stage1_13[60],stage1_12[138],stage1_11[140],stage1_10[143],stage1_9[222]}
   );
   gpc606_5 gpc460 (
      {stage0_9[378], stage0_9[379], stage0_9[380], stage0_9[381], stage0_9[382], stage0_9[383]},
      {stage0_11[366], stage0_11[367], stage0_11[368], stage0_11[369], stage0_11[370], stage0_11[371]},
      {stage1_13[61],stage1_12[139],stage1_11[141],stage1_10[144],stage1_9[223]}
   );
   gpc606_5 gpc461 (
      {stage0_9[384], stage0_9[385], stage0_9[386], stage0_9[387], stage0_9[388], stage0_9[389]},
      {stage0_11[372], stage0_11[373], stage0_11[374], stage0_11[375], stage0_11[376], stage0_11[377]},
      {stage1_13[62],stage1_12[140],stage1_11[142],stage1_10[145],stage1_9[224]}
   );
   gpc606_5 gpc462 (
      {stage0_9[390], stage0_9[391], stage0_9[392], stage0_9[393], stage0_9[394], stage0_9[395]},
      {stage0_11[378], stage0_11[379], stage0_11[380], stage0_11[381], stage0_11[382], stage0_11[383]},
      {stage1_13[63],stage1_12[141],stage1_11[143],stage1_10[146],stage1_9[225]}
   );
   gpc606_5 gpc463 (
      {stage0_9[396], stage0_9[397], stage0_9[398], stage0_9[399], stage0_9[400], stage0_9[401]},
      {stage0_11[384], stage0_11[385], stage0_11[386], stage0_11[387], stage0_11[388], stage0_11[389]},
      {stage1_13[64],stage1_12[142],stage1_11[144],stage1_10[147],stage1_9[226]}
   );
   gpc606_5 gpc464 (
      {stage0_9[402], stage0_9[403], stage0_9[404], stage0_9[405], stage0_9[406], stage0_9[407]},
      {stage0_11[390], stage0_11[391], stage0_11[392], stage0_11[393], stage0_11[394], stage0_11[395]},
      {stage1_13[65],stage1_12[143],stage1_11[145],stage1_10[148],stage1_9[227]}
   );
   gpc606_5 gpc465 (
      {stage0_9[408], stage0_9[409], stage0_9[410], stage0_9[411], stage0_9[412], stage0_9[413]},
      {stage0_11[396], stage0_11[397], stage0_11[398], stage0_11[399], stage0_11[400], stage0_11[401]},
      {stage1_13[66],stage1_12[144],stage1_11[146],stage1_10[149],stage1_9[228]}
   );
   gpc606_5 gpc466 (
      {stage0_9[414], stage0_9[415], stage0_9[416], stage0_9[417], stage0_9[418], stage0_9[419]},
      {stage0_11[402], stage0_11[403], stage0_11[404], stage0_11[405], stage0_11[406], stage0_11[407]},
      {stage1_13[67],stage1_12[145],stage1_11[147],stage1_10[150],stage1_9[229]}
   );
   gpc606_5 gpc467 (
      {stage0_9[420], stage0_9[421], stage0_9[422], stage0_9[423], stage0_9[424], stage0_9[425]},
      {stage0_11[408], stage0_11[409], stage0_11[410], stage0_11[411], stage0_11[412], stage0_11[413]},
      {stage1_13[68],stage1_12[146],stage1_11[148],stage1_10[151],stage1_9[230]}
   );
   gpc606_5 gpc468 (
      {stage0_9[426], stage0_9[427], stage0_9[428], stage0_9[429], stage0_9[430], stage0_9[431]},
      {stage0_11[414], stage0_11[415], stage0_11[416], stage0_11[417], stage0_11[418], stage0_11[419]},
      {stage1_13[69],stage1_12[147],stage1_11[149],stage1_10[152],stage1_9[231]}
   );
   gpc606_5 gpc469 (
      {stage0_9[432], stage0_9[433], stage0_9[434], stage0_9[435], stage0_9[436], stage0_9[437]},
      {stage0_11[420], stage0_11[421], stage0_11[422], stage0_11[423], stage0_11[424], stage0_11[425]},
      {stage1_13[70],stage1_12[148],stage1_11[150],stage1_10[153],stage1_9[232]}
   );
   gpc606_5 gpc470 (
      {stage0_9[438], stage0_9[439], stage0_9[440], stage0_9[441], stage0_9[442], stage0_9[443]},
      {stage0_11[426], stage0_11[427], stage0_11[428], stage0_11[429], stage0_11[430], stage0_11[431]},
      {stage1_13[71],stage1_12[149],stage1_11[151],stage1_10[154],stage1_9[233]}
   );
   gpc606_5 gpc471 (
      {stage0_9[444], stage0_9[445], stage0_9[446], stage0_9[447], stage0_9[448], stage0_9[449]},
      {stage0_11[432], stage0_11[433], stage0_11[434], stage0_11[435], stage0_11[436], stage0_11[437]},
      {stage1_13[72],stage1_12[150],stage1_11[152],stage1_10[155],stage1_9[234]}
   );
   gpc606_5 gpc472 (
      {stage0_9[450], stage0_9[451], stage0_9[452], stage0_9[453], stage0_9[454], stage0_9[455]},
      {stage0_11[438], stage0_11[439], stage0_11[440], stage0_11[441], stage0_11[442], stage0_11[443]},
      {stage1_13[73],stage1_12[151],stage1_11[153],stage1_10[156],stage1_9[235]}
   );
   gpc606_5 gpc473 (
      {stage0_9[456], stage0_9[457], stage0_9[458], stage0_9[459], stage0_9[460], stage0_9[461]},
      {stage0_11[444], stage0_11[445], stage0_11[446], stage0_11[447], stage0_11[448], stage0_11[449]},
      {stage1_13[74],stage1_12[152],stage1_11[154],stage1_10[157],stage1_9[236]}
   );
   gpc606_5 gpc474 (
      {stage0_9[462], stage0_9[463], stage0_9[464], stage0_9[465], stage0_9[466], stage0_9[467]},
      {stage0_11[450], stage0_11[451], stage0_11[452], stage0_11[453], stage0_11[454], stage0_11[455]},
      {stage1_13[75],stage1_12[153],stage1_11[155],stage1_10[158],stage1_9[237]}
   );
   gpc606_5 gpc475 (
      {stage0_9[468], stage0_9[469], stage0_9[470], stage0_9[471], stage0_9[472], stage0_9[473]},
      {stage0_11[456], stage0_11[457], stage0_11[458], stage0_11[459], stage0_11[460], stage0_11[461]},
      {stage1_13[76],stage1_12[154],stage1_11[156],stage1_10[159],stage1_9[238]}
   );
   gpc606_5 gpc476 (
      {stage0_9[474], stage0_9[475], stage0_9[476], stage0_9[477], stage0_9[478], stage0_9[479]},
      {stage0_11[462], stage0_11[463], stage0_11[464], stage0_11[465], stage0_11[466], stage0_11[467]},
      {stage1_13[77],stage1_12[155],stage1_11[157],stage1_10[160],stage1_9[239]}
   );
   gpc606_5 gpc477 (
      {stage0_9[480], stage0_9[481], stage0_9[482], stage0_9[483], stage0_9[484], stage0_9[485]},
      {stage0_11[468], stage0_11[469], stage0_11[470], stage0_11[471], stage0_11[472], stage0_11[473]},
      {stage1_13[78],stage1_12[156],stage1_11[158],stage1_10[161],stage1_9[240]}
   );
   gpc1_1 gpc478 (
      {stage0_2[447]},
      {stage1_2[159]}
   );
   gpc1_1 gpc479 (
      {stage0_2[448]},
      {stage1_2[160]}
   );
   gpc1_1 gpc480 (
      {stage0_2[449]},
      {stage1_2[161]}
   );
   gpc1_1 gpc481 (
      {stage0_2[450]},
      {stage1_2[162]}
   );
   gpc1_1 gpc482 (
      {stage0_2[451]},
      {stage1_2[163]}
   );
   gpc1_1 gpc483 (
      {stage0_2[452]},
      {stage1_2[164]}
   );
   gpc1_1 gpc484 (
      {stage0_2[453]},
      {stage1_2[165]}
   );
   gpc1_1 gpc485 (
      {stage0_2[454]},
      {stage1_2[166]}
   );
   gpc1_1 gpc486 (
      {stage0_2[455]},
      {stage1_2[167]}
   );
   gpc1_1 gpc487 (
      {stage0_2[456]},
      {stage1_2[168]}
   );
   gpc1_1 gpc488 (
      {stage0_2[457]},
      {stage1_2[169]}
   );
   gpc1_1 gpc489 (
      {stage0_2[458]},
      {stage1_2[170]}
   );
   gpc1_1 gpc490 (
      {stage0_2[459]},
      {stage1_2[171]}
   );
   gpc1_1 gpc491 (
      {stage0_2[460]},
      {stage1_2[172]}
   );
   gpc1_1 gpc492 (
      {stage0_2[461]},
      {stage1_2[173]}
   );
   gpc1_1 gpc493 (
      {stage0_2[462]},
      {stage1_2[174]}
   );
   gpc1_1 gpc494 (
      {stage0_2[463]},
      {stage1_2[175]}
   );
   gpc1_1 gpc495 (
      {stage0_2[464]},
      {stage1_2[176]}
   );
   gpc1_1 gpc496 (
      {stage0_2[465]},
      {stage1_2[177]}
   );
   gpc1_1 gpc497 (
      {stage0_2[466]},
      {stage1_2[178]}
   );
   gpc1_1 gpc498 (
      {stage0_2[467]},
      {stage1_2[179]}
   );
   gpc1_1 gpc499 (
      {stage0_2[468]},
      {stage1_2[180]}
   );
   gpc1_1 gpc500 (
      {stage0_2[469]},
      {stage1_2[181]}
   );
   gpc1_1 gpc501 (
      {stage0_2[470]},
      {stage1_2[182]}
   );
   gpc1_1 gpc502 (
      {stage0_2[471]},
      {stage1_2[183]}
   );
   gpc1_1 gpc503 (
      {stage0_2[472]},
      {stage1_2[184]}
   );
   gpc1_1 gpc504 (
      {stage0_2[473]},
      {stage1_2[185]}
   );
   gpc1_1 gpc505 (
      {stage0_2[474]},
      {stage1_2[186]}
   );
   gpc1_1 gpc506 (
      {stage0_2[475]},
      {stage1_2[187]}
   );
   gpc1_1 gpc507 (
      {stage0_2[476]},
      {stage1_2[188]}
   );
   gpc1_1 gpc508 (
      {stage0_2[477]},
      {stage1_2[189]}
   );
   gpc1_1 gpc509 (
      {stage0_2[478]},
      {stage1_2[190]}
   );
   gpc1_1 gpc510 (
      {stage0_2[479]},
      {stage1_2[191]}
   );
   gpc1_1 gpc511 (
      {stage0_2[480]},
      {stage1_2[192]}
   );
   gpc1_1 gpc512 (
      {stage0_2[481]},
      {stage1_2[193]}
   );
   gpc1_1 gpc513 (
      {stage0_2[482]},
      {stage1_2[194]}
   );
   gpc1_1 gpc514 (
      {stage0_2[483]},
      {stage1_2[195]}
   );
   gpc1_1 gpc515 (
      {stage0_2[484]},
      {stage1_2[196]}
   );
   gpc1_1 gpc516 (
      {stage0_2[485]},
      {stage1_2[197]}
   );
   gpc1_1 gpc517 (
      {stage0_3[450]},
      {stage1_3[160]}
   );
   gpc1_1 gpc518 (
      {stage0_3[451]},
      {stage1_3[161]}
   );
   gpc1_1 gpc519 (
      {stage0_3[452]},
      {stage1_3[162]}
   );
   gpc1_1 gpc520 (
      {stage0_3[453]},
      {stage1_3[163]}
   );
   gpc1_1 gpc521 (
      {stage0_3[454]},
      {stage1_3[164]}
   );
   gpc1_1 gpc522 (
      {stage0_3[455]},
      {stage1_3[165]}
   );
   gpc1_1 gpc523 (
      {stage0_3[456]},
      {stage1_3[166]}
   );
   gpc1_1 gpc524 (
      {stage0_3[457]},
      {stage1_3[167]}
   );
   gpc1_1 gpc525 (
      {stage0_3[458]},
      {stage1_3[168]}
   );
   gpc1_1 gpc526 (
      {stage0_3[459]},
      {stage1_3[169]}
   );
   gpc1_1 gpc527 (
      {stage0_3[460]},
      {stage1_3[170]}
   );
   gpc1_1 gpc528 (
      {stage0_3[461]},
      {stage1_3[171]}
   );
   gpc1_1 gpc529 (
      {stage0_3[462]},
      {stage1_3[172]}
   );
   gpc1_1 gpc530 (
      {stage0_3[463]},
      {stage1_3[173]}
   );
   gpc1_1 gpc531 (
      {stage0_3[464]},
      {stage1_3[174]}
   );
   gpc1_1 gpc532 (
      {stage0_3[465]},
      {stage1_3[175]}
   );
   gpc1_1 gpc533 (
      {stage0_3[466]},
      {stage1_3[176]}
   );
   gpc1_1 gpc534 (
      {stage0_3[467]},
      {stage1_3[177]}
   );
   gpc1_1 gpc535 (
      {stage0_3[468]},
      {stage1_3[178]}
   );
   gpc1_1 gpc536 (
      {stage0_3[469]},
      {stage1_3[179]}
   );
   gpc1_1 gpc537 (
      {stage0_3[470]},
      {stage1_3[180]}
   );
   gpc1_1 gpc538 (
      {stage0_3[471]},
      {stage1_3[181]}
   );
   gpc1_1 gpc539 (
      {stage0_3[472]},
      {stage1_3[182]}
   );
   gpc1_1 gpc540 (
      {stage0_3[473]},
      {stage1_3[183]}
   );
   gpc1_1 gpc541 (
      {stage0_3[474]},
      {stage1_3[184]}
   );
   gpc1_1 gpc542 (
      {stage0_3[475]},
      {stage1_3[185]}
   );
   gpc1_1 gpc543 (
      {stage0_3[476]},
      {stage1_3[186]}
   );
   gpc1_1 gpc544 (
      {stage0_3[477]},
      {stage1_3[187]}
   );
   gpc1_1 gpc545 (
      {stage0_3[478]},
      {stage1_3[188]}
   );
   gpc1_1 gpc546 (
      {stage0_3[479]},
      {stage1_3[189]}
   );
   gpc1_1 gpc547 (
      {stage0_3[480]},
      {stage1_3[190]}
   );
   gpc1_1 gpc548 (
      {stage0_3[481]},
      {stage1_3[191]}
   );
   gpc1_1 gpc549 (
      {stage0_3[482]},
      {stage1_3[192]}
   );
   gpc1_1 gpc550 (
      {stage0_3[483]},
      {stage1_3[193]}
   );
   gpc1_1 gpc551 (
      {stage0_3[484]},
      {stage1_3[194]}
   );
   gpc1_1 gpc552 (
      {stage0_3[485]},
      {stage1_3[195]}
   );
   gpc1_1 gpc553 (
      {stage0_4[481]},
      {stage1_4[236]}
   );
   gpc1_1 gpc554 (
      {stage0_4[482]},
      {stage1_4[237]}
   );
   gpc1_1 gpc555 (
      {stage0_4[483]},
      {stage1_4[238]}
   );
   gpc1_1 gpc556 (
      {stage0_4[484]},
      {stage1_4[239]}
   );
   gpc1_1 gpc557 (
      {stage0_4[485]},
      {stage1_4[240]}
   );
   gpc1_1 gpc558 (
      {stage0_6[480]},
      {stage1_6[164]}
   );
   gpc1_1 gpc559 (
      {stage0_6[481]},
      {stage1_6[165]}
   );
   gpc1_1 gpc560 (
      {stage0_6[482]},
      {stage1_6[166]}
   );
   gpc1_1 gpc561 (
      {stage0_6[483]},
      {stage1_6[167]}
   );
   gpc1_1 gpc562 (
      {stage0_6[484]},
      {stage1_6[168]}
   );
   gpc1_1 gpc563 (
      {stage0_6[485]},
      {stage1_6[169]}
   );
   gpc1_1 gpc564 (
      {stage0_10[468]},
      {stage1_10[162]}
   );
   gpc1_1 gpc565 (
      {stage0_10[469]},
      {stage1_10[163]}
   );
   gpc1_1 gpc566 (
      {stage0_10[470]},
      {stage1_10[164]}
   );
   gpc1_1 gpc567 (
      {stage0_10[471]},
      {stage1_10[165]}
   );
   gpc1_1 gpc568 (
      {stage0_10[472]},
      {stage1_10[166]}
   );
   gpc1_1 gpc569 (
      {stage0_10[473]},
      {stage1_10[167]}
   );
   gpc1_1 gpc570 (
      {stage0_10[474]},
      {stage1_10[168]}
   );
   gpc1_1 gpc571 (
      {stage0_10[475]},
      {stage1_10[169]}
   );
   gpc1_1 gpc572 (
      {stage0_10[476]},
      {stage1_10[170]}
   );
   gpc1_1 gpc573 (
      {stage0_10[477]},
      {stage1_10[171]}
   );
   gpc1_1 gpc574 (
      {stage0_10[478]},
      {stage1_10[172]}
   );
   gpc1_1 gpc575 (
      {stage0_10[479]},
      {stage1_10[173]}
   );
   gpc1_1 gpc576 (
      {stage0_10[480]},
      {stage1_10[174]}
   );
   gpc1_1 gpc577 (
      {stage0_10[481]},
      {stage1_10[175]}
   );
   gpc1_1 gpc578 (
      {stage0_10[482]},
      {stage1_10[176]}
   );
   gpc1_1 gpc579 (
      {stage0_10[483]},
      {stage1_10[177]}
   );
   gpc1_1 gpc580 (
      {stage0_10[484]},
      {stage1_10[178]}
   );
   gpc1_1 gpc581 (
      {stage0_10[485]},
      {stage1_10[179]}
   );
   gpc1_1 gpc582 (
      {stage0_11[474]},
      {stage1_11[159]}
   );
   gpc1_1 gpc583 (
      {stage0_11[475]},
      {stage1_11[160]}
   );
   gpc1_1 gpc584 (
      {stage0_11[476]},
      {stage1_11[161]}
   );
   gpc1_1 gpc585 (
      {stage0_11[477]},
      {stage1_11[162]}
   );
   gpc1_1 gpc586 (
      {stage0_11[478]},
      {stage1_11[163]}
   );
   gpc1_1 gpc587 (
      {stage0_11[479]},
      {stage1_11[164]}
   );
   gpc1_1 gpc588 (
      {stage0_11[480]},
      {stage1_11[165]}
   );
   gpc1_1 gpc589 (
      {stage0_11[481]},
      {stage1_11[166]}
   );
   gpc1_1 gpc590 (
      {stage0_11[482]},
      {stage1_11[167]}
   );
   gpc1_1 gpc591 (
      {stage0_11[483]},
      {stage1_11[168]}
   );
   gpc1_1 gpc592 (
      {stage0_11[484]},
      {stage1_11[169]}
   );
   gpc1_1 gpc593 (
      {stage0_11[485]},
      {stage1_11[170]}
   );
   gpc1163_5 gpc594 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc595 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc596 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc597 (
      {stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[3]},
      {stage1_3[3]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc598 (
      {stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[4]},
      {stage1_3[4]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc1163_5 gpc599 (
      {stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_2[5]},
      {stage1_3[5]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc1163_5 gpc600 (
      {stage1_0[18], stage1_0[19], stage1_0[20]},
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_2[6]},
      {stage1_3[6]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc1163_5 gpc601 (
      {stage1_0[21], stage1_0[22], stage1_0[23]},
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_2[7]},
      {stage1_3[7]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc1163_5 gpc602 (
      {stage1_0[24], stage1_0[25], stage1_0[26]},
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_2[8]},
      {stage1_3[8]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc1163_5 gpc603 (
      {stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59]},
      {stage1_2[9]},
      {stage1_3[9]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc1163_5 gpc604 (
      {stage1_0[30], stage1_0[31], stage1_0[32]},
      {stage1_1[60], stage1_1[61], stage1_1[62], stage1_1[63], stage1_1[64], stage1_1[65]},
      {stage1_2[10]},
      {stage1_3[10]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc1163_5 gpc605 (
      {stage1_0[33], stage1_0[34], stage1_0[35]},
      {stage1_1[66], stage1_1[67], stage1_1[68], stage1_1[69], stage1_1[70], stage1_1[71]},
      {stage1_2[11]},
      {stage1_3[11]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc1163_5 gpc606 (
      {stage1_0[36], stage1_0[37], stage1_0[38]},
      {stage1_1[72], stage1_1[73], stage1_1[74], stage1_1[75], stage1_1[76], stage1_1[77]},
      {stage1_2[12]},
      {stage1_3[12]},
      {stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12],stage2_0[12]}
   );
   gpc1163_5 gpc607 (
      {stage1_0[39], stage1_0[40], stage1_0[41]},
      {stage1_1[78], stage1_1[79], stage1_1[80], stage1_1[81], stage1_1[82], stage1_1[83]},
      {stage1_2[13]},
      {stage1_3[13]},
      {stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13],stage2_0[13]}
   );
   gpc1163_5 gpc608 (
      {stage1_0[42], stage1_0[43], stage1_0[44]},
      {stage1_1[84], stage1_1[85], stage1_1[86], stage1_1[87], stage1_1[88], stage1_1[89]},
      {stage1_2[14]},
      {stage1_3[14]},
      {stage2_4[14],stage2_3[14],stage2_2[14],stage2_1[14],stage2_0[14]}
   );
   gpc1163_5 gpc609 (
      {stage1_0[45], stage1_0[46], stage1_0[47]},
      {stage1_1[90], stage1_1[91], stage1_1[92], stage1_1[93], stage1_1[94], stage1_1[95]},
      {stage1_2[15]},
      {stage1_3[15]},
      {stage2_4[15],stage2_3[15],stage2_2[15],stage2_1[15],stage2_0[15]}
   );
   gpc1163_5 gpc610 (
      {stage1_0[48], stage1_0[49], stage1_0[50]},
      {stage1_1[96], stage1_1[97], stage1_1[98], stage1_1[99], stage1_1[100], stage1_1[101]},
      {stage1_2[16]},
      {stage1_3[16]},
      {stage2_4[16],stage2_3[16],stage2_2[16],stage2_1[16],stage2_0[16]}
   );
   gpc1163_5 gpc611 (
      {stage1_0[51], stage1_0[52], stage1_0[53]},
      {stage1_1[102], stage1_1[103], stage1_1[104], stage1_1[105], stage1_1[106], stage1_1[107]},
      {stage1_2[17]},
      {stage1_3[17]},
      {stage2_4[17],stage2_3[17],stage2_2[17],stage2_1[17],stage2_0[17]}
   );
   gpc1163_5 gpc612 (
      {stage1_0[54], stage1_0[55], stage1_0[56]},
      {stage1_1[108], stage1_1[109], stage1_1[110], stage1_1[111], stage1_1[112], stage1_1[113]},
      {stage1_2[18]},
      {stage1_3[18]},
      {stage2_4[18],stage2_3[18],stage2_2[18],stage2_1[18],stage2_0[18]}
   );
   gpc1163_5 gpc613 (
      {stage1_0[57], stage1_0[58], stage1_0[59]},
      {stage1_1[114], stage1_1[115], stage1_1[116], stage1_1[117], stage1_1[118], stage1_1[119]},
      {stage1_2[19]},
      {stage1_3[19]},
      {stage2_4[19],stage2_3[19],stage2_2[19],stage2_1[19],stage2_0[19]}
   );
   gpc606_5 gpc614 (
      {stage1_0[60], stage1_0[61], stage1_0[62], stage1_0[63], stage1_0[64], stage1_0[65]},
      {stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23], stage1_2[24], stage1_2[25]},
      {stage2_4[20],stage2_3[20],stage2_2[20],stage2_1[20],stage2_0[20]}
   );
   gpc606_5 gpc615 (
      {stage1_0[66], stage1_0[67], stage1_0[68], stage1_0[69], stage1_0[70], stage1_0[71]},
      {stage1_2[26], stage1_2[27], stage1_2[28], stage1_2[29], stage1_2[30], stage1_2[31]},
      {stage2_4[21],stage2_3[21],stage2_2[21],stage2_1[21],stage2_0[21]}
   );
   gpc606_5 gpc616 (
      {stage1_0[72], stage1_0[73], stage1_0[74], stage1_0[75], stage1_0[76], stage1_0[77]},
      {stage1_2[32], stage1_2[33], stage1_2[34], stage1_2[35], stage1_2[36], stage1_2[37]},
      {stage2_4[22],stage2_3[22],stage2_2[22],stage2_1[22],stage2_0[22]}
   );
   gpc606_5 gpc617 (
      {stage1_2[38], stage1_2[39], stage1_2[40], stage1_2[41], stage1_2[42], stage1_2[43]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[0],stage2_4[23],stage2_3[23],stage2_2[23]}
   );
   gpc606_5 gpc618 (
      {stage1_2[44], stage1_2[45], stage1_2[46], stage1_2[47], stage1_2[48], stage1_2[49]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[1],stage2_4[24],stage2_3[24],stage2_2[24]}
   );
   gpc606_5 gpc619 (
      {stage1_2[50], stage1_2[51], stage1_2[52], stage1_2[53], stage1_2[54], stage1_2[55]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[2],stage2_4[25],stage2_3[25],stage2_2[25]}
   );
   gpc606_5 gpc620 (
      {stage1_2[56], stage1_2[57], stage1_2[58], stage1_2[59], stage1_2[60], stage1_2[61]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[3],stage2_4[26],stage2_3[26],stage2_2[26]}
   );
   gpc606_5 gpc621 (
      {stage1_2[62], stage1_2[63], stage1_2[64], stage1_2[65], stage1_2[66], stage1_2[67]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[4],stage2_4[27],stage2_3[27],stage2_2[27]}
   );
   gpc615_5 gpc622 (
      {stage1_2[68], stage1_2[69], stage1_2[70], stage1_2[71], stage1_2[72]},
      {stage1_3[20]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[5],stage2_4[28],stage2_3[28],stage2_2[28]}
   );
   gpc615_5 gpc623 (
      {stage1_2[73], stage1_2[74], stage1_2[75], stage1_2[76], stage1_2[77]},
      {stage1_3[21]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[6],stage2_4[29],stage2_3[29],stage2_2[29]}
   );
   gpc615_5 gpc624 (
      {stage1_2[78], stage1_2[79], stage1_2[80], stage1_2[81], stage1_2[82]},
      {stage1_3[22]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[7],stage2_4[30],stage2_3[30],stage2_2[30]}
   );
   gpc615_5 gpc625 (
      {stage1_2[83], stage1_2[84], stage1_2[85], stage1_2[86], stage1_2[87]},
      {stage1_3[23]},
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage2_6[8],stage2_5[8],stage2_4[31],stage2_3[31],stage2_2[31]}
   );
   gpc615_5 gpc626 (
      {stage1_2[88], stage1_2[89], stage1_2[90], stage1_2[91], stage1_2[92]},
      {stage1_3[24]},
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage2_6[9],stage2_5[9],stage2_4[32],stage2_3[32],stage2_2[32]}
   );
   gpc615_5 gpc627 (
      {stage1_2[93], stage1_2[94], stage1_2[95], stage1_2[96], stage1_2[97]},
      {stage1_3[25]},
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage2_6[10],stage2_5[10],stage2_4[33],stage2_3[33],stage2_2[33]}
   );
   gpc615_5 gpc628 (
      {stage1_2[98], stage1_2[99], stage1_2[100], stage1_2[101], stage1_2[102]},
      {stage1_3[26]},
      {stage1_4[66], stage1_4[67], stage1_4[68], stage1_4[69], stage1_4[70], stage1_4[71]},
      {stage2_6[11],stage2_5[11],stage2_4[34],stage2_3[34],stage2_2[34]}
   );
   gpc615_5 gpc629 (
      {stage1_2[103], stage1_2[104], stage1_2[105], stage1_2[106], stage1_2[107]},
      {stage1_3[27]},
      {stage1_4[72], stage1_4[73], stage1_4[74], stage1_4[75], stage1_4[76], stage1_4[77]},
      {stage2_6[12],stage2_5[12],stage2_4[35],stage2_3[35],stage2_2[35]}
   );
   gpc615_5 gpc630 (
      {stage1_2[108], stage1_2[109], stage1_2[110], stage1_2[111], stage1_2[112]},
      {stage1_3[28]},
      {stage1_4[78], stage1_4[79], stage1_4[80], stage1_4[81], stage1_4[82], stage1_4[83]},
      {stage2_6[13],stage2_5[13],stage2_4[36],stage2_3[36],stage2_2[36]}
   );
   gpc615_5 gpc631 (
      {stage1_2[113], stage1_2[114], stage1_2[115], stage1_2[116], stage1_2[117]},
      {stage1_3[29]},
      {stage1_4[84], stage1_4[85], stage1_4[86], stage1_4[87], stage1_4[88], stage1_4[89]},
      {stage2_6[14],stage2_5[14],stage2_4[37],stage2_3[37],stage2_2[37]}
   );
   gpc615_5 gpc632 (
      {stage1_2[118], stage1_2[119], stage1_2[120], stage1_2[121], stage1_2[122]},
      {stage1_3[30]},
      {stage1_4[90], stage1_4[91], stage1_4[92], stage1_4[93], stage1_4[94], stage1_4[95]},
      {stage2_6[15],stage2_5[15],stage2_4[38],stage2_3[38],stage2_2[38]}
   );
   gpc615_5 gpc633 (
      {stage1_2[123], stage1_2[124], stage1_2[125], stage1_2[126], stage1_2[127]},
      {stage1_3[31]},
      {stage1_4[96], stage1_4[97], stage1_4[98], stage1_4[99], stage1_4[100], stage1_4[101]},
      {stage2_6[16],stage2_5[16],stage2_4[39],stage2_3[39],stage2_2[39]}
   );
   gpc615_5 gpc634 (
      {stage1_2[128], stage1_2[129], stage1_2[130], stage1_2[131], stage1_2[132]},
      {stage1_3[32]},
      {stage1_4[102], stage1_4[103], stage1_4[104], stage1_4[105], stage1_4[106], stage1_4[107]},
      {stage2_6[17],stage2_5[17],stage2_4[40],stage2_3[40],stage2_2[40]}
   );
   gpc615_5 gpc635 (
      {stage1_2[133], stage1_2[134], stage1_2[135], stage1_2[136], stage1_2[137]},
      {stage1_3[33]},
      {stage1_4[108], stage1_4[109], stage1_4[110], stage1_4[111], stage1_4[112], stage1_4[113]},
      {stage2_6[18],stage2_5[18],stage2_4[41],stage2_3[41],stage2_2[41]}
   );
   gpc615_5 gpc636 (
      {stage1_2[138], stage1_2[139], stage1_2[140], stage1_2[141], stage1_2[142]},
      {stage1_3[34]},
      {stage1_4[114], stage1_4[115], stage1_4[116], stage1_4[117], stage1_4[118], stage1_4[119]},
      {stage2_6[19],stage2_5[19],stage2_4[42],stage2_3[42],stage2_2[42]}
   );
   gpc615_5 gpc637 (
      {stage1_2[143], stage1_2[144], stage1_2[145], stage1_2[146], stage1_2[147]},
      {stage1_3[35]},
      {stage1_4[120], stage1_4[121], stage1_4[122], stage1_4[123], stage1_4[124], stage1_4[125]},
      {stage2_6[20],stage2_5[20],stage2_4[43],stage2_3[43],stage2_2[43]}
   );
   gpc615_5 gpc638 (
      {stage1_2[148], stage1_2[149], stage1_2[150], stage1_2[151], stage1_2[152]},
      {stage1_3[36]},
      {stage1_4[126], stage1_4[127], stage1_4[128], stage1_4[129], stage1_4[130], stage1_4[131]},
      {stage2_6[21],stage2_5[21],stage2_4[44],stage2_3[44],stage2_2[44]}
   );
   gpc615_5 gpc639 (
      {stage1_2[153], stage1_2[154], stage1_2[155], stage1_2[156], stage1_2[157]},
      {stage1_3[37]},
      {stage1_4[132], stage1_4[133], stage1_4[134], stage1_4[135], stage1_4[136], stage1_4[137]},
      {stage2_6[22],stage2_5[22],stage2_4[45],stage2_3[45],stage2_2[45]}
   );
   gpc615_5 gpc640 (
      {stage1_2[158], stage1_2[159], stage1_2[160], stage1_2[161], stage1_2[162]},
      {stage1_3[38]},
      {stage1_4[138], stage1_4[139], stage1_4[140], stage1_4[141], stage1_4[142], stage1_4[143]},
      {stage2_6[23],stage2_5[23],stage2_4[46],stage2_3[46],stage2_2[46]}
   );
   gpc615_5 gpc641 (
      {stage1_2[163], stage1_2[164], stage1_2[165], stage1_2[166], stage1_2[167]},
      {stage1_3[39]},
      {stage1_4[144], stage1_4[145], stage1_4[146], stage1_4[147], stage1_4[148], stage1_4[149]},
      {stage2_6[24],stage2_5[24],stage2_4[47],stage2_3[47],stage2_2[47]}
   );
   gpc615_5 gpc642 (
      {stage1_2[168], stage1_2[169], stage1_2[170], stage1_2[171], stage1_2[172]},
      {stage1_3[40]},
      {stage1_4[150], stage1_4[151], stage1_4[152], stage1_4[153], stage1_4[154], stage1_4[155]},
      {stage2_6[25],stage2_5[25],stage2_4[48],stage2_3[48],stage2_2[48]}
   );
   gpc615_5 gpc643 (
      {stage1_2[173], stage1_2[174], stage1_2[175], stage1_2[176], stage1_2[177]},
      {stage1_3[41]},
      {stage1_4[156], stage1_4[157], stage1_4[158], stage1_4[159], stage1_4[160], stage1_4[161]},
      {stage2_6[26],stage2_5[26],stage2_4[49],stage2_3[49],stage2_2[49]}
   );
   gpc615_5 gpc644 (
      {stage1_2[178], stage1_2[179], stage1_2[180], stage1_2[181], stage1_2[182]},
      {stage1_3[42]},
      {stage1_4[162], stage1_4[163], stage1_4[164], stage1_4[165], stage1_4[166], stage1_4[167]},
      {stage2_6[27],stage2_5[27],stage2_4[50],stage2_3[50],stage2_2[50]}
   );
   gpc615_5 gpc645 (
      {stage1_2[183], stage1_2[184], stage1_2[185], stage1_2[186], stage1_2[187]},
      {stage1_3[43]},
      {stage1_4[168], stage1_4[169], stage1_4[170], stage1_4[171], stage1_4[172], stage1_4[173]},
      {stage2_6[28],stage2_5[28],stage2_4[51],stage2_3[51],stage2_2[51]}
   );
   gpc615_5 gpc646 (
      {stage1_2[188], stage1_2[189], stage1_2[190], stage1_2[191], stage1_2[192]},
      {stage1_3[44]},
      {stage1_4[174], stage1_4[175], stage1_4[176], stage1_4[177], stage1_4[178], stage1_4[179]},
      {stage2_6[29],stage2_5[29],stage2_4[52],stage2_3[52],stage2_2[52]}
   );
   gpc615_5 gpc647 (
      {stage1_2[193], stage1_2[194], stage1_2[195], stage1_2[196], stage1_2[197]},
      {stage1_3[45]},
      {stage1_4[180], stage1_4[181], stage1_4[182], stage1_4[183], stage1_4[184], stage1_4[185]},
      {stage2_6[30],stage2_5[30],stage2_4[53],stage2_3[53],stage2_2[53]}
   );
   gpc615_5 gpc648 (
      {stage1_3[46], stage1_3[47], stage1_3[48], stage1_3[49], stage1_3[50]},
      {stage1_4[186]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[31],stage2_5[31],stage2_4[54],stage2_3[54]}
   );
   gpc615_5 gpc649 (
      {stage1_3[51], stage1_3[52], stage1_3[53], stage1_3[54], stage1_3[55]},
      {stage1_4[187]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[32],stage2_5[32],stage2_4[55],stage2_3[55]}
   );
   gpc615_5 gpc650 (
      {stage1_3[56], stage1_3[57], stage1_3[58], stage1_3[59], stage1_3[60]},
      {stage1_4[188]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[33],stage2_5[33],stage2_4[56],stage2_3[56]}
   );
   gpc615_5 gpc651 (
      {stage1_3[61], stage1_3[62], stage1_3[63], stage1_3[64], stage1_3[65]},
      {stage1_4[189]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[34],stage2_5[34],stage2_4[57],stage2_3[57]}
   );
   gpc615_5 gpc652 (
      {stage1_3[66], stage1_3[67], stage1_3[68], stage1_3[69], stage1_3[70]},
      {stage1_4[190]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[35],stage2_5[35],stage2_4[58],stage2_3[58]}
   );
   gpc615_5 gpc653 (
      {stage1_3[71], stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75]},
      {stage1_4[191]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[36],stage2_5[36],stage2_4[59],stage2_3[59]}
   );
   gpc615_5 gpc654 (
      {stage1_3[76], stage1_3[77], stage1_3[78], stage1_3[79], stage1_3[80]},
      {stage1_4[192]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[37],stage2_5[37],stage2_4[60],stage2_3[60]}
   );
   gpc615_5 gpc655 (
      {stage1_3[81], stage1_3[82], stage1_3[83], stage1_3[84], stage1_3[85]},
      {stage1_4[193]},
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage2_7[7],stage2_6[38],stage2_5[38],stage2_4[61],stage2_3[61]}
   );
   gpc615_5 gpc656 (
      {stage1_3[86], stage1_3[87], stage1_3[88], stage1_3[89], stage1_3[90]},
      {stage1_4[194]},
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage2_7[8],stage2_6[39],stage2_5[39],stage2_4[62],stage2_3[62]}
   );
   gpc615_5 gpc657 (
      {stage1_3[91], stage1_3[92], stage1_3[93], stage1_3[94], stage1_3[95]},
      {stage1_4[195]},
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage2_7[9],stage2_6[40],stage2_5[40],stage2_4[63],stage2_3[63]}
   );
   gpc615_5 gpc658 (
      {stage1_3[96], stage1_3[97], stage1_3[98], stage1_3[99], stage1_3[100]},
      {stage1_4[196]},
      {stage1_5[60], stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65]},
      {stage2_7[10],stage2_6[41],stage2_5[41],stage2_4[64],stage2_3[64]}
   );
   gpc615_5 gpc659 (
      {stage1_3[101], stage1_3[102], stage1_3[103], stage1_3[104], stage1_3[105]},
      {stage1_4[197]},
      {stage1_5[66], stage1_5[67], stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71]},
      {stage2_7[11],stage2_6[42],stage2_5[42],stage2_4[65],stage2_3[65]}
   );
   gpc615_5 gpc660 (
      {stage1_3[106], stage1_3[107], stage1_3[108], stage1_3[109], stage1_3[110]},
      {stage1_4[198]},
      {stage1_5[72], stage1_5[73], stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77]},
      {stage2_7[12],stage2_6[43],stage2_5[43],stage2_4[66],stage2_3[66]}
   );
   gpc615_5 gpc661 (
      {stage1_3[111], stage1_3[112], stage1_3[113], stage1_3[114], stage1_3[115]},
      {stage1_4[199]},
      {stage1_5[78], stage1_5[79], stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83]},
      {stage2_7[13],stage2_6[44],stage2_5[44],stage2_4[67],stage2_3[67]}
   );
   gpc615_5 gpc662 (
      {stage1_3[116], stage1_3[117], stage1_3[118], stage1_3[119], stage1_3[120]},
      {stage1_4[200]},
      {stage1_5[84], stage1_5[85], stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89]},
      {stage2_7[14],stage2_6[45],stage2_5[45],stage2_4[68],stage2_3[68]}
   );
   gpc615_5 gpc663 (
      {stage1_3[121], stage1_3[122], stage1_3[123], stage1_3[124], stage1_3[125]},
      {stage1_4[201]},
      {stage1_5[90], stage1_5[91], stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95]},
      {stage2_7[15],stage2_6[46],stage2_5[46],stage2_4[69],stage2_3[69]}
   );
   gpc615_5 gpc664 (
      {stage1_3[126], stage1_3[127], stage1_3[128], stage1_3[129], stage1_3[130]},
      {stage1_4[202]},
      {stage1_5[96], stage1_5[97], stage1_5[98], stage1_5[99], stage1_5[100], stage1_5[101]},
      {stage2_7[16],stage2_6[47],stage2_5[47],stage2_4[70],stage2_3[70]}
   );
   gpc615_5 gpc665 (
      {stage1_3[131], stage1_3[132], stage1_3[133], stage1_3[134], stage1_3[135]},
      {stage1_4[203]},
      {stage1_5[102], stage1_5[103], stage1_5[104], stage1_5[105], stage1_5[106], stage1_5[107]},
      {stage2_7[17],stage2_6[48],stage2_5[48],stage2_4[71],stage2_3[71]}
   );
   gpc615_5 gpc666 (
      {stage1_3[136], stage1_3[137], stage1_3[138], stage1_3[139], stage1_3[140]},
      {stage1_4[204]},
      {stage1_5[108], stage1_5[109], stage1_5[110], stage1_5[111], stage1_5[112], stage1_5[113]},
      {stage2_7[18],stage2_6[49],stage2_5[49],stage2_4[72],stage2_3[72]}
   );
   gpc615_5 gpc667 (
      {stage1_3[141], stage1_3[142], stage1_3[143], stage1_3[144], stage1_3[145]},
      {stage1_4[205]},
      {stage1_5[114], stage1_5[115], stage1_5[116], stage1_5[117], stage1_5[118], stage1_5[119]},
      {stage2_7[19],stage2_6[50],stage2_5[50],stage2_4[73],stage2_3[73]}
   );
   gpc615_5 gpc668 (
      {stage1_3[146], stage1_3[147], stage1_3[148], stage1_3[149], stage1_3[150]},
      {stage1_4[206]},
      {stage1_5[120], stage1_5[121], stage1_5[122], stage1_5[123], stage1_5[124], stage1_5[125]},
      {stage2_7[20],stage2_6[51],stage2_5[51],stage2_4[74],stage2_3[74]}
   );
   gpc615_5 gpc669 (
      {stage1_3[151], stage1_3[152], stage1_3[153], stage1_3[154], stage1_3[155]},
      {stage1_4[207]},
      {stage1_5[126], stage1_5[127], stage1_5[128], stage1_5[129], stage1_5[130], stage1_5[131]},
      {stage2_7[21],stage2_6[52],stage2_5[52],stage2_4[75],stage2_3[75]}
   );
   gpc615_5 gpc670 (
      {stage1_3[156], stage1_3[157], stage1_3[158], stage1_3[159], stage1_3[160]},
      {stage1_4[208]},
      {stage1_5[132], stage1_5[133], stage1_5[134], stage1_5[135], stage1_5[136], stage1_5[137]},
      {stage2_7[22],stage2_6[53],stage2_5[53],stage2_4[76],stage2_3[76]}
   );
   gpc615_5 gpc671 (
      {stage1_3[161], stage1_3[162], stage1_3[163], stage1_3[164], stage1_3[165]},
      {stage1_4[209]},
      {stage1_5[138], stage1_5[139], stage1_5[140], stage1_5[141], stage1_5[142], stage1_5[143]},
      {stage2_7[23],stage2_6[54],stage2_5[54],stage2_4[77],stage2_3[77]}
   );
   gpc615_5 gpc672 (
      {stage1_3[166], stage1_3[167], stage1_3[168], stage1_3[169], stage1_3[170]},
      {stage1_4[210]},
      {stage1_5[144], stage1_5[145], stage1_5[146], stage1_5[147], stage1_5[148], stage1_5[149]},
      {stage2_7[24],stage2_6[55],stage2_5[55],stage2_4[78],stage2_3[78]}
   );
   gpc615_5 gpc673 (
      {stage1_3[171], stage1_3[172], stage1_3[173], stage1_3[174], stage1_3[175]},
      {stage1_4[211]},
      {stage1_5[150], stage1_5[151], stage1_5[152], stage1_5[153], stage1_5[154], stage1_5[155]},
      {stage2_7[25],stage2_6[56],stage2_5[56],stage2_4[79],stage2_3[79]}
   );
   gpc615_5 gpc674 (
      {stage1_3[176], stage1_3[177], stage1_3[178], stage1_3[179], stage1_3[180]},
      {stage1_4[212]},
      {stage1_5[156], stage1_5[157], stage1_5[158], stage1_5[159], stage1_5[160], stage1_5[161]},
      {stage2_7[26],stage2_6[57],stage2_5[57],stage2_4[80],stage2_3[80]}
   );
   gpc615_5 gpc675 (
      {stage1_3[181], stage1_3[182], stage1_3[183], stage1_3[184], stage1_3[185]},
      {stage1_4[213]},
      {stage1_5[162], stage1_5[163], stage1_5[164], stage1_5[165], stage1_5[166], stage1_5[167]},
      {stage2_7[27],stage2_6[58],stage2_5[58],stage2_4[81],stage2_3[81]}
   );
   gpc615_5 gpc676 (
      {stage1_3[186], stage1_3[187], stage1_3[188], stage1_3[189], stage1_3[190]},
      {stage1_4[214]},
      {stage1_5[168], stage1_5[169], stage1_5[170], stage1_5[171], stage1_5[172], stage1_5[173]},
      {stage2_7[28],stage2_6[59],stage2_5[59],stage2_4[82],stage2_3[82]}
   );
   gpc615_5 gpc677 (
      {stage1_3[191], stage1_3[192], stage1_3[193], stage1_3[194], stage1_3[195]},
      {stage1_4[215]},
      {stage1_5[174], stage1_5[175], stage1_5[176], stage1_5[177], stage1_5[178], stage1_5[179]},
      {stage2_7[29],stage2_6[60],stage2_5[60],stage2_4[83],stage2_3[83]}
   );
   gpc606_5 gpc678 (
      {stage1_4[216], stage1_4[217], stage1_4[218], stage1_4[219], stage1_4[220], stage1_4[221]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[30],stage2_6[61],stage2_5[61],stage2_4[84]}
   );
   gpc606_5 gpc679 (
      {stage1_4[222], stage1_4[223], stage1_4[224], stage1_4[225], stage1_4[226], stage1_4[227]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[31],stage2_6[62],stage2_5[62],stage2_4[85]}
   );
   gpc606_5 gpc680 (
      {stage1_4[228], stage1_4[229], stage1_4[230], stage1_4[231], stage1_4[232], stage1_4[233]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[32],stage2_6[63],stage2_5[63],stage2_4[86]}
   );
   gpc606_5 gpc681 (
      {stage1_4[234], stage1_4[235], stage1_4[236], stage1_4[237], stage1_4[238], stage1_4[239]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[33],stage2_6[64],stage2_5[64],stage2_4[87]}
   );
   gpc606_5 gpc682 (
      {stage1_5[180], stage1_5[181], stage1_5[182], stage1_5[183], stage1_5[184], stage1_5[185]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[4],stage2_7[34],stage2_6[65],stage2_5[65]}
   );
   gpc606_5 gpc683 (
      {stage1_5[186], stage1_5[187], stage1_5[188], stage1_5[189], stage1_5[190], stage1_5[191]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[5],stage2_7[35],stage2_6[66],stage2_5[66]}
   );
   gpc606_5 gpc684 (
      {stage1_5[192], stage1_5[193], stage1_5[194], stage1_5[195], stage1_5[196], stage1_5[197]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[6],stage2_7[36],stage2_6[67],stage2_5[67]}
   );
   gpc606_5 gpc685 (
      {stage1_5[198], stage1_5[199], stage1_5[200], stage1_5[201], stage1_5[202], stage1_5[203]},
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage2_9[3],stage2_8[7],stage2_7[37],stage2_6[68],stage2_5[68]}
   );
   gpc606_5 gpc686 (
      {stage1_5[204], stage1_5[205], stage1_5[206], stage1_5[207], stage1_5[208], stage1_5[209]},
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29]},
      {stage2_9[4],stage2_8[8],stage2_7[38],stage2_6[69],stage2_5[69]}
   );
   gpc606_5 gpc687 (
      {stage1_5[210], stage1_5[211], stage1_5[212], stage1_5[213], stage1_5[214], stage1_5[215]},
      {stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35]},
      {stage2_9[5],stage2_8[9],stage2_7[39],stage2_6[70],stage2_5[70]}
   );
   gpc606_5 gpc688 (
      {stage1_5[216], stage1_5[217], stage1_5[218], stage1_5[219], stage1_5[220], stage1_5[221]},
      {stage1_7[36], stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage2_9[6],stage2_8[10],stage2_7[40],stage2_6[71],stage2_5[71]}
   );
   gpc606_5 gpc689 (
      {stage1_5[222], stage1_5[223], stage1_5[224], stage1_5[225], stage1_5[226], stage1_5[227]},
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47]},
      {stage2_9[7],stage2_8[11],stage2_7[41],stage2_6[72],stage2_5[72]}
   );
   gpc606_5 gpc690 (
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[8],stage2_8[12],stage2_7[42],stage2_6[73]}
   );
   gpc606_5 gpc691 (
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[9],stage2_8[13],stage2_7[43],stage2_6[74]}
   );
   gpc606_5 gpc692 (
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[10],stage2_8[14],stage2_7[44],stage2_6[75]}
   );
   gpc606_5 gpc693 (
      {stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[11],stage2_8[15],stage2_7[45],stage2_6[76]}
   );
   gpc606_5 gpc694 (
      {stage1_6[48], stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[12],stage2_8[16],stage2_7[46],stage2_6[77]}
   );
   gpc606_5 gpc695 (
      {stage1_6[54], stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[13],stage2_8[17],stage2_7[47],stage2_6[78]}
   );
   gpc606_5 gpc696 (
      {stage1_6[60], stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65]},
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage2_10[6],stage2_9[14],stage2_8[18],stage2_7[48],stage2_6[79]}
   );
   gpc606_5 gpc697 (
      {stage1_6[66], stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71]},
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage2_10[7],stage2_9[15],stage2_8[19],stage2_7[49],stage2_6[80]}
   );
   gpc606_5 gpc698 (
      {stage1_6[72], stage1_6[73], stage1_6[74], stage1_6[75], stage1_6[76], stage1_6[77]},
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage2_10[8],stage2_9[16],stage2_8[20],stage2_7[50],stage2_6[81]}
   );
   gpc606_5 gpc699 (
      {stage1_6[78], stage1_6[79], stage1_6[80], stage1_6[81], stage1_6[82], stage1_6[83]},
      {stage1_8[54], stage1_8[55], stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59]},
      {stage2_10[9],stage2_9[17],stage2_8[21],stage2_7[51],stage2_6[82]}
   );
   gpc606_5 gpc700 (
      {stage1_6[84], stage1_6[85], stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89]},
      {stage1_8[60], stage1_8[61], stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65]},
      {stage2_10[10],stage2_9[18],stage2_8[22],stage2_7[52],stage2_6[83]}
   );
   gpc606_5 gpc701 (
      {stage1_6[90], stage1_6[91], stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95]},
      {stage1_8[66], stage1_8[67], stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71]},
      {stage2_10[11],stage2_9[19],stage2_8[23],stage2_7[53],stage2_6[84]}
   );
   gpc606_5 gpc702 (
      {stage1_6[96], stage1_6[97], stage1_6[98], stage1_6[99], stage1_6[100], stage1_6[101]},
      {stage1_8[72], stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77]},
      {stage2_10[12],stage2_9[20],stage2_8[24],stage2_7[54],stage2_6[85]}
   );
   gpc606_5 gpc703 (
      {stage1_6[102], stage1_6[103], stage1_6[104], stage1_6[105], stage1_6[106], stage1_6[107]},
      {stage1_8[78], stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83]},
      {stage2_10[13],stage2_9[21],stage2_8[25],stage2_7[55],stage2_6[86]}
   );
   gpc606_5 gpc704 (
      {stage1_6[108], stage1_6[109], stage1_6[110], stage1_6[111], stage1_6[112], stage1_6[113]},
      {stage1_8[84], stage1_8[85], stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89]},
      {stage2_10[14],stage2_9[22],stage2_8[26],stage2_7[56],stage2_6[87]}
   );
   gpc606_5 gpc705 (
      {stage1_6[114], stage1_6[115], stage1_6[116], stage1_6[117], stage1_6[118], stage1_6[119]},
      {stage1_8[90], stage1_8[91], stage1_8[92], stage1_8[93], stage1_8[94], stage1_8[95]},
      {stage2_10[15],stage2_9[23],stage2_8[27],stage2_7[57],stage2_6[88]}
   );
   gpc606_5 gpc706 (
      {stage1_6[120], stage1_6[121], stage1_6[122], stage1_6[123], stage1_6[124], stage1_6[125]},
      {stage1_8[96], stage1_8[97], stage1_8[98], stage1_8[99], stage1_8[100], stage1_8[101]},
      {stage2_10[16],stage2_9[24],stage2_8[28],stage2_7[58],stage2_6[89]}
   );
   gpc606_5 gpc707 (
      {stage1_6[126], stage1_6[127], stage1_6[128], stage1_6[129], stage1_6[130], stage1_6[131]},
      {stage1_8[102], stage1_8[103], stage1_8[104], stage1_8[105], stage1_8[106], stage1_8[107]},
      {stage2_10[17],stage2_9[25],stage2_8[29],stage2_7[59],stage2_6[90]}
   );
   gpc606_5 gpc708 (
      {stage1_6[132], stage1_6[133], stage1_6[134], stage1_6[135], stage1_6[136], stage1_6[137]},
      {stage1_8[108], stage1_8[109], stage1_8[110], stage1_8[111], stage1_8[112], stage1_8[113]},
      {stage2_10[18],stage2_9[26],stage2_8[30],stage2_7[60],stage2_6[91]}
   );
   gpc606_5 gpc709 (
      {stage1_6[138], stage1_6[139], stage1_6[140], stage1_6[141], stage1_6[142], stage1_6[143]},
      {stage1_8[114], stage1_8[115], stage1_8[116], stage1_8[117], stage1_8[118], stage1_8[119]},
      {stage2_10[19],stage2_9[27],stage2_8[31],stage2_7[61],stage2_6[92]}
   );
   gpc606_5 gpc710 (
      {stage1_6[144], stage1_6[145], stage1_6[146], stage1_6[147], stage1_6[148], stage1_6[149]},
      {stage1_8[120], stage1_8[121], stage1_8[122], stage1_8[123], stage1_8[124], stage1_8[125]},
      {stage2_10[20],stage2_9[28],stage2_8[32],stage2_7[62],stage2_6[93]}
   );
   gpc615_5 gpc711 (
      {stage1_6[150], stage1_6[151], stage1_6[152], stage1_6[153], stage1_6[154]},
      {stage1_7[48]},
      {stage1_8[126], stage1_8[127], stage1_8[128], stage1_8[129], stage1_8[130], stage1_8[131]},
      {stage2_10[21],stage2_9[29],stage2_8[33],stage2_7[63],stage2_6[94]}
   );
   gpc615_5 gpc712 (
      {stage1_6[155], stage1_6[156], stage1_6[157], stage1_6[158], stage1_6[159]},
      {stage1_7[49]},
      {stage1_8[132], stage1_8[133], stage1_8[134], stage1_8[135], stage1_8[136], stage1_8[137]},
      {stage2_10[22],stage2_9[30],stage2_8[34],stage2_7[64],stage2_6[95]}
   );
   gpc615_5 gpc713 (
      {stage1_6[160], stage1_6[161], stage1_6[162], stage1_6[163], stage1_6[164]},
      {stage1_7[50]},
      {stage1_8[138], stage1_8[139], stage1_8[140], stage1_8[141], stage1_8[142], stage1_8[143]},
      {stage2_10[23],stage2_9[31],stage2_8[35],stage2_7[65],stage2_6[96]}
   );
   gpc615_5 gpc714 (
      {stage1_6[165], stage1_6[166], stage1_6[167], stage1_6[168], stage1_6[169]},
      {stage1_7[51]},
      {stage1_8[144], stage1_8[145], stage1_8[146], stage1_8[147], stage1_8[148], stage1_8[149]},
      {stage2_10[24],stage2_9[32],stage2_8[36],stage2_7[66],stage2_6[97]}
   );
   gpc615_5 gpc715 (
      {stage1_7[52], stage1_7[53], stage1_7[54], stage1_7[55], stage1_7[56]},
      {stage1_8[150]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[25],stage2_9[33],stage2_8[37],stage2_7[67]}
   );
   gpc615_5 gpc716 (
      {stage1_7[57], stage1_7[58], stage1_7[59], stage1_7[60], stage1_7[61]},
      {stage1_8[151]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[26],stage2_9[34],stage2_8[38],stage2_7[68]}
   );
   gpc615_5 gpc717 (
      {stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65], stage1_7[66]},
      {stage1_8[152]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[27],stage2_9[35],stage2_8[39],stage2_7[69]}
   );
   gpc615_5 gpc718 (
      {stage1_7[67], stage1_7[68], stage1_7[69], stage1_7[70], stage1_7[71]},
      {stage1_8[153]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[28],stage2_9[36],stage2_8[40],stage2_7[70]}
   );
   gpc615_5 gpc719 (
      {stage1_7[72], stage1_7[73], stage1_7[74], stage1_7[75], stage1_7[76]},
      {stage1_8[154]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[29],stage2_9[37],stage2_8[41],stage2_7[71]}
   );
   gpc615_5 gpc720 (
      {stage1_7[77], stage1_7[78], stage1_7[79], stage1_7[80], stage1_7[81]},
      {stage1_8[155]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[30],stage2_9[38],stage2_8[42],stage2_7[72]}
   );
   gpc615_5 gpc721 (
      {stage1_7[82], stage1_7[83], stage1_7[84], stage1_7[85], stage1_7[86]},
      {stage1_8[156]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[31],stage2_9[39],stage2_8[43],stage2_7[73]}
   );
   gpc615_5 gpc722 (
      {stage1_7[87], stage1_7[88], stage1_7[89], stage1_7[90], stage1_7[91]},
      {stage1_8[157]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[32],stage2_9[40],stage2_8[44],stage2_7[74]}
   );
   gpc615_5 gpc723 (
      {stage1_7[92], stage1_7[93], stage1_7[94], stage1_7[95], stage1_7[96]},
      {stage1_8[158]},
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage2_11[8],stage2_10[33],stage2_9[41],stage2_8[45],stage2_7[75]}
   );
   gpc615_5 gpc724 (
      {stage1_7[97], stage1_7[98], stage1_7[99], stage1_7[100], stage1_7[101]},
      {stage1_8[159]},
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage2_11[9],stage2_10[34],stage2_9[42],stage2_8[46],stage2_7[76]}
   );
   gpc615_5 gpc725 (
      {stage1_7[102], stage1_7[103], stage1_7[104], stage1_7[105], stage1_7[106]},
      {stage1_8[160]},
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage2_11[10],stage2_10[35],stage2_9[43],stage2_8[47],stage2_7[77]}
   );
   gpc615_5 gpc726 (
      {stage1_7[107], stage1_7[108], stage1_7[109], stage1_7[110], stage1_7[111]},
      {stage1_8[161]},
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage2_11[11],stage2_10[36],stage2_9[44],stage2_8[48],stage2_7[78]}
   );
   gpc615_5 gpc727 (
      {stage1_7[112], stage1_7[113], stage1_7[114], stage1_7[115], stage1_7[116]},
      {stage1_8[162]},
      {stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77]},
      {stage2_11[12],stage2_10[37],stage2_9[45],stage2_8[49],stage2_7[79]}
   );
   gpc615_5 gpc728 (
      {stage1_7[117], stage1_7[118], stage1_7[119], stage1_7[120], stage1_7[121]},
      {stage1_8[163]},
      {stage1_9[78], stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83]},
      {stage2_11[13],stage2_10[38],stage2_9[46],stage2_8[50],stage2_7[80]}
   );
   gpc615_5 gpc729 (
      {stage1_7[122], stage1_7[123], stage1_7[124], stage1_7[125], stage1_7[126]},
      {stage1_8[164]},
      {stage1_9[84], stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89]},
      {stage2_11[14],stage2_10[39],stage2_9[47],stage2_8[51],stage2_7[81]}
   );
   gpc615_5 gpc730 (
      {stage1_7[127], stage1_7[128], stage1_7[129], stage1_7[130], stage1_7[131]},
      {stage1_8[165]},
      {stage1_9[90], stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95]},
      {stage2_11[15],stage2_10[40],stage2_9[48],stage2_8[52],stage2_7[82]}
   );
   gpc615_5 gpc731 (
      {stage1_7[132], stage1_7[133], stage1_7[134], stage1_7[135], stage1_7[136]},
      {stage1_8[166]},
      {stage1_9[96], stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100], stage1_9[101]},
      {stage2_11[16],stage2_10[41],stage2_9[49],stage2_8[53],stage2_7[83]}
   );
   gpc615_5 gpc732 (
      {stage1_7[137], stage1_7[138], stage1_7[139], stage1_7[140], stage1_7[141]},
      {stage1_8[167]},
      {stage1_9[102], stage1_9[103], stage1_9[104], stage1_9[105], stage1_9[106], stage1_9[107]},
      {stage2_11[17],stage2_10[42],stage2_9[50],stage2_8[54],stage2_7[84]}
   );
   gpc615_5 gpc733 (
      {stage1_7[142], stage1_7[143], stage1_7[144], stage1_7[145], stage1_7[146]},
      {stage1_8[168]},
      {stage1_9[108], stage1_9[109], stage1_9[110], stage1_9[111], stage1_9[112], stage1_9[113]},
      {stage2_11[18],stage2_10[43],stage2_9[51],stage2_8[55],stage2_7[85]}
   );
   gpc615_5 gpc734 (
      {stage1_7[147], stage1_7[148], stage1_7[149], stage1_7[150], stage1_7[151]},
      {stage1_8[169]},
      {stage1_9[114], stage1_9[115], stage1_9[116], stage1_9[117], stage1_9[118], stage1_9[119]},
      {stage2_11[19],stage2_10[44],stage2_9[52],stage2_8[56],stage2_7[86]}
   );
   gpc615_5 gpc735 (
      {stage1_7[152], stage1_7[153], stage1_7[154], stage1_7[155], stage1_7[156]},
      {stage1_8[170]},
      {stage1_9[120], stage1_9[121], stage1_9[122], stage1_9[123], stage1_9[124], stage1_9[125]},
      {stage2_11[20],stage2_10[45],stage2_9[53],stage2_8[57],stage2_7[87]}
   );
   gpc615_5 gpc736 (
      {stage1_7[157], stage1_7[158], stage1_7[159], stage1_7[160], stage1_7[161]},
      {stage1_8[171]},
      {stage1_9[126], stage1_9[127], stage1_9[128], stage1_9[129], stage1_9[130], stage1_9[131]},
      {stage2_11[21],stage2_10[46],stage2_9[54],stage2_8[58],stage2_7[88]}
   );
   gpc606_5 gpc737 (
      {stage1_8[172], stage1_8[173], stage1_8[174], stage1_8[175], stage1_8[176], stage1_8[177]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[22],stage2_10[47],stage2_9[55],stage2_8[59]}
   );
   gpc606_5 gpc738 (
      {stage1_8[178], stage1_8[179], stage1_8[180], stage1_8[181], stage1_8[182], stage1_8[183]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[23],stage2_10[48],stage2_9[56],stage2_8[60]}
   );
   gpc606_5 gpc739 (
      {stage1_8[184], stage1_8[185], stage1_8[186], stage1_8[187], stage1_8[188], stage1_8[189]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[24],stage2_10[49],stage2_9[57],stage2_8[61]}
   );
   gpc606_5 gpc740 (
      {stage1_8[190], stage1_8[191], stage1_8[192], stage1_8[193], stage1_8[194], stage1_8[195]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[25],stage2_10[50],stage2_9[58],stage2_8[62]}
   );
   gpc606_5 gpc741 (
      {stage1_8[196], stage1_8[197], stage1_8[198], stage1_8[199], stage1_8[200], stage1_8[201]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[26],stage2_10[51],stage2_9[59],stage2_8[63]}
   );
   gpc606_5 gpc742 (
      {stage1_8[202], stage1_8[203], stage1_8[204], stage1_8[205], stage1_8[206], stage1_8[207]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[27],stage2_10[52],stage2_9[60],stage2_8[64]}
   );
   gpc606_5 gpc743 (
      {stage1_8[208], stage1_8[209], stage1_8[210], stage1_8[211], stage1_8[212], stage1_8[213]},
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage2_12[6],stage2_11[28],stage2_10[53],stage2_9[61],stage2_8[65]}
   );
   gpc615_5 gpc744 (
      {stage1_8[214], stage1_8[215], stage1_8[216], stage1_8[217], stage1_8[218]},
      {stage1_9[132]},
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage2_12[7],stage2_11[29],stage2_10[54],stage2_9[62],stage2_8[66]}
   );
   gpc615_5 gpc745 (
      {stage1_8[219], stage1_8[220], stage1_8[221], stage1_8[222], stage1_8[223]},
      {stage1_9[133]},
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage2_12[8],stage2_11[30],stage2_10[55],stage2_9[63],stage2_8[67]}
   );
   gpc615_5 gpc746 (
      {stage1_8[224], stage1_8[225], stage1_8[226], stage1_8[227], stage1_8[228]},
      {stage1_9[134]},
      {stage1_10[54], stage1_10[55], stage1_10[56], stage1_10[57], stage1_10[58], stage1_10[59]},
      {stage2_12[9],stage2_11[31],stage2_10[56],stage2_9[64],stage2_8[68]}
   );
   gpc615_5 gpc747 (
      {stage1_8[229], stage1_8[230], stage1_8[231], stage1_8[232], stage1_8[233]},
      {stage1_9[135]},
      {stage1_10[60], stage1_10[61], stage1_10[62], stage1_10[63], stage1_10[64], stage1_10[65]},
      {stage2_12[10],stage2_11[32],stage2_10[57],stage2_9[65],stage2_8[69]}
   );
   gpc615_5 gpc748 (
      {stage1_8[234], stage1_8[235], stage1_8[236], stage1_8[237], stage1_8[238]},
      {stage1_9[136]},
      {stage1_10[66], stage1_10[67], stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71]},
      {stage2_12[11],stage2_11[33],stage2_10[58],stage2_9[66],stage2_8[70]}
   );
   gpc606_5 gpc749 (
      {stage1_9[137], stage1_9[138], stage1_9[139], stage1_9[140], stage1_9[141], stage1_9[142]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[12],stage2_11[34],stage2_10[59],stage2_9[67]}
   );
   gpc606_5 gpc750 (
      {stage1_9[143], stage1_9[144], stage1_9[145], stage1_9[146], stage1_9[147], stage1_9[148]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[13],stage2_11[35],stage2_10[60],stage2_9[68]}
   );
   gpc606_5 gpc751 (
      {stage1_9[149], stage1_9[150], stage1_9[151], stage1_9[152], stage1_9[153], stage1_9[154]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[14],stage2_11[36],stage2_10[61],stage2_9[69]}
   );
   gpc606_5 gpc752 (
      {stage1_9[155], stage1_9[156], stage1_9[157], stage1_9[158], stage1_9[159], stage1_9[160]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[15],stage2_11[37],stage2_10[62],stage2_9[70]}
   );
   gpc606_5 gpc753 (
      {stage1_9[161], stage1_9[162], stage1_9[163], stage1_9[164], stage1_9[165], stage1_9[166]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[16],stage2_11[38],stage2_10[63],stage2_9[71]}
   );
   gpc606_5 gpc754 (
      {stage1_9[167], stage1_9[168], stage1_9[169], stage1_9[170], stage1_9[171], stage1_9[172]},
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage2_13[5],stage2_12[17],stage2_11[39],stage2_10[64],stage2_9[72]}
   );
   gpc606_5 gpc755 (
      {stage1_9[173], stage1_9[174], stage1_9[175], stage1_9[176], stage1_9[177], stage1_9[178]},
      {stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41]},
      {stage2_13[6],stage2_12[18],stage2_11[40],stage2_10[65],stage2_9[73]}
   );
   gpc615_5 gpc756 (
      {stage1_9[179], stage1_9[180], stage1_9[181], stage1_9[182], stage1_9[183]},
      {stage1_10[72]},
      {stage1_11[42], stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage2_13[7],stage2_12[19],stage2_11[41],stage2_10[66],stage2_9[74]}
   );
   gpc615_5 gpc757 (
      {stage1_9[184], stage1_9[185], stage1_9[186], stage1_9[187], stage1_9[188]},
      {stage1_10[73]},
      {stage1_11[48], stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage2_13[8],stage2_12[20],stage2_11[42],stage2_10[67],stage2_9[75]}
   );
   gpc615_5 gpc758 (
      {stage1_9[189], stage1_9[190], stage1_9[191], stage1_9[192], stage1_9[193]},
      {stage1_10[74]},
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58], stage1_11[59]},
      {stage2_13[9],stage2_12[21],stage2_11[43],stage2_10[68],stage2_9[76]}
   );
   gpc615_5 gpc759 (
      {stage1_9[194], stage1_9[195], stage1_9[196], stage1_9[197], stage1_9[198]},
      {stage1_10[75]},
      {stage1_11[60], stage1_11[61], stage1_11[62], stage1_11[63], stage1_11[64], stage1_11[65]},
      {stage2_13[10],stage2_12[22],stage2_11[44],stage2_10[69],stage2_9[77]}
   );
   gpc615_5 gpc760 (
      {stage1_9[199], stage1_9[200], stage1_9[201], stage1_9[202], stage1_9[203]},
      {stage1_10[76]},
      {stage1_11[66], stage1_11[67], stage1_11[68], stage1_11[69], stage1_11[70], stage1_11[71]},
      {stage2_13[11],stage2_12[23],stage2_11[45],stage2_10[70],stage2_9[78]}
   );
   gpc615_5 gpc761 (
      {stage1_9[204], stage1_9[205], stage1_9[206], stage1_9[207], stage1_9[208]},
      {stage1_10[77]},
      {stage1_11[72], stage1_11[73], stage1_11[74], stage1_11[75], stage1_11[76], stage1_11[77]},
      {stage2_13[12],stage2_12[24],stage2_11[46],stage2_10[71],stage2_9[79]}
   );
   gpc615_5 gpc762 (
      {stage1_9[209], stage1_9[210], stage1_9[211], stage1_9[212], stage1_9[213]},
      {stage1_10[78]},
      {stage1_11[78], stage1_11[79], stage1_11[80], stage1_11[81], stage1_11[82], stage1_11[83]},
      {stage2_13[13],stage2_12[25],stage2_11[47],stage2_10[72],stage2_9[80]}
   );
   gpc615_5 gpc763 (
      {stage1_9[214], stage1_9[215], stage1_9[216], stage1_9[217], stage1_9[218]},
      {stage1_10[79]},
      {stage1_11[84], stage1_11[85], stage1_11[86], stage1_11[87], stage1_11[88], stage1_11[89]},
      {stage2_13[14],stage2_12[26],stage2_11[48],stage2_10[73],stage2_9[81]}
   );
   gpc615_5 gpc764 (
      {stage1_9[219], stage1_9[220], stage1_9[221], stage1_9[222], stage1_9[223]},
      {stage1_10[80]},
      {stage1_11[90], stage1_11[91], stage1_11[92], stage1_11[93], stage1_11[94], stage1_11[95]},
      {stage2_13[15],stage2_12[27],stage2_11[49],stage2_10[74],stage2_9[82]}
   );
   gpc615_5 gpc765 (
      {stage1_9[224], stage1_9[225], stage1_9[226], stage1_9[227], stage1_9[228]},
      {stage1_10[81]},
      {stage1_11[96], stage1_11[97], stage1_11[98], stage1_11[99], stage1_11[100], stage1_11[101]},
      {stage2_13[16],stage2_12[28],stage2_11[50],stage2_10[75],stage2_9[83]}
   );
   gpc615_5 gpc766 (
      {stage1_9[229], stage1_9[230], stage1_9[231], stage1_9[232], stage1_9[233]},
      {stage1_10[82]},
      {stage1_11[102], stage1_11[103], stage1_11[104], stage1_11[105], stage1_11[106], stage1_11[107]},
      {stage2_13[17],stage2_12[29],stage2_11[51],stage2_10[76],stage2_9[84]}
   );
   gpc606_5 gpc767 (
      {stage1_10[83], stage1_10[84], stage1_10[85], stage1_10[86], stage1_10[87], stage1_10[88]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[18],stage2_12[30],stage2_11[52],stage2_10[77]}
   );
   gpc606_5 gpc768 (
      {stage1_10[89], stage1_10[90], stage1_10[91], stage1_10[92], stage1_10[93], stage1_10[94]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[19],stage2_12[31],stage2_11[53],stage2_10[78]}
   );
   gpc606_5 gpc769 (
      {stage1_10[95], stage1_10[96], stage1_10[97], stage1_10[98], stage1_10[99], stage1_10[100]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[20],stage2_12[32],stage2_11[54],stage2_10[79]}
   );
   gpc606_5 gpc770 (
      {stage1_10[101], stage1_10[102], stage1_10[103], stage1_10[104], stage1_10[105], stage1_10[106]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[21],stage2_12[33],stage2_11[55],stage2_10[80]}
   );
   gpc606_5 gpc771 (
      {stage1_10[107], stage1_10[108], stage1_10[109], stage1_10[110], stage1_10[111], stage1_10[112]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[22],stage2_12[34],stage2_11[56],stage2_10[81]}
   );
   gpc606_5 gpc772 (
      {stage1_10[113], stage1_10[114], stage1_10[115], stage1_10[116], stage1_10[117], stage1_10[118]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[23],stage2_12[35],stage2_11[57],stage2_10[82]}
   );
   gpc606_5 gpc773 (
      {stage1_10[119], stage1_10[120], stage1_10[121], stage1_10[122], stage1_10[123], stage1_10[124]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[24],stage2_12[36],stage2_11[58],stage2_10[83]}
   );
   gpc606_5 gpc774 (
      {stage1_10[125], stage1_10[126], stage1_10[127], stage1_10[128], stage1_10[129], stage1_10[130]},
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage2_14[7],stage2_13[25],stage2_12[37],stage2_11[59],stage2_10[84]}
   );
   gpc606_5 gpc775 (
      {stage1_10[131], stage1_10[132], stage1_10[133], stage1_10[134], stage1_10[135], stage1_10[136]},
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage2_14[8],stage2_13[26],stage2_12[38],stage2_11[60],stage2_10[85]}
   );
   gpc606_5 gpc776 (
      {stage1_10[137], stage1_10[138], stage1_10[139], stage1_10[140], stage1_10[141], stage1_10[142]},
      {stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage2_14[9],stage2_13[27],stage2_12[39],stage2_11[61],stage2_10[86]}
   );
   gpc606_5 gpc777 (
      {stage1_10[143], stage1_10[144], stage1_10[145], stage1_10[146], stage1_10[147], stage1_10[148]},
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64], stage1_12[65]},
      {stage2_14[10],stage2_13[28],stage2_12[40],stage2_11[62],stage2_10[87]}
   );
   gpc606_5 gpc778 (
      {stage1_10[149], stage1_10[150], stage1_10[151], stage1_10[152], stage1_10[153], stage1_10[154]},
      {stage1_12[66], stage1_12[67], stage1_12[68], stage1_12[69], stage1_12[70], stage1_12[71]},
      {stage2_14[11],stage2_13[29],stage2_12[41],stage2_11[63],stage2_10[88]}
   );
   gpc606_5 gpc779 (
      {stage1_10[155], stage1_10[156], stage1_10[157], stage1_10[158], stage1_10[159], stage1_10[160]},
      {stage1_12[72], stage1_12[73], stage1_12[74], stage1_12[75], stage1_12[76], stage1_12[77]},
      {stage2_14[12],stage2_13[30],stage2_12[42],stage2_11[64],stage2_10[89]}
   );
   gpc606_5 gpc780 (
      {stage1_10[161], stage1_10[162], stage1_10[163], stage1_10[164], stage1_10[165], stage1_10[166]},
      {stage1_12[78], stage1_12[79], stage1_12[80], stage1_12[81], stage1_12[82], stage1_12[83]},
      {stage2_14[13],stage2_13[31],stage2_12[43],stage2_11[65],stage2_10[90]}
   );
   gpc606_5 gpc781 (
      {stage1_10[167], stage1_10[168], stage1_10[169], stage1_10[170], stage1_10[171], stage1_10[172]},
      {stage1_12[84], stage1_12[85], stage1_12[86], stage1_12[87], stage1_12[88], stage1_12[89]},
      {stage2_14[14],stage2_13[32],stage2_12[44],stage2_11[66],stage2_10[91]}
   );
   gpc615_5 gpc782 (
      {stage1_11[108], stage1_11[109], stage1_11[110], stage1_11[111], stage1_11[112]},
      {stage1_12[90]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[15],stage2_13[33],stage2_12[45],stage2_11[67]}
   );
   gpc615_5 gpc783 (
      {stage1_11[113], stage1_11[114], stage1_11[115], stage1_11[116], stage1_11[117]},
      {stage1_12[91]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[16],stage2_13[34],stage2_12[46],stage2_11[68]}
   );
   gpc615_5 gpc784 (
      {stage1_11[118], stage1_11[119], stage1_11[120], stage1_11[121], stage1_11[122]},
      {stage1_12[92]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[17],stage2_13[35],stage2_12[47],stage2_11[69]}
   );
   gpc615_5 gpc785 (
      {stage1_11[123], stage1_11[124], stage1_11[125], stage1_11[126], stage1_11[127]},
      {stage1_12[93]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[18],stage2_13[36],stage2_12[48],stage2_11[70]}
   );
   gpc615_5 gpc786 (
      {stage1_11[128], stage1_11[129], stage1_11[130], stage1_11[131], stage1_11[132]},
      {stage1_12[94]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[19],stage2_13[37],stage2_12[49],stage2_11[71]}
   );
   gpc615_5 gpc787 (
      {stage1_11[133], stage1_11[134], stage1_11[135], stage1_11[136], stage1_11[137]},
      {stage1_12[95]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[20],stage2_13[38],stage2_12[50],stage2_11[72]}
   );
   gpc615_5 gpc788 (
      {stage1_11[138], stage1_11[139], stage1_11[140], stage1_11[141], stage1_11[142]},
      {stage1_12[96]},
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage2_15[6],stage2_14[21],stage2_13[39],stage2_12[51],stage2_11[73]}
   );
   gpc615_5 gpc789 (
      {stage1_11[143], stage1_11[144], stage1_11[145], stage1_11[146], stage1_11[147]},
      {stage1_12[97]},
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage2_15[7],stage2_14[22],stage2_13[40],stage2_12[52],stage2_11[74]}
   );
   gpc615_5 gpc790 (
      {stage1_11[148], stage1_11[149], stage1_11[150], stage1_11[151], stage1_11[152]},
      {stage1_12[98]},
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage2_15[8],stage2_14[23],stage2_13[41],stage2_12[53],stage2_11[75]}
   );
   gpc615_5 gpc791 (
      {stage1_11[153], stage1_11[154], stage1_11[155], stage1_11[156], stage1_11[157]},
      {stage1_12[99]},
      {stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59]},
      {stage2_15[9],stage2_14[24],stage2_13[42],stage2_12[54],stage2_11[76]}
   );
   gpc615_5 gpc792 (
      {stage1_11[158], stage1_11[159], stage1_11[160], stage1_11[161], stage1_11[162]},
      {stage1_12[100]},
      {stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage2_15[10],stage2_14[25],stage2_13[43],stage2_12[55],stage2_11[77]}
   );
   gpc615_5 gpc793 (
      {stage1_11[163], stage1_11[164], stage1_11[165], stage1_11[166], stage1_11[167]},
      {stage1_12[101]},
      {stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69], stage1_13[70], stage1_13[71]},
      {stage2_15[11],stage2_14[26],stage2_13[44],stage2_12[56],stage2_11[78]}
   );
   gpc1_1 gpc794 (
      {stage1_0[78]},
      {stage2_0[23]}
   );
   gpc1_1 gpc795 (
      {stage1_0[79]},
      {stage2_0[24]}
   );
   gpc1_1 gpc796 (
      {stage1_0[80]},
      {stage2_0[25]}
   );
   gpc1_1 gpc797 (
      {stage1_0[81]},
      {stage2_0[26]}
   );
   gpc1_1 gpc798 (
      {stage1_0[82]},
      {stage2_0[27]}
   );
   gpc1_1 gpc799 (
      {stage1_0[83]},
      {stage2_0[28]}
   );
   gpc1_1 gpc800 (
      {stage1_0[84]},
      {stage2_0[29]}
   );
   gpc1_1 gpc801 (
      {stage1_0[85]},
      {stage2_0[30]}
   );
   gpc1_1 gpc802 (
      {stage1_1[120]},
      {stage2_1[23]}
   );
   gpc1_1 gpc803 (
      {stage1_1[121]},
      {stage2_1[24]}
   );
   gpc1_1 gpc804 (
      {stage1_1[122]},
      {stage2_1[25]}
   );
   gpc1_1 gpc805 (
      {stage1_1[123]},
      {stage2_1[26]}
   );
   gpc1_1 gpc806 (
      {stage1_1[124]},
      {stage2_1[27]}
   );
   gpc1_1 gpc807 (
      {stage1_1[125]},
      {stage2_1[28]}
   );
   gpc1_1 gpc808 (
      {stage1_1[126]},
      {stage2_1[29]}
   );
   gpc1_1 gpc809 (
      {stage1_1[127]},
      {stage2_1[30]}
   );
   gpc1_1 gpc810 (
      {stage1_1[128]},
      {stage2_1[31]}
   );
   gpc1_1 gpc811 (
      {stage1_1[129]},
      {stage2_1[32]}
   );
   gpc1_1 gpc812 (
      {stage1_1[130]},
      {stage2_1[33]}
   );
   gpc1_1 gpc813 (
      {stage1_1[131]},
      {stage2_1[34]}
   );
   gpc1_1 gpc814 (
      {stage1_1[132]},
      {stage2_1[35]}
   );
   gpc1_1 gpc815 (
      {stage1_1[133]},
      {stage2_1[36]}
   );
   gpc1_1 gpc816 (
      {stage1_1[134]},
      {stage2_1[37]}
   );
   gpc1_1 gpc817 (
      {stage1_1[135]},
      {stage2_1[38]}
   );
   gpc1_1 gpc818 (
      {stage1_1[136]},
      {stage2_1[39]}
   );
   gpc1_1 gpc819 (
      {stage1_1[137]},
      {stage2_1[40]}
   );
   gpc1_1 gpc820 (
      {stage1_1[138]},
      {stage2_1[41]}
   );
   gpc1_1 gpc821 (
      {stage1_1[139]},
      {stage2_1[42]}
   );
   gpc1_1 gpc822 (
      {stage1_1[140]},
      {stage2_1[43]}
   );
   gpc1_1 gpc823 (
      {stage1_1[141]},
      {stage2_1[44]}
   );
   gpc1_1 gpc824 (
      {stage1_1[142]},
      {stage2_1[45]}
   );
   gpc1_1 gpc825 (
      {stage1_1[143]},
      {stage2_1[46]}
   );
   gpc1_1 gpc826 (
      {stage1_1[144]},
      {stage2_1[47]}
   );
   gpc1_1 gpc827 (
      {stage1_1[145]},
      {stage2_1[48]}
   );
   gpc1_1 gpc828 (
      {stage1_1[146]},
      {stage2_1[49]}
   );
   gpc1_1 gpc829 (
      {stage1_1[147]},
      {stage2_1[50]}
   );
   gpc1_1 gpc830 (
      {stage1_1[148]},
      {stage2_1[51]}
   );
   gpc1_1 gpc831 (
      {stage1_1[149]},
      {stage2_1[52]}
   );
   gpc1_1 gpc832 (
      {stage1_1[150]},
      {stage2_1[53]}
   );
   gpc1_1 gpc833 (
      {stage1_1[151]},
      {stage2_1[54]}
   );
   gpc1_1 gpc834 (
      {stage1_1[152]},
      {stage2_1[55]}
   );
   gpc1_1 gpc835 (
      {stage1_1[153]},
      {stage2_1[56]}
   );
   gpc1_1 gpc836 (
      {stage1_1[154]},
      {stage2_1[57]}
   );
   gpc1_1 gpc837 (
      {stage1_4[240]},
      {stage2_4[88]}
   );
   gpc1_1 gpc838 (
      {stage1_5[228]},
      {stage2_5[73]}
   );
   gpc1_1 gpc839 (
      {stage1_5[229]},
      {stage2_5[74]}
   );
   gpc1_1 gpc840 (
      {stage1_9[234]},
      {stage2_9[85]}
   );
   gpc1_1 gpc841 (
      {stage1_9[235]},
      {stage2_9[86]}
   );
   gpc1_1 gpc842 (
      {stage1_9[236]},
      {stage2_9[87]}
   );
   gpc1_1 gpc843 (
      {stage1_9[237]},
      {stage2_9[88]}
   );
   gpc1_1 gpc844 (
      {stage1_9[238]},
      {stage2_9[89]}
   );
   gpc1_1 gpc845 (
      {stage1_9[239]},
      {stage2_9[90]}
   );
   gpc1_1 gpc846 (
      {stage1_9[240]},
      {stage2_9[91]}
   );
   gpc1_1 gpc847 (
      {stage1_10[173]},
      {stage2_10[92]}
   );
   gpc1_1 gpc848 (
      {stage1_10[174]},
      {stage2_10[93]}
   );
   gpc1_1 gpc849 (
      {stage1_10[175]},
      {stage2_10[94]}
   );
   gpc1_1 gpc850 (
      {stage1_10[176]},
      {stage2_10[95]}
   );
   gpc1_1 gpc851 (
      {stage1_10[177]},
      {stage2_10[96]}
   );
   gpc1_1 gpc852 (
      {stage1_10[178]},
      {stage2_10[97]}
   );
   gpc1_1 gpc853 (
      {stage1_10[179]},
      {stage2_10[98]}
   );
   gpc1_1 gpc854 (
      {stage1_11[168]},
      {stage2_11[79]}
   );
   gpc1_1 gpc855 (
      {stage1_11[169]},
      {stage2_11[80]}
   );
   gpc1_1 gpc856 (
      {stage1_11[170]},
      {stage2_11[81]}
   );
   gpc1_1 gpc857 (
      {stage1_12[102]},
      {stage2_12[57]}
   );
   gpc1_1 gpc858 (
      {stage1_12[103]},
      {stage2_12[58]}
   );
   gpc1_1 gpc859 (
      {stage1_12[104]},
      {stage2_12[59]}
   );
   gpc1_1 gpc860 (
      {stage1_12[105]},
      {stage2_12[60]}
   );
   gpc1_1 gpc861 (
      {stage1_12[106]},
      {stage2_12[61]}
   );
   gpc1_1 gpc862 (
      {stage1_12[107]},
      {stage2_12[62]}
   );
   gpc1_1 gpc863 (
      {stage1_12[108]},
      {stage2_12[63]}
   );
   gpc1_1 gpc864 (
      {stage1_12[109]},
      {stage2_12[64]}
   );
   gpc1_1 gpc865 (
      {stage1_12[110]},
      {stage2_12[65]}
   );
   gpc1_1 gpc866 (
      {stage1_12[111]},
      {stage2_12[66]}
   );
   gpc1_1 gpc867 (
      {stage1_12[112]},
      {stage2_12[67]}
   );
   gpc1_1 gpc868 (
      {stage1_12[113]},
      {stage2_12[68]}
   );
   gpc1_1 gpc869 (
      {stage1_12[114]},
      {stage2_12[69]}
   );
   gpc1_1 gpc870 (
      {stage1_12[115]},
      {stage2_12[70]}
   );
   gpc1_1 gpc871 (
      {stage1_12[116]},
      {stage2_12[71]}
   );
   gpc1_1 gpc872 (
      {stage1_12[117]},
      {stage2_12[72]}
   );
   gpc1_1 gpc873 (
      {stage1_12[118]},
      {stage2_12[73]}
   );
   gpc1_1 gpc874 (
      {stage1_12[119]},
      {stage2_12[74]}
   );
   gpc1_1 gpc875 (
      {stage1_12[120]},
      {stage2_12[75]}
   );
   gpc1_1 gpc876 (
      {stage1_12[121]},
      {stage2_12[76]}
   );
   gpc1_1 gpc877 (
      {stage1_12[122]},
      {stage2_12[77]}
   );
   gpc1_1 gpc878 (
      {stage1_12[123]},
      {stage2_12[78]}
   );
   gpc1_1 gpc879 (
      {stage1_12[124]},
      {stage2_12[79]}
   );
   gpc1_1 gpc880 (
      {stage1_12[125]},
      {stage2_12[80]}
   );
   gpc1_1 gpc881 (
      {stage1_12[126]},
      {stage2_12[81]}
   );
   gpc1_1 gpc882 (
      {stage1_12[127]},
      {stage2_12[82]}
   );
   gpc1_1 gpc883 (
      {stage1_12[128]},
      {stage2_12[83]}
   );
   gpc1_1 gpc884 (
      {stage1_12[129]},
      {stage2_12[84]}
   );
   gpc1_1 gpc885 (
      {stage1_12[130]},
      {stage2_12[85]}
   );
   gpc1_1 gpc886 (
      {stage1_12[131]},
      {stage2_12[86]}
   );
   gpc1_1 gpc887 (
      {stage1_12[132]},
      {stage2_12[87]}
   );
   gpc1_1 gpc888 (
      {stage1_12[133]},
      {stage2_12[88]}
   );
   gpc1_1 gpc889 (
      {stage1_12[134]},
      {stage2_12[89]}
   );
   gpc1_1 gpc890 (
      {stage1_12[135]},
      {stage2_12[90]}
   );
   gpc1_1 gpc891 (
      {stage1_12[136]},
      {stage2_12[91]}
   );
   gpc1_1 gpc892 (
      {stage1_12[137]},
      {stage2_12[92]}
   );
   gpc1_1 gpc893 (
      {stage1_12[138]},
      {stage2_12[93]}
   );
   gpc1_1 gpc894 (
      {stage1_12[139]},
      {stage2_12[94]}
   );
   gpc1_1 gpc895 (
      {stage1_12[140]},
      {stage2_12[95]}
   );
   gpc1_1 gpc896 (
      {stage1_12[141]},
      {stage2_12[96]}
   );
   gpc1_1 gpc897 (
      {stage1_12[142]},
      {stage2_12[97]}
   );
   gpc1_1 gpc898 (
      {stage1_12[143]},
      {stage2_12[98]}
   );
   gpc1_1 gpc899 (
      {stage1_12[144]},
      {stage2_12[99]}
   );
   gpc1_1 gpc900 (
      {stage1_12[145]},
      {stage2_12[100]}
   );
   gpc1_1 gpc901 (
      {stage1_12[146]},
      {stage2_12[101]}
   );
   gpc1_1 gpc902 (
      {stage1_12[147]},
      {stage2_12[102]}
   );
   gpc1_1 gpc903 (
      {stage1_12[148]},
      {stage2_12[103]}
   );
   gpc1_1 gpc904 (
      {stage1_12[149]},
      {stage2_12[104]}
   );
   gpc1_1 gpc905 (
      {stage1_12[150]},
      {stage2_12[105]}
   );
   gpc1_1 gpc906 (
      {stage1_12[151]},
      {stage2_12[106]}
   );
   gpc1_1 gpc907 (
      {stage1_12[152]},
      {stage2_12[107]}
   );
   gpc1_1 gpc908 (
      {stage1_12[153]},
      {stage2_12[108]}
   );
   gpc1_1 gpc909 (
      {stage1_12[154]},
      {stage2_12[109]}
   );
   gpc1_1 gpc910 (
      {stage1_12[155]},
      {stage2_12[110]}
   );
   gpc1_1 gpc911 (
      {stage1_12[156]},
      {stage2_12[111]}
   );
   gpc1_1 gpc912 (
      {stage1_13[72]},
      {stage2_13[45]}
   );
   gpc1_1 gpc913 (
      {stage1_13[73]},
      {stage2_13[46]}
   );
   gpc1_1 gpc914 (
      {stage1_13[74]},
      {stage2_13[47]}
   );
   gpc1_1 gpc915 (
      {stage1_13[75]},
      {stage2_13[48]}
   );
   gpc1_1 gpc916 (
      {stage1_13[76]},
      {stage2_13[49]}
   );
   gpc1_1 gpc917 (
      {stage1_13[77]},
      {stage2_13[50]}
   );
   gpc1_1 gpc918 (
      {stage1_13[78]},
      {stage2_13[51]}
   );
   gpc1163_5 gpc919 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc920 (
      {stage2_0[3], stage2_0[4], stage2_0[5], stage2_0[6], stage2_0[7], stage2_0[8]},
      {stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc606_5 gpc921 (
      {stage2_0[9], stage2_0[10], stage2_0[11], stage2_0[12], stage2_0[13], stage2_0[14]},
      {stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11], stage2_2[12]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc606_5 gpc922 (
      {stage2_0[15], stage2_0[16], stage2_0[17], stage2_0[18], stage2_0[19], stage2_0[20]},
      {stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17], stage2_2[18]},
      {stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3],stage3_0[3]}
   );
   gpc606_5 gpc923 (
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5], stage2_3[6]},
      {stage3_5[0],stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4]}
   );
   gpc606_5 gpc924 (
      {stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15], stage2_1[16], stage2_1[17]},
      {stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11], stage2_3[12]},
      {stage3_5[1],stage3_4[5],stage3_3[5],stage3_2[5],stage3_1[5]}
   );
   gpc606_5 gpc925 (
      {stage2_1[18], stage2_1[19], stage2_1[20], stage2_1[21], stage2_1[22], stage2_1[23]},
      {stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17], stage2_3[18]},
      {stage3_5[2],stage3_4[6],stage3_3[6],stage3_2[6],stage3_1[6]}
   );
   gpc606_5 gpc926 (
      {stage2_1[24], stage2_1[25], stage2_1[26], stage2_1[27], stage2_1[28], stage2_1[29]},
      {stage2_3[19], stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23], stage2_3[24]},
      {stage3_5[3],stage3_4[7],stage3_3[7],stage3_2[7],stage3_1[7]}
   );
   gpc606_5 gpc927 (
      {stage2_1[30], stage2_1[31], stage2_1[32], stage2_1[33], stage2_1[34], stage2_1[35]},
      {stage2_3[25], stage2_3[26], stage2_3[27], stage2_3[28], stage2_3[29], stage2_3[30]},
      {stage3_5[4],stage3_4[8],stage3_3[8],stage3_2[8],stage3_1[8]}
   );
   gpc606_5 gpc928 (
      {stage2_1[36], stage2_1[37], stage2_1[38], stage2_1[39], stage2_1[40], stage2_1[41]},
      {stage2_3[31], stage2_3[32], stage2_3[33], stage2_3[34], stage2_3[35], stage2_3[36]},
      {stage3_5[5],stage3_4[9],stage3_3[9],stage3_2[9],stage3_1[9]}
   );
   gpc615_5 gpc929 (
      {stage2_2[19], stage2_2[20], stage2_2[21], stage2_2[22], stage2_2[23]},
      {stage2_3[37]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[6],stage3_4[10],stage3_3[10],stage3_2[10]}
   );
   gpc615_5 gpc930 (
      {stage2_2[24], stage2_2[25], stage2_2[26], stage2_2[27], stage2_2[28]},
      {stage2_3[38]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[7],stage3_4[11],stage3_3[11],stage3_2[11]}
   );
   gpc615_5 gpc931 (
      {stage2_2[29], stage2_2[30], stage2_2[31], stage2_2[32], stage2_2[33]},
      {stage2_3[39]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage3_6[2],stage3_5[8],stage3_4[12],stage3_3[12],stage3_2[12]}
   );
   gpc615_5 gpc932 (
      {stage2_2[34], stage2_2[35], stage2_2[36], stage2_2[37], stage2_2[38]},
      {stage2_3[40]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage3_6[3],stage3_5[9],stage3_4[13],stage3_3[13],stage3_2[13]}
   );
   gpc615_5 gpc933 (
      {stage2_2[39], stage2_2[40], stage2_2[41], stage2_2[42], stage2_2[43]},
      {stage2_3[41]},
      {stage2_4[24], stage2_4[25], stage2_4[26], stage2_4[27], stage2_4[28], stage2_4[29]},
      {stage3_6[4],stage3_5[10],stage3_4[14],stage3_3[14],stage3_2[14]}
   );
   gpc615_5 gpc934 (
      {stage2_2[44], stage2_2[45], stage2_2[46], stage2_2[47], stage2_2[48]},
      {stage2_3[42]},
      {stage2_4[30], stage2_4[31], stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35]},
      {stage3_6[5],stage3_5[11],stage3_4[15],stage3_3[15],stage3_2[15]}
   );
   gpc615_5 gpc935 (
      {stage2_2[49], stage2_2[50], stage2_2[51], stage2_2[52], stage2_2[53]},
      {stage2_3[43]},
      {stage2_4[36], stage2_4[37], stage2_4[38], stage2_4[39], stage2_4[40], stage2_4[41]},
      {stage3_6[6],stage3_5[12],stage3_4[16],stage3_3[16],stage3_2[16]}
   );
   gpc615_5 gpc936 (
      {stage2_3[44], stage2_3[45], stage2_3[46], stage2_3[47], stage2_3[48]},
      {stage2_4[42]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[7],stage3_5[13],stage3_4[17],stage3_3[17]}
   );
   gpc615_5 gpc937 (
      {stage2_3[49], stage2_3[50], stage2_3[51], stage2_3[52], stage2_3[53]},
      {stage2_4[43]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[8],stage3_5[14],stage3_4[18],stage3_3[18]}
   );
   gpc615_5 gpc938 (
      {stage2_3[54], stage2_3[55], stage2_3[56], stage2_3[57], stage2_3[58]},
      {stage2_4[44]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[9],stage3_5[15],stage3_4[19],stage3_3[19]}
   );
   gpc615_5 gpc939 (
      {stage2_3[59], stage2_3[60], stage2_3[61], stage2_3[62], stage2_3[63]},
      {stage2_4[45]},
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage3_7[3],stage3_6[10],stage3_5[16],stage3_4[20],stage3_3[20]}
   );
   gpc615_5 gpc940 (
      {stage2_3[64], stage2_3[65], stage2_3[66], stage2_3[67], stage2_3[68]},
      {stage2_4[46]},
      {stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29]},
      {stage3_7[4],stage3_6[11],stage3_5[17],stage3_4[21],stage3_3[21]}
   );
   gpc615_5 gpc941 (
      {stage2_3[69], stage2_3[70], stage2_3[71], stage2_3[72], stage2_3[73]},
      {stage2_4[47]},
      {stage2_5[30], stage2_5[31], stage2_5[32], stage2_5[33], stage2_5[34], stage2_5[35]},
      {stage3_7[5],stage3_6[12],stage3_5[18],stage3_4[22],stage3_3[22]}
   );
   gpc615_5 gpc942 (
      {stage2_3[74], stage2_3[75], stage2_3[76], stage2_3[77], stage2_3[78]},
      {stage2_4[48]},
      {stage2_5[36], stage2_5[37], stage2_5[38], stage2_5[39], stage2_5[40], stage2_5[41]},
      {stage3_7[6],stage3_6[13],stage3_5[19],stage3_4[23],stage3_3[23]}
   );
   gpc615_5 gpc943 (
      {stage2_3[79], stage2_3[80], stage2_3[81], stage2_3[82], stage2_3[83]},
      {stage2_4[49]},
      {stage2_5[42], stage2_5[43], stage2_5[44], stage2_5[45], stage2_5[46], stage2_5[47]},
      {stage3_7[7],stage3_6[14],stage3_5[20],stage3_4[24],stage3_3[24]}
   );
   gpc606_5 gpc944 (
      {stage2_4[50], stage2_4[51], stage2_4[52], stage2_4[53], stage2_4[54], stage2_4[55]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[8],stage3_6[15],stage3_5[21],stage3_4[25]}
   );
   gpc606_5 gpc945 (
      {stage2_4[56], stage2_4[57], stage2_4[58], stage2_4[59], stage2_4[60], stage2_4[61]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[9],stage3_6[16],stage3_5[22],stage3_4[26]}
   );
   gpc606_5 gpc946 (
      {stage2_4[62], stage2_4[63], stage2_4[64], stage2_4[65], stage2_4[66], stage2_4[67]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[10],stage3_6[17],stage3_5[23],stage3_4[27]}
   );
   gpc606_5 gpc947 (
      {stage2_4[68], stage2_4[69], stage2_4[70], stage2_4[71], stage2_4[72], stage2_4[73]},
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage3_8[3],stage3_7[11],stage3_6[18],stage3_5[24],stage3_4[28]}
   );
   gpc606_5 gpc948 (
      {stage2_4[74], stage2_4[75], stage2_4[76], stage2_4[77], stage2_4[78], stage2_4[79]},
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29]},
      {stage3_8[4],stage3_7[12],stage3_6[19],stage3_5[25],stage3_4[29]}
   );
   gpc606_5 gpc949 (
      {stage2_4[80], stage2_4[81], stage2_4[82], stage2_4[83], stage2_4[84], stage2_4[85]},
      {stage2_6[30], stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage3_8[5],stage3_7[13],stage3_6[20],stage3_5[26],stage3_4[30]}
   );
   gpc606_5 gpc950 (
      {stage2_5[48], stage2_5[49], stage2_5[50], stage2_5[51], stage2_5[52], stage2_5[53]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[6],stage3_7[14],stage3_6[21],stage3_5[27]}
   );
   gpc606_5 gpc951 (
      {stage2_5[54], stage2_5[55], stage2_5[56], stage2_5[57], stage2_5[58], stage2_5[59]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[7],stage3_7[15],stage3_6[22],stage3_5[28]}
   );
   gpc615_5 gpc952 (
      {stage2_5[60], stage2_5[61], stage2_5[62], stage2_5[63], stage2_5[64]},
      {stage2_6[36]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[8],stage3_7[16],stage3_6[23],stage3_5[29]}
   );
   gpc615_5 gpc953 (
      {stage2_5[65], stage2_5[66], stage2_5[67], stage2_5[68], stage2_5[69]},
      {stage2_6[37]},
      {stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage3_9[3],stage3_8[9],stage3_7[17],stage3_6[24],stage3_5[30]}
   );
   gpc615_5 gpc954 (
      {stage2_5[70], stage2_5[71], stage2_5[72], stage2_5[73], stage2_5[74]},
      {stage2_6[38]},
      {stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27], stage2_7[28], stage2_7[29]},
      {stage3_9[4],stage3_8[10],stage3_7[18],stage3_6[25],stage3_5[31]}
   );
   gpc615_5 gpc955 (
      {stage2_6[39], stage2_6[40], stage2_6[41], stage2_6[42], stage2_6[43]},
      {stage2_7[30]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[5],stage3_8[11],stage3_7[19],stage3_6[26]}
   );
   gpc615_5 gpc956 (
      {stage2_6[44], stage2_6[45], stage2_6[46], stage2_6[47], stage2_6[48]},
      {stage2_7[31]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[6],stage3_8[12],stage3_7[20],stage3_6[27]}
   );
   gpc615_5 gpc957 (
      {stage2_6[49], stage2_6[50], stage2_6[51], stage2_6[52], stage2_6[53]},
      {stage2_7[32]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[7],stage3_8[13],stage3_7[21],stage3_6[28]}
   );
   gpc615_5 gpc958 (
      {stage2_6[54], stage2_6[55], stage2_6[56], stage2_6[57], stage2_6[58]},
      {stage2_7[33]},
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23]},
      {stage3_10[3],stage3_9[8],stage3_8[14],stage3_7[22],stage3_6[29]}
   );
   gpc615_5 gpc959 (
      {stage2_6[59], stage2_6[60], stage2_6[61], stage2_6[62], stage2_6[63]},
      {stage2_7[34]},
      {stage2_8[24], stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29]},
      {stage3_10[4],stage3_9[9],stage3_8[15],stage3_7[23],stage3_6[30]}
   );
   gpc615_5 gpc960 (
      {stage2_6[64], stage2_6[65], stage2_6[66], stage2_6[67], stage2_6[68]},
      {stage2_7[35]},
      {stage2_8[30], stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35]},
      {stage3_10[5],stage3_9[10],stage3_8[16],stage3_7[24],stage3_6[31]}
   );
   gpc615_5 gpc961 (
      {stage2_6[69], stage2_6[70], stage2_6[71], stage2_6[72], stage2_6[73]},
      {stage2_7[36]},
      {stage2_8[36], stage2_8[37], stage2_8[38], stage2_8[39], stage2_8[40], stage2_8[41]},
      {stage3_10[6],stage3_9[11],stage3_8[17],stage3_7[25],stage3_6[32]}
   );
   gpc615_5 gpc962 (
      {stage2_6[74], stage2_6[75], stage2_6[76], stage2_6[77], stage2_6[78]},
      {stage2_7[37]},
      {stage2_8[42], stage2_8[43], stage2_8[44], stage2_8[45], stage2_8[46], stage2_8[47]},
      {stage3_10[7],stage3_9[12],stage3_8[18],stage3_7[26],stage3_6[33]}
   );
   gpc615_5 gpc963 (
      {stage2_6[79], stage2_6[80], stage2_6[81], stage2_6[82], stage2_6[83]},
      {stage2_7[38]},
      {stage2_8[48], stage2_8[49], stage2_8[50], stage2_8[51], stage2_8[52], stage2_8[53]},
      {stage3_10[8],stage3_9[13],stage3_8[19],stage3_7[27],stage3_6[34]}
   );
   gpc615_5 gpc964 (
      {stage2_6[84], stage2_6[85], stage2_6[86], stage2_6[87], stage2_6[88]},
      {stage2_7[39]},
      {stage2_8[54], stage2_8[55], stage2_8[56], stage2_8[57], stage2_8[58], stage2_8[59]},
      {stage3_10[9],stage3_9[14],stage3_8[20],stage3_7[28],stage3_6[35]}
   );
   gpc606_5 gpc965 (
      {stage2_7[40], stage2_7[41], stage2_7[42], stage2_7[43], stage2_7[44], stage2_7[45]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[10],stage3_9[15],stage3_8[21],stage3_7[29]}
   );
   gpc606_5 gpc966 (
      {stage2_7[46], stage2_7[47], stage2_7[48], stage2_7[49], stage2_7[50], stage2_7[51]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[11],stage3_9[16],stage3_8[22],stage3_7[30]}
   );
   gpc606_5 gpc967 (
      {stage2_7[52], stage2_7[53], stage2_7[54], stage2_7[55], stage2_7[56], stage2_7[57]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[12],stage3_9[17],stage3_8[23],stage3_7[31]}
   );
   gpc606_5 gpc968 (
      {stage2_7[58], stage2_7[59], stage2_7[60], stage2_7[61], stage2_7[62], stage2_7[63]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[13],stage3_9[18],stage3_8[24],stage3_7[32]}
   );
   gpc615_5 gpc969 (
      {stage2_7[64], stage2_7[65], stage2_7[66], stage2_7[67], stage2_7[68]},
      {stage2_8[60]},
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage3_11[4],stage3_10[14],stage3_9[19],stage3_8[25],stage3_7[33]}
   );
   gpc615_5 gpc970 (
      {stage2_7[69], stage2_7[70], stage2_7[71], stage2_7[72], stage2_7[73]},
      {stage2_8[61]},
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage3_11[5],stage3_10[15],stage3_9[20],stage3_8[26],stage3_7[34]}
   );
   gpc615_5 gpc971 (
      {stage2_7[74], stage2_7[75], stage2_7[76], stage2_7[77], stage2_7[78]},
      {stage2_8[62]},
      {stage2_9[36], stage2_9[37], stage2_9[38], stage2_9[39], stage2_9[40], stage2_9[41]},
      {stage3_11[6],stage3_10[16],stage3_9[21],stage3_8[27],stage3_7[35]}
   );
   gpc615_5 gpc972 (
      {stage2_7[79], stage2_7[80], stage2_7[81], stage2_7[82], stage2_7[83]},
      {stage2_8[63]},
      {stage2_9[42], stage2_9[43], stage2_9[44], stage2_9[45], stage2_9[46], stage2_9[47]},
      {stage3_11[7],stage3_10[17],stage3_9[22],stage3_8[28],stage3_7[36]}
   );
   gpc615_5 gpc973 (
      {stage2_7[84], stage2_7[85], stage2_7[86], stage2_7[87], stage2_7[88]},
      {stage2_8[64]},
      {stage2_9[48], stage2_9[49], stage2_9[50], stage2_9[51], stage2_9[52], stage2_9[53]},
      {stage3_11[8],stage3_10[18],stage3_9[23],stage3_8[29],stage3_7[37]}
   );
   gpc606_5 gpc974 (
      {stage2_8[65], stage2_8[66], stage2_8[67], stage2_8[68], stage2_8[69], stage2_8[70]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[9],stage3_10[19],stage3_9[24],stage3_8[30]}
   );
   gpc1163_5 gpc975 (
      {stage2_9[54], stage2_9[55], stage2_9[56]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage2_11[0]},
      {stage2_12[0]},
      {stage3_13[0],stage3_12[1],stage3_11[10],stage3_10[20],stage3_9[25]}
   );
   gpc1163_5 gpc976 (
      {stage2_9[57], stage2_9[58], stage2_9[59]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage2_11[1]},
      {stage2_12[1]},
      {stage3_13[1],stage3_12[2],stage3_11[11],stage3_10[21],stage3_9[26]}
   );
   gpc1163_5 gpc977 (
      {stage2_9[60], stage2_9[61], stage2_9[62]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage2_11[2]},
      {stage2_12[2]},
      {stage3_13[2],stage3_12[3],stage3_11[12],stage3_10[22],stage3_9[27]}
   );
   gpc1163_5 gpc978 (
      {stage2_9[63], stage2_9[64], stage2_9[65]},
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage2_11[3]},
      {stage2_12[3]},
      {stage3_13[3],stage3_12[4],stage3_11[13],stage3_10[23],stage3_9[28]}
   );
   gpc615_5 gpc979 (
      {stage2_9[66], stage2_9[67], stage2_9[68], stage2_9[69], stage2_9[70]},
      {stage2_10[30]},
      {stage2_11[4], stage2_11[5], stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9]},
      {stage3_13[4],stage3_12[5],stage3_11[14],stage3_10[24],stage3_9[29]}
   );
   gpc615_5 gpc980 (
      {stage2_9[71], stage2_9[72], stage2_9[73], stage2_9[74], stage2_9[75]},
      {stage2_10[31]},
      {stage2_11[10], stage2_11[11], stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15]},
      {stage3_13[5],stage3_12[6],stage3_11[15],stage3_10[25],stage3_9[30]}
   );
   gpc615_5 gpc981 (
      {stage2_9[76], stage2_9[77], stage2_9[78], stage2_9[79], stage2_9[80]},
      {stage2_10[32]},
      {stage2_11[16], stage2_11[17], stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21]},
      {stage3_13[6],stage3_12[7],stage3_11[16],stage3_10[26],stage3_9[31]}
   );
   gpc606_5 gpc982 (
      {stage2_10[33], stage2_10[34], stage2_10[35], stage2_10[36], stage2_10[37], stage2_10[38]},
      {stage2_12[4], stage2_12[5], stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9]},
      {stage3_14[0],stage3_13[7],stage3_12[8],stage3_11[17],stage3_10[27]}
   );
   gpc606_5 gpc983 (
      {stage2_10[39], stage2_10[40], stage2_10[41], stage2_10[42], stage2_10[43], stage2_10[44]},
      {stage2_12[10], stage2_12[11], stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15]},
      {stage3_14[1],stage3_13[8],stage3_12[9],stage3_11[18],stage3_10[28]}
   );
   gpc606_5 gpc984 (
      {stage2_10[45], stage2_10[46], stage2_10[47], stage2_10[48], stage2_10[49], stage2_10[50]},
      {stage2_12[16], stage2_12[17], stage2_12[18], stage2_12[19], stage2_12[20], stage2_12[21]},
      {stage3_14[2],stage3_13[9],stage3_12[10],stage3_11[19],stage3_10[29]}
   );
   gpc606_5 gpc985 (
      {stage2_10[51], stage2_10[52], stage2_10[53], stage2_10[54], stage2_10[55], stage2_10[56]},
      {stage2_12[22], stage2_12[23], stage2_12[24], stage2_12[25], stage2_12[26], stage2_12[27]},
      {stage3_14[3],stage3_13[10],stage3_12[11],stage3_11[20],stage3_10[30]}
   );
   gpc606_5 gpc986 (
      {stage2_10[57], stage2_10[58], stage2_10[59], stage2_10[60], stage2_10[61], stage2_10[62]},
      {stage2_12[28], stage2_12[29], stage2_12[30], stage2_12[31], stage2_12[32], stage2_12[33]},
      {stage3_14[4],stage3_13[11],stage3_12[12],stage3_11[21],stage3_10[31]}
   );
   gpc606_5 gpc987 (
      {stage2_10[63], stage2_10[64], stage2_10[65], stage2_10[66], stage2_10[67], stage2_10[68]},
      {stage2_12[34], stage2_12[35], stage2_12[36], stage2_12[37], stage2_12[38], stage2_12[39]},
      {stage3_14[5],stage3_13[12],stage3_12[13],stage3_11[22],stage3_10[32]}
   );
   gpc606_5 gpc988 (
      {stage2_10[69], stage2_10[70], stage2_10[71], stage2_10[72], stage2_10[73], stage2_10[74]},
      {stage2_12[40], stage2_12[41], stage2_12[42], stage2_12[43], stage2_12[44], stage2_12[45]},
      {stage3_14[6],stage3_13[13],stage3_12[14],stage3_11[23],stage3_10[33]}
   );
   gpc606_5 gpc989 (
      {stage2_10[75], stage2_10[76], stage2_10[77], stage2_10[78], stage2_10[79], stage2_10[80]},
      {stage2_12[46], stage2_12[47], stage2_12[48], stage2_12[49], stage2_12[50], stage2_12[51]},
      {stage3_14[7],stage3_13[14],stage3_12[15],stage3_11[24],stage3_10[34]}
   );
   gpc606_5 gpc990 (
      {stage2_10[81], stage2_10[82], stage2_10[83], stage2_10[84], stage2_10[85], stage2_10[86]},
      {stage2_12[52], stage2_12[53], stage2_12[54], stage2_12[55], stage2_12[56], stage2_12[57]},
      {stage3_14[8],stage3_13[15],stage3_12[16],stage3_11[25],stage3_10[35]}
   );
   gpc606_5 gpc991 (
      {stage2_10[87], stage2_10[88], stage2_10[89], stage2_10[90], stage2_10[91], stage2_10[92]},
      {stage2_12[58], stage2_12[59], stage2_12[60], stage2_12[61], stage2_12[62], stage2_12[63]},
      {stage3_14[9],stage3_13[16],stage3_12[17],stage3_11[26],stage3_10[36]}
   );
   gpc606_5 gpc992 (
      {stage2_10[93], stage2_10[94], stage2_10[95], stage2_10[96], stage2_10[97], stage2_10[98]},
      {stage2_12[64], stage2_12[65], stage2_12[66], stage2_12[67], stage2_12[68], stage2_12[69]},
      {stage3_14[10],stage3_13[17],stage3_12[18],stage3_11[27],stage3_10[37]}
   );
   gpc606_5 gpc993 (
      {stage2_11[22], stage2_11[23], stage2_11[24], stage2_11[25], stage2_11[26], stage2_11[27]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[11],stage3_13[18],stage3_12[19],stage3_11[28]}
   );
   gpc606_5 gpc994 (
      {stage2_11[28], stage2_11[29], stage2_11[30], stage2_11[31], stage2_11[32], stage2_11[33]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[12],stage3_13[19],stage3_12[20],stage3_11[29]}
   );
   gpc606_5 gpc995 (
      {stage2_11[34], stage2_11[35], stage2_11[36], stage2_11[37], stage2_11[38], stage2_11[39]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[13],stage3_13[20],stage3_12[21],stage3_11[30]}
   );
   gpc606_5 gpc996 (
      {stage2_11[40], stage2_11[41], stage2_11[42], stage2_11[43], stage2_11[44], stage2_11[45]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[14],stage3_13[21],stage3_12[22],stage3_11[31]}
   );
   gpc606_5 gpc997 (
      {stage2_11[46], stage2_11[47], stage2_11[48], stage2_11[49], stage2_11[50], stage2_11[51]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[15],stage3_13[22],stage3_12[23],stage3_11[32]}
   );
   gpc606_5 gpc998 (
      {stage2_11[52], stage2_11[53], stage2_11[54], stage2_11[55], stage2_11[56], stage2_11[57]},
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage3_15[5],stage3_14[16],stage3_13[23],stage3_12[24],stage3_11[33]}
   );
   gpc615_5 gpc999 (
      {stage2_11[58], stage2_11[59], stage2_11[60], stage2_11[61], stage2_11[62]},
      {stage2_12[70]},
      {stage2_13[36], stage2_13[37], stage2_13[38], stage2_13[39], stage2_13[40], stage2_13[41]},
      {stage3_15[6],stage3_14[17],stage3_13[24],stage3_12[25],stage3_11[34]}
   );
   gpc606_5 gpc1000 (
      {stage2_12[71], stage2_12[72], stage2_12[73], stage2_12[74], stage2_12[75], stage2_12[76]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[7],stage3_14[18],stage3_13[25],stage3_12[26]}
   );
   gpc606_5 gpc1001 (
      {stage2_12[77], stage2_12[78], stage2_12[79], stage2_12[80], stage2_12[81], stage2_12[82]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[8],stage3_14[19],stage3_13[26],stage3_12[27]}
   );
   gpc606_5 gpc1002 (
      {stage2_12[83], stage2_12[84], stage2_12[85], stage2_12[86], stage2_12[87], stage2_12[88]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[9],stage3_14[20],stage3_13[27],stage3_12[28]}
   );
   gpc606_5 gpc1003 (
      {stage2_12[89], stage2_12[90], stage2_12[91], stage2_12[92], stage2_12[93], stage2_12[94]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[10],stage3_14[21],stage3_13[28],stage3_12[29]}
   );
   gpc606_5 gpc1004 (
      {stage2_13[42], stage2_13[43], stage2_13[44], stage2_13[45], stage2_13[46], stage2_13[47]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[4],stage3_15[11],stage3_14[22],stage3_13[29]}
   );
   gpc1_1 gpc1005 (
      {stage2_0[21]},
      {stage3_0[4]}
   );
   gpc1_1 gpc1006 (
      {stage2_0[22]},
      {stage3_0[5]}
   );
   gpc1_1 gpc1007 (
      {stage2_0[23]},
      {stage3_0[6]}
   );
   gpc1_1 gpc1008 (
      {stage2_0[24]},
      {stage3_0[7]}
   );
   gpc1_1 gpc1009 (
      {stage2_0[25]},
      {stage3_0[8]}
   );
   gpc1_1 gpc1010 (
      {stage2_0[26]},
      {stage3_0[9]}
   );
   gpc1_1 gpc1011 (
      {stage2_0[27]},
      {stage3_0[10]}
   );
   gpc1_1 gpc1012 (
      {stage2_0[28]},
      {stage3_0[11]}
   );
   gpc1_1 gpc1013 (
      {stage2_0[29]},
      {stage3_0[12]}
   );
   gpc1_1 gpc1014 (
      {stage2_0[30]},
      {stage3_0[13]}
   );
   gpc1_1 gpc1015 (
      {stage2_1[42]},
      {stage3_1[10]}
   );
   gpc1_1 gpc1016 (
      {stage2_1[43]},
      {stage3_1[11]}
   );
   gpc1_1 gpc1017 (
      {stage2_1[44]},
      {stage3_1[12]}
   );
   gpc1_1 gpc1018 (
      {stage2_1[45]},
      {stage3_1[13]}
   );
   gpc1_1 gpc1019 (
      {stage2_1[46]},
      {stage3_1[14]}
   );
   gpc1_1 gpc1020 (
      {stage2_1[47]},
      {stage3_1[15]}
   );
   gpc1_1 gpc1021 (
      {stage2_1[48]},
      {stage3_1[16]}
   );
   gpc1_1 gpc1022 (
      {stage2_1[49]},
      {stage3_1[17]}
   );
   gpc1_1 gpc1023 (
      {stage2_1[50]},
      {stage3_1[18]}
   );
   gpc1_1 gpc1024 (
      {stage2_1[51]},
      {stage3_1[19]}
   );
   gpc1_1 gpc1025 (
      {stage2_1[52]},
      {stage3_1[20]}
   );
   gpc1_1 gpc1026 (
      {stage2_1[53]},
      {stage3_1[21]}
   );
   gpc1_1 gpc1027 (
      {stage2_1[54]},
      {stage3_1[22]}
   );
   gpc1_1 gpc1028 (
      {stage2_1[55]},
      {stage3_1[23]}
   );
   gpc1_1 gpc1029 (
      {stage2_1[56]},
      {stage3_1[24]}
   );
   gpc1_1 gpc1030 (
      {stage2_1[57]},
      {stage3_1[25]}
   );
   gpc1_1 gpc1031 (
      {stage2_4[86]},
      {stage3_4[31]}
   );
   gpc1_1 gpc1032 (
      {stage2_4[87]},
      {stage3_4[32]}
   );
   gpc1_1 gpc1033 (
      {stage2_4[88]},
      {stage3_4[33]}
   );
   gpc1_1 gpc1034 (
      {stage2_6[89]},
      {stage3_6[36]}
   );
   gpc1_1 gpc1035 (
      {stage2_6[90]},
      {stage3_6[37]}
   );
   gpc1_1 gpc1036 (
      {stage2_6[91]},
      {stage3_6[38]}
   );
   gpc1_1 gpc1037 (
      {stage2_6[92]},
      {stage3_6[39]}
   );
   gpc1_1 gpc1038 (
      {stage2_6[93]},
      {stage3_6[40]}
   );
   gpc1_1 gpc1039 (
      {stage2_6[94]},
      {stage3_6[41]}
   );
   gpc1_1 gpc1040 (
      {stage2_6[95]},
      {stage3_6[42]}
   );
   gpc1_1 gpc1041 (
      {stage2_6[96]},
      {stage3_6[43]}
   );
   gpc1_1 gpc1042 (
      {stage2_6[97]},
      {stage3_6[44]}
   );
   gpc1_1 gpc1043 (
      {stage2_9[81]},
      {stage3_9[32]}
   );
   gpc1_1 gpc1044 (
      {stage2_9[82]},
      {stage3_9[33]}
   );
   gpc1_1 gpc1045 (
      {stage2_9[83]},
      {stage3_9[34]}
   );
   gpc1_1 gpc1046 (
      {stage2_9[84]},
      {stage3_9[35]}
   );
   gpc1_1 gpc1047 (
      {stage2_9[85]},
      {stage3_9[36]}
   );
   gpc1_1 gpc1048 (
      {stage2_9[86]},
      {stage3_9[37]}
   );
   gpc1_1 gpc1049 (
      {stage2_9[87]},
      {stage3_9[38]}
   );
   gpc1_1 gpc1050 (
      {stage2_9[88]},
      {stage3_9[39]}
   );
   gpc1_1 gpc1051 (
      {stage2_9[89]},
      {stage3_9[40]}
   );
   gpc1_1 gpc1052 (
      {stage2_9[90]},
      {stage3_9[41]}
   );
   gpc1_1 gpc1053 (
      {stage2_9[91]},
      {stage3_9[42]}
   );
   gpc1_1 gpc1054 (
      {stage2_11[63]},
      {stage3_11[35]}
   );
   gpc1_1 gpc1055 (
      {stage2_11[64]},
      {stage3_11[36]}
   );
   gpc1_1 gpc1056 (
      {stage2_11[65]},
      {stage3_11[37]}
   );
   gpc1_1 gpc1057 (
      {stage2_11[66]},
      {stage3_11[38]}
   );
   gpc1_1 gpc1058 (
      {stage2_11[67]},
      {stage3_11[39]}
   );
   gpc1_1 gpc1059 (
      {stage2_11[68]},
      {stage3_11[40]}
   );
   gpc1_1 gpc1060 (
      {stage2_11[69]},
      {stage3_11[41]}
   );
   gpc1_1 gpc1061 (
      {stage2_11[70]},
      {stage3_11[42]}
   );
   gpc1_1 gpc1062 (
      {stage2_11[71]},
      {stage3_11[43]}
   );
   gpc1_1 gpc1063 (
      {stage2_11[72]},
      {stage3_11[44]}
   );
   gpc1_1 gpc1064 (
      {stage2_11[73]},
      {stage3_11[45]}
   );
   gpc1_1 gpc1065 (
      {stage2_11[74]},
      {stage3_11[46]}
   );
   gpc1_1 gpc1066 (
      {stage2_11[75]},
      {stage3_11[47]}
   );
   gpc1_1 gpc1067 (
      {stage2_11[76]},
      {stage3_11[48]}
   );
   gpc1_1 gpc1068 (
      {stage2_11[77]},
      {stage3_11[49]}
   );
   gpc1_1 gpc1069 (
      {stage2_11[78]},
      {stage3_11[50]}
   );
   gpc1_1 gpc1070 (
      {stage2_11[79]},
      {stage3_11[51]}
   );
   gpc1_1 gpc1071 (
      {stage2_11[80]},
      {stage3_11[52]}
   );
   gpc1_1 gpc1072 (
      {stage2_11[81]},
      {stage3_11[53]}
   );
   gpc1_1 gpc1073 (
      {stage2_12[95]},
      {stage3_12[30]}
   );
   gpc1_1 gpc1074 (
      {stage2_12[96]},
      {stage3_12[31]}
   );
   gpc1_1 gpc1075 (
      {stage2_12[97]},
      {stage3_12[32]}
   );
   gpc1_1 gpc1076 (
      {stage2_12[98]},
      {stage3_12[33]}
   );
   gpc1_1 gpc1077 (
      {stage2_12[99]},
      {stage3_12[34]}
   );
   gpc1_1 gpc1078 (
      {stage2_12[100]},
      {stage3_12[35]}
   );
   gpc1_1 gpc1079 (
      {stage2_12[101]},
      {stage3_12[36]}
   );
   gpc1_1 gpc1080 (
      {stage2_12[102]},
      {stage3_12[37]}
   );
   gpc1_1 gpc1081 (
      {stage2_12[103]},
      {stage3_12[38]}
   );
   gpc1_1 gpc1082 (
      {stage2_12[104]},
      {stage3_12[39]}
   );
   gpc1_1 gpc1083 (
      {stage2_12[105]},
      {stage3_12[40]}
   );
   gpc1_1 gpc1084 (
      {stage2_12[106]},
      {stage3_12[41]}
   );
   gpc1_1 gpc1085 (
      {stage2_12[107]},
      {stage3_12[42]}
   );
   gpc1_1 gpc1086 (
      {stage2_12[108]},
      {stage3_12[43]}
   );
   gpc1_1 gpc1087 (
      {stage2_12[109]},
      {stage3_12[44]}
   );
   gpc1_1 gpc1088 (
      {stage2_12[110]},
      {stage3_12[45]}
   );
   gpc1_1 gpc1089 (
      {stage2_12[111]},
      {stage3_12[46]}
   );
   gpc1_1 gpc1090 (
      {stage2_13[48]},
      {stage3_13[30]}
   );
   gpc1_1 gpc1091 (
      {stage2_13[49]},
      {stage3_13[31]}
   );
   gpc1_1 gpc1092 (
      {stage2_13[50]},
      {stage3_13[32]}
   );
   gpc1_1 gpc1093 (
      {stage2_13[51]},
      {stage3_13[33]}
   );
   gpc1_1 gpc1094 (
      {stage2_14[24]},
      {stage3_14[23]}
   );
   gpc1_1 gpc1095 (
      {stage2_14[25]},
      {stage3_14[24]}
   );
   gpc1_1 gpc1096 (
      {stage2_14[26]},
      {stage3_14[25]}
   );
   gpc1_1 gpc1097 (
      {stage2_15[6]},
      {stage3_15[12]}
   );
   gpc1_1 gpc1098 (
      {stage2_15[7]},
      {stage3_15[13]}
   );
   gpc1_1 gpc1099 (
      {stage2_15[8]},
      {stage3_15[14]}
   );
   gpc1_1 gpc1100 (
      {stage2_15[9]},
      {stage3_15[15]}
   );
   gpc1_1 gpc1101 (
      {stage2_15[10]},
      {stage3_15[16]}
   );
   gpc1_1 gpc1102 (
      {stage2_15[11]},
      {stage3_15[17]}
   );
   gpc606_5 gpc1103 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc606_5 gpc1104 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc606_5 gpc1105 (
      {stage3_1[6], stage3_1[7], stage3_1[8], stage3_1[9], stage3_1[10], stage3_1[11]},
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage4_5[1],stage4_4[2],stage4_3[2],stage4_2[2],stage4_1[2]}
   );
   gpc606_5 gpc1106 (
      {stage3_1[12], stage3_1[13], stage3_1[14], stage3_1[15], stage3_1[16], stage3_1[17]},
      {stage3_3[12], stage3_3[13], stage3_3[14], stage3_3[15], stage3_3[16], stage3_3[17]},
      {stage4_5[2],stage4_4[3],stage4_3[3],stage4_2[3],stage4_1[3]}
   );
   gpc615_5 gpc1107 (
      {stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9], stage3_2[10]},
      {stage3_3[18]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[3],stage4_4[4],stage4_3[4],stage4_2[4]}
   );
   gpc615_5 gpc1108 (
      {stage3_2[11], stage3_2[12], stage3_2[13], stage3_2[14], stage3_2[15]},
      {stage3_3[19]},
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage4_6[1],stage4_5[4],stage4_4[5],stage4_3[5],stage4_2[5]}
   );
   gpc615_5 gpc1109 (
      {stage3_3[20], stage3_3[21], stage3_3[22], stage3_3[23], stage3_3[24]},
      {stage3_4[12]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[2],stage4_5[5],stage4_4[6],stage4_3[6]}
   );
   gpc606_5 gpc1110 (
      {stage3_4[13], stage3_4[14], stage3_4[15], stage3_4[16], stage3_4[17], stage3_4[18]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[1],stage4_6[3],stage4_5[6],stage4_4[7]}
   );
   gpc606_5 gpc1111 (
      {stage3_4[19], stage3_4[20], stage3_4[21], stage3_4[22], stage3_4[23], stage3_4[24]},
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10], stage3_6[11]},
      {stage4_8[1],stage4_7[2],stage4_6[4],stage4_5[7],stage4_4[8]}
   );
   gpc606_5 gpc1112 (
      {stage3_4[25], stage3_4[26], stage3_4[27], stage3_4[28], stage3_4[29], stage3_4[30]},
      {stage3_6[12], stage3_6[13], stage3_6[14], stage3_6[15], stage3_6[16], stage3_6[17]},
      {stage4_8[2],stage4_7[3],stage4_6[5],stage4_5[8],stage4_4[9]}
   );
   gpc606_5 gpc1113 (
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[3],stage4_7[4],stage4_6[6],stage4_5[9]}
   );
   gpc606_5 gpc1114 (
      {stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17]},
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage4_9[1],stage4_8[4],stage4_7[5],stage4_6[7],stage4_5[10]}
   );
   gpc606_5 gpc1115 (
      {stage3_5[18], stage3_5[19], stage3_5[20], stage3_5[21], stage3_5[22], stage3_5[23]},
      {stage3_7[12], stage3_7[13], stage3_7[14], stage3_7[15], stage3_7[16], stage3_7[17]},
      {stage4_9[2],stage4_8[5],stage4_7[6],stage4_6[8],stage4_5[11]}
   );
   gpc606_5 gpc1116 (
      {stage3_5[24], stage3_5[25], stage3_5[26], stage3_5[27], stage3_5[28], stage3_5[29]},
      {stage3_7[18], stage3_7[19], stage3_7[20], stage3_7[21], stage3_7[22], stage3_7[23]},
      {stage4_9[3],stage4_8[6],stage4_7[7],stage4_6[9],stage4_5[12]}
   );
   gpc606_5 gpc1117 (
      {stage3_6[18], stage3_6[19], stage3_6[20], stage3_6[21], stage3_6[22], stage3_6[23]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[4],stage4_8[7],stage4_7[8],stage4_6[10]}
   );
   gpc615_5 gpc1118 (
      {stage3_6[24], stage3_6[25], stage3_6[26], stage3_6[27], stage3_6[28]},
      {stage3_7[24]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[5],stage4_8[8],stage4_7[9],stage4_6[11]}
   );
   gpc615_5 gpc1119 (
      {stage3_6[29], stage3_6[30], stage3_6[31], stage3_6[32], stage3_6[33]},
      {stage3_7[25]},
      {stage3_8[12], stage3_8[13], stage3_8[14], stage3_8[15], stage3_8[16], stage3_8[17]},
      {stage4_10[2],stage4_9[6],stage4_8[9],stage4_7[10],stage4_6[12]}
   );
   gpc615_5 gpc1120 (
      {stage3_6[34], stage3_6[35], stage3_6[36], stage3_6[37], stage3_6[38]},
      {stage3_7[26]},
      {stage3_8[18], stage3_8[19], stage3_8[20], stage3_8[21], stage3_8[22], stage3_8[23]},
      {stage4_10[3],stage4_9[7],stage4_8[10],stage4_7[11],stage4_6[13]}
   );
   gpc615_5 gpc1121 (
      {stage3_6[39], stage3_6[40], stage3_6[41], stage3_6[42], stage3_6[43]},
      {stage3_7[27]},
      {stage3_8[24], stage3_8[25], stage3_8[26], stage3_8[27], stage3_8[28], stage3_8[29]},
      {stage4_10[4],stage4_9[8],stage4_8[11],stage4_7[12],stage4_6[14]}
   );
   gpc615_5 gpc1122 (
      {stage3_7[28], stage3_7[29], stage3_7[30], stage3_7[31], stage3_7[32]},
      {stage3_8[30]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[5],stage4_9[9],stage4_8[12],stage4_7[13]}
   );
   gpc606_5 gpc1123 (
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[0],stage4_11[1],stage4_10[6],stage4_9[10]}
   );
   gpc606_5 gpc1124 (
      {stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15], stage3_9[16], stage3_9[17]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[1],stage4_11[2],stage4_10[7],stage4_9[11]}
   );
   gpc606_5 gpc1125 (
      {stage3_9[18], stage3_9[19], stage3_9[20], stage3_9[21], stage3_9[22], stage3_9[23]},
      {stage3_11[12], stage3_11[13], stage3_11[14], stage3_11[15], stage3_11[16], stage3_11[17]},
      {stage4_13[2],stage4_12[2],stage4_11[3],stage4_10[8],stage4_9[12]}
   );
   gpc606_5 gpc1126 (
      {stage3_9[24], stage3_9[25], stage3_9[26], stage3_9[27], stage3_9[28], stage3_9[29]},
      {stage3_11[18], stage3_11[19], stage3_11[20], stage3_11[21], stage3_11[22], stage3_11[23]},
      {stage4_13[3],stage4_12[3],stage4_11[4],stage4_10[9],stage4_9[13]}
   );
   gpc606_5 gpc1127 (
      {stage3_9[30], stage3_9[31], stage3_9[32], stage3_9[33], stage3_9[34], stage3_9[35]},
      {stage3_11[24], stage3_11[25], stage3_11[26], stage3_11[27], stage3_11[28], stage3_11[29]},
      {stage4_13[4],stage4_12[4],stage4_11[5],stage4_10[10],stage4_9[14]}
   );
   gpc606_5 gpc1128 (
      {stage3_9[36], stage3_9[37], stage3_9[38], stage3_9[39], stage3_9[40], stage3_9[41]},
      {stage3_11[30], stage3_11[31], stage3_11[32], stage3_11[33], stage3_11[34], stage3_11[35]},
      {stage4_13[5],stage4_12[5],stage4_11[6],stage4_10[11],stage4_9[15]}
   );
   gpc2135_5 gpc1129 (
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4]},
      {stage3_11[36], stage3_11[37], stage3_11[38]},
      {stage3_12[0]},
      {stage3_13[0], stage3_13[1]},
      {stage4_14[0],stage4_13[6],stage4_12[6],stage4_11[7],stage4_10[12]}
   );
   gpc2135_5 gpc1130 (
      {stage3_10[5], stage3_10[6], stage3_10[7], stage3_10[8], stage3_10[9]},
      {stage3_11[39], stage3_11[40], stage3_11[41]},
      {stage3_12[1]},
      {stage3_13[2], stage3_13[3]},
      {stage4_14[1],stage4_13[7],stage4_12[7],stage4_11[8],stage4_10[13]}
   );
   gpc2135_5 gpc1131 (
      {stage3_10[10], stage3_10[11], stage3_10[12], stage3_10[13], stage3_10[14]},
      {stage3_11[42], stage3_11[43], stage3_11[44]},
      {stage3_12[2]},
      {stage3_13[4], stage3_13[5]},
      {stage4_14[2],stage4_13[8],stage4_12[8],stage4_11[9],stage4_10[14]}
   );
   gpc2135_5 gpc1132 (
      {stage3_10[15], stage3_10[16], stage3_10[17], stage3_10[18], stage3_10[19]},
      {stage3_11[45], stage3_11[46], stage3_11[47]},
      {stage3_12[3]},
      {stage3_13[6], stage3_13[7]},
      {stage4_14[3],stage4_13[9],stage4_12[9],stage4_11[10],stage4_10[15]}
   );
   gpc606_5 gpc1133 (
      {stage3_10[20], stage3_10[21], stage3_10[22], stage3_10[23], stage3_10[24], stage3_10[25]},
      {stage3_12[4], stage3_12[5], stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9]},
      {stage4_14[4],stage4_13[10],stage4_12[10],stage4_11[11],stage4_10[16]}
   );
   gpc606_5 gpc1134 (
      {stage3_10[26], stage3_10[27], stage3_10[28], stage3_10[29], stage3_10[30], stage3_10[31]},
      {stage3_12[10], stage3_12[11], stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15]},
      {stage4_14[5],stage4_13[11],stage4_12[11],stage4_11[12],stage4_10[17]}
   );
   gpc606_5 gpc1135 (
      {stage3_10[32], stage3_10[33], stage3_10[34], stage3_10[35], stage3_10[36], stage3_10[37]},
      {stage3_12[16], stage3_12[17], stage3_12[18], stage3_12[19], stage3_12[20], stage3_12[21]},
      {stage4_14[6],stage4_13[12],stage4_12[12],stage4_11[13],stage4_10[18]}
   );
   gpc615_5 gpc1136 (
      {stage3_11[48], stage3_11[49], stage3_11[50], stage3_11[51], stage3_11[52]},
      {stage3_12[22]},
      {stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11], stage3_13[12], stage3_13[13]},
      {stage4_15[0],stage4_14[7],stage4_13[13],stage4_12[13],stage4_11[14]}
   );
   gpc606_5 gpc1137 (
      {stage3_12[23], stage3_12[24], stage3_12[25], stage3_12[26], stage3_12[27], stage3_12[28]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[1],stage4_14[8],stage4_13[14],stage4_12[14]}
   );
   gpc606_5 gpc1138 (
      {stage3_12[29], stage3_12[30], stage3_12[31], stage3_12[32], stage3_12[33], stage3_12[34]},
      {stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10], stage3_14[11]},
      {stage4_16[1],stage4_15[2],stage4_14[9],stage4_13[15],stage4_12[15]}
   );
   gpc606_5 gpc1139 (
      {stage3_12[35], stage3_12[36], stage3_12[37], stage3_12[38], stage3_12[39], stage3_12[40]},
      {stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15], stage3_14[16], stage3_14[17]},
      {stage4_16[2],stage4_15[3],stage4_14[10],stage4_13[16],stage4_12[16]}
   );
   gpc606_5 gpc1140 (
      {stage3_12[41], stage3_12[42], stage3_12[43], stage3_12[44], stage3_12[45], stage3_12[46]},
      {stage3_14[18], stage3_14[19], stage3_14[20], stage3_14[21], stage3_14[22], stage3_14[23]},
      {stage4_16[3],stage4_15[4],stage4_14[11],stage4_13[17],stage4_12[17]}
   );
   gpc606_5 gpc1141 (
      {stage3_13[14], stage3_13[15], stage3_13[16], stage3_13[17], stage3_13[18], stage3_13[19]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[4],stage4_15[5],stage4_14[12],stage4_13[18]}
   );
   gpc606_5 gpc1142 (
      {stage3_13[20], stage3_13[21], stage3_13[22], stage3_13[23], stage3_13[24], stage3_13[25]},
      {stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11]},
      {stage4_17[1],stage4_16[5],stage4_15[6],stage4_14[13],stage4_13[19]}
   );
   gpc606_5 gpc1143 (
      {stage3_13[26], stage3_13[27], stage3_13[28], stage3_13[29], stage3_13[30], stage3_13[31]},
      {stage3_15[12], stage3_15[13], stage3_15[14], stage3_15[15], stage3_15[16], stage3_15[17]},
      {stage4_17[2],stage4_16[6],stage4_15[7],stage4_14[14],stage4_13[20]}
   );
   gpc1_1 gpc1144 (
      {stage3_0[6]},
      {stage4_0[1]}
   );
   gpc1_1 gpc1145 (
      {stage3_0[7]},
      {stage4_0[2]}
   );
   gpc1_1 gpc1146 (
      {stage3_0[8]},
      {stage4_0[3]}
   );
   gpc1_1 gpc1147 (
      {stage3_0[9]},
      {stage4_0[4]}
   );
   gpc1_1 gpc1148 (
      {stage3_0[10]},
      {stage4_0[5]}
   );
   gpc1_1 gpc1149 (
      {stage3_0[11]},
      {stage4_0[6]}
   );
   gpc1_1 gpc1150 (
      {stage3_0[12]},
      {stage4_0[7]}
   );
   gpc1_1 gpc1151 (
      {stage3_0[13]},
      {stage4_0[8]}
   );
   gpc1_1 gpc1152 (
      {stage3_1[18]},
      {stage4_1[4]}
   );
   gpc1_1 gpc1153 (
      {stage3_1[19]},
      {stage4_1[5]}
   );
   gpc1_1 gpc1154 (
      {stage3_1[20]},
      {stage4_1[6]}
   );
   gpc1_1 gpc1155 (
      {stage3_1[21]},
      {stage4_1[7]}
   );
   gpc1_1 gpc1156 (
      {stage3_1[22]},
      {stage4_1[8]}
   );
   gpc1_1 gpc1157 (
      {stage3_1[23]},
      {stage4_1[9]}
   );
   gpc1_1 gpc1158 (
      {stage3_1[24]},
      {stage4_1[10]}
   );
   gpc1_1 gpc1159 (
      {stage3_1[25]},
      {stage4_1[11]}
   );
   gpc1_1 gpc1160 (
      {stage3_2[16]},
      {stage4_2[6]}
   );
   gpc1_1 gpc1161 (
      {stage3_4[31]},
      {stage4_4[10]}
   );
   gpc1_1 gpc1162 (
      {stage3_4[32]},
      {stage4_4[11]}
   );
   gpc1_1 gpc1163 (
      {stage3_4[33]},
      {stage4_4[12]}
   );
   gpc1_1 gpc1164 (
      {stage3_5[30]},
      {stage4_5[13]}
   );
   gpc1_1 gpc1165 (
      {stage3_5[31]},
      {stage4_5[14]}
   );
   gpc1_1 gpc1166 (
      {stage3_6[44]},
      {stage4_6[15]}
   );
   gpc1_1 gpc1167 (
      {stage3_7[33]},
      {stage4_7[14]}
   );
   gpc1_1 gpc1168 (
      {stage3_7[34]},
      {stage4_7[15]}
   );
   gpc1_1 gpc1169 (
      {stage3_7[35]},
      {stage4_7[16]}
   );
   gpc1_1 gpc1170 (
      {stage3_7[36]},
      {stage4_7[17]}
   );
   gpc1_1 gpc1171 (
      {stage3_7[37]},
      {stage4_7[18]}
   );
   gpc1_1 gpc1172 (
      {stage3_9[42]},
      {stage4_9[16]}
   );
   gpc1_1 gpc1173 (
      {stage3_11[53]},
      {stage4_11[15]}
   );
   gpc1_1 gpc1174 (
      {stage3_13[32]},
      {stage4_13[21]}
   );
   gpc1_1 gpc1175 (
      {stage3_13[33]},
      {stage4_13[22]}
   );
   gpc1_1 gpc1176 (
      {stage3_14[24]},
      {stage4_14[15]}
   );
   gpc1_1 gpc1177 (
      {stage3_14[25]},
      {stage4_14[16]}
   );
   gpc1_1 gpc1178 (
      {stage3_16[0]},
      {stage4_16[7]}
   );
   gpc1_1 gpc1179 (
      {stage3_16[1]},
      {stage4_16[8]}
   );
   gpc1_1 gpc1180 (
      {stage3_16[2]},
      {stage4_16[9]}
   );
   gpc1_1 gpc1181 (
      {stage3_16[3]},
      {stage4_16[10]}
   );
   gpc1_1 gpc1182 (
      {stage3_16[4]},
      {stage4_16[11]}
   );
   gpc1_1 gpc1183 (
      {stage3_17[0]},
      {stage4_17[3]}
   );
   gpc1163_5 gpc1184 (
      {stage4_0[0], stage4_0[1], stage4_0[2]},
      {stage4_1[0], stage4_1[1], stage4_1[2], stage4_1[3], stage4_1[4], stage4_1[5]},
      {stage4_2[0]},
      {stage4_3[0]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc623_5 gpc1185 (
      {stage4_2[1], stage4_2[2], stage4_2[3]},
      {stage4_3[1], stage4_3[2]},
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5]},
      {stage5_6[0],stage5_5[0],stage5_4[1],stage5_3[1],stage5_2[1]}
   );
   gpc606_5 gpc1186 (
      {stage4_4[6], stage4_4[7], stage4_4[8], stage4_4[9], stage4_4[10], stage4_4[11]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage5_8[0],stage5_7[0],stage5_6[1],stage5_5[1],stage5_4[2]}
   );
   gpc615_5 gpc1187 (
      {stage4_5[0], stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4]},
      {stage4_6[6]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5]},
      {stage5_9[0],stage5_8[1],stage5_7[1],stage5_6[2],stage5_5[2]}
   );
   gpc615_5 gpc1188 (
      {stage4_5[5], stage4_5[6], stage4_5[7], stage4_5[8], stage4_5[9]},
      {stage4_6[7]},
      {stage4_7[6], stage4_7[7], stage4_7[8], stage4_7[9], stage4_7[10], stage4_7[11]},
      {stage5_9[1],stage5_8[2],stage5_7[2],stage5_6[3],stage5_5[3]}
   );
   gpc615_5 gpc1189 (
      {stage4_5[10], stage4_5[11], stage4_5[12], stage4_5[13], stage4_5[14]},
      {stage4_6[8]},
      {stage4_7[12], stage4_7[13], stage4_7[14], stage4_7[15], stage4_7[16], stage4_7[17]},
      {stage5_9[2],stage5_8[3],stage5_7[3],stage5_6[4],stage5_5[4]}
   );
   gpc606_5 gpc1190 (
      {stage4_6[9], stage4_6[10], stage4_6[11], stage4_6[12], stage4_6[13], stage4_6[14]},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage5_10[0],stage5_9[3],stage5_8[4],stage5_7[4],stage5_6[5]}
   );
   gpc2135_5 gpc1191 (
      {stage4_9[0], stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4]},
      {stage4_10[0], stage4_10[1], stage4_10[2]},
      {stage4_11[0]},
      {stage4_12[0], stage4_12[1]},
      {stage5_13[0],stage5_12[0],stage5_11[0],stage5_10[1],stage5_9[4]}
   );
   gpc2135_5 gpc1192 (
      {stage4_9[5], stage4_9[6], stage4_9[7], stage4_9[8], stage4_9[9]},
      {stage4_10[3], stage4_10[4], stage4_10[5]},
      {stage4_11[1]},
      {stage4_12[2], stage4_12[3]},
      {stage5_13[1],stage5_12[1],stage5_11[1],stage5_10[2],stage5_9[5]}
   );
   gpc7_3 gpc1193 (
      {stage4_9[10], stage4_9[11], stage4_9[12], stage4_9[13], stage4_9[14], stage4_9[15], stage4_9[16]},
      {stage5_11[2],stage5_10[3],stage5_9[6]}
   );
   gpc2135_5 gpc1194 (
      {stage4_10[6], stage4_10[7], stage4_10[8], stage4_10[9], stage4_10[10]},
      {stage4_11[2], stage4_11[3], stage4_11[4]},
      {stage4_12[4]},
      {stage4_13[0], stage4_13[1]},
      {stage5_14[0],stage5_13[2],stage5_12[2],stage5_11[3],stage5_10[4]}
   );
   gpc606_5 gpc1195 (
      {stage4_10[11], stage4_10[12], stage4_10[13], stage4_10[14], stage4_10[15], stage4_10[16]},
      {stage4_12[5], stage4_12[6], stage4_12[7], stage4_12[8], stage4_12[9], stage4_12[10]},
      {stage5_14[1],stage5_13[3],stage5_12[3],stage5_11[4],stage5_10[5]}
   );
   gpc615_5 gpc1196 (
      {stage4_11[5], stage4_11[6], stage4_11[7], stage4_11[8], stage4_11[9]},
      {stage4_12[11]},
      {stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5], stage4_13[6], stage4_13[7]},
      {stage5_15[0],stage5_14[2],stage5_13[4],stage5_12[4],stage5_11[5]}
   );
   gpc615_5 gpc1197 (
      {stage4_11[10], stage4_11[11], stage4_11[12], stage4_11[13], stage4_11[14]},
      {stage4_12[12]},
      {stage4_13[8], stage4_13[9], stage4_13[10], stage4_13[11], stage4_13[12], stage4_13[13]},
      {stage5_15[1],stage5_14[3],stage5_13[5],stage5_12[5],stage5_11[6]}
   );
   gpc606_5 gpc1198 (
      {stage4_12[13], stage4_12[14], stage4_12[15], stage4_12[16], stage4_12[17], 1'b0},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[2],stage5_14[4],stage5_13[6],stage5_12[6]}
   );
   gpc606_5 gpc1199 (
      {stage4_13[14], stage4_13[15], stage4_13[16], stage4_13[17], stage4_13[18], stage4_13[19]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5]},
      {stage5_17[0],stage5_16[1],stage5_15[3],stage5_14[5],stage5_13[7]}
   );
   gpc606_5 gpc1200 (
      {stage4_14[6], stage4_14[7], stage4_14[8], stage4_14[9], stage4_14[10], stage4_14[11]},
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage5_18[0],stage5_17[1],stage5_16[2],stage5_15[4],stage5_14[6]}
   );
   gpc615_5 gpc1201 (
      {stage4_14[12], stage4_14[13], stage4_14[14], stage4_14[15], stage4_14[16]},
      {stage4_15[6]},
      {stage4_16[6], stage4_16[7], stage4_16[8], stage4_16[9], stage4_16[10], stage4_16[11]},
      {stage5_18[1],stage5_17[2],stage5_16[3],stage5_15[5],stage5_14[7]}
   );
   gpc1_1 gpc1202 (
      {stage4_0[3]},
      {stage5_0[1]}
   );
   gpc1_1 gpc1203 (
      {stage4_0[4]},
      {stage5_0[2]}
   );
   gpc1_1 gpc1204 (
      {stage4_0[5]},
      {stage5_0[3]}
   );
   gpc1_1 gpc1205 (
      {stage4_0[6]},
      {stage5_0[4]}
   );
   gpc1_1 gpc1206 (
      {stage4_0[7]},
      {stage5_0[5]}
   );
   gpc1_1 gpc1207 (
      {stage4_0[8]},
      {stage5_0[6]}
   );
   gpc1_1 gpc1208 (
      {stage4_1[6]},
      {stage5_1[1]}
   );
   gpc1_1 gpc1209 (
      {stage4_1[7]},
      {stage5_1[2]}
   );
   gpc1_1 gpc1210 (
      {stage4_1[8]},
      {stage5_1[3]}
   );
   gpc1_1 gpc1211 (
      {stage4_1[9]},
      {stage5_1[4]}
   );
   gpc1_1 gpc1212 (
      {stage4_1[10]},
      {stage5_1[5]}
   );
   gpc1_1 gpc1213 (
      {stage4_1[11]},
      {stage5_1[6]}
   );
   gpc1_1 gpc1214 (
      {stage4_2[4]},
      {stage5_2[2]}
   );
   gpc1_1 gpc1215 (
      {stage4_2[5]},
      {stage5_2[3]}
   );
   gpc1_1 gpc1216 (
      {stage4_2[6]},
      {stage5_2[4]}
   );
   gpc1_1 gpc1217 (
      {stage4_3[3]},
      {stage5_3[2]}
   );
   gpc1_1 gpc1218 (
      {stage4_3[4]},
      {stage5_3[3]}
   );
   gpc1_1 gpc1219 (
      {stage4_3[5]},
      {stage5_3[4]}
   );
   gpc1_1 gpc1220 (
      {stage4_3[6]},
      {stage5_3[5]}
   );
   gpc1_1 gpc1221 (
      {stage4_4[12]},
      {stage5_4[3]}
   );
   gpc1_1 gpc1222 (
      {stage4_6[15]},
      {stage5_6[6]}
   );
   gpc1_1 gpc1223 (
      {stage4_7[18]},
      {stage5_7[5]}
   );
   gpc1_1 gpc1224 (
      {stage4_8[6]},
      {stage5_8[5]}
   );
   gpc1_1 gpc1225 (
      {stage4_8[7]},
      {stage5_8[6]}
   );
   gpc1_1 gpc1226 (
      {stage4_8[8]},
      {stage5_8[7]}
   );
   gpc1_1 gpc1227 (
      {stage4_8[9]},
      {stage5_8[8]}
   );
   gpc1_1 gpc1228 (
      {stage4_8[10]},
      {stage5_8[9]}
   );
   gpc1_1 gpc1229 (
      {stage4_8[11]},
      {stage5_8[10]}
   );
   gpc1_1 gpc1230 (
      {stage4_8[12]},
      {stage5_8[11]}
   );
   gpc1_1 gpc1231 (
      {stage4_10[17]},
      {stage5_10[6]}
   );
   gpc1_1 gpc1232 (
      {stage4_10[18]},
      {stage5_10[7]}
   );
   gpc1_1 gpc1233 (
      {stage4_11[15]},
      {stage5_11[7]}
   );
   gpc1_1 gpc1234 (
      {stage4_13[20]},
      {stage5_13[8]}
   );
   gpc1_1 gpc1235 (
      {stage4_13[21]},
      {stage5_13[9]}
   );
   gpc1_1 gpc1236 (
      {stage4_13[22]},
      {stage5_13[10]}
   );
   gpc1_1 gpc1237 (
      {stage4_15[7]},
      {stage5_15[6]}
   );
   gpc1_1 gpc1238 (
      {stage4_17[0]},
      {stage5_17[3]}
   );
   gpc1_1 gpc1239 (
      {stage4_17[1]},
      {stage5_17[4]}
   );
   gpc1_1 gpc1240 (
      {stage4_17[2]},
      {stage5_17[5]}
   );
   gpc1_1 gpc1241 (
      {stage4_17[3]},
      {stage5_17[6]}
   );
   gpc117_4 gpc1242 (
      {stage5_0[0], stage5_0[1], stage5_0[2], stage5_0[3], stage5_0[4], stage5_0[5], stage5_0[6]},
      {stage5_1[0]},
      {stage5_2[0]},
      {stage6_3[0],stage6_2[0],stage6_1[0],stage6_0[0]}
   );
   gpc215_4 gpc1243 (
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4]},
      {stage5_6[0]},
      {stage5_7[0], stage5_7[1]},
      {stage6_8[0],stage6_7[0],stage6_6[0],stage6_5[0]}
   );
   gpc615_5 gpc1244 (
      {stage5_6[1], stage5_6[2], stage5_6[3], stage5_6[4], stage5_6[5]},
      {stage5_7[2]},
      {stage5_8[0], stage5_8[1], stage5_8[2], stage5_8[3], stage5_8[4], stage5_8[5]},
      {stage6_10[0],stage6_9[0],stage6_8[1],stage6_7[1],stage6_6[1]}
   );
   gpc623_5 gpc1245 (
      {stage5_7[3], stage5_7[4], stage5_7[5]},
      {stage5_8[6], stage5_8[7]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3], stage5_9[4], stage5_9[5]},
      {stage6_11[0],stage6_10[1],stage6_9[1],stage6_8[2],stage6_7[2]}
   );
   gpc1163_5 gpc1246 (
      {stage5_10[0], stage5_10[1], stage5_10[2]},
      {stage5_11[0], stage5_11[1], stage5_11[2], stage5_11[3], stage5_11[4], stage5_11[5]},
      {stage5_12[0]},
      {stage5_13[0]},
      {stage6_14[0],stage6_13[0],stage6_12[0],stage6_11[1],stage6_10[2]}
   );
   gpc615_5 gpc1247 (
      {stage5_10[3], stage5_10[4], stage5_10[5], stage5_10[6], stage5_10[7]},
      {stage5_11[6]},
      {stage5_12[1], stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5], stage5_12[6]},
      {stage6_14[1],stage6_13[1],stage6_12[1],stage6_11[2],stage6_10[3]}
   );
   gpc1163_5 gpc1248 (
      {stage5_13[1], stage5_13[2], stage5_13[3]},
      {stage5_14[0], stage5_14[1], stage5_14[2], stage5_14[3], stage5_14[4], stage5_14[5]},
      {stage5_15[0]},
      {stage5_16[0]},
      {stage6_17[0],stage6_16[0],stage6_15[0],stage6_14[2],stage6_13[2]}
   );
   gpc615_5 gpc1249 (
      {stage5_13[4], stage5_13[5], stage5_13[6], stage5_13[7], stage5_13[8]},
      {stage5_14[6]},
      {stage5_15[1], stage5_15[2], stage5_15[3], stage5_15[4], stage5_15[5], stage5_15[6]},
      {stage6_17[1],stage6_16[1],stage6_15[1],stage6_14[3],stage6_13[3]}
   );
   gpc1163_5 gpc1250 (
      {stage5_16[1], stage5_16[2], stage5_16[3]},
      {stage5_17[0], stage5_17[1], stage5_17[2], stage5_17[3], stage5_17[4], stage5_17[5]},
      {stage5_18[0]},
      {1'b0},
      {stage6_20[0],stage6_19[0],stage6_18[0],stage6_17[2],stage6_16[2]}
   );
   gpc1_1 gpc1251 (
      {stage5_1[1]},
      {stage6_1[1]}
   );
   gpc1_1 gpc1252 (
      {stage5_1[2]},
      {stage6_1[2]}
   );
   gpc1_1 gpc1253 (
      {stage5_1[3]},
      {stage6_1[3]}
   );
   gpc1_1 gpc1254 (
      {stage5_1[4]},
      {stage6_1[4]}
   );
   gpc1_1 gpc1255 (
      {stage5_1[5]},
      {stage6_1[5]}
   );
   gpc1_1 gpc1256 (
      {stage5_1[6]},
      {stage6_1[6]}
   );
   gpc1_1 gpc1257 (
      {stage5_2[1]},
      {stage6_2[1]}
   );
   gpc1_1 gpc1258 (
      {stage5_2[2]},
      {stage6_2[2]}
   );
   gpc1_1 gpc1259 (
      {stage5_2[3]},
      {stage6_2[3]}
   );
   gpc1_1 gpc1260 (
      {stage5_2[4]},
      {stage6_2[4]}
   );
   gpc1_1 gpc1261 (
      {stage5_3[0]},
      {stage6_3[1]}
   );
   gpc1_1 gpc1262 (
      {stage5_3[1]},
      {stage6_3[2]}
   );
   gpc1_1 gpc1263 (
      {stage5_3[2]},
      {stage6_3[3]}
   );
   gpc1_1 gpc1264 (
      {stage5_3[3]},
      {stage6_3[4]}
   );
   gpc1_1 gpc1265 (
      {stage5_3[4]},
      {stage6_3[5]}
   );
   gpc1_1 gpc1266 (
      {stage5_3[5]},
      {stage6_3[6]}
   );
   gpc1_1 gpc1267 (
      {stage5_4[0]},
      {stage6_4[0]}
   );
   gpc1_1 gpc1268 (
      {stage5_4[1]},
      {stage6_4[1]}
   );
   gpc1_1 gpc1269 (
      {stage5_4[2]},
      {stage6_4[2]}
   );
   gpc1_1 gpc1270 (
      {stage5_4[3]},
      {stage6_4[3]}
   );
   gpc1_1 gpc1271 (
      {stage5_6[6]},
      {stage6_6[2]}
   );
   gpc1_1 gpc1272 (
      {stage5_8[8]},
      {stage6_8[3]}
   );
   gpc1_1 gpc1273 (
      {stage5_8[9]},
      {stage6_8[4]}
   );
   gpc1_1 gpc1274 (
      {stage5_8[10]},
      {stage6_8[5]}
   );
   gpc1_1 gpc1275 (
      {stage5_8[11]},
      {stage6_8[6]}
   );
   gpc1_1 gpc1276 (
      {stage5_9[6]},
      {stage6_9[2]}
   );
   gpc1_1 gpc1277 (
      {stage5_11[7]},
      {stage6_11[3]}
   );
   gpc1_1 gpc1278 (
      {stage5_13[9]},
      {stage6_13[4]}
   );
   gpc1_1 gpc1279 (
      {stage5_13[10]},
      {stage6_13[5]}
   );
   gpc1_1 gpc1280 (
      {stage5_14[7]},
      {stage6_14[4]}
   );
   gpc1_1 gpc1281 (
      {stage5_17[6]},
      {stage6_17[3]}
   );
   gpc1_1 gpc1282 (
      {stage5_18[1]},
      {stage6_18[1]}
   );
   gpc606_5 gpc1283 (
      {stage6_1[0], stage6_1[1], stage6_1[2], stage6_1[3], stage6_1[4], stage6_1[5]},
      {stage6_3[0], stage6_3[1], stage6_3[2], stage6_3[3], stage6_3[4], stage6_3[5]},
      {stage7_5[0],stage7_4[0],stage7_3[0],stage7_2[0],stage7_1[0]}
   );
   gpc1415_5 gpc1284 (
      {stage6_2[0], stage6_2[1], stage6_2[2], stage6_2[3], stage6_2[4]},
      {stage6_3[6]},
      {stage6_4[0], stage6_4[1], stage6_4[2], stage6_4[3]},
      {stage6_5[0]},
      {stage7_6[0],stage7_5[1],stage7_4[1],stage7_3[1],stage7_2[1]}
   );
   gpc623_5 gpc1285 (
      {stage6_6[0], stage6_6[1], stage6_6[2]},
      {stage6_7[0], stage6_7[1]},
      {stage6_8[0], stage6_8[1], stage6_8[2], stage6_8[3], stage6_8[4], stage6_8[5]},
      {stage7_10[0],stage7_9[0],stage7_8[0],stage7_7[0],stage7_6[1]}
   );
   gpc1343_5 gpc1286 (
      {stage6_9[0], stage6_9[1], stage6_9[2]},
      {stage6_10[0], stage6_10[1], stage6_10[2], stage6_10[3]},
      {stage6_11[0], stage6_11[1], stage6_11[2]},
      {stage6_12[0]},
      {stage7_13[0],stage7_12[0],stage7_11[0],stage7_10[1],stage7_9[1]}
   );
   gpc207_4 gpc1287 (
      {stage6_13[0], stage6_13[1], stage6_13[2], stage6_13[3], stage6_13[4], stage6_13[5], 1'b0},
      {stage6_15[0], stage6_15[1]},
      {stage7_16[0],stage7_15[0],stage7_14[0],stage7_13[1]}
   );
   gpc1406_5 gpc1288 (
      {stage6_14[0], stage6_14[1], stage6_14[2], stage6_14[3], stage6_14[4], 1'b0},
      {stage6_16[0], stage6_16[1], stage6_16[2], 1'b0},
      {stage6_17[0]},
      {stage7_18[0],stage7_17[0],stage7_16[1],stage7_15[1],stage7_14[1]}
   );
   gpc135_4 gpc1289 (
      {stage6_17[1], stage6_17[2], stage6_17[3], 1'b0, 1'b0},
      {stage6_18[0], stage6_18[1], 1'b0},
      {stage6_19[0]},
      {stage7_20[0],stage7_19[0],stage7_18[1],stage7_17[1]}
   );
   gpc1_1 gpc1290 (
      {stage6_0[0]},
      {stage7_0[0]}
   );
   gpc1_1 gpc1291 (
      {stage6_1[6]},
      {stage7_1[1]}
   );
   gpc1_1 gpc1292 (
      {stage6_7[2]},
      {stage7_7[1]}
   );
   gpc1_1 gpc1293 (
      {stage6_8[6]},
      {stage7_8[1]}
   );
   gpc1_1 gpc1294 (
      {stage6_11[3]},
      {stage7_11[1]}
   );
   gpc1_1 gpc1295 (
      {stage6_12[1]},
      {stage7_12[1]}
   );
   gpc1_1 gpc1296 (
      {stage6_20[0]},
      {stage7_20[1]}
   );
endmodule
module rowadder2_1_21(input [20:0] src0, input [20:0] src1, output [21:0] dst0);
    wire [20:0] gene;
    wire [20:0] prop;
    wire [23:0] out;
    wire [23:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_19_gene (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(gene[19])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_19_prop (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(prop[19])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_20_gene (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(gene[20])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_20_prop (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(prop[20])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    CARRY4 carry4_23_20 (
        .CO(carryout[23:20]),
        .O(out[23:20]),
        .CI(carryout[19]),
        .CYINIT(1'h0),
        .DI({3'h0, gene[20:20]}),
        .S({3'h0, prop[20:20]})
    );
    assign dst0 = {carryout[20], out[20:0]};
endmodule


module testbench();
    reg [485:0] src0;
    reg [485:0] src1;
    reg [485:0] src2;
    reg [485:0] src3;
    reg [485:0] src4;
    reg [485:0] src5;
    reg [485:0] src6;
    reg [485:0] src7;
    reg [485:0] src8;
    reg [485:0] src9;
    reg [485:0] src10;
    reg [485:0] src11;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [20:0] srcsum;
    wire [20:0] dstsum;
    wire test;
    compressor2_1_486_12 compressor2_1_486_12(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255] + src0[256] + src0[257] + src0[258] + src0[259] + src0[260] + src0[261] + src0[262] + src0[263] + src0[264] + src0[265] + src0[266] + src0[267] + src0[268] + src0[269] + src0[270] + src0[271] + src0[272] + src0[273] + src0[274] + src0[275] + src0[276] + src0[277] + src0[278] + src0[279] + src0[280] + src0[281] + src0[282] + src0[283] + src0[284] + src0[285] + src0[286] + src0[287] + src0[288] + src0[289] + src0[290] + src0[291] + src0[292] + src0[293] + src0[294] + src0[295] + src0[296] + src0[297] + src0[298] + src0[299] + src0[300] + src0[301] + src0[302] + src0[303] + src0[304] + src0[305] + src0[306] + src0[307] + src0[308] + src0[309] + src0[310] + src0[311] + src0[312] + src0[313] + src0[314] + src0[315] + src0[316] + src0[317] + src0[318] + src0[319] + src0[320] + src0[321] + src0[322] + src0[323] + src0[324] + src0[325] + src0[326] + src0[327] + src0[328] + src0[329] + src0[330] + src0[331] + src0[332] + src0[333] + src0[334] + src0[335] + src0[336] + src0[337] + src0[338] + src0[339] + src0[340] + src0[341] + src0[342] + src0[343] + src0[344] + src0[345] + src0[346] + src0[347] + src0[348] + src0[349] + src0[350] + src0[351] + src0[352] + src0[353] + src0[354] + src0[355] + src0[356] + src0[357] + src0[358] + src0[359] + src0[360] + src0[361] + src0[362] + src0[363] + src0[364] + src0[365] + src0[366] + src0[367] + src0[368] + src0[369] + src0[370] + src0[371] + src0[372] + src0[373] + src0[374] + src0[375] + src0[376] + src0[377] + src0[378] + src0[379] + src0[380] + src0[381] + src0[382] + src0[383] + src0[384] + src0[385] + src0[386] + src0[387] + src0[388] + src0[389] + src0[390] + src0[391] + src0[392] + src0[393] + src0[394] + src0[395] + src0[396] + src0[397] + src0[398] + src0[399] + src0[400] + src0[401] + src0[402] + src0[403] + src0[404] + src0[405] + src0[406] + src0[407] + src0[408] + src0[409] + src0[410] + src0[411] + src0[412] + src0[413] + src0[414] + src0[415] + src0[416] + src0[417] + src0[418] + src0[419] + src0[420] + src0[421] + src0[422] + src0[423] + src0[424] + src0[425] + src0[426] + src0[427] + src0[428] + src0[429] + src0[430] + src0[431] + src0[432] + src0[433] + src0[434] + src0[435] + src0[436] + src0[437] + src0[438] + src0[439] + src0[440] + src0[441] + src0[442] + src0[443] + src0[444] + src0[445] + src0[446] + src0[447] + src0[448] + src0[449] + src0[450] + src0[451] + src0[452] + src0[453] + src0[454] + src0[455] + src0[456] + src0[457] + src0[458] + src0[459] + src0[460] + src0[461] + src0[462] + src0[463] + src0[464] + src0[465] + src0[466] + src0[467] + src0[468] + src0[469] + src0[470] + src0[471] + src0[472] + src0[473] + src0[474] + src0[475] + src0[476] + src0[477] + src0[478] + src0[479] + src0[480] + src0[481] + src0[482] + src0[483] + src0[484] + src0[485])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255] + src1[256] + src1[257] + src1[258] + src1[259] + src1[260] + src1[261] + src1[262] + src1[263] + src1[264] + src1[265] + src1[266] + src1[267] + src1[268] + src1[269] + src1[270] + src1[271] + src1[272] + src1[273] + src1[274] + src1[275] + src1[276] + src1[277] + src1[278] + src1[279] + src1[280] + src1[281] + src1[282] + src1[283] + src1[284] + src1[285] + src1[286] + src1[287] + src1[288] + src1[289] + src1[290] + src1[291] + src1[292] + src1[293] + src1[294] + src1[295] + src1[296] + src1[297] + src1[298] + src1[299] + src1[300] + src1[301] + src1[302] + src1[303] + src1[304] + src1[305] + src1[306] + src1[307] + src1[308] + src1[309] + src1[310] + src1[311] + src1[312] + src1[313] + src1[314] + src1[315] + src1[316] + src1[317] + src1[318] + src1[319] + src1[320] + src1[321] + src1[322] + src1[323] + src1[324] + src1[325] + src1[326] + src1[327] + src1[328] + src1[329] + src1[330] + src1[331] + src1[332] + src1[333] + src1[334] + src1[335] + src1[336] + src1[337] + src1[338] + src1[339] + src1[340] + src1[341] + src1[342] + src1[343] + src1[344] + src1[345] + src1[346] + src1[347] + src1[348] + src1[349] + src1[350] + src1[351] + src1[352] + src1[353] + src1[354] + src1[355] + src1[356] + src1[357] + src1[358] + src1[359] + src1[360] + src1[361] + src1[362] + src1[363] + src1[364] + src1[365] + src1[366] + src1[367] + src1[368] + src1[369] + src1[370] + src1[371] + src1[372] + src1[373] + src1[374] + src1[375] + src1[376] + src1[377] + src1[378] + src1[379] + src1[380] + src1[381] + src1[382] + src1[383] + src1[384] + src1[385] + src1[386] + src1[387] + src1[388] + src1[389] + src1[390] + src1[391] + src1[392] + src1[393] + src1[394] + src1[395] + src1[396] + src1[397] + src1[398] + src1[399] + src1[400] + src1[401] + src1[402] + src1[403] + src1[404] + src1[405] + src1[406] + src1[407] + src1[408] + src1[409] + src1[410] + src1[411] + src1[412] + src1[413] + src1[414] + src1[415] + src1[416] + src1[417] + src1[418] + src1[419] + src1[420] + src1[421] + src1[422] + src1[423] + src1[424] + src1[425] + src1[426] + src1[427] + src1[428] + src1[429] + src1[430] + src1[431] + src1[432] + src1[433] + src1[434] + src1[435] + src1[436] + src1[437] + src1[438] + src1[439] + src1[440] + src1[441] + src1[442] + src1[443] + src1[444] + src1[445] + src1[446] + src1[447] + src1[448] + src1[449] + src1[450] + src1[451] + src1[452] + src1[453] + src1[454] + src1[455] + src1[456] + src1[457] + src1[458] + src1[459] + src1[460] + src1[461] + src1[462] + src1[463] + src1[464] + src1[465] + src1[466] + src1[467] + src1[468] + src1[469] + src1[470] + src1[471] + src1[472] + src1[473] + src1[474] + src1[475] + src1[476] + src1[477] + src1[478] + src1[479] + src1[480] + src1[481] + src1[482] + src1[483] + src1[484] + src1[485])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255] + src2[256] + src2[257] + src2[258] + src2[259] + src2[260] + src2[261] + src2[262] + src2[263] + src2[264] + src2[265] + src2[266] + src2[267] + src2[268] + src2[269] + src2[270] + src2[271] + src2[272] + src2[273] + src2[274] + src2[275] + src2[276] + src2[277] + src2[278] + src2[279] + src2[280] + src2[281] + src2[282] + src2[283] + src2[284] + src2[285] + src2[286] + src2[287] + src2[288] + src2[289] + src2[290] + src2[291] + src2[292] + src2[293] + src2[294] + src2[295] + src2[296] + src2[297] + src2[298] + src2[299] + src2[300] + src2[301] + src2[302] + src2[303] + src2[304] + src2[305] + src2[306] + src2[307] + src2[308] + src2[309] + src2[310] + src2[311] + src2[312] + src2[313] + src2[314] + src2[315] + src2[316] + src2[317] + src2[318] + src2[319] + src2[320] + src2[321] + src2[322] + src2[323] + src2[324] + src2[325] + src2[326] + src2[327] + src2[328] + src2[329] + src2[330] + src2[331] + src2[332] + src2[333] + src2[334] + src2[335] + src2[336] + src2[337] + src2[338] + src2[339] + src2[340] + src2[341] + src2[342] + src2[343] + src2[344] + src2[345] + src2[346] + src2[347] + src2[348] + src2[349] + src2[350] + src2[351] + src2[352] + src2[353] + src2[354] + src2[355] + src2[356] + src2[357] + src2[358] + src2[359] + src2[360] + src2[361] + src2[362] + src2[363] + src2[364] + src2[365] + src2[366] + src2[367] + src2[368] + src2[369] + src2[370] + src2[371] + src2[372] + src2[373] + src2[374] + src2[375] + src2[376] + src2[377] + src2[378] + src2[379] + src2[380] + src2[381] + src2[382] + src2[383] + src2[384] + src2[385] + src2[386] + src2[387] + src2[388] + src2[389] + src2[390] + src2[391] + src2[392] + src2[393] + src2[394] + src2[395] + src2[396] + src2[397] + src2[398] + src2[399] + src2[400] + src2[401] + src2[402] + src2[403] + src2[404] + src2[405] + src2[406] + src2[407] + src2[408] + src2[409] + src2[410] + src2[411] + src2[412] + src2[413] + src2[414] + src2[415] + src2[416] + src2[417] + src2[418] + src2[419] + src2[420] + src2[421] + src2[422] + src2[423] + src2[424] + src2[425] + src2[426] + src2[427] + src2[428] + src2[429] + src2[430] + src2[431] + src2[432] + src2[433] + src2[434] + src2[435] + src2[436] + src2[437] + src2[438] + src2[439] + src2[440] + src2[441] + src2[442] + src2[443] + src2[444] + src2[445] + src2[446] + src2[447] + src2[448] + src2[449] + src2[450] + src2[451] + src2[452] + src2[453] + src2[454] + src2[455] + src2[456] + src2[457] + src2[458] + src2[459] + src2[460] + src2[461] + src2[462] + src2[463] + src2[464] + src2[465] + src2[466] + src2[467] + src2[468] + src2[469] + src2[470] + src2[471] + src2[472] + src2[473] + src2[474] + src2[475] + src2[476] + src2[477] + src2[478] + src2[479] + src2[480] + src2[481] + src2[482] + src2[483] + src2[484] + src2[485])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255] + src3[256] + src3[257] + src3[258] + src3[259] + src3[260] + src3[261] + src3[262] + src3[263] + src3[264] + src3[265] + src3[266] + src3[267] + src3[268] + src3[269] + src3[270] + src3[271] + src3[272] + src3[273] + src3[274] + src3[275] + src3[276] + src3[277] + src3[278] + src3[279] + src3[280] + src3[281] + src3[282] + src3[283] + src3[284] + src3[285] + src3[286] + src3[287] + src3[288] + src3[289] + src3[290] + src3[291] + src3[292] + src3[293] + src3[294] + src3[295] + src3[296] + src3[297] + src3[298] + src3[299] + src3[300] + src3[301] + src3[302] + src3[303] + src3[304] + src3[305] + src3[306] + src3[307] + src3[308] + src3[309] + src3[310] + src3[311] + src3[312] + src3[313] + src3[314] + src3[315] + src3[316] + src3[317] + src3[318] + src3[319] + src3[320] + src3[321] + src3[322] + src3[323] + src3[324] + src3[325] + src3[326] + src3[327] + src3[328] + src3[329] + src3[330] + src3[331] + src3[332] + src3[333] + src3[334] + src3[335] + src3[336] + src3[337] + src3[338] + src3[339] + src3[340] + src3[341] + src3[342] + src3[343] + src3[344] + src3[345] + src3[346] + src3[347] + src3[348] + src3[349] + src3[350] + src3[351] + src3[352] + src3[353] + src3[354] + src3[355] + src3[356] + src3[357] + src3[358] + src3[359] + src3[360] + src3[361] + src3[362] + src3[363] + src3[364] + src3[365] + src3[366] + src3[367] + src3[368] + src3[369] + src3[370] + src3[371] + src3[372] + src3[373] + src3[374] + src3[375] + src3[376] + src3[377] + src3[378] + src3[379] + src3[380] + src3[381] + src3[382] + src3[383] + src3[384] + src3[385] + src3[386] + src3[387] + src3[388] + src3[389] + src3[390] + src3[391] + src3[392] + src3[393] + src3[394] + src3[395] + src3[396] + src3[397] + src3[398] + src3[399] + src3[400] + src3[401] + src3[402] + src3[403] + src3[404] + src3[405] + src3[406] + src3[407] + src3[408] + src3[409] + src3[410] + src3[411] + src3[412] + src3[413] + src3[414] + src3[415] + src3[416] + src3[417] + src3[418] + src3[419] + src3[420] + src3[421] + src3[422] + src3[423] + src3[424] + src3[425] + src3[426] + src3[427] + src3[428] + src3[429] + src3[430] + src3[431] + src3[432] + src3[433] + src3[434] + src3[435] + src3[436] + src3[437] + src3[438] + src3[439] + src3[440] + src3[441] + src3[442] + src3[443] + src3[444] + src3[445] + src3[446] + src3[447] + src3[448] + src3[449] + src3[450] + src3[451] + src3[452] + src3[453] + src3[454] + src3[455] + src3[456] + src3[457] + src3[458] + src3[459] + src3[460] + src3[461] + src3[462] + src3[463] + src3[464] + src3[465] + src3[466] + src3[467] + src3[468] + src3[469] + src3[470] + src3[471] + src3[472] + src3[473] + src3[474] + src3[475] + src3[476] + src3[477] + src3[478] + src3[479] + src3[480] + src3[481] + src3[482] + src3[483] + src3[484] + src3[485])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255] + src4[256] + src4[257] + src4[258] + src4[259] + src4[260] + src4[261] + src4[262] + src4[263] + src4[264] + src4[265] + src4[266] + src4[267] + src4[268] + src4[269] + src4[270] + src4[271] + src4[272] + src4[273] + src4[274] + src4[275] + src4[276] + src4[277] + src4[278] + src4[279] + src4[280] + src4[281] + src4[282] + src4[283] + src4[284] + src4[285] + src4[286] + src4[287] + src4[288] + src4[289] + src4[290] + src4[291] + src4[292] + src4[293] + src4[294] + src4[295] + src4[296] + src4[297] + src4[298] + src4[299] + src4[300] + src4[301] + src4[302] + src4[303] + src4[304] + src4[305] + src4[306] + src4[307] + src4[308] + src4[309] + src4[310] + src4[311] + src4[312] + src4[313] + src4[314] + src4[315] + src4[316] + src4[317] + src4[318] + src4[319] + src4[320] + src4[321] + src4[322] + src4[323] + src4[324] + src4[325] + src4[326] + src4[327] + src4[328] + src4[329] + src4[330] + src4[331] + src4[332] + src4[333] + src4[334] + src4[335] + src4[336] + src4[337] + src4[338] + src4[339] + src4[340] + src4[341] + src4[342] + src4[343] + src4[344] + src4[345] + src4[346] + src4[347] + src4[348] + src4[349] + src4[350] + src4[351] + src4[352] + src4[353] + src4[354] + src4[355] + src4[356] + src4[357] + src4[358] + src4[359] + src4[360] + src4[361] + src4[362] + src4[363] + src4[364] + src4[365] + src4[366] + src4[367] + src4[368] + src4[369] + src4[370] + src4[371] + src4[372] + src4[373] + src4[374] + src4[375] + src4[376] + src4[377] + src4[378] + src4[379] + src4[380] + src4[381] + src4[382] + src4[383] + src4[384] + src4[385] + src4[386] + src4[387] + src4[388] + src4[389] + src4[390] + src4[391] + src4[392] + src4[393] + src4[394] + src4[395] + src4[396] + src4[397] + src4[398] + src4[399] + src4[400] + src4[401] + src4[402] + src4[403] + src4[404] + src4[405] + src4[406] + src4[407] + src4[408] + src4[409] + src4[410] + src4[411] + src4[412] + src4[413] + src4[414] + src4[415] + src4[416] + src4[417] + src4[418] + src4[419] + src4[420] + src4[421] + src4[422] + src4[423] + src4[424] + src4[425] + src4[426] + src4[427] + src4[428] + src4[429] + src4[430] + src4[431] + src4[432] + src4[433] + src4[434] + src4[435] + src4[436] + src4[437] + src4[438] + src4[439] + src4[440] + src4[441] + src4[442] + src4[443] + src4[444] + src4[445] + src4[446] + src4[447] + src4[448] + src4[449] + src4[450] + src4[451] + src4[452] + src4[453] + src4[454] + src4[455] + src4[456] + src4[457] + src4[458] + src4[459] + src4[460] + src4[461] + src4[462] + src4[463] + src4[464] + src4[465] + src4[466] + src4[467] + src4[468] + src4[469] + src4[470] + src4[471] + src4[472] + src4[473] + src4[474] + src4[475] + src4[476] + src4[477] + src4[478] + src4[479] + src4[480] + src4[481] + src4[482] + src4[483] + src4[484] + src4[485])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255] + src5[256] + src5[257] + src5[258] + src5[259] + src5[260] + src5[261] + src5[262] + src5[263] + src5[264] + src5[265] + src5[266] + src5[267] + src5[268] + src5[269] + src5[270] + src5[271] + src5[272] + src5[273] + src5[274] + src5[275] + src5[276] + src5[277] + src5[278] + src5[279] + src5[280] + src5[281] + src5[282] + src5[283] + src5[284] + src5[285] + src5[286] + src5[287] + src5[288] + src5[289] + src5[290] + src5[291] + src5[292] + src5[293] + src5[294] + src5[295] + src5[296] + src5[297] + src5[298] + src5[299] + src5[300] + src5[301] + src5[302] + src5[303] + src5[304] + src5[305] + src5[306] + src5[307] + src5[308] + src5[309] + src5[310] + src5[311] + src5[312] + src5[313] + src5[314] + src5[315] + src5[316] + src5[317] + src5[318] + src5[319] + src5[320] + src5[321] + src5[322] + src5[323] + src5[324] + src5[325] + src5[326] + src5[327] + src5[328] + src5[329] + src5[330] + src5[331] + src5[332] + src5[333] + src5[334] + src5[335] + src5[336] + src5[337] + src5[338] + src5[339] + src5[340] + src5[341] + src5[342] + src5[343] + src5[344] + src5[345] + src5[346] + src5[347] + src5[348] + src5[349] + src5[350] + src5[351] + src5[352] + src5[353] + src5[354] + src5[355] + src5[356] + src5[357] + src5[358] + src5[359] + src5[360] + src5[361] + src5[362] + src5[363] + src5[364] + src5[365] + src5[366] + src5[367] + src5[368] + src5[369] + src5[370] + src5[371] + src5[372] + src5[373] + src5[374] + src5[375] + src5[376] + src5[377] + src5[378] + src5[379] + src5[380] + src5[381] + src5[382] + src5[383] + src5[384] + src5[385] + src5[386] + src5[387] + src5[388] + src5[389] + src5[390] + src5[391] + src5[392] + src5[393] + src5[394] + src5[395] + src5[396] + src5[397] + src5[398] + src5[399] + src5[400] + src5[401] + src5[402] + src5[403] + src5[404] + src5[405] + src5[406] + src5[407] + src5[408] + src5[409] + src5[410] + src5[411] + src5[412] + src5[413] + src5[414] + src5[415] + src5[416] + src5[417] + src5[418] + src5[419] + src5[420] + src5[421] + src5[422] + src5[423] + src5[424] + src5[425] + src5[426] + src5[427] + src5[428] + src5[429] + src5[430] + src5[431] + src5[432] + src5[433] + src5[434] + src5[435] + src5[436] + src5[437] + src5[438] + src5[439] + src5[440] + src5[441] + src5[442] + src5[443] + src5[444] + src5[445] + src5[446] + src5[447] + src5[448] + src5[449] + src5[450] + src5[451] + src5[452] + src5[453] + src5[454] + src5[455] + src5[456] + src5[457] + src5[458] + src5[459] + src5[460] + src5[461] + src5[462] + src5[463] + src5[464] + src5[465] + src5[466] + src5[467] + src5[468] + src5[469] + src5[470] + src5[471] + src5[472] + src5[473] + src5[474] + src5[475] + src5[476] + src5[477] + src5[478] + src5[479] + src5[480] + src5[481] + src5[482] + src5[483] + src5[484] + src5[485])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255] + src6[256] + src6[257] + src6[258] + src6[259] + src6[260] + src6[261] + src6[262] + src6[263] + src6[264] + src6[265] + src6[266] + src6[267] + src6[268] + src6[269] + src6[270] + src6[271] + src6[272] + src6[273] + src6[274] + src6[275] + src6[276] + src6[277] + src6[278] + src6[279] + src6[280] + src6[281] + src6[282] + src6[283] + src6[284] + src6[285] + src6[286] + src6[287] + src6[288] + src6[289] + src6[290] + src6[291] + src6[292] + src6[293] + src6[294] + src6[295] + src6[296] + src6[297] + src6[298] + src6[299] + src6[300] + src6[301] + src6[302] + src6[303] + src6[304] + src6[305] + src6[306] + src6[307] + src6[308] + src6[309] + src6[310] + src6[311] + src6[312] + src6[313] + src6[314] + src6[315] + src6[316] + src6[317] + src6[318] + src6[319] + src6[320] + src6[321] + src6[322] + src6[323] + src6[324] + src6[325] + src6[326] + src6[327] + src6[328] + src6[329] + src6[330] + src6[331] + src6[332] + src6[333] + src6[334] + src6[335] + src6[336] + src6[337] + src6[338] + src6[339] + src6[340] + src6[341] + src6[342] + src6[343] + src6[344] + src6[345] + src6[346] + src6[347] + src6[348] + src6[349] + src6[350] + src6[351] + src6[352] + src6[353] + src6[354] + src6[355] + src6[356] + src6[357] + src6[358] + src6[359] + src6[360] + src6[361] + src6[362] + src6[363] + src6[364] + src6[365] + src6[366] + src6[367] + src6[368] + src6[369] + src6[370] + src6[371] + src6[372] + src6[373] + src6[374] + src6[375] + src6[376] + src6[377] + src6[378] + src6[379] + src6[380] + src6[381] + src6[382] + src6[383] + src6[384] + src6[385] + src6[386] + src6[387] + src6[388] + src6[389] + src6[390] + src6[391] + src6[392] + src6[393] + src6[394] + src6[395] + src6[396] + src6[397] + src6[398] + src6[399] + src6[400] + src6[401] + src6[402] + src6[403] + src6[404] + src6[405] + src6[406] + src6[407] + src6[408] + src6[409] + src6[410] + src6[411] + src6[412] + src6[413] + src6[414] + src6[415] + src6[416] + src6[417] + src6[418] + src6[419] + src6[420] + src6[421] + src6[422] + src6[423] + src6[424] + src6[425] + src6[426] + src6[427] + src6[428] + src6[429] + src6[430] + src6[431] + src6[432] + src6[433] + src6[434] + src6[435] + src6[436] + src6[437] + src6[438] + src6[439] + src6[440] + src6[441] + src6[442] + src6[443] + src6[444] + src6[445] + src6[446] + src6[447] + src6[448] + src6[449] + src6[450] + src6[451] + src6[452] + src6[453] + src6[454] + src6[455] + src6[456] + src6[457] + src6[458] + src6[459] + src6[460] + src6[461] + src6[462] + src6[463] + src6[464] + src6[465] + src6[466] + src6[467] + src6[468] + src6[469] + src6[470] + src6[471] + src6[472] + src6[473] + src6[474] + src6[475] + src6[476] + src6[477] + src6[478] + src6[479] + src6[480] + src6[481] + src6[482] + src6[483] + src6[484] + src6[485])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255] + src7[256] + src7[257] + src7[258] + src7[259] + src7[260] + src7[261] + src7[262] + src7[263] + src7[264] + src7[265] + src7[266] + src7[267] + src7[268] + src7[269] + src7[270] + src7[271] + src7[272] + src7[273] + src7[274] + src7[275] + src7[276] + src7[277] + src7[278] + src7[279] + src7[280] + src7[281] + src7[282] + src7[283] + src7[284] + src7[285] + src7[286] + src7[287] + src7[288] + src7[289] + src7[290] + src7[291] + src7[292] + src7[293] + src7[294] + src7[295] + src7[296] + src7[297] + src7[298] + src7[299] + src7[300] + src7[301] + src7[302] + src7[303] + src7[304] + src7[305] + src7[306] + src7[307] + src7[308] + src7[309] + src7[310] + src7[311] + src7[312] + src7[313] + src7[314] + src7[315] + src7[316] + src7[317] + src7[318] + src7[319] + src7[320] + src7[321] + src7[322] + src7[323] + src7[324] + src7[325] + src7[326] + src7[327] + src7[328] + src7[329] + src7[330] + src7[331] + src7[332] + src7[333] + src7[334] + src7[335] + src7[336] + src7[337] + src7[338] + src7[339] + src7[340] + src7[341] + src7[342] + src7[343] + src7[344] + src7[345] + src7[346] + src7[347] + src7[348] + src7[349] + src7[350] + src7[351] + src7[352] + src7[353] + src7[354] + src7[355] + src7[356] + src7[357] + src7[358] + src7[359] + src7[360] + src7[361] + src7[362] + src7[363] + src7[364] + src7[365] + src7[366] + src7[367] + src7[368] + src7[369] + src7[370] + src7[371] + src7[372] + src7[373] + src7[374] + src7[375] + src7[376] + src7[377] + src7[378] + src7[379] + src7[380] + src7[381] + src7[382] + src7[383] + src7[384] + src7[385] + src7[386] + src7[387] + src7[388] + src7[389] + src7[390] + src7[391] + src7[392] + src7[393] + src7[394] + src7[395] + src7[396] + src7[397] + src7[398] + src7[399] + src7[400] + src7[401] + src7[402] + src7[403] + src7[404] + src7[405] + src7[406] + src7[407] + src7[408] + src7[409] + src7[410] + src7[411] + src7[412] + src7[413] + src7[414] + src7[415] + src7[416] + src7[417] + src7[418] + src7[419] + src7[420] + src7[421] + src7[422] + src7[423] + src7[424] + src7[425] + src7[426] + src7[427] + src7[428] + src7[429] + src7[430] + src7[431] + src7[432] + src7[433] + src7[434] + src7[435] + src7[436] + src7[437] + src7[438] + src7[439] + src7[440] + src7[441] + src7[442] + src7[443] + src7[444] + src7[445] + src7[446] + src7[447] + src7[448] + src7[449] + src7[450] + src7[451] + src7[452] + src7[453] + src7[454] + src7[455] + src7[456] + src7[457] + src7[458] + src7[459] + src7[460] + src7[461] + src7[462] + src7[463] + src7[464] + src7[465] + src7[466] + src7[467] + src7[468] + src7[469] + src7[470] + src7[471] + src7[472] + src7[473] + src7[474] + src7[475] + src7[476] + src7[477] + src7[478] + src7[479] + src7[480] + src7[481] + src7[482] + src7[483] + src7[484] + src7[485])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255] + src8[256] + src8[257] + src8[258] + src8[259] + src8[260] + src8[261] + src8[262] + src8[263] + src8[264] + src8[265] + src8[266] + src8[267] + src8[268] + src8[269] + src8[270] + src8[271] + src8[272] + src8[273] + src8[274] + src8[275] + src8[276] + src8[277] + src8[278] + src8[279] + src8[280] + src8[281] + src8[282] + src8[283] + src8[284] + src8[285] + src8[286] + src8[287] + src8[288] + src8[289] + src8[290] + src8[291] + src8[292] + src8[293] + src8[294] + src8[295] + src8[296] + src8[297] + src8[298] + src8[299] + src8[300] + src8[301] + src8[302] + src8[303] + src8[304] + src8[305] + src8[306] + src8[307] + src8[308] + src8[309] + src8[310] + src8[311] + src8[312] + src8[313] + src8[314] + src8[315] + src8[316] + src8[317] + src8[318] + src8[319] + src8[320] + src8[321] + src8[322] + src8[323] + src8[324] + src8[325] + src8[326] + src8[327] + src8[328] + src8[329] + src8[330] + src8[331] + src8[332] + src8[333] + src8[334] + src8[335] + src8[336] + src8[337] + src8[338] + src8[339] + src8[340] + src8[341] + src8[342] + src8[343] + src8[344] + src8[345] + src8[346] + src8[347] + src8[348] + src8[349] + src8[350] + src8[351] + src8[352] + src8[353] + src8[354] + src8[355] + src8[356] + src8[357] + src8[358] + src8[359] + src8[360] + src8[361] + src8[362] + src8[363] + src8[364] + src8[365] + src8[366] + src8[367] + src8[368] + src8[369] + src8[370] + src8[371] + src8[372] + src8[373] + src8[374] + src8[375] + src8[376] + src8[377] + src8[378] + src8[379] + src8[380] + src8[381] + src8[382] + src8[383] + src8[384] + src8[385] + src8[386] + src8[387] + src8[388] + src8[389] + src8[390] + src8[391] + src8[392] + src8[393] + src8[394] + src8[395] + src8[396] + src8[397] + src8[398] + src8[399] + src8[400] + src8[401] + src8[402] + src8[403] + src8[404] + src8[405] + src8[406] + src8[407] + src8[408] + src8[409] + src8[410] + src8[411] + src8[412] + src8[413] + src8[414] + src8[415] + src8[416] + src8[417] + src8[418] + src8[419] + src8[420] + src8[421] + src8[422] + src8[423] + src8[424] + src8[425] + src8[426] + src8[427] + src8[428] + src8[429] + src8[430] + src8[431] + src8[432] + src8[433] + src8[434] + src8[435] + src8[436] + src8[437] + src8[438] + src8[439] + src8[440] + src8[441] + src8[442] + src8[443] + src8[444] + src8[445] + src8[446] + src8[447] + src8[448] + src8[449] + src8[450] + src8[451] + src8[452] + src8[453] + src8[454] + src8[455] + src8[456] + src8[457] + src8[458] + src8[459] + src8[460] + src8[461] + src8[462] + src8[463] + src8[464] + src8[465] + src8[466] + src8[467] + src8[468] + src8[469] + src8[470] + src8[471] + src8[472] + src8[473] + src8[474] + src8[475] + src8[476] + src8[477] + src8[478] + src8[479] + src8[480] + src8[481] + src8[482] + src8[483] + src8[484] + src8[485])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255] + src9[256] + src9[257] + src9[258] + src9[259] + src9[260] + src9[261] + src9[262] + src9[263] + src9[264] + src9[265] + src9[266] + src9[267] + src9[268] + src9[269] + src9[270] + src9[271] + src9[272] + src9[273] + src9[274] + src9[275] + src9[276] + src9[277] + src9[278] + src9[279] + src9[280] + src9[281] + src9[282] + src9[283] + src9[284] + src9[285] + src9[286] + src9[287] + src9[288] + src9[289] + src9[290] + src9[291] + src9[292] + src9[293] + src9[294] + src9[295] + src9[296] + src9[297] + src9[298] + src9[299] + src9[300] + src9[301] + src9[302] + src9[303] + src9[304] + src9[305] + src9[306] + src9[307] + src9[308] + src9[309] + src9[310] + src9[311] + src9[312] + src9[313] + src9[314] + src9[315] + src9[316] + src9[317] + src9[318] + src9[319] + src9[320] + src9[321] + src9[322] + src9[323] + src9[324] + src9[325] + src9[326] + src9[327] + src9[328] + src9[329] + src9[330] + src9[331] + src9[332] + src9[333] + src9[334] + src9[335] + src9[336] + src9[337] + src9[338] + src9[339] + src9[340] + src9[341] + src9[342] + src9[343] + src9[344] + src9[345] + src9[346] + src9[347] + src9[348] + src9[349] + src9[350] + src9[351] + src9[352] + src9[353] + src9[354] + src9[355] + src9[356] + src9[357] + src9[358] + src9[359] + src9[360] + src9[361] + src9[362] + src9[363] + src9[364] + src9[365] + src9[366] + src9[367] + src9[368] + src9[369] + src9[370] + src9[371] + src9[372] + src9[373] + src9[374] + src9[375] + src9[376] + src9[377] + src9[378] + src9[379] + src9[380] + src9[381] + src9[382] + src9[383] + src9[384] + src9[385] + src9[386] + src9[387] + src9[388] + src9[389] + src9[390] + src9[391] + src9[392] + src9[393] + src9[394] + src9[395] + src9[396] + src9[397] + src9[398] + src9[399] + src9[400] + src9[401] + src9[402] + src9[403] + src9[404] + src9[405] + src9[406] + src9[407] + src9[408] + src9[409] + src9[410] + src9[411] + src9[412] + src9[413] + src9[414] + src9[415] + src9[416] + src9[417] + src9[418] + src9[419] + src9[420] + src9[421] + src9[422] + src9[423] + src9[424] + src9[425] + src9[426] + src9[427] + src9[428] + src9[429] + src9[430] + src9[431] + src9[432] + src9[433] + src9[434] + src9[435] + src9[436] + src9[437] + src9[438] + src9[439] + src9[440] + src9[441] + src9[442] + src9[443] + src9[444] + src9[445] + src9[446] + src9[447] + src9[448] + src9[449] + src9[450] + src9[451] + src9[452] + src9[453] + src9[454] + src9[455] + src9[456] + src9[457] + src9[458] + src9[459] + src9[460] + src9[461] + src9[462] + src9[463] + src9[464] + src9[465] + src9[466] + src9[467] + src9[468] + src9[469] + src9[470] + src9[471] + src9[472] + src9[473] + src9[474] + src9[475] + src9[476] + src9[477] + src9[478] + src9[479] + src9[480] + src9[481] + src9[482] + src9[483] + src9[484] + src9[485])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255] + src10[256] + src10[257] + src10[258] + src10[259] + src10[260] + src10[261] + src10[262] + src10[263] + src10[264] + src10[265] + src10[266] + src10[267] + src10[268] + src10[269] + src10[270] + src10[271] + src10[272] + src10[273] + src10[274] + src10[275] + src10[276] + src10[277] + src10[278] + src10[279] + src10[280] + src10[281] + src10[282] + src10[283] + src10[284] + src10[285] + src10[286] + src10[287] + src10[288] + src10[289] + src10[290] + src10[291] + src10[292] + src10[293] + src10[294] + src10[295] + src10[296] + src10[297] + src10[298] + src10[299] + src10[300] + src10[301] + src10[302] + src10[303] + src10[304] + src10[305] + src10[306] + src10[307] + src10[308] + src10[309] + src10[310] + src10[311] + src10[312] + src10[313] + src10[314] + src10[315] + src10[316] + src10[317] + src10[318] + src10[319] + src10[320] + src10[321] + src10[322] + src10[323] + src10[324] + src10[325] + src10[326] + src10[327] + src10[328] + src10[329] + src10[330] + src10[331] + src10[332] + src10[333] + src10[334] + src10[335] + src10[336] + src10[337] + src10[338] + src10[339] + src10[340] + src10[341] + src10[342] + src10[343] + src10[344] + src10[345] + src10[346] + src10[347] + src10[348] + src10[349] + src10[350] + src10[351] + src10[352] + src10[353] + src10[354] + src10[355] + src10[356] + src10[357] + src10[358] + src10[359] + src10[360] + src10[361] + src10[362] + src10[363] + src10[364] + src10[365] + src10[366] + src10[367] + src10[368] + src10[369] + src10[370] + src10[371] + src10[372] + src10[373] + src10[374] + src10[375] + src10[376] + src10[377] + src10[378] + src10[379] + src10[380] + src10[381] + src10[382] + src10[383] + src10[384] + src10[385] + src10[386] + src10[387] + src10[388] + src10[389] + src10[390] + src10[391] + src10[392] + src10[393] + src10[394] + src10[395] + src10[396] + src10[397] + src10[398] + src10[399] + src10[400] + src10[401] + src10[402] + src10[403] + src10[404] + src10[405] + src10[406] + src10[407] + src10[408] + src10[409] + src10[410] + src10[411] + src10[412] + src10[413] + src10[414] + src10[415] + src10[416] + src10[417] + src10[418] + src10[419] + src10[420] + src10[421] + src10[422] + src10[423] + src10[424] + src10[425] + src10[426] + src10[427] + src10[428] + src10[429] + src10[430] + src10[431] + src10[432] + src10[433] + src10[434] + src10[435] + src10[436] + src10[437] + src10[438] + src10[439] + src10[440] + src10[441] + src10[442] + src10[443] + src10[444] + src10[445] + src10[446] + src10[447] + src10[448] + src10[449] + src10[450] + src10[451] + src10[452] + src10[453] + src10[454] + src10[455] + src10[456] + src10[457] + src10[458] + src10[459] + src10[460] + src10[461] + src10[462] + src10[463] + src10[464] + src10[465] + src10[466] + src10[467] + src10[468] + src10[469] + src10[470] + src10[471] + src10[472] + src10[473] + src10[474] + src10[475] + src10[476] + src10[477] + src10[478] + src10[479] + src10[480] + src10[481] + src10[482] + src10[483] + src10[484] + src10[485])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255] + src11[256] + src11[257] + src11[258] + src11[259] + src11[260] + src11[261] + src11[262] + src11[263] + src11[264] + src11[265] + src11[266] + src11[267] + src11[268] + src11[269] + src11[270] + src11[271] + src11[272] + src11[273] + src11[274] + src11[275] + src11[276] + src11[277] + src11[278] + src11[279] + src11[280] + src11[281] + src11[282] + src11[283] + src11[284] + src11[285] + src11[286] + src11[287] + src11[288] + src11[289] + src11[290] + src11[291] + src11[292] + src11[293] + src11[294] + src11[295] + src11[296] + src11[297] + src11[298] + src11[299] + src11[300] + src11[301] + src11[302] + src11[303] + src11[304] + src11[305] + src11[306] + src11[307] + src11[308] + src11[309] + src11[310] + src11[311] + src11[312] + src11[313] + src11[314] + src11[315] + src11[316] + src11[317] + src11[318] + src11[319] + src11[320] + src11[321] + src11[322] + src11[323] + src11[324] + src11[325] + src11[326] + src11[327] + src11[328] + src11[329] + src11[330] + src11[331] + src11[332] + src11[333] + src11[334] + src11[335] + src11[336] + src11[337] + src11[338] + src11[339] + src11[340] + src11[341] + src11[342] + src11[343] + src11[344] + src11[345] + src11[346] + src11[347] + src11[348] + src11[349] + src11[350] + src11[351] + src11[352] + src11[353] + src11[354] + src11[355] + src11[356] + src11[357] + src11[358] + src11[359] + src11[360] + src11[361] + src11[362] + src11[363] + src11[364] + src11[365] + src11[366] + src11[367] + src11[368] + src11[369] + src11[370] + src11[371] + src11[372] + src11[373] + src11[374] + src11[375] + src11[376] + src11[377] + src11[378] + src11[379] + src11[380] + src11[381] + src11[382] + src11[383] + src11[384] + src11[385] + src11[386] + src11[387] + src11[388] + src11[389] + src11[390] + src11[391] + src11[392] + src11[393] + src11[394] + src11[395] + src11[396] + src11[397] + src11[398] + src11[399] + src11[400] + src11[401] + src11[402] + src11[403] + src11[404] + src11[405] + src11[406] + src11[407] + src11[408] + src11[409] + src11[410] + src11[411] + src11[412] + src11[413] + src11[414] + src11[415] + src11[416] + src11[417] + src11[418] + src11[419] + src11[420] + src11[421] + src11[422] + src11[423] + src11[424] + src11[425] + src11[426] + src11[427] + src11[428] + src11[429] + src11[430] + src11[431] + src11[432] + src11[433] + src11[434] + src11[435] + src11[436] + src11[437] + src11[438] + src11[439] + src11[440] + src11[441] + src11[442] + src11[443] + src11[444] + src11[445] + src11[446] + src11[447] + src11[448] + src11[449] + src11[450] + src11[451] + src11[452] + src11[453] + src11[454] + src11[455] + src11[456] + src11[457] + src11[458] + src11[459] + src11[460] + src11[461] + src11[462] + src11[463] + src11[464] + src11[465] + src11[466] + src11[467] + src11[468] + src11[469] + src11[470] + src11[471] + src11[472] + src11[473] + src11[474] + src11[475] + src11[476] + src11[477] + src11[478] + src11[479] + src11[480] + src11[481] + src11[482] + src11[483] + src11[484] + src11[485])<<11);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hcd20e48d0da7ee6764e8531ad7599a10236672f0356c5fce70250d46519859678d365483c971c3decdc04a2c6507e86394312bf377207c1cebf4eaa4c02d02980207bad070da5db648da0b2138dd2640f8e87add7e4c864b8abf4229d6e2146e57cc249639d85242775c9467132cfd21fe3a2a767d99d82c4034744fbbb04fce7a2009e303dabfc055df2863237eb95650f486c88dcec09f4bfeb73c8af402102c538e5fdbde4c107f94e28f31f1e3bb52af9dee804fa69c1034eb9694f04c493ed96030d9a6e25989b66e7190aa6a189d0b5e00bef36229469bf3a14f4063534f8e737bd041374b82dfdeb8e0d88584bed8b137835d4e91186a0b544dccb84e7df61930153999352619b46f31c1d3a9522cde7ca9da5474506d31229c25122bb57e0ce07bc1b2e27179876fec10bea639b0c41b022e77b86a7552b125618a47bc8e97491155317af9f166723ac25768670af13b2eeae32b186c1f943c6e359c0c6c528a94c0197b8e9c9ef955641ae38be74e18a2a03100e82acd0c26b8ccbb8ad3bd469938f0ea91c35268338c1421635de47271fc117a6736f56d91b074fecb0717005e5a6fbdad68e486b308ef47fb8bb2f25250953b0bf3c026427272d8a1818c04a91e2b5e835f973b863deda7c84828bf90fe03273d056d204645afe2cfed91229e8e47bd4b3c1126452db2c813c4c34c5dabd876d13fe0fa21805026c4753b600881388fc7f5449aeed7735c4660726cfaef39e93c6a40dd70a69c98af076e7d83df1874d96e8ba5e7a58f1d48e28c0019c2bc9b83b5521190e011296d25d6d51d7580a2a7bc8f25503aa607325204cccfc253dabc25388d61dd4acc0240c003a010f354a795cd48ca526ff07f4ad9fb29989b6fe792130eaec077b407f56a8df4f3773185fcb17b17225e1df10525778e82fa82610915573331b4239390c25730886376eb5debfe031038ff78c22fc66fd32e240e63854da3289a3024c87ec322df203595033e0f842d075ac9df5000093bad8e07;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'haac899394c10706748bd986387e8756e4fd7b2c248a022deb593664bdc399b3dcde993c50a068449b75df8f8d83a950116cac64f1bec869b04c618e496fc6c92906232ee8cc60fde9bf9291ab215d4e6417b07b1d0c6b68ecff05ec8c40744f85ba2386d527b66f2a8bdd04a3d1016a8a26570f12da1aa85aa1ae5e774a9af37b8ba9c7aced7a7a1d5fd69d6dbba04241c45a78f89237f32f0e98bee465b43cca97ac955e9a203a33dcbab317bf6f4bb036df288d58cd518e0db3b62d020e420716cd3a009eedabbe3d292dd43051f3b22fde6f4c56d9787619ae170e279c5e642306acff95c9dca1759714632f5b5f6ac0a06666d6b512c8815839b7162c6651e648554927d51ce4596ed4cec95c47609ed2113522d040901a4b5dffde4136a34a4693bfee79fe808de20fd209caa6cab1c97a489697cda67e5b129dd8bafb77e2f51af37b4ec085dbcdd83bf6b72a8698b121790ef7c3d7524f96fa25495f4b6d978cab75687405ad1640403ef6fcfbfaf5365de132d65b3d681f3cc354be0ad8da6b047110fa214e7e7e810b738ad9bacdce08f48701696c7f7b76c3bbfec1466bd46db4c48e31de2c690b6688b546d8808424821a1b2b0d2539d22b2998d2ef015828848f211f1eec790917b04c5c1f8707189a551d44c30761bf29e22955b4eba778f8edd6051ca99e1a05679fd203f448dee2be49c750e8a48b84064349e97cab85f52b30122a6468edc68a07ea7cfdbe17838acbb21a1684afbc75d5fe70d2ff270bdfbd084666a9de06bf27372b6300b9bd9aea9a96c8e446942d42605e944c3282e0e3f7d1b523cb0678b694ac80ab2b65e86630d0019acdd1beb7c9a952fb1b9b6230ca5a7242206b720311f6764f6fb85f58ee7b7c90b5c67d8d1881958b97b834009631ab70fdd5f6e113611f5de5e612414f92c263c0a6befc6e769c411fb0236e4bcf1c8b231ebe415090e7ee6aecf4a8b37f3cd9cf35d64eb060cded65350f03f4e573febd13c11b6dd3ea85ea0e42a35f3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h3556de12cc5021ccebe0ecbbd8fef506eb575efc382b1aa310648f6a8372d8f16b59928c46cfedf436a0912d36e453ee40f3468c61443a94756a28d28f2a243e38721d215715af1e5a557d7f261715dc17b4fd8a33e2382dd2d7daecaa4d66b87857526cbc74baf2f3ca2d0828cec2a8fda5fedd92733a49a509983a69d485a4fe9c3dd130f2f1a03d84571a23df0faf08b943fec38628775bd88adee9e0ef270f7b99474fb8bb2276e29dde2b0932d35dca8f3c902626f5279dadd7c4ebb384aab4a34beb4d0e9f913adfc35f21db982f0ac3e671b7f0597066b3f4cdd0a3eb8f72e1f6dd7adeb7ed681508e0a61ea4e2f7c73ba8f99d578420691133b5a64f2b61322f76ecd1a4d973550e70c55e1a2616a06570a20ad887f32188cb810578430ba99d42036b461933af58da5456217b9661cd5f7ccc0f6067dfee803637b508d9c75ba3023380cbad4485bfd01cc93af10db2db08af08c7dfa17de33088720423450c026a1ce40926f71b184dd3da37d0d1416cbc9dca3014503a5bcc1e76768cd1953659567839472bce1cc845eb27ea3de93b3f848312c40f89e7f6ba203264e0acf1fdd321ca79951c8e9ee29e7e4977861a2488391211e5b9bb145cfbcb8004b4677d698b26825da042d061965578430bd4bff808a4dd15f32d797257fc67e8e27320e74995c017554414109e6a170dfd8be713de3c77fe136e8995e435eb2198737af3d78955414817be9d444a1d5502f65240a6a93f4179f9af383edc7e5969f71df472c76dacfee1758cdc6e8fa0241db447fa10893f3f80757baf20a589d774ad6f53960860aea78e11728a495f6013fcd4c42858ca480cc26908c0ab17b190f8eaa283e9ed79d18bdcbe87632e851b45ffb383c5920223631fbc034e96967f0c190ce1f09357f3dc6b6d3f9b8fc61473ce6d079741a2d63502333fed2a6786ae1c77943a15c1f12a68c7d0c1b1ede103278f5d418c87570d316d5329ecec3cfc0e151489070d1228542f1dc70c00076237df25;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h6d8b6bfee89ce4089247980b20ed154eb0fe76935cb2f0277b760258387e27a1f2fc6c4485ce92b942ea0a69c7407c78f12b5a456cc873fbb1b8e2ac654346259a2b3cd9bd8029dfc6c64e18c7b4422a11c8d266bcacb506651fc6749b635ee8d8bf74e74b3a978dc8a119e3cbd0d8c07f9025aef7b330eec8db023948c3a7a94370e931c62144dfe2e64f7baf04e5ed8383cd377e61c9f98aec8659e9e982eca1f96f92d6a9c22b323dfedda07b040188a6314c3eba1ce39ec868890a59eeac0ff9daa0f88a68659d5812096250bcd5f16ddcef25386312ad88fb7f7bb418318121366a5a008f7f13f84172f8e2a4bdb981b0918b17548c204ad04ee70f7bb1afa1f7f145ed2b8eeb12291583afe305e2e9378f75f5b2e2e11d0d8df86f9b78b7c30261c96aa1a5bfe385c39aa8cea1a4307b25de8afcf06d77fd367be799e119685175814dcceecfa06413fd853e792c0cbb5d3dd6c2a3c33648de3c8a701efa1ef3c906d0123d654d389328d2d1afb08fe08cf1469ded9d3343bf120cb1ab7407bcc1b5dab52c394c056c390b19d12da32c3d36254ebcae8adc1e85c574026199e691377822eb7165afd7f8f384ce50019abe022c6d7d38ea168047ddf381e4101028bafd1cb62ebbf709dafa0dc9b3d46f9fbfed1880f9498805f0840139a02f678651b23763385be5470ba61ac6e84612d4f20842b40c56d0c75e80fab2e07611d5c19418a69432d012fac8490db0ce44479da552412ad9c42c1f9481cb7c56d9999c30c4f277a20f5d01245ad4b924e27cda368130d56741b819cefca4661c18fccaa47ca97c7d28a0ff178128a8634b66c9676ae8c92f0fc8cb354f09c03a753518b7e80434ac8e82c7a11f64e1f263d02644e82c788059285f504a92a637c43e5102e508c8377079e22fc05d635db68cd53ad50056cd1d8e15d9efcbb67ea2372650b4c05e08f45a834f6da37e8763f03366f98309a5a368c74b80bfc263b81f122f58ccdb0a023a9fd7c9864ecfaf0213d8a79439;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'ha62844d64140bc0d244e004a9a08f658986f161072d6a669eba57d15d88b984332b989ee2eb599d31e4017b1317f58466196dc6a267133c4f6436a038745e1fe1a7a52159ac32853a55b74f315a3339e1ff1295a78794b5c13b84f14df81a582a56712bbae33304ab50284b6b3140ea628ac0915753825c54167f1e21fe4a794e56f87ab5660fe5ca9d09a7e72c71d4dcd0807c3eb6c7f7df5933ecd1cb42229a24130b3c4e53c7ed516992fc3451c458731bc2a40fb652aa27c92f054f57d2f4d0223e18010100994fd0f9ecd3aa70a1bf300d5d3859b849b2f7cd496861439a405fbb6dbb25bc6c6eecf53e42c92c42d04a3719381adfc8cb243ff9d8994e20555e2c9450eae74eb40184564933177ec62d15a05af1e820d0405b3a44524eddf0a67512de5e31a618cfc32d51dc23332b84088af0725f3d0bf4ac7311b5699d809336510533043028e75a77ef4752735f4c174cc8ab24fd406857616c5510a3e5a32e4bb4cd6a5be55e20855022a77b6b0be957396406510e428161ba0e9b378ef49291bb16d90cc0377a1e435a537a440ca5f829eb0c1ff5ae1b3e7959037e68a14c5424095a88c238a5d25de17d9442c30c42e7a8ae73fdb25789f7cae8bfce24bef34911b12f9c6513a4a6941539916ba1119e9ef10b84e4bbaac38a6071baedf926c0e9ccfd748bf777ecaf19857943d76c07c41cde57c3c653979d7c1d811e0eb34d28051ff2f7ca48afbd088e23d68c27b131f95ef065cc55d97d7350ac2b25f2739f1351f67d23a2d4b0eac0282a9d6c73d9ba67e435e2225223bbb090cd6d0c45a6a763c9ed1dad434fb5a73e9d0f7ca4d200637b466d288e289ac81de50b098f05c801e794f01220c1b0ef51c446ee82d453c24619513c317a2ae37402ae01f44ecaea12e24b9cbdd35ff41dc83d6ed079128fb50760bf3408a62f5798069b71742c2ac362c163cbb1f707a7d3ec1f64294378309a20cc6e530cae1b7e5d1763b2cad07fa9f3dcdf9d1c2a0e5c33404f2cf825e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h7e9e0ba49b5ffa520925d759ec537bd5a370b640cdef4b5289094cc9df91cb5a829f33197d3819fd5771227e6b082f0c5bac5505f26e0da8f8276f14f10301452d74e28cf80b45331d166edcf4691d65d322db4091927bb087b09a51c269fc9cfc590df0cef42494b06c61edcfb8f7b581075a424465576f345366b3b10d2a0ce1dc2edfa26747b4132b3eb7b250af7c3e3defb048cb3ccf4f8cc4d552142574b6d019b33f1887b03b20345f0fd48d2a1061326a13a2a22f8d2b3cf67d3a5cb04471ba4b7fd33efd8dc04d1cc6e898c99322897a23668333e25715860a6eb50f44e7b92c48eea7fb115e9b4f83e554240b3034b6c9d675b48eba9f6c21488c60ffaf0f7718da6f90f871b3a44abd1446fd82cf2e4a575f6e6ff5d89e6fd7f6278b522f6643016a4b7f5b14e14ab23ffc6424a0b21774285652ae2ecdac7ddb3944320ed03618d07c434b04fc036a43ddbd0db1a9a8df12787cae39c216621388dd4cca339ece58be6b7349f295167e4c5ffa054fea22be72db3d59c5bed5e6beb477ec27a5b6e1eaf0b43c806a11dd66789f18cadaf3dff26b6b6d23f141bcea2357fd79dc199877ae7f6a6e997528741aad36e9944080dfb51935e5f90442bd3a58893a93fa24bd69a2179b619e1b309e3bf699607f3189b06e2cc2a23a85e691000ac0d4e259e0b973c7389cf8256d07b369507d4564c0bcaf7ddae1eeb7d2e37ccae900b856783e1ffe37944f38b327278d27c98acae0c676d87f3a2d59cbd2eed1810e90c8d8d4f781b387ae55f89189aee470d6255a4a55118eecf1a587d62cd7977713003b7b439cf76a0702c5c2a5a2dc6fe46e89e67ce1ea0ccb3c55a94135bf4f6738f07511fb5cab726f07f705654c8e297e159833e756feb57d1191244a49e002160541d033fccb8a42bc26d5e0407cd5f1b2520b0520af97a6af4ce3b2e855e0f0dfedceb76a3701c9340a90ad3ddef5ccb471b56f4b6adc5a0e17ec9373781d52a00782288d92015f392587b87dc7618023c1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hbb4d3411670414d9c884c656555f75a10b7fcd245357b927237749d7a990fe58a4d06c496249bbbd386bcd858b65edb2670f8ee05efc4d3a9e17f0dc4b73688f4810c10c6baafddd323ff8919fd784477d700d3310b771169e71a0e823abe598cafbc08cd560313adb1c8c3aab34558dc3c82ae7ada7459e7cbf47fa7d71e8cdcc199cc67b21267178f5db2109509eded23f54b482f94a1b8e08e86eabbf237e7aba79a17c93809ffcf589d361d40e20fbd5008cf3c85a22bb03e06692f191dad515496798c58486a09b3e1400cf4c996d6f32c4403f996e3898ffadfc314ffc7ac2062a3eecc57e6f6e6cf9282a9b707e0a9b3c60620129be485ec118a21d71ef03e452c50f12563875d7e9fe4cb6eac278d2177c13f01f1fe57f6a4a2fc7053a51a42544c8c57eab941c223889df687126aff2f52ff2e44b5359e774a3aed0e80dcf5965c218ee139461bc9a8f082c76ba7334fdffdfbcba9fd99f9e788750ccb7ff4a748bf4d0c67d08dc6804ce30f8d58e2ce7f270ecd1ef34db8176d625465848455b348215b4948708dc7fa6fe45bef59d288c812c0dc73d29c5d2120529f42d11393316a21bf387126ff5d09c24b74f1259a77b22fcf4eb3afa4cd834b954d2bf59d2c76d5643fc1edb954f82089ca784267dd097b668a9ae1ebd593c4bde229a328c253a3359af99939062dad370c9a6ee481ac0eeeaa0edd4d261414abe1455b0c205b3c7f8a04bf449f69f0015d514eeea30095dcb4df2744d575be82af41cf0b4c5ee6fc8012e6e9a5a499d2521837fe25492cb728638e3ed0189eb864da37a32f7b15af836eafcba769f9e722a16819703cea2002c3014342c89826f6488fdd9efc368cd1f1bb3d3b8757c59bbfd50b5e6f608e2a451add38c8a877e6fbcbab3a393ba445f16c7a82020ba7fa9f8e54b3f53a7c672ed93cac96a9afbf95e256a1b85d312f39700cb17f3312c185e8c6d54fc08424ed2a7376326bd60347dfafc9ddc5c5931093f9f15623dbc43c21a692a22c3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h455dbda3efa1ddb161ac918c85090c6a68c94ce516fa9dbf7d06b35ed0b0aa07f06e143f4eed972ca1a141093284333644f338c2b3ce65332520c954d30915fe8818b2cff0b50f554c2626d0b709ae4821d07b40b76b286979de7caaddf00bf8292aaf1a31880e9f69a60b36ed48f0d182ae5f90834274fdf56fa9e2f91974faaf9f6e0ab281f946897b077d3eaad96a96c4b9e05fe182899b1a31cdc448744bcc26e17649568b349797d56ddf4a5bb6fc28918bd7a7b4b672d6a63cced2f3b1378649e39981b66841353d5913d61941785f133aef73dd709fa90462c70b3e49622fc6f3650488ce038d586ec84577cb0853543b48993265117fb8a344bee01321560dbc79cf77c12de2bfec9a0b8ecc5d53e17e00f51f3e32e13b64034020b7bb2ece0ab7e727153c2295f70a2dab0c35dba8d22de0a070fb4a424c0a73bcd57d2d397d8e614517b5c07ccdb66ef1868fc8eaf1936ac638db78aa51871245f0709135547f749d007b594c6dde34354822e3e8b15b19b60544d2ae1440645acddfde871dfda2aefedcfc0ffd46b77f905d3e33924330302335655d883530b8e0965cc2dc3822544e02319c966715770711f36cb2f6c0a0573b25a22080bfc612f4d2b4676154da642366f8ea554465e424a0bc1fa976ac0b11354dd43bf105421a84175edefb99609df203d53dda0d7e7244322cfc92d3ca85d06e8dc815631dc17199f8be37d8fd93aed8f840108b32b03204e2745fb73d93927bbee638b121f2d70790ffee95c4b7e27480c29301a5100c589f58fe018f870e3a84e858f1de3ca23d9b108e89daad9383bfc6c1cc2e39e840ca18537bee3010e6cc794679e1a1ecdd109b302a4d8f7d68d33613a9256033ddc5798fdf2eaaf710a0ceaee7d9a96954c4e46683bfa762c7b152edd605252acd89b981aa26baabf6c04f69f02384cf97fd868eae2efe6617125d27ff2c9232fa9ce6cdff0e230f7ed49486d2ee0799b751dc4d1b0bfb2efba2030920a55e9bf81cce9b70809a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hffe550570e188037ec8994627bcdd90a711ad5731c88b26cf310df0948e9de81ac8e6661ac36e366917382d718a68d9d1f20800224de7b727d2c85f60cae9bd321ca801a2c122ee7965ccc81bc8f157c331aec4b7b2f2def5e393b5350078e7ea169271ab9edae85c49db4778647b507b72854469778f6080285aba6927ff6c4fbb907ce452fb8d8c0688753411cb00f17dfc9a5fd6dfbd1d0631451aff6957da3d17c2fe509d9120a0970286df606291ad448c799d2cd6d9ca837370abf67a86f4a10f75435d7c5bd24a295e75484da650ea08d8bffa37e0f902ec5fff1c126699d1211c53e3d576f144b477b58c8c73d2a2c37a5148fbdbbef78fdb5fff74d525b8c5bd9dd8c269b64deca0dd834aca6e374ae07b1abe461749fa443ddd7d7993336572506f3ae04a82ee0d33e90ad9f4c3aa6d3787119e0a0f3ee5d91ee0ff300a9888a1f4574c78d3cab15fa1cbc08647658222aa6bb4ac57413356237d7a7d9706785ed11413ec59e66021bedf050c423ca049eb497cf46bf4a1cdbb0854a6bc113fcc90cb9003c918980c76cdf3ba382442dc34f7b9c6e4c5a437794ba06b8e19928e42d2cb623566c850d92d4413a4ec81e4040801d2f752a32b695215b1cd7803bf2e34e61ae48e97a7d50a6a8a88aa224c2bf35cb678dcdcf518cf8e9cc3e25bd1ebbc19c213aa02cd85cc8c61262d9c5e4f22260584e35f7dbcfa3c28534086a7c64c3795f71c7a3d3c870ed09ed55e6f8cf158977041b4d1daa8825e835807ac31c803bf5f2f0414a2dfe5965e11a0cc88ab61faf973ca52cdc3049c2c582bdfeceb843fc50be904e2169ba2786a3a9804e42bb05136b866c1f342430db7ff6a4af068e7a205184479575e6ae935e4452e41716cdae261abdfdedff164ddc642f2918d318e0772f33f87b602b0360629920aabd2bc7a21ef114c0e6e110e019ea1a70c08fe2a4ae72c75d6f51fb828666badbc2808844a3e141da24ef340542ccf6107eee5c83fd387917388ce8146480f9d42;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h7a1ba12d390921215d115729c37f888418c1766b809e72df30e324e567b7378465f6b29469ce6719b5b2fcf890d8af395b3672956ce36a23fb4d324fa48111d973b77b690a5e89499fe01b8fd8c25364c27a0494aed47e3066ee8688d9b357a0e0c3c1af70e4efd51fe044feda15d8e72463e91b89c0113ba652b7574d8a081c16b5362b45bec2a6b6475acfafb634843ae6190866fce7fbdfb6f8e2e079cd4adfc9ed8272ad46e71d2ef02a356a8c1fe0484f2e001adaacb9d411a4f560b40ea22708e7b17b3f8260e41f2abe37add8c4c7296f3c3f92c315f42f206a86397a7e1a8ff42b6976dfeab9844a4b0393546176bfd05abaf998e75f8cb0f85d3c7b5867706af9439b9228ca6bf9a2d6fae88fabfaf178072f95687d7cf221dfa55232f050b65c88f92b1fcba4c3d7fe1606fe4da0c16caa91c32a51e665a7e91a0d15837e67257e3bdf82cf3424799d92efe7cf1aa4e2166b6ab4264e29e2ea1c9086d3d41ef56f7b0a9011092723820d19f4ae13f18a269a1041da8ae59e5d5753e961d975d713042d985f57a64304917b798d8d14af254680164adda91b3beb4c6e978fbaa9454d4c02cfb1f87b71d0a222f9ac413a928bb30b78a7594ee18d524cf548e5226abc88106960340702d0cd0492cf96b33c517770c9f6716d1a9f87ca65d67e9b5671431c4b44bd324563ce32d891eb55a2e7f1451f8881b4f30e707077b57b38d6db0956c54aad4e7b40d0355279f1ee2776075755da6e59cca68e384b971e319cea16c31ac72fc3f14641571364a19265e7713ae0be399b1fa1c9d322c33788b4f045d5c0b9330985514df32cb792d6fd691f03a83db48e212e845dd1ecf921dd3c1a1e64813ff072b9f910f5a134be0cbebea1b6813813b817fb8e78525e2094b204a1458aa9d6996b70d51b73c27cbee794e6edfaa297da72914ffeeb98e90fd4c33132bafc4dd49381a5c92ecdec7791a77169e248317000dfdf6becf2b2d469e371f8855cfe2106512efb0e5dd88b48dfb1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h2db0aa88e177e040113cd2bec70a8b95a9e5b9b1fe9ab34d0535db8e237ce5e4dd34e546efeefc01774c8869a6eb1345346775f8607894caca2d0a550f40d74dc6de465b790dea15bcc8c32a9581a9612eb93e1dc371f8b5d4703e2b07fbd9384305443262040170d7e5bc68e8a2ddf435b0fc3c5e68f5b742b6853559cd31222eeb167cab7b3045b7199d4c5b01043d75e4f33af73fc6154a4515dd16596b530950bfff1d17b5a36f0187837dcf47897d607e2e9ea68b7f97480a434cd9523aa1cc931ffdbd45ced1bb49a7ba14a6e3dbf663ee72221f2f16207fd976293219a433a0f0835e2f05f2aa968b37de4f13965b879591ea0fcca7994eea86036e35515783bef2cde35f12e557b298ebb356067233a024c10f2e963f3947a5ade5db121bee92aa05fc62bc8e3797a00ede8c3475a07274ec8598284ef1046dc1774db78f6e134f0548380debb73d7454d797d9ca09ddfb7133679f93242162e8de99eaa28ae323b57a1a3f76da068818e8cd5e5a2337b369d22729be6c409529855bbbb1b77be87764ad088574d9fcceafbdb467aaccb1434987e9e68f549dda9e3d7608c199bd1e17721dfef85802f9b30104aeaeba0d46d3743c2009f5bdaf94890e8652f1a0139a7228d0c57d47f46edadd4f11465b3d00fdc326f9b84051c4ab072ea03be575cecf6cefd0708552404aa43e58dc56d02ca6a75fe705bcae8726de8bc2564fa8be36ab4020a50275cd429fc96c8f06d5db4b861f7a9de58d8b92e2e3b64ca62c07d59f2b199db23776e39d41a430293a42c00627cca544037d1c671728eb8a4278185b207073600811a63d23d03c49e70039eef5390b3c57e8a143fc828e370f07639e574afecce5d2c94d2ddf6f13ea5a7f44fa27048578c9370691e91e5892d139ad541e94d0337e181e15999356e736930aa1fa4da8b9df33764ad4ae05f72a79b0ec7b5b393bdd1b1c8949ececd1339d243b57d3988da0bb7b71c068bfd9c1941fffd94fcdd8e412984a841576241ca75;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h9005b3297f3e77b1d5df8fa4def793261688abaa9df6fb5af45f12e0d802c948ab53d438f3286ff8187429e766bbc20bce9ed87ff1ce2f6087358fa2e9cd006038ae86d91c75d3f82f1712c812aaac09d5e33f9bd78b5fbc0ecb53a98ef84897e28194158d5f0f0ea65af4f582fd969b71571bed6f468587e45cc0971f75c8075834a806d9cbc91960677fdaea10a59ac926a9b92c9082afa89b2d4f28579c181178a0b56eeddd79840c3ad65d57125dbb16f313fda407035531679eb1c86f618cc5b2271f94f635c0bdb6b5b237ac7e76eae7f9d5c5f7a46297fef44116a5c276ab83ce416df8d54147623c530972171ba55eaf70886bd96828c9e3cfff18c699dd0f8c36acebe749771a1832698ad992b2106c77d112c25872cf7630b940cdcaad20f442b900c380e86c1b6e100deb908b94d166e3a8b81524e58c4a1979c26cb51080b1f24c3e2981eaeb158be35a82baee69853bc5b9f79095906e8572d4606a3af3545e94b6574c3b8cfb9dfee17b8c1748adbab7e6ef21e71e0c69c37e251d3e69b435315eb2958641e6619438fac30113e6beada0707d78d56bdfecce07166fd9e99c69b6450b1503a3063a94960d69243c0bf1eccb81283b3c8886722b983a8ac9482f477bf04ecc85f7ca8583f7d0cb81a89e19277302ef04e853178efe9846e94c4557eda096b49ea9086fb29d5c0611388948687df8ea2431fc1cdc27069f5c9c437ce85d6c33ebbc024160812d05fd5783fd48b6cd4c8ca22d608f658171a6d0217a89f439f7c45e7959b0a572d4919a872237671b0225f6c8aced6ae0b5dcd66d37ec231598f18d50d8137ac9809e333ea7b46d07623b0644d1b9a3d269311f2795fc1e5437a2460954f741be5aafa1c9e68b864137c9810d00c336f71dbe339e5c277a659b23143a030819dc618aed3bf37889e0416dc9207ca8b7f332d621b591ad18b60f3d83333a3e477ab4846247610895bd9b971a5bbb2ffac42c0287fdea1ea04fd9b6c791ceefc16e91d97c1b2699;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h5c169e92fe78f142688b90fe08a7b480e90274804482eed7bb3c753fd338b91caabe1204542aff94760bf93e74a34b6560d9b9f86a46d5030ca553068a1f60586dc25f08bffded65b0a1633f19d9ecab7ef683f04567a070d3d90f5f58cd26b2dd54692d2056ad404bc264e17664d246014ef3e4bb961708c4f8805d7749dcb4c242563ed2cc4273e9f68fe67b0a1c21a9a9da5b4422a8fb967a71ffc0bd1027e5890bc675e2b2b75a57e6e9a0bc01d41ad902a3427b3ef542ec49dbb60c0650fc13ee940cd7fc181b0dbaf7ab81aa500d406563b047b2c501c982d518b2c728ba08828c7e7a33e5096356849f8c35c9f7faf7111ecd211bd1dab92237e92909f406c40ae39e2960d61f25b9a35373e1815865ccb4a0ad8fc547027a4bdb6fd64c12cecb67546fd442d1aa819f29170725581f6f1034a9e940363f6619344a6242cdf07ac34a5fde68ac8f01daf61d6ddc88eaefef025bf16f1695ec41d3570eb3384fa5f5b8d6676f2fb569cb6a034056442e6347978d5557b4799d8fd31fac8db40e3cc0dbfb173e75d7d0e095a2d366f0f9745a8512717de3e27bc25f33b4559381316e1145993cefbd59b66062c9d4dbc8ed606a5851f3074b864bf4a47c2a8d98c202945f7d3c1c449d6c6c9253b3777d91472c2deafd2ee34ea637f03e798c95f4ceffc68647856f5d73d1651cde2c1312252c913e5635d936cf232c5430d1b0493f812ec77925ea80b03017b0a792628674c7771f24596366b878f236c9c0671a23344e26676a51cfd92c93457db4e16d53911abc56e9c5f0f35aad746f7dd903cb89d8ad83998cc2ed3e510100040f46bee31edf3b196490a5ffa72c21f14b1d3161319373cb40c0c11ea571f4159186cae676b6c10fdd4bde9c7ad33ecf896a38a925417b4428736a3a904417664c63b7e6c112ff6002d9aa6b0de4538a982c0ce6d89a3d228718ebcf5fdc30f51d0bf66dafc6e88bb79ee1c11207d5bffade3d4e8e9cd86be90fa9ac2ba9183e800334a32c4462;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hde9890d71098385dfd69925018eae14c999bac452ed3441254b3fe330febd09af49decf861f2a689cb0a1175ba6920811bdff579082ae681420c8070e10e729b9a1e9fee71dfa7df6c4900704f006d98f8af182b6ce78ff2d5df93aaaec0851dd8f9f8956cd5d0afea7e699725afbf90537f5a6e5381ff787393fa63b2b9f7981f385e4c998a707cb43266780f26d491aa2c1eeb96b2ef252b6fcf4e5759e70d05f4307422f49fca98e8aa8652f27b6648d59afd1b1990fb5daf2023d1738653d08c0f149752256e769b9e8fe3b747f462cc324dd85c4a7832652f2ba948fbc0ac2b9babaf07257bc2f561f7179c137f7882b8c948ca1d02630ba6591612ec37d2e7b2900b58ece1fb449c8c9c8d9f5f12f728634cc2953123f17554e2a60e0f83f00dd4341d99f975d19a622bf748d6a386b595eb86d51a2becdabea6e97507e857304d36854aac9ccd095597e0acee772688f93e711cae276291e84e2bd1108235b0080502bf996a8d90a56f40d6e756377a15c3bfef9190d91183fa33952cd63e902fb51710165e6414bff0dcbb465b3262e91373732c8ec63aa42557d022af9f1fa604180faa175f80c7812edd36df6cb91b2e83601fb03d93dc36f481c1855a667be4b73815229ef743ece46f93ff47431c25c8c6b92d9f78ddc2c2070c4b8f7de4f5a71f579b38c05cf4e185a5397045ed73b0ed9563b8298c7af11d74886065b0f749c5528059e6647dc5d99ab5e5f1be504eb39fcaafdca1ead3cb502cfee686578ac53dfd33db1f46378dd33c4b4e4c0060a9a0136994dfa6d0f16fe9ec5ae90ae55491f955e3afb87a26bf54a9b786429458c64f368125b27b555015cacf62aa19199d5346dd933270d27c2a1c1c17e17f47488f8c3ed4991380b8f4ebc6e924633609542813fc25923054f0d7157ee2ee52c0091e81dd069ee2ff160e408d75bb3731a21ccf550196b291f8d73187660ad2e4a48217ac5d5c11ac0d7fe4785ae41f9595ef1cce02444d39fc6f5647a9c5ee554;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h9c8b9a1972a19bf94d3d22bddb16652c4812cba2cf1265da7fdfdd37c87c8fb9f0f7442029f8b31b8bf4ef9cab1eccb729fe662ca8fef2db248df80503c8ecf1861d9cc340f69ba8c71ae28d5b76254cae4f60ec5b40d398fbd9e3c4a49e6871a5b4ebba16a6366745dda5b0db159df6ce64a71cd7f5fba65e141718098b4667ff88d07a26df0c43859b57a0eb29bbffcce564013813d88160ec1b533400e6c7fedf0718a87ecd6475b345895748f07d6b2e0836b6f2112c0505fd66acd2a8a0a58b2371e127803d89cc9068e5893ce3f55fcf38a1dc7f371af7911fbddf55c00b0912b3278440280fb28c847c357d8c4a241fa88f5d136437dd7567ae6fe7a71df83d859be1268bf267258d09b5b8dbdbd84498ffa44eb08a9088e122eae985904e6ca5a5e8b24cc0e67caa81e4f504524d520835b40883739b17022826315d95d7b29c9ef2112fd3f2c191c975dab10d5a93a141d38232ed8cf85b485ccb30606ad0557057cefc7f00304cfbb422253ef2438cda42b053ada7e432fb5d5fc0c70a9fbacf3f2a2e35672902b54435dc585e2975df941f8ae6844bedc1e47fd490930443530e4453972542836af886c7f98ff19c8365b1712b61977143afab9bf3575e1f90c9d72a4b0e0282dff7bf940c58c8d2cca230dc04749f07b8e56ae250c510bb8fc0903270d1ecdf4c3c0f40ce69548b80444817091a391c5fce71dd7f11c2c2f1f12a1d2e0621be6c713522c5383e7c3411c430622a75b02408c4c4dea09082aede18f2e6d803ae5c09770ed5c6c1c9cb96516a8ef664f7d0b8b8039fb03c4dd08ff8f040e9f494919ce9c4ba813b1c78e399009b0fe177c15635d0a599830ecbdcd718d137e4ed3a74f1e017f33cb0da0100d479c45406f34fffbce2e588cb7496e215d28fef4b1e40ec8c64984aa2c705ff74698e3a78cb6c483e5a3371f217de64f4c0448b7484e07f803d8d454585e2a7b7efe436daade46fb86c8d58a31eb9f33eba8cc1823986a2c8c4f3eae620e6e20275;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h57aaf521e8f76a1a71edb5efb1b7e406e4c77329d60d137eead77f4a8472164850d5e77a4b0f8057fd867b23c0c3e1fee8c09cb52a55a52224d6ee6da158271d098fc3bac8ac7a4d79acf8f695680b1055eebb440db977ebe45e1983f15eef5052c405e339723bba8d0b4236b83afeb8fe374d12a6145f09cc721c3a4c2b0267bdc12245fd87a88e2ec85f10103ac18507b2d4216799fddfdef27c55fa9c13c6c44e68332170854c2d6c7ec37d0dcf6d49a7fdca3554af5b5ea88b1044c2e288ecfd2ca2dadf8fe765a1ebf74c5c22b98ab5d4c7e52dcc3de8d7fab4972580574213d56188ec28566d650b4920b4e3e832e05eccf4a9bd06590c376f3c8158c8fbd95b4a32b07095b3f82c64c4da197f749be895d714d07b6fa8b9c38c9892b5e32e7185d595fe2304f8994c93cde24fac0ab1c4989cf0e9632a358b666b22e54b83b423f8079f2d3a319f3a903198f4a63ef86e732c6bf116d2a545d51ad904782556765fa2b95307c9ddd2de0e61ab1a548fa7ea4b50d021381468ebca375926c89cdab87b9bfbba27b87cd123c6134af235ea314d6b482353b78b2f71372f4314da24e7425843842d8934742449dfc848beb80f80df6dcf1a7726cecc46c36f8445d6585b55e8d7f03f4b956d721b01bd5f47b9f7979b7d6d172045bab3b1f394ec17a3bec70ee8b8f379f6259f80f3429d47e5041510498422961e733ec2aad175d1c7816b47346381eb299fc54a8e845728a757e176b113dde671ed885b37284980940d5a37d9baecbfc96b353d2a038d31fb6f45981f5359003f7b4f2603e8f4cb128b95e19efa193d10074c2406d214bf70dbba3bb7680c2de4bc77fd466a7dbcd8c817d3fba04c2e8700d20b5a3b7bb7063da68176d0d8dc4f8f27d44b1f8a26696d21272251de3db14b39b1f54fcbf9ee074193212c99701636bd2b036070563fccd5dcf6766fe0b240e5e47d25fb886a019f329601c9d96ef08b7727b372ce20aba7a9667fee6c3039e159dde8cf2cc56a9dd6a0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hd18313c80ad19570dc92fa8941bd0d5d8e60e2f242304834255431716f3e8bb5a061d94a2ff48b6fdca323157f74f94fed4fe71f9481e6d0053dfc73e9a18230353a60ef808fcf2dbd86947c7ae9757817ce32e5ded5b0d3100564ba776691957c42b725808e5ef882d3fb3ce5c88de1c718a60821812b77864e0e98d77069ddf88fead964535d7fe6525ef948cb9594e33332783a5612c803a7cd9c246bc68f06c9b9acdd9e1950ca18406e2fa56b356b2690e5674f64b914d807325a02494a12c8174fb4073f1061f24a9c47d4f5335a4398df04bf91813c556f2237bd24cfd443e6141aac3ce8d69fb4528e48134e7ceeec376a6fcd553619352b7337de0b5968783e63f49312745e6249ea1303b3f8cca545602b8717d485c00a25fcb13f03421ded9c3eb07a25ada6b64cf600df9981882c2e7e5b234d0472a0753d8a6d976a0ff026c9049747d8bcb3e5a0d5bf39626a26025b40984cb38bd8c3be3b67b171ba146d277f9726de27b9dfa3d749896d7f3d132e9afd8f5064396aa2b188173b623efc190673b46d683369c685ca08ff81e48c6574f955d0a91b9554c8965e944016094cfd095b5a8962969a584943b4d199bf3ffbff97c5bd95d34f536c748f2994dfafa113c68615659d389767132e6ab5cbe2f0c1735a6e7f064f56cc32db84b375cddeb6435351542df442e8810f62d1f2cb9bd72ef10970eb84b37e8dd45fdeb389f4bf6328193160b2459bb1d9b1a79b4afe2e9d3f7255cd50bf62af861090c919fba3e3aadb81e84bb76ecfbdb2f0adc5ef79ad27772cfb2e205b19b2ba9f190be15306d23b788d565a13361333164bd4e5764fe2c51e3981bce324f700bb649c03c93cb2bf9f80324689de446d3a22a04706980d191847f90218d4354c9193af083f34dfac09fcac3d9343bca3057ee59e1527f7793a9452c30726ca526f7c50e0340876f9fd170d44ef5eb851a2818f33f30552e5c31434c0245d41e9b9ae0c6df79327bf60c3738090980d8d6b283fdfd73;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hc53012d843a326dca78f7e1b51b23d645ab85d58639c439c188b369c291c18d4c6147b7bc30c6674a46c2871224d7104cecfc14faf8dd00832359685df9467e96504bc4e7f38d2c12ea307d91c5de78af3abcb331ad71bc55014ddcddd7d9011f80b7df3713d9762c667301c83e8a35eaaae705b46b22ed70990fb45ae2dc5b582c6311cb6a16b4ddca6f41f8b9a1d24bc248f38859907e2db0ee14b1fa35ba7e0cc39d9c1fb6dd3578dcc30506b40b653c13e8c62c7ed2e07b2dff06a338d6de5a802e406a6171c8559f42e783aa3763d2757b5583f1be8cc148f49ca843a5142c555003641d5fea5fb81ea4f532c214f0be1183a0f016005754b7750d4333fed4d000486ed5114766b8e013d608a2f29d518f8468b07e998b6f487857a138ecfad2b32ed8fa718d9a42289a1bcc35c787924befe6b2cc3336c807c308da9e6f21fa49a4cd06ee10609bec0562b8c94622f80f84c736d1c5ef01261bc96e18349ee4bb5ed7feb3fe6302f943c93decef18853e6c3a95526101e649078e6491e33776c6c5f23ada001b2e3e33d00927e7a1163755777f52cc0fe5e56a04d76c4fc3f70856ddf2bb51c059e79011de72dd56f8329e134d9d63f6fdbcf53da3579f8dc7509d8b0a69d32c22845c1faf25add073db08f8391fb36dde6cfe6969cc8cf39f1400c89cf31df0fcaddd15a267151b312aea31a27c305580813df23a8b2818ce359b8bea0749138c735917582c89c42dd6eb361738de9c149a1f80e174db9b71370433d83c5a0d3e5607482e7c6a62a190c35df3eeb7c9324e9dbf706480620092ca09f55ddbc3139d8d545150f6b051a6fced28c3fb6d60556087eb161ce996756767dda45a4a6425ee1e336ca837d4d9541daaf43f24e5855a4915ce9573198628f51b515b3b1efc7d48f906393efb8a068bc5043cebfaff3cd204e407f0c497db0e29094c21c0e2e8046ea638661b461db8b06e926e241d801e83e11b6b4d0c773f6171fa94bf17e8695593bb99a05d4ffb93474a5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h6abef856cf57a4ad080f68e2b707d708c6090ba6cd4a2c05997f31114bc6fa00ba739bf27464b938978d5507b8337a762b0b2723a736da78fa5f335e7dafcf193248b2095a8fec0cf88330e8cac8fb2895de7db0b54a2422c5777060b7f0af81bf7b39a12f630ffff6bebb1fd6ace913c97557902a19c2389ef260d5c5eaec2fc33dcc9552e9effc54901e8c2add6324dd2c1c857c2b60c522295e2cea72b3ede674ff37165a3e6718c67d0f1cc0f9ea7b788b7dedb1f7a78e7ed46bff9b0ad64a09bb72ec67f336939f68727f3747ad35bda32bbcf2206fda65b08d099b142f94ac3dd46742e772f8a383857649f11856204d5c908bd3dfc0660d066d584d2be2a4cc6574c9dc85335c8087761ddf836835864b3227d519491d93c2f4e230035c1e94bfe36ea7bcc38056a9b891f002081fa33bccf9aa72284122f2d589893a9ea93129ab68e6de19df724635f068af6a69bf46da246cbc4e6666f0660847a9c2f6ba6d76bee1ce4302a89c365ff16d68385ab63bdaa07d61a8a29b240bb894d29461b904e0965ff4b9c8705f39aa278b299c491072c6be2c9f722d131f0c6440f9e3a01f3041ff91c4ff003309c73cc9f10c71aeebf9dc6a648ce0b726f9f616af0b540ffe4948585507833b5dab9f8028744f240f15748004af129ad16d21019733d6d54dce6c4a27638bbd8fa60768f76c00fb8bd5a7dbcf795b2f637c520490fb3fd3c5e61b6c023542efa2649f30ba5282bc68decd32f39dea05e5db2ed0f8a93002865b7d0eca2678086a9da1ce92e5089a3f254749c5265046b27d4d68a7ed801fd7ceb1e18035686b2ce660af9688269361f15dcae3d30c6c19c0c947bfec932046f135c8ce48ac8bdee45fef0953e2277709872503b16761e57728db34b07b2cc24f4c577a0abf218d9af8200f2ea5322d698511a3b4002c0ee0d8b6de77f029a845b6b5602ee5cf0eeea3f8d5a86558e5b15a8d41d1cb5e328ed1348738b3ab882721a9fe8c71ff446c1ac5827d0dd90d002cde;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'he34cecec995a01643c4a53f0af31f3b1df915d9ae658ec8e7ec28494f1463dd558217298c68309cb8eee13faaa51988680c3db992371d2d6a50498fb06d95779d99f72c0184799c5da9cf3ffb25d56ece3f9f964818c45fa99b1717a28dea12f57c8f6644c68beda704f81d3c8243c46799d3c7430bdcc156034f8b568601b1a955f6beffe046c3f388114cb1524ae901bae69e5a03554b93012a2bf9842abc9e9233fcece1a1f81eb33faf23a5428f0130b316003040eb750d926197c61a77048e44a06d0bb28f9cd8961c710ab5a0d37fd3865583cbd8cc498c5d562697c413119184136c1b47bb6ba6ff6c8486e0ad98d06169094a2244722c8e02cb79b03079aa8622a74b332f12cfb2d0d09e11074c856b095ad2264985ca1578b12a8d240d2187c7bcbf7e216b5c69aa4e5b6dce3e80b0012a0e9b283b045eaef1d0c729e75b19409329fdc999fb7b643ecda510b9efc10aa5be9f33017e9c69d031897d83970097da568fa5899405f71cb589ab3870f97eeb9156192d4bad8fbbecd54bfcbc875b581198b9a2e401c202e616612a350ebe29f5e7dcf1c65322a6cd9ad7731ac2358150645956f1618e18929228dfd1fce6e5d98e9ad7af5ba817c9c826b582ad6998263ae2eb7f3031338d06e28ad684e078886951be93656dd465001d4b8f247165a9f86bce48a08435c6b86ef6c903eff4368e77b8b50d57bed9e53e50474be1d5ee677d3a937ffe60abe8ed46ecbd6010b0c6e70c78380d03f67c2f012de92e3768c0e5b1522ccd8024fd469b4c9b1638c46566f264c7907166ae604137e9e2a942ddd75d2801a0ac182cf73e5c473b6b26547d0ed074017cc60061628db1829f31fbe6e044af29b4b73b6ed7393ef39a4f09946473b15dfa535ffbe9785d49135c51f4e441323a2de9fd1d6393ce8081840a56b5a5d4fbe886c8d96de0775a2ad70a3770c2e5a26acd1591591df32bafaf51617a1dce0c45536bf6f662f3764a5d0a711cdcc22f1c3e7fe99715a8a6ebacb5e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h532b1db588243818e09bbf77b26f7e4cb2b4c875c7219e4d4bc3daf4a88d5fcc15fae4e50ab95ad97783cd224e4ef531280f446fec74fca3bee90bbdf5fa1e883fdd40214c24f17af09acb233f092142fd73801f1e8c4429cfa02d74249e6db0f445b612d799837dd694931afe9525d7dea066c82b891cb7976fa1868c6ff0cf9513690187aa76c9f18370212c5bdd586520b864f1c9e98ea7b2c9409d48c92c761b3479d892ecc90d5cfd4d082b043b01de9152c8cf1bc0d702d379cff92af85ae693b13a051a015832cc5791e9e966ee5684a0faefadd9b16dcbc3885e93ebccd4de58ae7033c3c71ecf13a7211c0371c16deb624b48e7b92f284b0dae91e9a2a2006f8d1f87d86934c79d5229eeb04f2faaf89534856569ad1ce646bf129f6714baa0d042d63659b5438255087cd6d6026325000d3d90507eef9ef68192c72e8e16b760866348378d3b109b1ec914161a3cc8e8bbaed677bcf95864fdcecba4a96a1396ebc332c1d5684294147f31e82f2027f0779231f1ae4bab526ecbd15874ea44d2c98fe98d05b83b9d229a0772a233fc092277fc906b961b3130ca29817d2ef64a12c886f3f35982a28d7269c96de9200b863e7aca48c3c2557bdeca50df801014f6ea76f04b162ae69af6b378c478e4067740a134501bc656b2034aafeea6d87b31a5306aeec1a5feeecaba42e99aa7dcdc86b01b0342357609fb0ef838ba634f7da9996f3a9ec52035359ae9b0d86d7271673639dff92bd26af7b7934b8827c4dc985bdf76ddbb2442cc102b6ab7be6aca09de791b2f1461de2d20a310d7cce6e3b2d8352627c6393cb4a0eac82aa24493947cb968bbd537ef9f5fcf34b9de0fbeb07e31f6ecf24d5e32acc7a2dd3a6ea83ea2df49e8533fa0e35f7919be8a84a74a1ce7a99afc5797b66040affcf6d72ffce4c2e8dfb518538385b802074d2e1ff5988d4236a215192abe8532049d87de33efcdba7c5aadb9831cc53a2795f28f824ffb8d9d0be07ff149fb0a34476258854ef5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h7e5a312af2f56258fb92533892709b3d721f12fc598fb9f56a6bceaa95dce64165a1cf0180a58e53a5d6445a99a3174c5fad0de4fb71cadcdbda0d751df2bac8918ababba22a05659ed326b835f139ada6ccc6d7030e84e934eb64cdf0e24e00122b40cf24111921f8801aa2afb026ce0ebe01bc44c80ae5bcbb9200d62f764734b90ce2ba15f94ec1f43f2e5a764eb3afb9bf39b1c5d213f5da00c81c017695d780ac3b9b0aa56d2cc3311aadeee8245fefafb371186bbccabc83965348fc6fc0886630f90aa5b21dbdf6a30f73a710581ae0d58b74612ea2e0d2acb13b12ecc9116de15d32d3fa3fd03a5bfc4e536c7863cb726b566e6f7c7b022136c79ae093b0e47845cb90204b6a8b036070b83fdaf120892d8bab34f161f1fb12ebb0e095467ad3b12f554ace443cdad31d37889eb6842b0e37e18b08a693fc2394cb5ea3db432a5a452db08af835d33293276b3769bd1605153607c325632ba74adb213b128e693eed7ec64527311d9a2a8b8e1d71069ba2480ae3e57a4299e27c1f66d2eb1dc38c5519a944720f23cb0f4dc46653aaa5f467e812761165e81eefa51169767d88f02721089a8ff3b2476ad1ffade3dc4076431e901d0eead1b08b6deae777e84dfb5bc44bf694ac47011070e87ff68ceabc75bbe17d691b6c587f52163bc25f9592a40211bf50696c5d3535fd0dbd858c12eb62de1e44a8dac837079404fda2c572254ec71013790e24afc6e98189b162fa113da882114e6833caf14a10376cf374a08467e75cc8d9ce9dc01234c3004a0a8d4f068152749e1b53bcaaee9e52bdac9d3b8e634d092db4faee2f74006bbc81a01c4669c5f1cfdd7a092fb0c8d78a60a65b99771211ac8ef6834f2e5889ec69a42d760e7c44e9dc964439e5ee25d39da942d93a80ed2919ce327137d24d6d0968dae0f70a5d80720c8fd1cad805501d27adb391289fac29863e81e71ad915916e64af111ceed62d131cb96e89d052861b3ecb7ba4565d0007978b2c8723a7d0ce713a8a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hecec0bdac630ef9767de658e71f41af7b11fd0d2934232f829ab0d814824311bf3cdd290a06ddbbce5cb85d0d17742c32cdd15be4057346415a3f9542bbefb737119abd0bc04dd3b20a4420790762ce0ddbd6867c6632aab0bdcfb982ab425519edbec07033f07891a7b7dc47f5418ba2bec8e052f76676e389b95fec6ed9a9313907c4c9c0b1bb6223749b56a6fb8a0826f4d2f3b22b78f193fc6e5ef57fa8948d368f679857d88e3a8dadaec8d043d3b8399e589af0cc0cd652ed7ca6500b2bd780e74bd64be01b1f0fb7ffbdfb0290d41f291342b55d97907fcba9aef73a423c159890da5d02073bc06b55f9cb2358052641032a3c1ff7211935df043966bfb0ad2fa3c7dd8948fbca2cd4219d96f975a9b1d1ea5bd619f17b608aba03fc9c3a7efcdd20a1270f130d66e80ffa71b339414d8aa5a3c6813188977449140db234d5ad5ab30f6a75ab00ad392e2cc291989cb7e34ed7162911691223e5877dff2b72c0e726d27eae57483bdfd34ac17545c91f19bca98de79182a29966387bc81e065e08443b42f505b6d5527e93d096bb7805ec8302b836b1a4664a021e321bb1f2b0807e85ad1387075fdb3bbde5a2badfed0fc1790f2da9aef04e10ddbb240553e3e7a612d3ab8d2cb39ba188e1ec5b33fa519f1e98c11e37e95089cd54deee596683fd0297b5fdd9f58079ace154ebc8f26d1ca9b234f76b4d400d344a215782e5998aad41a70f01c9b9d6b994944601979780c9fdad8dfefb047edbdda0fea628a67057468cb63d157a4e99c0c3d9ad7a213782111408c86e55a0a7d1a96e695a86c4f4974c2d76249c000b4554adbf5d370f93a0af922231ddeeb20bb6abac7ba42a0e18897c94c4b196a75bc560eebb442c361e1c340041e56977d863353d298f995a7870b36ae5a8ca3a64dea475c398572d95de62c0f75b1e2afedb52b26b51578edf36c181d6467bed5db35b8cc0cc87b262afb67a4426c61574eb9df116eb00558fd71dad13ffe16a5bc55aa1552f1a4166716;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h91cefe970ca70fb5396c73eba8bbbbde813c947d5d19e2cd523d38a9076d2f0470615a324c1269bb82236bd4c5549fae40fb96024cbc01cd443817ce7ed83c2755dc3679545446db852eb0edc52ce0f37565c0f2d23bb1becb5c998145e857d85a15cfc776e96fab8333712c970e8417e9f613765cbafd3d612fe0b9cd42155b3f8061fa9cac2b63b1320957e3c6ea2a75f09ccc2c4c7767824823e0561d6c61fb065d876fe4f9a60df29994da069d08bf1ff2afcf5a65fac905ff4eae7daf02e43c5b644178a8f204465d36e0a57aa0660411ab20f98ce2e969904d6448aca16c8bd516410929a781d86ef20e84bfeaa688ffb84a94ce26c317ca9813175b3f280fd1e824b0cd1f21f06da4723b502fec97a39b822da9b66a22ab65d7facd23985bb7bbae321bb69311494fa67024e661120860e3e2d2d622889538583991561c26a801ded6332d37ee3510fec714c3f824484b3e2ec21610fdb2a075b909250dc2dd2e5509931863d82fe5e4b32b18bca545523685158d745726a2502ae1ffa5132164d06eae8fed5d92f8d80003bf062e5b0c78a9b3e577a8cad710553a7e9e8d9edef3425d099387664544c976ed03d089bdbe6a60db0de79382f29e796bff743485b81c5d259f4c2ef4d95ec5aec6aa173c209b53badd01a395b1c96871921f93f1c6dd2414b9eba642f5f9074b08a01644607ff34b85011b7809fd951d3bb5391c94b8dfaad0343b9ce5b54cfa9e1362cf76cacc16612f5bcc1ba249a5e57d5963f134436a57d189d378f084541545bc6b38e2a4af9183f71a1956dde74c31076de4f6c4066032a42b16d0cd239f64630023e6e9bdf42ad5efcf646c37546a22ffdf5496d719736e4f47b40ec3b68385c6ae3911a9f5d3105c83557a470ffb0ae2d66df67df34399182dbfc16ef3b7f092e9dd6eb755c78b25a49cfd28cc6b11f05eddb0f0159537544432e951546ecd8596490cb5e35e7db499292de1a5d4a991243356be4dcbfd2cf4898c378a9ee2e1e2cfd2a77c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h6d24d3e7883701154d2de443ecf98e765d8d28801365cfadc5e961b0320c9a22a5c780aa7438c757f0fffebf0010f8890e4840432a766f914fe87d9be3923f13a3b745057911458b52de9a3d63c4fd10892f3a99cc7c12aa026e0c1d606d3af966ba89a445db88d865b37ce0e67fc55957371f4bd5d37e1376a18cf4f3fb482fb6bed3c426a70608e0565be3c32abfb88de05a6e870b84c93b2cbd1df144eddcb6ebd3e0bf34835d332aa8f13673d9adce97bc24dba93673a2ec63b27c5e7022823f0c09e87ea9dc2731f0a6be02c3f7b951835daf762ae617ab7fb8bcf6b5aa4b22c3d281f08041ba84bc2a28d3f4879ef0980d777688d34981621f2b80471c3480f66abef6b740e6f76d053861a717aa9efc9021ba209683b4c753a2b8c831b0de4f481fe890fbbbd0f540ca149ef534aae5b65e227f4ae4c774cb4b0d827f04dd7c2251bef48e5383b1f02eb0e8a28a6d85e1635d7bedff096d6a91779fadfbd4a003e432384676f13aae9e2a3151eeca4120c462913925ac66c0845d69ff26c816652f2b88f7abe207f13e88891ca1d1d37ad50bc162c99b9e29c5bc9972a1448db2795aa47cc033621748f08b31200c57b237d87592d88b52ddf757d70e6e588efb0b3d06dc695618a4462c966908587d1b217bc7e5b4ef955c1cb8ed34c0c35c3a48e4e01d413f4eccbc40764c2fb0d156e5454c24731f95bb190ac5eca45611216660123a5dd98c7e54764647a1b46e79297b1e2de6609bc2e6c31ad979668f4adeeb42b379ffd6e90448a81e62a6a787ad94331777d89851cff6b348fb3657d869ecc7732020d6e54bc5e58f7db86a6a5c62a7c36a89cbe5a058e3dbc62db586cb458d8bf1d74e68480cf7656035b3d97770c3504d16af960caac4a43040928f4e1d7cedcec5fe79bbc8e0eb307950ca00deb914c06304b8db59d166bfd7d06a5f43c21555558beac595942ac698198e28850bc42db36423141afa5178643ecac0e91a297055f888e3781ab9a42f0a3d09191881ab;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h6d8d4c79bed0108d004f3b189daa29baf8908fca43363e79b44e150c791676b6d07bc1c252b7ffeda067de014a731b2399d6b2bd1e95e228a43922082fcf8c04edb069d04fe29cf6dc6319da418b8aa92bce60302ad3870859a24e070c796a95ee0d94ab735d3158ab5aa3e1858294a6e597fa0403be085c49eded6836ec97eb82e35ed869d5a775e331d434d9e1818a8fd94adf0ca611d2a755eaad36576324c03e321080606d9bbd65a4dd3619c38e5e185240149a5996a39e5821d76367a05dd44dec3f9d0240ed9437dc07bebbe0361d2b0bacc0394b7424c894275a74580d2ba7edd2f225b90245af1f663aee210e821f8e8e97d0642c1e9c143884270761f132c587e098b034d7851f1fae5b0fb8a61c2f11a7702073d547ecb97507b93039446f816b2b11496e971831af36442251e6c8b413a8976fbaf12473c2cb0618b114500509a65cdc153cbedb399c4c1be883ba2898833b1501f226bf76cc7ab2ee351851c71c45599f4d799604c946c8dd13ab5eb2fcee7e45f456ea2771887037c2ef57f7ea7fcc0d814665c7ddeb93e76af29a802a2d872a90e682c5547f325c3141ec2c4a32df99e0a27abd563931f08f46c413a915a85d17b8232443ba174110d0e138956764b8a4909bc9f70ad157db69c1b117d759b6e4fef16525dec771ec6c5c8447c122ad3d6b7723a17197918a27e4365f1b5e53b87c4a2b739b42f6dd0db6323e21f8185a2d414059616850fc0717a454fa618bdb0387b0fa2b792248247d48b7442c8b72df025efa9100bc4a297ef85d1e3276db1a58052bcc456e114827de5cfc644e484b0e0ade64fbc07068ebde8501167144105ada39dabf68a17281886a30e0826b7aec1337c5736b93e73e53191f04e28b2df15310a9a4bd42846a7cadc5e52a22747fe08ddab6d2741254e39a5186a681a65c36ef42684dfb8ed7fb76045b424117d68fd761e10036d60e224e025096286339d50af2cca549796dcb5299d51a026e4346b06e8a6c71915d3004805b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h88a97c374bf403d5b005bb0129e4864c142c24fe249bd13ed451d545524e17e73d4df0b6af0b0045a3194644cba199d8fbf4a3302d1c1b05f261ed2bdbdb083357c7d22c202028b838e70530f64d21b3c4953626a9ec998e0acf4e5a04ab8bdeae8d23e1638d4c71bccec42911f814e463a3031da72f3ccbff8d43b53877ba73e80c21753880b1016e0f94048326568e079b3bbe2d13ae3442baf14777739fa6297b4a71ddb28568cdc3f98f52d9fbbe6c6578a26dfe0dd0ccaeedb738aef0262c8f391554a8500bdada457c0dfb7afcd5abca3abf3548da2e17fda5a23d303f254f239a3221177fd7d3939226dccd3c13d65385f71d9a357f5c31fc7e061e2480a5e8a80d589a6d4a506b7ca719c7ee80da121f428995aaeeb74a6f89c83770bf00ef1333bd6bee5c0dee48710daf30caa811465bd7079bc39179b0f24a5395498956e476d4a37ccb0432b645f34614ca7f0a4516d25d736a4829a6485d05aa8d944e18223758f43f9a1391fff42c4ef8b1c28c43cf8dbf1b60fe96c085248b7340e21ceea8d9e686b7770c36acccc155d2326b6dc8cfa40ca47be9ddb3fd3b22a21f03ed1733f9ab92419d81c2b98a83bb3f4d9a7b1417e19b22450d69dcf89f9fa1b7d82cef307748956406999ea322c79a9265a35c0e82b1cb1624e760ebc2b5c8754f481b466d9d0adeeab01a0b63c3016a70c3bfc76f212a07c1858f576d636c124282cfa8aa42a603ff31656bea8115e5ad5429fe01ab9033d156bfca71d6fae236926d10603c56c5da0f6c72223ea1751bfe6309f1c0593237d2837c7d45d9208f44c4606e3ceeb8af36ec1524ba144eba229ad91452376547df6a91dd13c8dc4ba9903cb48d261d5d9e7f751ea3c0c2d14ba2e3247844733fe41cc643cd5449c1c28fb2f927178229a8ed6950181f9f0269a749a37ca78b32075073a6c75caabeb5ef95313b3399f43dc88e6111ffcb5a7df5100bd4e0bc713f7f82569c306f2cf92d7c316eacba20930b51987b00d435e83b13cb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h119923a01398738054f253c744f18cc50882c969f72d782ba73d813ddeb9b395705d2f1d44206dec195e98c487fce4029ee1158e2a5899da762075f3b7c37271ccb6f1e8e8851decfbca6a38ed0c6ca813e9d8ab838a24600888acf9bd4e01fb1d29a1e9bbaba023b800705ae3b1df4ccbdb0ce897a0248d17ef1251eb546fa664f8926c2b47fc3869cde7d1f45e6011ec7d476a2030af20eab22eea8e285bfbdff2d1a7fa035838ef1677206876337c755e8d38b29a018980e14eeb58670a6a14526a859efa3a46c14c7567c83e480cec989249c1233aa90b636a5c12b0ba69fa268a16b57512513ebf8a1a9d5d255961bdf92e4f4224670432765e3ab50ca1e4e904c7a4cee30cfee7f5b36e373485d41133da03f8354d05083d5865ebda58b6c9cc50cf3b6e2e402f039137d147178a5bcfcaa04663a7d40a2a4d0db4053a6c8d1b1abc2fcaaac56a5d6328dfcad6bb288124448ec3850320cec61066005a6937a1e94130d3748acbaf5b8333f57dd4a94c436f5e24315cb127ea3d71be8828256fcf0c768519457b2a1e5b2176c69ad47de99f314c59cf20386cc0ed4f2b0d53a2d14419c794bf17e5b865dcebab2b40e0b59a8253c6dee8b2d549532f52431f10f237f2fcc7da630b54916577ac4a5a77f9660fccd26d7e1562c850aa2fd5165c2b6efdb724f68f6dff2a90f9fd977e9eb1bb28f38b96e7fbcc44124bcda1c60c9d2654a6cb2fbfbc36b00a0f0023fd92c1f13033b9773326503aba197511d977975875b9b9f57002911b40256134c716f46a77d8a162d347830ddc03dd0b355baf13f62c48df3cf76b40c04022ec7af708ff77dfcf6625334a22876d8ce6819daf4bbeb94b18611cfaa91dc4e36c15c5fa28a42ed4b8d0a7639d422d755bf55cd6574d98f7596bd05c041edfbe246cb94faa511bf170a344168cfafd4bca01aed27bd6fb39e75d6b1bd6c6b7b5e1fa5790a6c9cad5221af451971fbea56324812b1be945f8fa5e368dc35656d71e28ae10de485286b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h8bf4c59ec594d7e65508536ccb9f86a2140a8b58e45f98cb8553840c7dbcd8a67952b7fcfecad1792c021490a3468f9609061442d50ec09c9167de25317c6c5b4d0fbde5c8af403591873a283d93803e56b128292bb98d8143bb6ea8d0de8e583386df112fed9e0ce46abf79f0ee2f6f701ae6fd7afaf2eb5288a203fb2366a117ab3592896b01d5f25227b1d27a56e33861f1fb41a612fae39b592155ea007832b51d55391105c8812b09fb2186d303e09c5895f71f5e8c98c8c638b0f26d2035ee93f9e3b7e1ec2e69bcd750a1dbbbbb5abe58861d76dd94a32a9dcf5c5162fd65d1b097a84df91ae616cc741aa262e8e3ed417b450ce2006f8b77ffaa0bd4b7f3f66e00e1309fddc032422a3b937df841c5ba7e624eaf425b6f9bebd4780720504d7c267ce5c3af6c39b04c4a1c4028a009e3c19a971ddfb50488929b647962036a3978569f7df44e223cca79eb6e464f19a21b9de0a973bbe91e6c2d0b2ec593c1bbef2b35ecef1b86d2ec8b0593549da762fdb83064b53103d02c7f1fa871f244c757c9edb5fb3bf7261bdb75e6461f807069835f6d06105ab7086ec6a7234ab143cd492c3d4fa85bab53d55ff76fa5fce6e60a223c602f948e4f53397f098223e1321b49cc764d6a3f7c1a9f80b796001fc5a574ec6fd62952598971d43cee676c1ba798b57b0d8f80e5e2b65cd98a52732e2314d3f83315703d93f9f9650bf1c9cabc782159a9510cad3736374332bbb46e66a5aeae769e84b9906a6c8c2fd4973eaaf1f4fd79954a63c734d0eb85a18174fbedccd5f0dd7b93905b03b8e8b45fb3aae4911820fb739d9f4b12df9d6caa57d0cbf9c3bc128aa23e8ad4d8f1aa79926362512c1221b0e6966c49d1c1ebf84f2a4c67a651ab795b8c5138665619709c3ad6bc21ee1d2158f9835b86a8a03e9755031043dc9aa566e509202d3effe2809ecf738c5522f2512059ae52ec304f0355f66742e4e349036f244795fa452a123b13f976728c06dbfe9a71ba7c64fd719f80dc61;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hde4d12e434dd9518dd08f4c7f1f928139e0b6907f6113b5939684a4b1560983d863ecf138abf7a364ef6a1212864f52d27d0dc25e21b117d9dd98ddbc8383e506b997ca604e98e640fc8e6dd09a8c686fd371cdf41c90ae18b5ac70f10e67e2544baba6fd4a098747b804b4c82f042e4311b1ad5385113c31f394b64666f7b517308b513a90b0ce82f5497b6dac0ac7c732551616ecf0c6dfb3b3ea203130c4f13ebdca0cf2f032004954d52925f423e02cc163ed486ea155a04eb3b270eeb76f648403e82d4c77bf9da04f0cda01965b310d4e57c416ce016d20b390eb1a447cd5bcfb592bc05fc3ea87797d302db2e71804cb46bc271842710b876f0db3e6e9ea5f0bb60b1a3a78d005ede879ae1044c35ade55bbb0cb1a1cb5690a8c7e724c76751ad28ef01573bc59a7b25cced27fa57887486fec026527628953be12b15b8d89d0d5b3dd94f372536e877e83272aee31b344efbefafae2375b86b729fc8b07894131898f4cc9344931bf47b51189157b85a966960c63242feef8c34094eb9331a8dd35435057785418225c172e0e64a081e251e398d000e02b35eeab8fd84191e4c00786d3872bdeefdff3e1ec6caa94bfa18784776b4087e3a561f6de8ac53634f0d7596c2f9ecabaab16e18377e608cde468093d91afe9fb4a639d6226785829a491044f67a654f79db0bf1238dbdd48594ac6ba31a3639689a9221458d2b22fce3814da225544d9a88fa53787712f55c952dde68d6699af490f8080ed76ae6ae64befec85ff07d2af16d3fb5c680640d6d980e151b1f60a66a157754a8524d60a9156dc52c1f1857380170f21def1544462880b281b71341a3c97ba8824fa7e48f9064f3b1ff128258493a4b02b3d5bb11645bb9b6a1df8e00e815381dd0c6ca8f5c90728279b92986b8cbed9c6e95d2ec641c8521343f3c6cef78c4707f3220d90343e35aaf7f0ec31fb3098f25853827da9871966c7fff784c341d22ed658d559c9ace7defa99a63b6e00560ecc5f0535e0158c4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h8e00bce2f9d446c865d1215297bd75ad56ff3aa9d84491e63ab682a24de80dcecadcfb5c70bf82cb4e154484603d4b43c006aa5717e488a326b671017d2ed0675b01caace9b8543308fa8c44223180fbbd5dc215929639940f3d6611104b978a13a206690303210caa55918baa7cd0aa9591af9693a221014f4e8ddd731659a25bd728142a55054d04439e0d9af3217d12eaa2b041557b58a9481466e278f6471b459b3b7084241358817c13e3ee99b89ca213e69f5a328c17b494a312a0804d15a331e416cea7aa1fbf109fb44fac83a4c19832bf14d94355a71dceff5659debd0afcf2e590b2856aadbd9332cb938d444f20f90427197075b6476a7982081f7fcd6001a0cb58f0b84f9e867967b952ff0d20151cf9eea7833859bc913c670ae2f395ba4433a7288b497ccef6cb2fb3b0fe24d4ef4756d1b7c3d0e353cfd948fc2aed66e89d7c158bfe29947be3f6d053068b8c6c6043cbe7f43e034ae27d487f0a9d5682a019d9fb5db6bb45d6c45b12947437cc7e86472aca44e9420285cd21e6780a7dde13c698d4dcef62b1766e4400a37a3d021f54ad5e2ea6b264183fa8c1327b6d2c73e42c00955ac03d13eb00c6cacdef22c93e7a12b6986c33d6885e389493a534b8414aa16e7fa25b410bb2e3234329a1bd4666d56b25c8a70456e87dcc0d5b1d96136d17fa5565f3e62eda35c790b79afffcf054a026cd7dbec8ba24d31a7aa20adfb4de6e54db9893a7a9ade1000578976bdd1dd5930568ce0633857af894f8086baa3873e289c84615351d29f92f4a7756f103a1228f3833f6fce80b386b77125f3fd89f054672be21564e4a5903eb903a96cc8da70cfbd3d04a316aecde4c6fe95b0d0ee2c4d4b2696731668263dc73ac1c4b1136a3b5e6cc8a80c4652492f62497a418b1451906df5decd56c3cdcb4be161945fe4e7e1e04168dbb51866cf189fb4e83539fd869df7f342764dbf238265c7cf0381ff211cc14159d29fc52f01d0a69e79fbe2e481dd05224f9ab90136191;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hcf1b1cdd3d4bf3c70eef41dc55c80df60ef1b46de689cc51bc88c687b61b4006ff6fff253ba722637a002a4176d01b42c7141b0087448faae7f4e0eebbe6350fb3b2d77711c2a0fb791912ef593ec246f8be66db71f22013fb4831771143e7cf55bbbd94410e93de8136a965f76520f8749bde18f0338b03955f30df86670933cdf55a9e72e3faed7aa41ad74ded41fd4845d7840bce3a5e682a2759d23cb2ed4cc71230074171e9d727ceb88d625c0c215760e43da63ccafbb7c5b40d9a8e09f578739c89cb6a86a992a4b24ac31a39464171d435119df1f0e2326445942a6ee1cbc3cbe85b592c04d24621bc35d0870372301d56825ac28c8ff4e37f93eccb4fb085628bb14b18d76283cfdbd55dec709f708605fb29525d7a832a8d9a9ae63f1f5dbc80a32d0fa2760c275914d1fb44358690bac9230b6741d8e2de4fd4020276d9bbbe38667cb9a453a803830b0f47a7c9d447d00c4639d35dd0012625061ed8922be45133e9e393bd247ba63ca755862acd788f68b56c2e759dc2f4278b688884de83ce74c800f622d6cc67638eb01fd5ce6f125368b84e9b2f8888151f91c296eab0cc49c645d49d1c399357e980070b0ce1ee3cda1890be0354497a0f8f11c948b63f5c53da04ff5bd7caa10ef9f677f3907b66277fa09a3cb84594a97f62db17636ca2b5881d13f909689070d816f61107f328f9c401a82fce01ec509af5e033125a819551471ab299158f7b74184ff7515f3ba17116391496b97b93eb6459365cb8f1ad3f9c1d1f3589df58f6f81f54b241e062e43a6ad4051e7df270282571f95ad15ac28210c8e98697760b2d5dfe1543dc3b14fa28d07017cec0d24bbb8d0e8214cce1c568a5e562e1c254480044466ea6676efeee3339581b21796520cc2383600fd11b423567b4b0931536d6aa8cd2156884fe5a93c7aa32732fd2f34aa482206f222d41f826c57fdcb806e28c114cba6eaf2591e091440f988b066ae79781d1b91786f472840fc3c5bb842cb6592652e65c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h492fab61d11543fcab8716e531fd81ee2b3eb73da51153b2d3038cd547e8ba6d68033f89073e92263caecc8f74e0a7601ab7e49ec405b9dc842f0315724d62ad993bfe1a306385c7badee39b73428b02439c1efb3222269c6625e5badeeb56479ff33801001e3dc6ea3a4a454314f7f4f0eed4f2a2c736f7a63addeb8534474d89d00de67983ea8228e8a617197236c05a7b8f1f7c8faabb26bc367a919616f68ed5066658fdf953efedb242021fbed3340a92439bee4708c27ed9fe5a3a2f6bee4dd8133a7e69e67b894d62df2803702e3d85a10f4688d522ce289713b6d2c6c3bd5e45767b2b283915ae583dd4877524bf012682919ea919676d9da6da5beb7c88e95dbe7ef89bbcf0670650dc59d7e176681bb1d88b50531c4484909fb8491649bc9aad56e62aafaa62dc402e183a47c56de9e5146d33ac2b974b50670de449f32aa0a5085ada2f7477773963a067c3393d1c6460fac577bee36f39f15a13ce15fccee8188d0ee2ce0ce2761b162247564b67155415f157edd178472c0c489f144158fe933c09e92892863e568cd430ffa12a32ea76cf7c1b713b31bf4e895c9378f5e8e1d061374599cc8a97d635dc41bca2196c3bce92720792ab0a2879591e90c71351531702bb8dc64b0fbec920ecb012ee6ec88303ca0a4cb6eb21740f89efff96eb1206fc039fa04800be037700135e31707a1ecd7a2a13e0c2a332fd6b778aec0e8c7890d543ace4477004fd196f4616f981dcc7578d47b5e2846505a1e59a29986b9704ef94cc3d1acdae9cd19519f43fa012ac7754f2832306fff0c3dd86042b6bf5e8940c6bcc8c31a6038a1559a7d9f86be5984bdf323ef7918d17b36ebd8e5bdd8215cde875738afc2ce4e32065252480a665a2f35f9ab8218a0739435436b6aa176ddd08c468477975ef9f18d1319bd4f3e0f41b5af37b7d404b53eb8b5ce2e4101cd8a90377184d1ec11af8d07d743b756188e59b30258b6a6e72c9d8cc95374932657f8b6a7d6fccf6b8dd0731737fdc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h18264a0a94b56149d1af07e1c3b19f3588e792127370d2bc656d971b19bb27ca09c29e794d1272a0337ea2ab60322c76c7b516e2233c3780bd3ca27ee5eff7b8eae83d02b150da1652e87756954a76336d306afd480cf33608b512157ddc2f399346ce8cafe2233e8b08696591aef4ea6f11c846ede5357673f5d0e45ef6484deeef756f5c7661387b2de28529144bc6e9c32d8c162240330cdf97a80667feb975aad4ae75aeec468e769b206942e0c6352633458bfb1361db96a55b85532489e7156e2d662193d0e1bff78e766f85cfb86329cd424c530a1e474a6f5ee49e0797e2d5071cf6d08f5e0003cb5f0e0051e9460d02da5917bf528f2cd52d2b1bdaec64a710492ea88b88344c782454d877f80a3313b6f18096cba30a8af4c1e9c50a91236a9b96d8a9b549a927a245da2dfa82b5a0301b2e5bddeefe4ff934d0cbdee1bbfd04dbb8a9cc14472702ed0cb618ccb8467dbe1759fc558676e00062b931655d246cf4d7b5cdff9c59cade3dc8d8670226d9cbba282defd02dba0aa463c322587dfde0c046b674f3103a4b81d1fbd61fbb8255898a6b9f4da884c7d44fda30f7a2664059f1b26b3d1a26d5af3b166d5dd65fddce2cf9857f8f581ea93df04d6f99e841ef7c872033b511950cf1fe2696cdf9179ad34edf044375cc5e6c6c22e25799c68280b2cbe7cce121b50cb88f5e902efcdae53198520da2e43615d6eafff3881cf7a8b9ee315330579255ae385437b608410f675f259899a8fcf572682959c1aeb519282d43d91d7cbb5a13a24423cf425851ee4c24708ca6b90a3c607012ab0265862878a1151c2c46c647375871dff540e1eb053df1a8f8bfc6601693328ac775241afa747f72164a634aa4e7e77791fceece1d586bf18353c314c68a0358325a2335afc368f39b78e6a30e4ded4ecf49e7bf15041d8ff31e8254233bdf2e986804d178a9052664668455b0700366f844c01a550820b953acab8a3fb55a53957b53b2654406bc74324101c6711cb4f613acc3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h22a6862aca5c3700b2dbcb5c48eee0e544e510fce37b5f5817cc99e55a1591442817896c7805c14f2fa31322d442d6e5a8578b5f025c5c0378faaad5fea2fb3bbe4c1e35e433f34263c66faab7d665031a360bc9bb661c0822f890492d4f9afb72e603bf7e3f9a81441f318edefbd53c7c38b087493d2104859effe225e4ef8c9f8e7a34f544556c570b4d322e5fdf8b9aa1cdf7c5c34513935f5a585e01f78c44187caf188884f5b656ac124bb200d5b1e758e3beb6a3c6ba44f8c0a59fa51febba04c80f636157b7385e9a0300e2a1b20d18fd51b59332c156fcfce1b089be6025bef3f94629ec539d73396d31458aed406402e9d5389338d4742d9518e84001800437ac374c3ec7ad04828710e5b48894ba8db6155fab3aba06816c294f6df7997401efce64933fdccb63de16dc30c1817dcbee0b5770dff7b8021e2d27f596afc32f0abc4961bb2c230c19b770c97981c9b19ef5aad87cd6560dad4a8ab8fc91410da3a56c19d7872772824939f140af0a007a62e5ef7316928bcf01e5a1990988a62f086f8a4629662817b89cc2e80e35fecf4f98fb6f7bbeb8b0400546617da94b23e3322a1eb771a52f5ea6362684578e2562893b96ed18491a41dafdac1e63b95770303175deeade21e5c001f0873329022f68767cccf4d405c36484bc00f10b8a7617bf3f1edf924ba114542b9647f3f51b175bd7f359cecf8a8ff34a6cdf99e7c0f909bef214759b2c3645429df03186d266ef2d709307dfb3a67173698661a8e7e3c7898ba383d9b17610a94c6b63d8ed08de2dbafc2b2d14f2dbb31d57fb27e3e324551b7fdd6d728f6a6c8c5e685f4914f66315e556000fb0b3bc125d202dad9f33bb9f0ebec7c621e20fdf20e884b9484c154bc29a2a1fb8c3e9e889e7ec38b36d41ac741936b2a08dc273a62ff19cc4ed232509202331ac9ac862b580649f5c38fca468faf90363fd0bf2f3fcb803cfd7f1e418cc798dc0456b5ad5bfa013b66d68615de3636be79ad543a566de82f5831f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hee664b67f40bc9e5abf21f2fa19031363e26595b118250bbac4959c04eb96629562cb2f87ac0c10898db3c4a5611b5f6e5f2f6f969ea70fd0de5733d3457a9675f9afe5f96f3360be0f1bffddc5fb4654dd38121304ef33ac5032af04fd6c02e36c3b74c10d2faa91a9fbe8dc304f7eeb85f1c450bc11e7e0579c3b7dac90f1580293330e31410332620bf1b68c4291fbd8b9a4c114e87ea7c497b1f405069c08e00d0e81c70c51f7b60f67ae35bdffcc00e9fbb704347edb02c3d3243623f5ec3eb1107ef2d6b5673710831e31160969e290f5b94dbebaab523facd459c68719df6a87ddb8bf41bbc81dc55797ce2709cc1d72332ff3c40201f5a4599ae2d08257973b1134b0e2990b27d19f3610bc69eae8ac0b947abacf0f1f7b28b07b9e5bb9bab1f9bb8069e0933efe229f5e2f2c87ec9056f877fc3de6448c146afa25ea312863576cf455c90531df5d7079de30ccbfa3c9900587573914899c8affcdc1e4e36b27b034eb27733c965658546d572e0ec2a744fa9cea174394f34855e6e043b272fc0a26c5119ae90abc8119869312109401a053e276ed12c01be0d0b4a7a712cfd544a90bd771630856eb0fb1e7304204f65a08ca922677920e772b0451824179b65ac9bd065733d9bdf47e80366200dafee02bed7268d8b61859c101084913b978fb90bd08ec9978d71b5d3180e078ed60a34d5dcf0accc63bdacd81040cd1662719d6fb303e9ca9cbac8e411788ca4e4199e592174edf58cf20b7cf35bc1d83aae696f6dfb0be096eaaec743e739eeeebedf7d0860b0b6502b01d8a430bf892151a0b5ed5e606981bcc2b7e3c0d1064ce25e3a3bc3d1e6fc3d49836d78b93cdf5272b9f575a908443ce65088dcc2db2c69ef0593268650a4d4e6ed49afbabe7a45122c274c47f4886c7cded427a232f3bd64dbb6a40385468a5b57fa282468122ff98de621ebff84f542f6bb425f11711bae2aae50c7c065c3921be07664a61a47f5fb8948a7a8d3513b615ed1e71e5f8e08174b2b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hb59b487a006e32d971a885f7d82c53d1a7dfefdeb9cda61ff0cf2ccf3961b74a7ecb24031cd0371da5375548abbf0186ce6a6e597dd50531101d7b6d0265a883ccdf64c1ef33ccfacab48acd6c8afba0d2bb8fcc0822a62e79b04f698320aa76d541cfd8d2ad14d79ff5e355211faffbefbad91a84db2b5c633d98b6c703948df04f3632fff332f4ecdffed89a59416e7c4c7a9207c7e29322a76d8063f0d787976541fe52380f0cb7defba6979b7f028470b793fb17ea04d0abc11c1ea350601a8993a77e776dac0d1b1ee93bd53d6c1e9b2ccd43a41233bc427d8ccc3ca1b82ef5c25973ac91668c91c5f021cdecf4e636ca87c14c58fae80877cf9993ff679d80a0a207f06af9374491a7472b34e035912b4bbaa849ef4f8cc9ea70d68cf9b217b1a48555ad0585de4c983c5d0fee0db8815916ec1b4a873dc9c028406bfe30235c14b1dd599e376e6baaa52ddca35850243a07b93461ad01207d575da11b99126024679104f8c357328acafd6a5fc698e88329bcfeeb25ed3039745ab4ae6563ce967439716b97fdb79bc83acedcb478b29eeac7e5d2a60db2e312bb335718d321c59b15a0426d39cb0754c64bfbf858d5f9dad7b04aa72cf854fcd802eb9c40b60bf7a435e6e3aa8aae7b123e1d2bf501f30a42929070dbedc2ebfaab597fcfb88b5010882801a71fb5c9bddd252c02c9f9b38ba13329494587502a2a4ca7ae5315cc954ecdbf5ed4e9652df840bd29640e917714bb4348be83bf0ac43fbab07423076f66561afa2e11c7f7f736427e0f9f04aab3d64c9e766d44f89b19ec03028311c8fe36aacf2b2742af88af286781dedfc8bbdc1ac74ec09fa41672936e5181bec7221d056d090499ed1e89636a55dd975a27043245a04237044d3f58290d003a03514a46ba7c4d6f4509c99ad1be5e335812ac1e1c45b8f2adb92a8571489a2f1eaa03545db05aae75c8bba32ed7d40c85e8632aa69eb733f8b71e03a22764ecb160c350969b5c5c3881b799d27f64bbfbb5e0b7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h13a08dc86de63f889d205cb2adf32881a4cdfeb3ea2cefc404054e5c11269a01fd70743899ad0a624e805c127142a0630325d40d554d32134cc6d1f880abc30d97cd8ba89b82d43ad869a58a12ccad58575809bb22227065f541feca892ef7c76dd1ba0265ab5604c9521de24f5946bd2e804920adb2764dc4a8a77f9a6fea79e3a38b874f97c98bc85880a950f0cdd55b1bf869e357787a07152e94565242e76dedc5397a40ce2402eec5d3d3096bc049d44721f5c983d3fb8e2ffddd7631683dda6c59c254b11a96b690c947d43f65183ea53aed5268a5505790c0be18dac96db301079552511152547cbd59454f41d4272bf05cbd8b1117d8d190e90addf072e7f2ee3b2d4a994286d50129d93a418948bcfe6bc5e50f858da6ad015b691bf4e16d34a38fc149e49a7c77d47e61760c8725006b8e24c5473443f41cb10efc0f2131f6657f3c5980974bfff5d1d58c1e77001aedb3bf54bb95ddd7bf9e6cdb7806e3d23fa1d365a9eb09bccd5f308f386107c528618ed101dbffa7570df9bfc63ba1430aa77344875386482048abba439eba727449fd40f5c51554fe6d77f7fcc4b6b86afcc973ad07b21cb443309da5193becfa9780a0ed9f848682516af7fc929ccd1f5fc0ccd67a1fb6dbae5cd20c3c1ee8d8a3a2ccfe00e69bdef701669510bea7583eab11bde2a09e7a43f8c5f2726da4c00702711e54985b502eb6d8f83aca891eed6af0751ccb59955bbde054a8de15e13c12efc349e0c35dbf1b74ce1e61637c03246b16a89e6b8b664cc5603125f254c9452a772fde80451269212ba6364ed7e0d745929deed36eb877a4cf84cab8af93392c1b788cdf1f6cc2340709f90789a17870e033462980c5b77caaf71f236b0b7c83f3186c29a16560eda1df2fe8629ff16bb255075cc51c48c3fd701ddc128e8313268e90dfdf627e5ef467c8a432d2ba0f36fd7190d8675314cba9b14674d44345071f61f208f4af3e676f12d1ce2bb34a581bbe915e4d56d6ebed4c48ca3572955b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h7f8e6aec8b6a4b4298fb052b457ff2a902baa37bbf35f9e5d6e3cc0bc881d182b57b44bd067c82b91289a26d337634b8272646829527d4eb59375608e78ffc6f0f6c9b2f9715b69a31246ab5de58f9f13b8e2cfdc90cb4e7437432cd84ff5e6ff0d298b07713f855da7cb46ef8bdce162eb5fbed0bb6bbae9166ea4106cff947a74dcf2f0a186f5a031b49f54f5d52ef2b19be6fa67499d2e85e3773b1c0dd46fbf463f80325416a376ef50374f03c7f1e61cdc3802cfbff7f3524df400e41d969d3b9ea90337e25cf1777c3bc3ffd68b7ece27844e7dabad9c555dad25d6ff0060c5bf095d8261ae567c7eab1cdc5fe08fd21c47661fd9263301388b555b1b50b3c600eee2eaee708ba2bd1ee737e6a66f6a9e3700f6c90eecf81ef2b990bc045bb1d320a53b653a155eaaa2d67cd6bb2ab4e6d78d6b13587ab18c26f8e477d23f1bd146fa767a22f5dbc96a87ae5bc9fa2060cc552d98532da6eef39b19f15e93f2aa1f4f38e07e5789253c662627c2ea95486899d57672ba00b902f31b5a0a4470c13c52d41901ca2bb59ae9258e6db923b235f51727f4632b93869718f1aa3a1caa2634639b63271a13675077dafb63fcbb28bdea5fe8f4ba90b620b27edcea1c1c947ad06106f8cbeb76388b1094b71da01819e6c430c11723a71cd99f5076d6bb4a720b06c0ef12b87befe6447baa8004faa0d2de00f96c177507583bd10b365d50c4c56931ef889bf69eeb29f13316930ef536926c505bbe5372940e495910084909c40d9787320a058eda82850ef04e9ed7fe86ea0e32cac2d4d8c0b886df27f897e60fd9ed8e4080a76d38448a970600560894160d9ff71c49b0fd60c26bddcbe7d7c77382b570bd9014184f5d2dd5dc486f1f6a83ca470fe94f57b5e5934e581c5dbd46e27e34f2f7c45cf21bc8260c5a3982acc47c81ea4f5884124e39a4a2f30fbca94f1cda6a58c3cdeeaf4dbca342a344912d14dc0814a1f2da532cfe3ea6eba295e44091daeb0435339a1484691441211d8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h1a5af09c362f81b82c223cc9231831d1e7780e9363a29e5c52575739ec66fd8fd044db862a942bda313a74a4594e5553957ffe8aef1924f29e96ad2fdeaa36dc5b6f0ee122c43d81230399efd1f59b38faa8ff342d22c514daf530321d3238c402ca71c267eebd6c61e6c394800c5d778c708422476137248a43587ea377071e0298222ab5480f76d99cac7be1bb576877cb2ab73b9c442e1b6bace4263d144526ca9a7916db54dbc00efbe481c05c3e36af8990f502122325cfc74b09305b32695880af9368c9ac81b433b54e76f336f11c4ad9fb9d643f18680632daf4d850cb6654f667c98a77c5174a5e0780c2c8ea408e80e08587ca8ce1d44ef4d1c25599e23992fa7db6731c96da9e3e318282e68284e405706ef7384c41598f475ba0031dbce1f072ef7dabfb6538ec9f7194eea2f6ccfcfff7f1eb515dd945a61a3fff9d4112bc87e7b5f0265c40e67a4d9600e74e9c4be641f4f1c14be44892e162aa6e161f292193a0a235dbe3d6a7c4e9ab7c159907bcb4d69d6bac093069051202be062ba03218e2a9316839ebbc3a3d1c4ed0805207caade705dc166362fe2e95bc7480916bf4691249f32e1c4ed41dd627dfa27754bab4750aaec6a9bcf226b819a5a66ae44f71267c91ddd319e42910c29903a8c7f0b98ba9656318cc4c95643418fc64d64854795ef8046c88aa9c75939cf456497c637f4dd8ff54952253876c96f2b835ae66bd06c41151e7b4491062d403e060517ba48d9b7b8721752c8e61f1e28c038ddbbb40734558bdcd067b503a594868dc446c6e7076ffcb52b1322cad4f37bca09b94de5bf6fbedf1602c18a151edab18c4584fc78003d75e5262e3851f84d0c4827104e9f9c78fec38a8449a78e2d6c51fd0c2df3cef9734913e8bf99e1288693930333a748cc42c8bf78decb47b022391b7389fc41909a687bf3b7af12b9eb0e65b14a3d30b98350913f28f5dd0acf637ca67c479cf10e9d8bdb8fd8bd2d6c5e3e65f8f1618478d5e85bcb6835d2fe27c04;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h8400ac7e4ebced0460493cec204c4b10fac63665edef735b263ed91fade7f6dfd8286e610b1813e1c5462e6412914c80dfe17b16d6eac5fae00bba6eae5ce35b83f1885d88296c06f38c1503da09ee75b713e47fdf823343c8916bc2db10b51eac25f5cb84a62baf7f775ebef7159761ba50aed8b24a72e9a9d5079a8095145caafa4ff7ea2cfb95d3ecda8efe2131c802bfb07c7fc1ec8dbc847d9b63793e5a4da286ce55c0faae8b6d87f72ce419e7987c007eea575c87e26c9dd72ca67642a7069f579dff611a720de5691034925133e8e0d7f0dfde4bc4410b66a73c1f17db4dab0347025a5688fc999e94af243d0bae779f496bbaba0f9bea4d984052b588e39796c524e62c351cec3e31010d08d37ac7a2afbe2de022adac7ff070dc0d527e766808016af7887ea9f55a87a656f2d7c2ac30b411d816f4f463f52e0ff388b1ae43298e71b8add2f1fbb7d8e678633e765ec5f286dc2c3f6abaea8d0410ede272452efdaaef06051db853d7065a687d27a5a85f57a42c2348781820b86b88af5f00ef7610ac5ba78c4d3428bcfd33b16f24ce5f8265b7f41a63f1955ad3bff54f943346ab16591ad611b7a7f266363924f752300ac64cc516c512773e35a2fa82acdb820bf0f617c8a034521b343efa2428b56d28f8565391fcff5c2a28b74a0716f7450781c3254c97995e5e129d8ed90f26e89c2e15bb98c9185a3c3901bf7fb6f03c8eb683de7887f629dddcfe9122ba99186a206a8fd482ac99b5b406050f2cbdfeb85796f3e51c99521218ab88de9191ec2c5d4102311c89fb602a8f66b000d11884f9b6b808e8efd9ca04bcc86e49dafe5371f5a66cac6966e0cc9dc4600fba59d1be31884b1e3decf1ceaf81935b65af16795d9e3028c2987aaef1aa9b564df5568da448ec30ac861e1081a2756ab15b420bc69a0ba9d9afca8f353d68c312f575cf01fd05541c7b87b6d0f9b42601b02a2a97d009c22e9a7b3a9cc748f69b05a2e75854b3995e1920790686f226ddaf3c80f0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h6244856f790152e5674e3f22d6f8c1d56538dfc8e473abc63b708c89f5d46af739c3bcb467ada910df3b6c4e81424310322433db0f867ce754e8c52a18be6fdd207f6f434b66057e4380850bee2cf787b1519d493e1154903e4d50f6652c2fa8822c2ede40402774142e80870190bc573816f71c85bf9375c6ffab78da2b522b0ecd2191281b7754868fb46fc7b0054bfe8a764f56f18573c2f9879e634bbae0d006144e7bb7919de57086fde9c8dc26fc70614b4f825079bdebc88893058cdefa4d1f5cdfe2bc97f1af4a9f9e335d9e3ed932f0317d993d417afa2e7b278cece0a0c73f90285eeb16c22f8b1ac89143a0ed75c5301363016df3e1cc67ff0d2c97d882efba0a995f93bfeb736f2ba020d57be7b6a41db9300ffcd0448f5cf760825417abc16db4f933677b9b2cd4e85155ed44ba1233326551de96fca0c6d69232f2ca87d9219bb882272b9a984002e82bbb3eeaa4572233f6d8d7ae913595f060fd6656adeb78fefb5fdd9e3cfd7db0d5a8a6274ce44cb67b12baa061d7ea5c58b76a28324185f54632b955f0c20a97bb61a6db4804027304f6f12c9cb158344cb5087e8034488a7079beb71c0db64d11728dee320e641b50560d5403237121d024d3c10001249928cac21ac4d0d8d3cc439c9efbda09ddb43e17be4f21a08845bed018d1298eccb497c4c501ea8b261f932173227aff5c9a153abf05c12c0221c85318ffb29ba1b222ae9d3b4bf57d17d85fb4180951d59031138f1897efc02da03f44aa6da263adf6871b09b833459df7358b92a2ab3e5b34ddd889a1777c4a9c901a8efb916dbaccfef6cc832fd92e45984c5ee5c3971396978087b8b80fb95475d102eaa452de51e2c47406b7069ca7e0bb64a048ed1c1a37da84609d0fdb000a885966ffdb8c4be3bd9f38fab93bb42010a683a2435bc07235b59e60055a616858094973e470b9f456d3d4c73a71bba1db72fcc3cb7afe44d12f7076c2f7eca9173a13fc1703ca45a35f93917f147a56c5d5aea54186;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h83f8fd0b862ed9e5deb554c8d0f12fecb89a38a6bf487f7d74760575c4e19da861d712140aa307a2ae5e689bb8e94e4d54d5c22874874770c63263e2a1f85d807427730d2c8d44dc47d0f025ca96fc3540f68f5f412883da72c6e450c0fbc5cfcf463c2d0a22c24b03e83de4daf835b8223cafc6ee50c5022bcd25122dff39c2617fcf55d94806e3604e028820f540535a38a1f5ba917bfaa0e7fff0beaee85cfc8bc38f5833452fd67dd71d69cd0a00b315d5a561417f33907d0d0c94469274470e2597dcade25ae8dc7b49ef8cd9355c1bf80b6bb0c6bfaeae47ce75d798198c99c1125f1ebcd7fed348735ffce5fbaa3984ee44b4916859e55c6b3684b2c634813332ac101a6388c018521f4387b3a854f76f731769e7283309e4574f914ff493fa7faf1be9794d0e28fdaef2c1ffd009f44de13641579454c1526b583d535d9c381676095c1f4d8b2f7c0833ff1ffc549b5047f50a5f2eaa0b8bd1e901af79e419dfa452a20859f4f01ef03d83560a86f2b9afcf64bed221769e85a1f52ebdfc546ca5ad69d5b95844a2d682b07d6af4c8aaa52fe0a32357e6052c07f0a289517a273399952d28dc00b7e455feb64008922cf10538b32a2f9a9eca77a205c2b765133d5c6eb6abbf89fe73e45cf7e75c5054f901cc806c76e4299ac90919b20000273837c749b706bb60776f40269acee8a72120ab35dfbfb77591e77d7f4cede72fac2ccdcd21532700f9860e422ca62d848bdb57b23bba54c6f06281b542ea5760f0446955e269f1bf80a8dd8048f281f2e9aafa8a5f0bd153c9e3aa6d5073eb63d131ab6dac907d539f9ee57b7525e66e5778b5396bf7b218203d6f8a033c58fc662537da1493c1f3bd76b61e812ed46ab81cb55dc78bc1c1284b02b645c77fcbe2bc7cf776a9de843d4672ece14db5ec7af72b550fdbf04b6652f7ceeac269c2d45bdb3a6a30097b02ed1e1197f4c837fd707a31325059b7fbc61fb51e4d9a4ed1fa34dea4e78a694403870e1ec3b2368191c81239;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h53c54f2ee0d810cc83d1ef9ffed9142ecbe900b8289cdd357c6090628e15373aa5e5f676d8fedb518067b53c784653c625f0a1ee72f3543db4cc0e17a95d0db447bfab3f3ca277fc05c8b9f3821811483c1b2367f8a6b84a103dd590115889cee7ff95745dde446f9db921d75cb076ef765ba2c31a60b659410ebe6e9379dcb0249f856b988ef76a1115cb355ca69e9d9c1fdff7df29721e09eb55453259069ff9e138f8c718b5dea8385dd3410f27b125527ebf285be48cd4cf96cadec5f761c1c8aeab23cc50f8f2ea3716e217fd2cca6a553cc90ea16722291137bae4525644aa3d02dac2c60dd599ea6661e17b8136b9d18bfab72b80d28601839e17fa0806195c257f70e410f6c9e7b0d03da23b921763de476cca1b9af9adf714c4409c92de6433394f57d8bcdcfcc0adc0be09834c6e86a3d0bc19cd52ec47f80d640e47d42cc31260bd62e640ec8895b3032228527da947fbbe88297aafb556d925e7fb77b1716c239952399c27499b0d1cd178b05a0a8332a55825e3856d2f3633e975853bf79f1acbc8b60ca8c30522a54b3a37db9ac7db9e70b516487bd14c8b47151dee53df3eb33010398360bb162c6b0e212926979db83a4d956aee5655423e0d2033edd0c74c0916a6ce5304d26d35938e2604e3c77db543dbb009e7bb51e1cb36554ca27d272f8d17e35dc15099ea51dc7ec0e6d626ea5a9626190815f789148ec2e7c43d8204839caafce51af54a91039f6883567c1584271661157dae2717d7c1224163df3133c4beaef3ef4539f57ee2ed37a9d10bf714c210ac6eea08172edbe33e55a58dc586d9126266f94db8ce5d508c609338dc60c29ffab6dd4e01a349643e67b51ba9ee821c98a1eb77f5c1620794a700178a6f7a16c87de08c4ba1d97a215ef28bbdb0e980e98858142458b4b91fce93fc850ca393b958a88de731839fd553664d69063ca4899bed06b3b8a0b147838a3a92f96fa8105ba73560c24fc70d7a8adca3bb95497aeac980703f52e44db89d520d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h9b821821c34c2a9afe529a843ece43fa0231c5ef37d9d7af33eddc3f2f9fb083ab7cad31cffa9502faca5ab3a9a783b6456b2d87a1f15acc5a1945475bb491a8347ab3046abb4611079e4985eb2e9f5cd6b26f2dcef56a28f312a2033e811a030f7d2c03157fcccc06eb08cb3bceeeb489ae0fec3e9f2403a27f328b9ff8d79e7e71f1c69c2a6ba37bd87e4d81cb1995b5408f0ff5e85eed975e7e1bf05cd0b07eadf09befef52853d8c6d946d3957a3f9b124c5b6bf90bbf3f2f7ba4c100cd696fe686f2cca42c03efcae80a88bf0a12a06b15b5b0581e252f41410a8cab6b6aded3de843763303c54161a970fffb6c98c834ab3a98bf1a5053c8d1eec0f66f0e9e4761a07a998f3a8023d1a741ed7d3cedb4405e76ca48ce563352f9ab3c3e561497ec4124128afc9ed77d11e5426d9aaa4fcc1a971f2dd336e3a2e386413de5e01fc1147460aa68f01963454ff5b3f8508af5c098d314e326579698f5b58e47a442b706b98f66bd3b0e42fff6e78cfbd43cc7675f3c74af8ea7fb260af27b7babc52b8806481fedad2da755644fef529456a92fa98aca55f4a1aab4dfef51a3b1e16b31888daf583c3cf972b129031951b6d65b9e12a9ae93e03ca6ce0848406277c6fe33dc2c8b1c2d680d96b6afb2b58c84a8340f2e4332120b856ea55f049a8128f0692ae994655500a556650f010e9e7877367af27381babcf6d868e6295c05c3c194d7f5d84ffae4ad907ea34f28e1bf2f373bcbd34bc03d94d89ce33228f4271bf12c4966fbdc4f6dab4cbfe27764ed3ea2cadb82c020821abe3aa9fd42751fdebee17e913b8201f1a5b6c0ec1e47f6f38847b9cc78a30cf1708f023b9ce82cc07103908a35000ef3c5ef88672462e6466cddffeacfaf7a0580e0132c966d86e8d4deb09c71f9b81bcf22b6f8504b05345e7e6a3489f986c29aa5caa70c8ba0c4d48fa2ebaa4378316327c26724950faf97d06ecb1a79bc75b139a9cffaa29214154f268594177d010798a7d4f2487ca119f0074b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hc94fcbe6a34bff0b63caaa2a8d4a6621736c56a0191bd491ea71475546494884adf7bbdec26d16c60d1427fe4335e22bb2b53a1d7ce4ad960b247db61e7254b72473119677e7bfe14adf1e48ca3211ecd6853d1677c1b5e8e0009b89bcbacf5d6b5e0b94bb59628910148484dd8fe4c00e2df1e3253c346d89dac4c450c4582d313e351078561e9a21c585298fde893e543392f464fdc73abb066c925fb168905ccc32e18ccc7be5df11debce412bc736960f18960ae4aeb9d784a5c19171363b9c879d6913d951b2a6ce2d75859148a042ce146b9c2a72d916218ee468c0be4595efe6e2e268beda07e84bb925529869663b7d0dc953a33c926b4932d70bd2ea1751d33dd4826eb70b63fa09e4dcca99999ecbfc74c2ce1b82b0c57fc628aa46ffffd9c81c998641d775c4ad4325ab831227308cfd8d50ae9c57f3911a4f48c0b985c173968972b7c963389acf1e45424266018d8e3857b09ea7359ef9cd9e1a967b713d2f88221b56e75cfcbecfe06a245b0db41185b510320a9e3e6083951bdb5eea261a8c75b0d6800ef7bcb68dd84b405ef320133ad5254c4931bcc22ad09ee8a9cbc50217ee0abed42bf31ae4ec3337eba6f90c28ddddf56ed060004d681cfedc9380f638f197ecb05832ca50c225a668c05471c6c7d2efe990125b021d192a57a8e0df9213a45dc3b908bf2a0a366b79460dce8897428a5e414e66b6ddf675d61ab30047ff73f5dbb9f1877906fd6b4e078e8175022408b8c5825cfb2ac71250aeb85d6bddf32242f044fceb7dd9c0c7262ef6452935133185590ff57d423fe6b2fa8ddb77729710aa2d0080028de1185fbc685445909b8ca2253d94576ad3bb37f036750d38741fe74e9d2547a826e3a60e059b312728c5dcf5d19c9e2af5241f8cd72128e3fddec6adc90015e18e02b87b48686c9269b1d66a044c0850771361a9befbb89974f18c4f08d6fc18c30a4e8062b2b1658da8e77b779fc843f8392e4e6ef29ea6072402768f591d2539b7832dfc1b92c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h3db25a3ec633d76b4d7c4f1aa8151722624eaa90d7b4f2bc4317489f8956bf14f587db5ca1e310ae26e2d3332e260aac980b2478227c43564fba507f09499f7d295f0d8d14cf28ee54e52a99e37704af135b798e1b42eb67028250da241ff2191b7b555e95c335db40d2698ce58505de4dd20c520f0059915dfec06b4cf47db713782f6f3ac9ab258352b4552383973843cbda41d6f8e255641cba15fe99989e028cd8f8deb2953a0ea5bc1ea0d79733d88848cc46631948bf8587f3146b774c6c298e255d5e707e8931eb4a859e39154628b02b24a3de1dc37f1b6df057b961fd242f4d33ed6ad3d5143c5f7168ba08976748a353d0d18c5b7ea79259bb9fd470f20e605e9cd39704619755a7242804ce6f5d8d3566ccdb46b477ffc33f4e74643146f4385e7daa1ac9517758aea207980aa2c667b410e706d9e268d34abd26b7e5e501fa53e5fac0256195e5068a1be884122add1abf60bd3ec5bb83e46f2079453201c31178644343e32b2052912e2fdb9134b00a3e21e7c5e62e364dc1e8d61449f3e8b3ac79196038f10c3b0269021ad28f12c198000be014720b482a540686fe0c41f38d91f4ab21f6043fa4e651fe9f3c08c0a9634b7817cbd320346f1b0057ffbf8d31dcf005bb3ec35f35f6a332b844a8c67f7ba6c91f59780aac6877f270b74ed2bc48d8fcec15e62f42824c3cf5dc221eeb79c9c98f0e70ddcd74e7a6dd66ce824d8b9c739fcd221fe0ea8ec465e060414d12d857ee1e6b88bf86b795d9bf930fb029c320d34b47e1ac163b4dbd3fc7b23d5531a8b7cd3234bc7a9e5745195910cd395083b9042a4351f7e0d1e5fd556df75fe6afa12938f013e0b082aa428f1afe0441b236253fa5f54224bceaa8ea393d1bed62f65a0edcce5980d1fe80b6e2bbac43ef012eedfd96186bc36d0cdfdc3e543d190dbafa668b8f5304b16d524bd23b20584345167a76ce8512fb70d7f54ae7f68ebae091bbb2e6496885eed5ff907d35a20c90a950718c1065c0e0c7ca67a940;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hd00ff8d815315e2cd6c197cfb165ae87dc8b98ae8f26f3521c9df765b679f40e8a045142142e0b85642754c37b4c87ef24228e7480d92b9e885e5772255d29b0ed23efe8b96bd7a61051da4c3e38ad62a0b547e0733e98b3a573dcbe43b2a7ec3f8f232b39bc8d6fa0dc68b27b9f85b0e2fc84b5bb200ce24c6a9eebad5207a838892ef1d69d8e2a9b80390c870515a7a80fa616729d80faef9a23fa1c3da0e38395fd93eebec3ba7a6d3846a20871a14d549075420a1e8ee53e96804fdd8a6e2e8ec2c4926182887378cc94f3c11c4bb0d62c5c62cf9c925e854cd4e0d694acd7192309c9958c99edab183c1954265e9c81dbb3e7595162f8153bb11bfa73ad87d88cff5a2efe392210566c2a4a9e5953df4568472953cba90da8a43338a95c743b86cc248bdde3e8450ba8adc5473ef4aba02dc2da80f08bccb706e1b548456259d9ceebc3f7de74ecca9304c56750693a3bcc57e2e8e7ce37567d068b9a67ff17cd5b0cbfc7779e3307ed875d13095f2c18eececb103e4aeaa466d24330e6f1e65252134a26aad82faa63c53ac0cb28b06680e5ffdd98e7eb623a17010ef4b12c79840efb2f2901bdcf59261deddd2dc5cad47e6e33865cd410ce78da135b7c12b0969a10bf9694a08750633ea4be411332864c52c22cb9d8f455b26879ad8bf7da020ace0aa2b3f07e3b90e2197b8ff380bc9c746c830c2af2234d5ba11a43ac4e6422984cca7a07184731d235d19ab55d5850a7f401ce227ed80296015e66181cf065e4aa72e65c6c11540cb1fd8a14b6352ae23f1be8f23a63cba47ce1e5b446e923b2407a31ab1793b46fa717bd8b909362b325ca93959e70d3d41fc0898eb696bbab3b2bb44fe89148f5241cb8c2c52dcdd10e672b6e557e40404f4573c96a69f88a29cb6e31abe2cb4581685600ab6d203ce5221391d426f282367781ff64bf56ad5930caaa026b310af40d3b9d5dabdac0a071e5f3d7fac82983541e99457909e461cb218138961531fa4bfa1d863419354e7885;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hbbacf5c9943ac042839e1f77921e331be38918aba53fe3028e0ee7577d832ba56b62bbd2201a930b2ca73a873ed0727ea61c66dae378fc7e9880fecc514e4cecc9e27a7817ce185bb5ec99bae868ed922ffbaa51a41cb6c9eea152bb1f13c313b779c425649146e78a24a625c1f08df843f84d94456af56aa6bb08d3351ce83842acde7934d5db4d76ee7da274c1ae4abd18e5a389bc50f681288b4210b55b5dee1f00cbf8f637b19cf29094e72c52ae681ccc9964b630229481fdb6f1c328e12226605af3b422b4e43e093f13208e449c84bec2996652b1eab03bdeac906ea554e69600f0937359892243e7718fa34212e640bba20b367d9da18ff1979996beda127d0af8b676cb71822c378032843f044b2a800b13270c49d153f5e138d7c4c489259259610540dc7670fa7a0a7ab9e8e0de00ba7c5a19e35adeefc69fc52303914019d838f21ab2117063f2e19a089fd4382bd9fe7ecbd5eba8430b7813347b7edfffda6e1ad3351b5c35b44eb39074f4a3f5b62662f4df5d0cd30adcf297b37f01c621298a98e07833d3109e01f98898b40c4cc8ee18f6499215fbf0d459e843b163cf2ef4fd418152f3034af55d273a7ec21b1c257f88bd094596cac2b09f0b68816f4aa09fb1728878c0827bf4dab1c7af0705e38b79268308437659e75d6f59935c23e0fb626ccc16853bae67f3c4ada8269dd7ccfb77a3ed0abce2602f31574a7e5ec1ed74c70f1c5ceb92d3aad90c1710b73fd1d03432988fb2918ec0ba4d82e6102797d9972764021245136e333283136b026af05e841d8f123476d0a2a32ce4238f739d860a95646a74ea167eca8d24842d73758d0c8ef91ff881fe282a05a4dc73b040c767358dcd3b39f7f0360811c7b0a8256711804eb872fea3fdc1776f36690948624b75d46c604c7c1299ed4bbe72aacc4fdc0a824d00037a66fa814904d42f66467898c41a71832deef6dac1bfacf325121b60b89c799ff40e00229ff9bc54d7f55f726044c49aeb1d3295bef1ee8714;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hfb07af9c6efd67764f5861b3e4c7e90d61e32606c075d67ad43b0d0e05774fbcd4f1a519330ae9a21a0eb46097798e17feff93f05b63e37eba0d4ce878d0f7a311542219c972230aeb4fc18aa3c9e7eb5cbc2fecb8222b30a93d0b5c130c509a42fd163e88729f2a496c01e0bc1050ab750f1c9ffcca753d28e42e8ba57854c10e6cf3e24db70b347fffc76282c4225434ec9facf8d9b60c68e78d51074b5332845b129cfd6a16de21cab7b35cea66c32f480e641a581d43ddb9090865d92b8d8dbb74618c7cfbe595c9f4a103d683f96b4559989a6146104503abcb6b8652631412e2bd6b3e90f30c1b00168ed33dc6e86c0573669d1fc431f3bbdfc8f9ae68041c932994028dfbf92b381d8fff46070dad66a3519f53b5b34457995823ffd72168997f81e9c88f20406290820045e7f5e00e0bd5f8c2b28c13dd9fd8373924941de1417db116d9c6b686fb303b716a1580d640832a31579acba19c62c7f8238d278081ce4583eeea6c2145736a3ce469959242987be7a0245eae4d42502a5b5e2a97fabc3b87e2411b35ca29a380a3643631e9d5d813351f0a49d877a0628e91d3571733d2d389971da18cf91995c74a5701931cadf98d3bc1da0ed0f888a451ea078d1fbab3dae89f7d1fbad449ce926f6cf054c4561e1811ad4e81107b0611ae206be1c8dbba3a3e15b43415d818ea95c47769003f29a7b18b083ae235124d99190aced20ca2460b85b3467b7d5aeecd9ce4c72112711a1e4e0a34cdec07a2ea7a040bf16b3b1ccafb5c997a5e5e4d5ef3d92741158bbb06503522a5d1ea5699814a1ec852b9923bcde5c6839d5c9189cc28192676cc2af5dd312861f2cd12fa17b287f2af803da6d00d92942eea924c61a09966bce9078058765e74c965809376e75ee2a39e1dc442d63f9c5def3da0ab0255778ce4b9679422f6cab658a5b6dc76b018a7b1f3578f6cb1a8a2692246dc794b1584759343ccc7a601af3c399206a70362285c76678633b55f3f556252837351b974cae7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hdfe79516c3906c359e1240ab38eca907d02c10cc8e2bbfd0b92b247b81c38af60bd8ad4c5d0c2c526f24838d9179d6ddf9650d0924ccd8576a83862dd70b11d35fe070c2b400c05ec313f94df36a676850783c6251097b9c96b43060e06c99d5d1231bad0bef2abf2626d7a7c49e956c2e5e5d67db44d4fbf6b4beb557fc3296d8a0bd57878bcee12515559830c8df298f4a9a9d571aaedf4b2c3fd589f928fb13b10a90aa80ad1a8a88b813c4919135a5a0275e719023d4b11c3515ab7658f17a3ca9f9f72962f7642d9c67af3b2468e7d853f181219f08bd39589c4c81a22421c52379299964d03e6a7198ddc77ce676b9860e61b8c952046c9f426f0edeb401ccf746c22a0d3bb24929c1af9f8642ca09cd38ccfc90014cd3e6b0a04d10354e15473cba97e8986b305e2e86333a37963853d066b9e6f916658a371ee093602262f95e2717bd476c06c6397fe11e622c1681da66ef72ccd7367ec7cc92df29c0ee0cfddcb96d744b520287f156867bf02d10266c52b4698aa6a12dae6c594f622a6f858a545b16845699e3275ee52be4b3da71ca61b29092d0a1550040413bf41f1ff806a022c62b6d23f02c904687b34ad11cc8f00dd535987602b50774a1c7a8ca96f428d62ef58270ade737023c177cd82800c25da6d81ed00d02a1086e6206ca6cc0150c8bd6e5bdf9fbf4fb8674c3dd5bc7e263450d66e8eaf647daf27540c14ed819d4e2d5f3127d9ed8a1348109147fcea48816d56b47239dc33de164a17ddeb090734c0b2ce5876a2a634eb709f6d0bd408f9b867e755948fae0d6a9c24598af0cc824c6ef443f981ae7206481a66962c415c8f79f2fefcbc81b7bca4f142f24335ca5484bea26e7f88ad797cee0300b448248347dd4fc4cc981958b7cbd30147ce566cadbb604d793d1d0781762b5844a63954549d35bc156aec98c22709db7c8aafcd410cc439ad4364bb7cd1c9cc51fd8c9fd2b9a243f3d38e98823bcac8ed52e8154eadb90a5912fa71eedae572df207e36e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'ha941ce4bdec9f549877b8c1a19b202d8564400567a51c98829f0372f46481c4edfccfdf4e5c5488b57e79cf6b4a02d763e38cbba4009fa6ddd6dddef337db00a6ce5b7de04d75d44797af4b1695e79c03f0da4c310175ee25fea9934812d733b2dfe1a4e5c7058a4d62334ff30652612971a53e284fa6a1d60bd71a37f8218d7f1a01ad9524d3ae7256b541d79fbb939543738250d3b7b7f8cc1f83dee1ecb2624fd5e3c0dfda45287d8e37c00e06a50e65cf06a5075d9afefddc3177b9cbc0207960d91b689b992b766e7d3f0000a1233b198aa1a3607a01b3d0ba6e84ad94f1c6a4ddf3a9a50e557cdaeaccfd807562ec3fa6254f8857d6afb0df41fe3f1ebe7b96ca9cbd2c0b06a4bc3fd27d516767172a1381c112285a81f60feddf0c6648d272755d56bd8e3430a3e29f34334f14f7e50baad6762e167d13da026c284abfe7784b49a712c64fe85c0d8658c49d2ea123935b03bc6433eaadd753f8d86d3776df74e799690d8bdd19e3b38d663638779da019a894b79f8f096bf3b0fa392d5d46292e22ede2ff00197c9993f5c40d7944a6cfce18554ecbce7ec280b9fe3f197ef9ee91722abf3d86373abf2967821d012d5630d1c6c917eaba4768ca5bfdb0027e0e628e26d500a6cfe3e1aabc1ac78f711f681104e2daf4d1ca2d476365f7613665928beb5b7e97612b199810e9ee059b4117d55ded025d8b639f5020b836ee909bd090bd6fe490bd193d2f761eaf980bd96cb5c29ee52cae8d5891b2fd3c368d920dca2fac3e8c9901d202451de67a23ca7e245d3b87ce06f955f2ccbb739c572dac51c792db9afca57eaa6e5e1810e1461ac53396267cb9ec30b992c676ff5987c9b22b2a93d0fd5d3dac1d069d51b5e79b227f6f0d5da12d55d16dc172f844b0651d96db9b6b1992de2bfcd0355976c691a8445022daeae3d1298fe042639bd0f36670672bd88093892ab4bc4709140bb679bc5c38088ccde5f0e47894cb76d6510d2b4958e95aae7d1771d846193fa7070cf7814;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h7c705707ba8f39a7e4c91966f1775837488ac39166f2df2055ee313601ccfc4ecdb7ca271c0d97be1694ae6e591ce574f912cd6acab2a047282b967b375c3f5f805bf0f9e6ae0f5dbc577365cf54d0d9f4d30d6fc9292e7c258449115e3d25471131434136223817fd5c3c8e4582aba6c8f5b7414b878a6bd2390f88794f9c868f50708cbddec9c0e77dacead8fa10673b6569de07335d07d695787fef2dd7af2c7c82c1b7a1fcc2272b22d0e719f67ef2d881788d2741d51ab328ac35df26e2fd6c5d96ec960ca940ce092d64126fad67445e3d916ca3fb452382611cd493486996533b3addd4b183ef645b96b62a0d1240a166864eb186d9220f52e2e73123d1b54340958a77f15e5d79de4bee07fe3fb7bef056b66cd367ff7ab4d6399fc712d4cc4f6de21ab9247084df5b4d28eaf7ff05af17dc90db13f442d45b903bd6e08cf8cfa6faa0f934657c619c7477f0412a37db6d30a01b49dd9f632490a1171e8f5acfd76e937e560195829d21909794286c38ce0b0576567db9b6add2207213f4f4960c13d140c011583b86cf7304b768d02071a6d8a57045d0366befe78970994a60253285143d833fdcfd9656276101333b9486f9648c9acdf1c69fe520ab8077fe9fd4b67c75aae8387ca979e38070eb0e43910fd9cb330cce59da56d499be67be1959cfe3024a81b3b9935d56fa40b6ec930715dbd936fef28e8cdfe5afa16a2e09c71292e982cb66ee23b3589f45b11b107b725892bad5d76b276b63f450ec29e10d6155d32902dc655d3c35160792776a82f4e89bf174e8e3dbb02ff49fdcdc4a915e419fb475d3218f8a1d0d8c1dae242570fb51eb3023a78b6e8d1bdebab0e6c5f0b6377838ba38b19c52c933e3897aa65726a5b69507367313b261b144fc5466647e05c1d4d2992d039cd14fcb5d640e1f50422b5b957da6ffc8843846fab9d8244d1d5dec08a6fe98b612ebec996a5b64bbd39ee482b0a9f3d5f34b2a0821b509df11ad057f64e05c275c6cac2321e99fbc5c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hbed3ed27d4ec8eba461940b4a2446e813e5b7e4986426ea2763be1c3c1a95f59c39d928dffdf3cdd29dfd450ae31af6bb12ce14a38253cecd7ddc93bed2d905651aa5d647665ca4f7ab795ad5247382263522bd1870c39892ebbcc5f01a8edbf2ef959b559deec6ddcdab7987aee5adfc58d624a065aa2594b01e0d00074d4e66682054fe003df8619dd8a28b34ec8fe9a9076e4a907c907b7d616400b9114f7a7be7745019f2b5e180d116b53841a76cc7bc2bfe4d65833224df2afb9b90969b5e02ad645d2feb6a5f89e3868530d5f6741f4f27a63313ae8e5a904a7d1367a20d84631ba8e84ede6b0fd9922d3f3d1be21b5ac50d9f09b02868a01f38673918771e5dd61ae542c47f61f079fb6f72235cbbce871d0b615583612cc65f84644914e7188c54bff15b6374b1994ed6ed37e39deadedfdc8633ef0f59e69356ab978226dd727844b2cb0b6a877127f6058f2766282a862d404c92b6f6b38cd01ff776efff72b72423dbaf73cc81554625a27f461b80e8f66d24d67005f609dec41ee8ab5fa91fbd721bce9dc417ce694a110428262e34216785dbfcb5385596161389ebec2e9b76d2f048a876fd84ded5030ff16eb836c0c0fd0ba0b81a677bc3536e36bbebb209e9cfddd9061217e6423f86df4821e2326f219709544caabea52a3776368fa031286d613d35e8fb0aff4b73dbccd81945532298309879ffaf298e32e1b8f49fee2b9a96c5d1f26e581c2e982966cd5fae7a25e578473dd85d6505ebf1878174b29e1908d3a565671adc7ba8120c112e49f4b151ab47619112f00d8a9e429d4e3ed3285ff38cebc010a8f4e1cb4283ecb284a4a610b2fb67ce0ffc3047d96b9ff6fcc2b3ebe5baeb3bf69e1451bbc9d8af282a0007c455c7ab93d311a7d591ef0b93b36c0d0d4dc99650a0f89ab2739be4a72ae410961fbd1bf49eab0cef7ee5960698a3b45b04221be34fe06471ebb325b24b4f226cf448073247e01f210002456a69ccbd9488e06fc538e8342b05918f47c3a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h2f1544e6d05db8748fbd52ec7f2d8c35b0d53904ae26bcb95cf353e2c5726a9c3a3012933da8c8a329a859743b84dbfce08f7a863a443ca7719dc1295f356315973fe92da5aeacc27f25efb81dbde1bbc4868d5381ec248ce11932bc002d543e617e81268296fb5afe41febb2d475de2fceed26978b6c844d3c63c4120a17a8fc29481b07e18dfb3f41eaa74c057bf373032fd40c72f3b3c85da5d6962e949164aad355c6084fd1371b6e6e10d73576cf0c5fbe62b0f5697a2caaccbef316c8395c3ff1139447bc48660e3641c8d2fc1010f73c20ec61637057120c6686443fa181966dc4a5d8f9d6b618dd3f2f4cdfeecdb892d3cd44d4cf785dec9124425ff42ac875f8bec5cb6e12150df693b3e200fdfd6d2eb7b4782cb1840cf119070f0e637a965c23eac6d04dcbec776726b1761512e0f42f894f95aa8d53076d6c3f8aac4a7096d68ac60f09a0fe152ee2dcc03f41fcee0be62af87c65f01eadbd7013c3e6201e38f3a7adc44ef653499ea19a1adbabc01e7c48da6b406340f73c15459a9d8811a9825502314bd485b64b9d2749e4e6443450d82f3f4ff460d318ed829dd50927c81f6c27c742c65595e438d3c3c94281c544b05ccb2813439e888d4369aac43d20f8d94953851b8845075386c8f9af4de8521526302f37c1b1e384a7df76ca6ec87f92e765892b395eed6a74c2e341b1098e853db90192b00da8ef682148f77bc1fbbc8ad6e5e99ef36216a20d65d3f1084fc14eb1d12a81e6153e210c8d9535ab7a9d2acd8f5a21ef920a96ccba9af5f7d55303a01b2d5b3f2561e71adc45830839b9e9351ff67c48f0ca27ed167472776fecec9bfafcb999acc3f3b35c7e0f5ca82e42fb765db46499c028c61ffc1a0289805efb80aa97a569e5eb9493741a307d4a4ad5fd095f153d0d2844dd9dcd8f1b8bbc906a6207dd0609be4a32243d05bc268624d7388866c8a17293b300a202fc89d696cf028a0cbe0e3e19ec9320619b42b2824446364fe1535419a72c8c2f096d87e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h75e0fbaae80b7c90a46450b802e2a4a6886ef1693aa7d2f616f69ffe246730946f0c340f9af4f9baf72e8657a5eb53ef002ac65ea17aa08fdee25c7b9f402f981ddf9fcb5fc9515153c366c28c05dc1e7e9b88e14516c1d27eed690e4720c2248d43fdf34c6d784620cc63b85be1739a98f58637a2945769b5d134803d3e1ec1912280ac713e64045462f0cf08e053e3261f597741db430175abfa36bb0922ac9c2131f246fb0ce9275fb9120ecaa6cc5e38e43c8bdfc29d5524a26fcb4734bc9aac4c109fa94004cf04ad1cefcae10813046a58e443e1e1b3137c78d437f4a23fb99594f64b81bb62c0605d18c5c876df2ec23d3222b0666c65f889ddeaf87392fa144c20b5205949b623ff4d4f952506559ae605105ae1da620c05193c9c6387be02e46a019df1b321ddb50da402401114b3665db567481c0cd6a8abc5ca03a8053053cbaed9b63ba50f109d4e96aab96745a4c9cea4b7c2168350eed90d369f1e3664afc27791ee2d7daa1018d2d0bf90c0bc9abd11c7651c59b8138ec1f8a81bb219101c3d42c970ebad300ed7edb19562ba69aaeeab6ac3e598c985f9fba7b42bee4413430858ea7ae2cab174724fa1c8aa4e1cc9b48776a61ae5853121ad65c8aebbc2aeeaecc77bceafb76951b4f88aa163bceb5d887dbc32f3f3e00dabf28dd7860a9cfa01401501121fd6a0dcac5f81316711ca27846bdb6d305b27850eb622c9b1f3f1c1a4924f64383c0a70ea56d5bc045aa1f47838467b6b83ae5ccb25e09a1f292f144973fc168b2cea4804d8e6ac38cefb0debc7053b25809eafc556be9c6c07debe6d2ab17fdf77afe8129c8016ec9a613174b4e610fc2263131c48b890a9a24f74eaf9f02af5f940f84121067d88de762e4b8c8871e914f28d306deee2399b68d0e3cccac73fd5eedae2cf455c38ba08ef9e1a4091e27111645848102750621d9095a0d92001044abb6b7181a4a701d7b096f0428e5c6eea598de69dacf1640dc4d4071e01b572ce55243aa3fffa63b527;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h876f1b13c924ce8e80e43a6c7c26b6635e4730918ea4898ce45f6d2ff17bdfbb2f715b586fd923bb03ddb9f5a445e91a6c4904a1ba1771e53d42afc61809cdfc038f94c0e702b4f521ca75f082f34436b340f472401ab4e7e39b6323a80ff78a2ae6ab80623cd6fc18566b8a86d5dda38ac38b2c11ae5f4ca7b17f88fd4a6f7ab1b43a1f90976ef06b0501d514d45e9ee7e933c78f9126d197df4dca6ac759f608b2d5f9eb77a9178a841964a717c5b2e7b4dcfef2b67090d31b5113ae430816c21cf12f4ae89dfa74a2b7fcecbfbd5739041e8a57e6f843cf9292f3dae2e085436a98a348dbb30a0ed4b8cf9e758bc6a2e1bda002e52ce9607e27791d0fae76215447291c8c526532cd435ce9962947b24be9b91fee0a266aa889a2537c96f1cef3eefd2cfc968fc44ac6adda19444dc1d162c053db13489faff7f696565daf1e4a9adfb44f37d7fecc23022958ba00c51b31a5bb7de87e8a1a76ab7f9952f7bbd799f231df0d2cd4d1fcdd2d099af8a721778ec359ea3d88001a380bfb882c2e94213ad04a913560be027f75a85d0fd5815bd14bea326d12a99ed3c2f3254a23644d0c1f0d9b4939bcf73b76025342885b1744b06994f3d48206518135b98b916700eeab157079471d2aa78aae35cdece68016d5821fd781b4091f555c08ce7a713f35053ff1b564317ee41c54a8ebfd01a82f81f4e770639f3e0fb964c864cd5f6a5fc7a1c49c976e5b053d1033a9b86ef2b9f4fab2cf1f38a5ac3f60255d6746dbd870a139a10cb2b91cf20491cc210b30ca83e78cc53a55e680ab89f13f032d1a1ea72c3c3cb40df3e48eeeae7acc743344a2a979594a3fde6fd2457b13f5234ff792f7ff2b3d1c387b2a8bf2177734353d8517279cc31721b8dd2eabc445f2268165f747a81a4772b0c2081c3dc0bc60c605a2e9c4456c46dd3ec662734a7ba544566726095ea11bfa9d2cc3a86033cafa04b72159bd72547ca6d7aef1d944143d177b5565cda60a537042fc19f0cba1fc3a44de94c4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hf6c19f801e78a26337ea249d74cfebfdaf412174f099663c14cf2b8a32a893e6d992b08f192cd1ad33fda7437bff60aa9e5bed9663f6498e3d9781602577f292fc1a7a32cf73f74f084fa978067edd2cc068c582bbd743857e4300572613c206bcc297fbb32803f1adc5f6f4067f82bc3bc82c0ceb5b055942513fe765493a93a4779214ef9152a559e4dc0b53c818fb4fbf069e52b5610e5a0757ab9e90f0b79c589fb0f89a67e13d1811109db46fbc28d803cada5510c340023f8e1f5099e3906a0369d4b3844b9c2ec31f1a2ce60be212c71d2b98abd0b526dc5511cb6217c03f180284c2ff4761cfedfff9f22ed4754bc6e78cc502caaa781dd6b96a559e9bb94563e801fff061cfec303070670d56f50d12d2ac1168b41619ed0084b72e25c5691fba50c7d166c8575ca216af048458ebabfee7f1e4aa0a3fe676757456905066e2506db42b238d0b91a9d6514cd0cb9f9b05ac93ed78b6615bd4fd0388e31930ceb61397393d3c6030fc8642124cfcc03b18d2a362e66959b0181a31cb62c7a8ac49d95ff9a053e53a92547b6b23f27285218643866bebe41ae08c03e7eb4f65ebd56dd7f94cd93ed907c9bc9f94ae623fe7895fc87ec1fa39a7f928cb83455d468f7e3e1e46479d6eca323c6261486b74ae5dad54626c91fcd7b753e858b14c5aa48889359c7b7bcdcaefc3cdefe1ca760fc16ff2902dfa09e688d5cd0f7ea153d35abc48c9867ddbcb9a071d7d9cd210385f680492bce126f563a8718dbb8100505c6052035b66895ac92bde36efd20d4e2e4b3d1ae03e8c88795540c3d55572ce4c9e5c114b44719b09e1e2c1c36465385a0025cf41280710e2f114981ab32f35fad53cc37824835dd63816eb16914a4c45d5b964efd3b0c3bb00c5a8c48bede4c7c101d86be43c9eb4b506e97480ed20bebfaf862a59c3da4529a11c79b5828e391e01e54a3b9b51b6d46d50c6d76311bad78ec04c19343e407ffe5924146fb86055f56dc355721822b8b5de412c5587ace9a336;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h7a85fbad4846cf4d435a7744e7ab0229632eecb08ba3b0dc0e8afe1f170ee39739a24308caa606366d7db5319f96ab1c6a3868f61fe78459ff3e60c484299b93e27864aa7091e09e29101e624ca9cc8454399331e29ec8332f8d5c80baa3d606b796c5dda3d9774953c3ea6b718f1abfc1babfc1fb1e2a2b789ff27428d8955187a656deaccf1fe95facbfe7b608465a2609f99850ca54d0e2dbcf92b3c59b0dcb48064fcc3b30de66a35390fce066238134706887c2645ed7e90e40b1ba28188cfa5b3050baa433f086c6d3d10c793c0a811480d3f3bdf2d06be13b3c559b91d020773a4d39818395f4c7519600d929d950c3ef4d09d25356569775e9e4e0e051776446d3594c1c60e4a9dfc7002441468a2f08f7752654988bfa295871c8667b987bb0a18ad167b8b199c21434db0fc0adbe8f9d2b011158f81b37f24194e97bc703eb524f924d7bdb06bb3e6a85903b325b1f63ad934fa2da3cc1297f9fd79760c6dcd841c2d523fba2708fb40b0fa3a8dbb0f587a0ef268bf809828115b1407cd68d1a2e827dae7532663600f8c9134551e226469fab4e29b349496627d4b9d25ff8cb30c554a30e94ec930e12036c29e4107caff038983c77475e0e1610e8cb9b9fd611ae56cbbac663350a3d74819d8815f464e8360912d6d1fb1bdfab0ec9c482ea28f6e147d96bd1856eeceff5d853f2ece69611ca0000871f9a30a9a6d0686e8197d14790343d987a280c2dfbf2a1e63901ec8dcd7316d9881cb0ae620825922ca07c247cb49c350af776ac4b40d1e855aa3837ff400fd9942ba2bc28e3612c0244ccb877d2c6c7ed83be099d8a2fa8523421f21090e8e823c9cd1d561c7a464dd961eb68f4379453c47f88e3ce531d8c27aeef81c5ac6f74911c147902966d7ecb01a57fd27742e74c8054d1e1d31b025fc1e17b878d9b77e902437bcaa14c10662afd847dc3e0935c2181581cc5f12fc73d278e6fd0d98a5bb36b3d7bdae9564fdeb95bd5b44b1f790193280318c86eb56b9c6f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h4fdde32f7e71b1be67748fe312f31faab05c5de96377947de8886dab87219212df2d1b222f140652a5f82b1a3aeda2fdcaa426cd0996862be2d5244016828a701cd7dc106aa163b29655a511e671fc2af846c3705e0cf002246ef7469a8e8534043b82583e302a670d6e9a1d2e2a0c0397154379ec2e51ded8a0a53b6294ee275ed2e7694b424c13447db7475ef988104e37786f327885fc82f54e9b027822e6cc0c4abb95fe86fda169e2184c398e8257802511ef6fc03460e156414fa7601256d317aa321ae04e6661b76bda8267b172fa380abed539d7ea6bc306b8f9318466fd8dbafa102dc88e2a8a711b88d1be80935b1069835a161929722098b26cf8b87f9ae8d65c20005e87dcc567bff4cc582ab18fccd85d82d72104963e781a88f7dbb05a27093c9386f259ff5a6a35e875d2ff891d6f277679cf4e8a6cf65aeb86633bab58cf4577169b42117d7134195bd258e3e316964bbcc749794bfaf26f97f93ccd62d829ad25e16dc5b9cc732e7531c8c44f8ac71788b47e5337c446bcd243cc0da31c50660e552ab2437747af65dae3d812fab2fe22f81a55082f2f50792b88c1c76a1765697ca5e78b24e298a3ef5887fc8083e7927e66acc56c7c1d0073de1ff1991ef5ce522beec6aa558fb59530c6be4b257889491ac9de5fbed9a8be5481cb5d6e8db7aa1f83434be28bd42643d75dc067827a9e2d53099cb74f5c81d05ec22957be7abc40aa33b988de6c5defeba7266ac3f557dcba4df3db9b0757908174bc9f2f6ee5cff0544ecb314fc6f49cc94eb692a6011b06ce624f2e396a77ddd9ae6436a8096dc7da318636ab039932f7238dfd07166374946aa4053c44168c247baa737b5ea51c7f3154c189ceb6fa4fc2bd21122e361d8ca05f3dcf87e4815f3d0f5bc27ef0c890e57e48570d8068b7efee6d06c7f6e7a7f76634e030bf0a9e6c0b1b62266dbe25891d976c0b0da424eb43537a85b08eea2cd80e02923ac28248e6bd49f4fbfc91cf11672a2962d63258066950;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'ha92b09a8a0cf9f396822af47eac5f7a695faca5d3848d5d50fe59531aff81bc659d84f639e082be25ed98eca1c8345c30e027f9afb7161b730a3c2b9931455edf08a89c8cb8ac90040d8fc931fefcda55e9b0d1e36755f1fd1aef2140c16a73bba202d17c5fd0cdcbc38b2eba8334d65708cb9526e3d8cbf655712f4dab13df6dd38957fdcbe836fb3b35c4448bc2bd59c87f06cd8b669a416f277069809a0ad373954a8a96a4803bf474037d239d8dfe757d12e1b0e35bc567634928802467617661572575e3285061b92d11a4666ac1698d4f827210e99e095ed03c16cc087eaed021f241ce273506b71dbe302e3d7a4f57701b7b7134075dafcd9da00be2a9bae3659402cf6ac92c60fb3a2426e4848328239ca31b4250584921f886a7560a8cb56bba7aad19fa3270d3d0b132511b16b6ca8e215b24cf8a00edcf6d46117a4c1c7665fdf7864c7208d66960af05d623e4674fecd6efe5c5fc5aaccddea41cd73dcf3408029a369575f357929cf27f56152e58aa6809ef0a11a99f3d9b097620bb5529f0004450054125db3d9fd735abacec1958319632f8dfbb862edb656ec905f75cf20e4ef953e53066fb9526beafb414a25aab88ca41bfb4a19a8248721a9dfaa846ded1b5ec531b0f5f40d8b46f88a81cd857d243a1448a4c84fdac907376f8aecc466efefea61d94dca611b2f55e1be0b80094216c53c3ad06d4d78d4b90f233e087995f7f766481870e8c4f1131be56b8bfa7507339b334ede160e6e6b14a96c8b712a6e23a06daf9ff9ae7019868f0988c21c15b186b61718749a01f0f2d6e7c747d4772a706edac3b900304755f16ec3f8fb2535e0fd938d4549857b5613053372b6ae0e3bb74c46a7ac8e2a3e2873610eead43f784bfbbdc1fa6f5296e061d194ff543bb7e9a6d44fc3f58e35d6f572714307d9cfdeeec7366b363d050f7f392f6860bae6b7e20476e6d4ee440235107f090e7c290f9dfe68fa0c91fc9c7eb3c2316fb9586938b4dec1c1273f2be3263473e4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hc2d3d9357a53dde4ffff0cb5af361c710c1d2e68e123441f8440edc7740ede152277c3c50413bf6c3d4a2a1bd3a0e6775a147ee88b3c02aa26376292be6d39f05a7c534bbc5240555a72c5f9ef56f0cd6c8ac89fa0f92035082e4d2de5349752d046e4f529dbefa98ab0eb84f8ec57cae0540057074b6073bb4d5ea0bc6e6cec9d73a87dbe5ea1327a4bc7257031526f2ed8412315bb0538fbdcc1229f2931e6619a0b3ddf6757b2a4626746bc5d83641aca0a78232a42d763f45385a720ba72e27b28fef2c84031ca1e4df3c6de3a8628bfad296835a18dad349cc898dbe230306a8dcadb94c8954262150908f8f0a7e0af3a3d0ab0027c9b80285c0258f2ae2e0ef311ca118e35e51bcafd061e127af0b00e17ceee6341ccebac54452e14ec5d5af228a99b0ad3041457fe65c8c085fdea3e66ca351101f141e746cf8a100ae89934d9142c4ea49f89d09f7034fbd2114a18f748de7f202b63d31ebc08bd8624f7af69f4e5b73e8c6b2c8a3f8c2c8d6eeda8c190ce04e75dba854ba534c18c34de72c233ddb14e22afcb6ae72b819549c803836efe01151aa6e06a8d168fc61e7bdb68537d2ef514769d173a932214fa7f75b2813662bf50ae6f973e6f3432a11ddfddb83d582e1eb35ca99c31b42e6939c4e8dc28fcd21545a2f95424f1794a772fdced2cafcbd32a984eabeeab35fde5cc87b4f9646974a264cec397c14fd53ff7f58672d92d866a5e83b9c815790d1a4cd629f0ed9a19ebb3ed6913baeb8a39c93594e129c59108b12d28470fcf6fbc7ac619f70448371e954801e310ee4424864c917b31e9d63ddcc0ff438ddd1a629c5d3d90080b8be7df52311025677282463f115454aa8dfffb64634db41b8457781178f7fe7a988e60cbd0cc06cbd74078482f6273316350899c0c4cd34edbfda61492749278e4d722d43bcf672708903a22a35e32b2a56e27b574b4f4ac9a78bb2344145df8696ebf9b309b675c4c41b292b86d1e789771458ec2e21c19075f6aaf4a405cba0f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h8c4631d2220592134519b723408e45d18d5b07685247b5581f68e188b41955e32891bec8fd88fe54af9e8e80d1bc4fac13be27920dcaaad4952566fe450f4c631343833cd6f1152316c7b6a9c00c7f5c9befcd6c35b8e77114cfead7ae7ac0ddd9e52c9b694a6bb2da2928eeb199372621dca69d72e05e082a0c470a91ceeb6f54a501de5e6b0f8c471e35d8173622ea5eba2c4643746e70101dad4ee638c4e9564d8d17a8119cf735f7d63e572d0a8d43adcb4d55bf3a6624156e39ee5dfb5265525c2a8502aa1713efab872154a80c06b47d84c6e2456fdbcbe154ad706addb7a13d9b795153d3c01a2bc1ebaf3ca466101e4ce16f9148d69188fa3ddcec15d0f56039d01c4f7492d0f3439cd2fff4a794442e56ad5b9d58575ec60f137b60eb59b6eed1ac797e1eaca22d20c9e0bfbfcbd5b1825b00c86db28bb31599ef74b1a9fd888a85a5d72623d13187cf4598a327efc78c14c5fe1f30ec21d53425503ad0613f1dfe4967bf53642fca0a95a9490555157c1ac146fd38530b7ea89595d8ec926f00feb1fdf451cab9e871852737f26be54dce82c48be924c02898cb55d8e748be4588ba34144535ddfc7c1d3d55087214d51ff3348c87ec9a3e08a55cc108ad25b0b0cca7696ca02d3f7af0ffe3d7a8c5d81a995702f70778161e24249ab83ae13474a0ca2f0821f0da0caec101989ed0c22dec1850641ad030cdb8a50a5c37d41ac24c8277c94903011861127b5fc32f150f8cecd96be1cb046d68e08881e8fb3d057af1f0b2bbc46b47a5256a4d0d2a82c57a5f8ec50e1c485dff495a369ec239a40691dcc96e54412af4bb42751057f9129d6380594ef9af95090e1ee86566fe78e14569e5fa8c0ea3725ab64c824829a3a10cdf94ae417756536bb0f1d82831a251656b93d07b10826e7bd69b4e160644ebb2ca592910c200d5cf6dd5332fe8cc88f37522c4d066446aabf544490c9a9a6d393c737fb0fb04692806c0c41ea220485f88ec7e4ecf40f13d37a2f5c6df3b2a48d6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hfde97505fb479aed5401f149d817cb3906291405fcd3c54d69dadb914137a24835286bcf657be6e2244ac5bb4be33cb5fed7a8dea15359465850ebcc4dc77beac4bdd103f45925c1fc6c6b3be567e174d002da95702e27effe2bc95bec6aa62677e2a64bbf0e73d346bada9ea44010023e62a4891673d1091786596e7ed5e1f5b2c9c161889fa1af55e97069c4996a37381d2397a24f376803aa1c1ee861c0738912f8846ea46ea07c258fb21301eddf62a3159f2dce7dc2e0d93c8cff102146da90003cf7c03d8432d0f2c47b4edda2de6a970b7a6ceaf5e9eec401df8cd0646a65799a2b74592846e6939a77dc620ab4a9337a10560528e0a7419c8dee97437b724abb8bcf3b22c09ccb92fbd373092e121392f58ba7d2f2417eb125e3cd0a251d5cfed14244b6dacf58c74a156f30175e3402919cefc9ebad330364a7f42571748401ccb1a2a4307a01d3504e77560bac57a807b78db9c00c4705c2f9ed186bca1b7e580656901d8575e1e3220d47ce85f333b20702d5bf5036e7f5d1ad950cb0ed644a0ae88a4983ccfb94823a584097b2c8f47c9e72c12aead4fd5d72ca9d4c93a4bed3ff11884471224293cfc7a390af52db617c1773304d89e4cb61e847121daf7aa8bce54e28a3d0f2d4cec6de667932ea92c2fdd29eac0e134004b5aa8f6897b36a541b2eac6e755473ed8d6f293ebbab85e236310a8cf32663372237d32fb94f3736f782e540e1e9ae7bbb692e223b32f828f8f8fbf3262cee29729694923335201c895f858aca773cc918e0654ae4395476559a29f6cb412fd37bae4457e09332d875f8069b63466428e3c6824d89557d1440d905cdfec23500e3df57bf16edbb462194e5bb6b97f664c136a1e33b4d6116fc74032b2a2367ce815fd3bc8fd8c7545600f8112c4fdd3fba72aa22b9ac805a30d17de08e659f8d443eceaeef31f9f4d8d6131674a683983cb5da90f8a97d16812dfd8374bcfcd1824fb26ff7638e9ef3c5ca627dd5b13836529a0d077439afe2ca;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h9af4c489dd83cec6afc1a336a30725f04442155f20542a38d2bd96c651e4f997f972b63842fb2e59210d43368c2bc9f9bbe6e300f39c05d008852fb3135fda7a458240dccc205c998071fb0b77aaf6c305ef3493a816e143417e13895f3317c41becbf4a5aadbdc616c79429b4c7f3c53639ecb28db9c9494ce6261e5710fe36ee462f3bc6e3ad53925c3df14a201614785779059178d20118863b3b536f774f6628c562a1ad90ba28bbef5cb1281f388cda6d8d6e1c8f36ab55012baad4aba56d3f3805a095a59883dbe0a732f10bfc704b80a6c32215d24464ad934ee40521bd814a2123a8f6f52ac0a06b5ddf550440026e22ff2892f3735779efaa8ab3902bb4fe6ba419c693dc9876ba0342ed1c055b40cb68fe57a3ef522bcc1f2ddd64fdf08df5931f620ecc9e84f34e4e9cb916aedf40693e481bcec027d9f59c04ba34d5f057696f14f8709e4f9bd2042551614dedb9d1158c493e85fdc225472c7a03647eaa1eae0b64dfcf66f36a6ac0fe5491a94476cb400024faa071ef3877996d2c7f8fdf30880812117ffeeec4868768214326c4c8e39af8e89f4b4ec3608559c3d6d7db1ba17a7856c505b13900c6d15b565f8f41f131b6c495c2f2c4df72af7f4a50e4f2a3db98460950e0d8697afaf09034ef41c0620460f4000e0d65f12daa69b616b8672920842b714673280f5c21b5824cdb2b36616562d4335b06074ca91c065e67d27d6a2838d1d24fef2d2f61a4fee61cc8511f1a6aa5dddf1d08c58bcdc07b55b3a64067664b35da0987d39d67031117b92d4cda85f49c368ae3002e81749b61f962e5a17b5495bc99fe078158f735353408569ce491c1624c1f9a0a4a447fba8ac2b5010aae3e8e5addd4ea74c6f60fa1bd8681ba5f81c2695343bd23864ce132818622885fd6cf8f38db083f0a3fa181294571449a3f97ebe40df204f0f2aa9ca2453fe142c8653a22ba8191f1485beccad9c92a5907fa91a5ef3e7b6c9cb1c37e33ec0fa13ffc0508e01b9911e8d1db5a6d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'haadce4f365bb0b6f6cbf7c2f74166acbcdae6db1180ad3f580f6c34ec6e726d419676190803d319646bcd0cf4168221ef313dbb26fc90983b21fc9e05af6492341657228b51fdbf45ca65275dfa085968184ad8219cb6bda31939f536b4f5666aeab10d587c26d43a538bbf7f34dbd694ed8e8a51fd318adb4c8b172bdc35807f9ac00a9a9a1cd404e62079f6df535b26522d5aa2bc1cf3a8fd73433eb9970c14e5e4dabd68e27aa58c1f88b6e3fe12fbb4ace1d6e0520068307380721eaa7110cf68f93ac0e03e70f6e02b7fe687cfe01d74547c28a5c5be6351121cc32449b2e0df9225d4a08a2f9a12de1d2d326ea53786ccd34467976a8f98153ba14986a533d1a9dd102febcb187b41251fb3665ea6e0e14ef09f249ca01dc0f191b90b12fb659c091db01282a32ac5b28ef4ceaaaedec35442b9e759173f9279b60b2c44fad65d9a5a422f8537d9dde54925c25490032720dcd4356c203dc5bb95254b0a98e5c65f05b750eda6f5597fad30f71147b138be28ea51a960315c4b3da81283f751911fef14995be8c543d73c565be5881b5e77e1d15f91c4a4f95bc7e6aaa665b4846c15f9783a4f54ad5122ac91352214d93454044a1187dcc4516928ff47e5bfcc3d3144bd5bc0a0ea515750896dd95a40393a123c34b7d5b576a632c1cca1b2f5a32c4098fe5b56b20a2977a0fee6282d4b33805c831ef3d8d96c3526e76cd92f9c3d56b331bca454a43674630f9ec3b41f88a35295f210d87162fcd52af198388583c7600eb566f6825f173327384939f282a0cfd28894221af03408424548ebf9904e7a2aa98c8e0e33f11fa7440ede695b66316c7d88e963b8fbba1f4bdf3cbfbcecf7117b404aa6e7bc92168561c047f5b032db6d3101e705f5a99fc58ef629314f1d48e8f4331620153f528b9480257072925c3da3ca27f2d86d467abd2e5cac6bd63b4107521cedb623fcf4b28468b16f87462946a18b10dfa4044986b6c91e2f2adf9141b613107db9ccaa7563fe802d3ea9a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h9df2676c0a458108448c2f6a6a4ac92f369403c252225d1e17f7f453fc449c705cc143d0abda8a88986a416658d065943ebaa14d6b5165e66388cf7845f695cbfbea9b2456a8749bcdf481e81df263d15b4d1a516431c6cc452f53755971041fdffb14f093c80474504a24fa22c53cc9f7505072b98a2202c2d3ae096cf16e0259800e375ab95a21c1849d487361078ab46099a0a891c51da5f903a2847e2801a4d8ad9dc76b228aa543e7830d32cf9cbe3a3c3034c53f335d7fd9f1adbcd6f3b65e7849169446b1e4da8c066ea7e84c815d4e2269d3243cd8d3588d724d15d0a3a5038e4f7c72e1b7b83d48b432ad33e795981854a60389060508130356eb18f61e2f8c57b45463759714ac9c13da20e1d52518b2fce9967013ec3a2e0c3fe5b728de70f45734b2a8a0b1103a3c8141efa5d7c6142e4912b3b97ce2a60cdd8aac99e35f579e6c963c895970d510e2d18b22329a569b8090becfe47b704d4e899825f41f274715b1c9d4b5baeadd9ea2d1d24e97655785feb9b6f61acea94e8aa066477225649ed465742958b3caf6343400e87a6e3266d83e02ee82df27ae8ceab3c859f39667c381e2e5559a2569a019984a9309802291ea605ff53a9fc28908fef7f3e189285518e2400447c73bd8fec06364686d41704678f3ceed81a1e4a010614666dd209d2cbbe2134d0f0d1ebf1a7147eefab4d8d55c3ea9353b35208b1416e16b6799d33f1762fb565776b6d181ed8b4bcce41533ccc431afa47d849468cf4fbb9bc0da242740704fca3442085e2b0a0b5e8af6718f3c3a58be884a4bc7e5bd3f0b50dd9a3c823abf55cda6763cfe725a48b60831cc66298f90ab507990ee266129039f313548e14e0e61b6c4efa3ba1a3ec5f02bc41a086dd1f9e9bf33185c6a0c3a56b5d1989c908974463f0763f0229541e36122afb35b10c31fd113ba11c9d539615a8249b4e311f8457f8cda2b54d62e99cfea8b40850ec32a91ce652b110d6cc82b494ab8808de1a9e2145f7abb4afc2923;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h49c161b893a787ac62243b43506abed7b739ba25058f48277920a116758459c05477b6e475deefc610c9b78991febff8a092463a0ce2291959f402d710abbdd53256427a6c6b4e01a86463266c4e1cdb0defaf613db23dbb0a2c491b0e2f4461476766da2133b056e686679c13721d8756d1f264fee112213579dfd11e991c7ea2251848649edfcfaeff20650951bd621c6cbe0411ffb14b1ba7a1f2b15ff5eb928eea97a83d52202efef67b4c3c4e153b548661b5fa2bf35cca740a2763eb9a107a0feb40804cadade48b588d8e16c0e9aff8e6c2577c466ea140298ba12198509a20b308d44b0badc402a02c3c88d4afcd70e984ff6d1fd9961beb4242448d74637655a8dfa8fa1fa9369fc7787b80cc8cb55d9aa84334255bd05bc737eecb08299b8f057cf1966983cb31fda2a60cd9b420a2260ece056a66dd0c4a790089419815751155710c45a063bb46aa6e261ea18fe6cf04ddd9852035faccbed1ba8aaf94bd5bd869f396ea97ae91c2ec54ecb986f761574cd01acb78d31352f082d9dd7ab575c041514574210021d7a8af4b66e63de0c0a3deb6bd91ab564169545e17b0bfc84af2053fbd4fe5cc90bf3ad06765b2c4bab7dcce4ad73a7e68cbc9268ab32820f2049fe36c92e57f32de0ab52b0a847e758bbc764b1d9a296a2d0e91a10371fc4f066fca35bf2222115ecf777f165e3100aa96bbc1bc39f207f0c77fc5031d07933ff99d9fb20bb655623786675bf5f5135b3072df2053a2d95d6b0e0885edfe6fb4de45c79d59170d1ee0f230c5cd746ca3f62fc819c67e13abf493f9c91b8cc519e6a08c7604f0a66e84078552ecba9a9a1f6f2d8cb2e259190969998a4dddc1f6eab1baf5f56e1069bd1f704f816959c90ab109e349cecbba48a99bbf0a42fc74e60810832fd7457123786d31fc43f01da854cb3f15758f07159672323505bd8fcf9fd4c8025baa85ddc226cadea6308197b077f259d6f94dcd52cd5b74145c325c5ddee5fb2a8cb8b4817c398d6f59af0d47;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h1c33063497128faa9b00a2622b7942ad23bdafa094a764246a7e2e7e3a50fe330941bba19a93468430571abcb92d8cf5d468e8abbe7f267cd3f42366c053231e4361fe81cd9ae0f4a85ce9f585242fe00b8fd109f8b65c7992dc258f10ce514e2e1195944ef707f5b9d8bb53378193504d4fd21bec3201725cb22767469dbe215a158f81559197539451043ff177567fecbf0e36482099af0a90a7445918ae658711c0c177e2618dfbb40fbcb3632e7dfef1e683a6af2ee96ad56dc89995c0d85ccfd0b96e035ac3e8d08bfc9f7b96e7bc001c04f8e3070a7eacdb5da8d6ed8b7f890b8d95ad260018c3492d7845cc93bbb7afb300b386ad67bd802f3bf6cfbd6f4cbac13c9494ee442eff38bd2752fee901dd96b9cc70faca3dacd39a990d1e668ca6f29aa654304349760808b56ee4063d58ab68ab080d691b9be94f91f48cec6d8d29990820ce7e742e7da69f4baf5505dc494546d972443b80f6a5368b4961dcc0b2e82a26c1d5af55cbc253d186f52d4c4574ca772285120eda69759751da29dd3d4a4257bd5217beed2684804332174fb4fe4375eea296e17b58cae6a69ddab64fe320ab0567269fb3b9a9cf98db9be756da5f2e6f60b80ee9ce31286893cc0a29da8ab5f3efd8a81e4fa89161110eaa2def35e244c192ee56009b3c599140cce98188e3bc2e25305f47bdeb82f90678b3bed4094003a4ed8f0789f11eb3aa920ae059b310e5069da93866bce521083403327ed85b862911e7814cedf87344ed160ac7e20a06f08c28d49b4bcfd65c1deb1326cebbdae3166236aae19271db54db27614ec81b6cb82ff8d49731a5917d7e3a07e9aae99dd6b21c26ccc750776e06757f7a120be2d78632c795afb0740dff2ce47d68977baec45a534d579aeb8894b56c5dfde7d6258a3787be4b482375ccec0cc1a2b74da4754c9b993c5d4e4630f08b63f5c74f81ec3539847e24f603db1ab349dc8d55c9230bdd8c43f085ff11477130af2b1a86f198c0cb04eeaa81dce25b81dd8f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hef4c026a735bdd0ab8a222b6d0f7d40c72bb7016578dfa63cffa03da7595892a9682028a275ee4b90e12b8b183e994bafd2b16b28b2bc857a8eedc36b2e0de08a843d9ed34debc3d6d507ec6902dfdc1bbeebf7b4378cbebdb707ddf2b45ab7a7b3f219ac4166ddee76d4ebd7cff7ae88896d34d3a0de3faf92fb82dd521485343c29acfbb586226cce131d473de90a3556aef08e83c90fab78dfb3801fc579fbed8f54b462014ec2579d65d7b7e1d7e5babef69dac819784125fb0c00e2ef532c581f6279e9db7357200b85b97c84df7b769d9d124aecf179dfbc4e96fdf4b8c45029a4cba53f5f91c150e0fc57ca40a2d301c392850d8e64d0428802169c69d4efa5b525803868812ec8340cf2bae948f3fd12673a66e90d702982842c70cd661b10ae58e38801618be4d1add95b9e31406de430bf3e893e0950e9f352ce379c445565f2280806ee7f665ed96bf8a68db16971f3b502f86d5ce3d34db0143a1376ae81e7287c5bc1ea71488addf181dca4eda5316ec644239f2b7aef8c1f39b11a86ff576e82ad635cbb63fe1c2ab14aa6f806f3d9304c1660f9e3b70133575ea003e8fc61e70d6432bb4ba7e9e381c0a2419c4f7f7a01d5cc77ebe1df889b0dccfa74b6f9fa3875d6edcd15fb062bfb02802de8b65e485feae0053431487ee4fd8e6017597c0ae7a1f53d17868f9dc1c18dacaca4261bc167fab8228a022dece9595cf23b7612a455015e0b95d1db7ae2974f5e908143f5716f432bf8f18c26eef464137968c87cf3d84433e5a03a9a25fa998c3c9b3c314bc8efb13738695bc83223890afa9dc4dcf247b6d7983c5e40072d35ba5faa5d32e3757c47e8c8c51c963de33c44d5bc19cb6ccfd6ffd3a028b1a8c00d290dd4e61db86369387593659d1598996fbb4fd60dee1221707ecd8624659bfe22c74c0e54c77e7d2322a87d95d7d24d792aa06285a9f5ecf558f82d27605bbb992ea031fabaa64cddc79c5433937468533548b5080f26713e1b4475840d1c8a950e76;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h4039efac1a6aa5e2fdf35e35d1e402637382a9daf0d9045affb2428317d445f2062e704ae1a051a13dbeaf6492a7e2e881c90a5961eef924c1266720ed66b1670a17ed7dbcda20e81854e050a533b2e933c0bfd1cfb42c15abee778ed2f4fdcfe8fc3602f148886d6822d020b15d3f2a40755b3e6d8e3297857879d79a690ba97c64064c3bebf1f98243351ae3a01a0dcd0fdc56dc9366c469f0fc88664a44a629f96788149d61fa65b8fb31a6ab08607fca8be67a4f44b0d21914f11c60d267b706edfb7f42789225770f4ed8fae26dbf4cdbadb06f08d117130502d2a2309c91f23310a93d071bf1e238844e9ff50534887803330b30f2a178365ae7d4ccee6360447e8cbbecf4ba8ddb864bb869415ed1dc975ed43dec69476ef6a2057714eac55e2b39a587460dc8a0f5d6d1127c67331d62437fcd81ca6e4cfa5b3ddde4fd35279233e25976733578de437c12b08726504a36d1edf92e71a9b0cc39191b0ea5f5af211f1b5c17c9f07a05638f38a6c2db0b08ef230d957101e68ce6404d7e69a820e8d609c415657feaf00aeee57ae1600265e7a99e6314d127e4b5b6d922811c5e3f6ab20e2f6a57214c6ab38589e0594ae76afb1fb03a0dcc9301ecc1abd54be4d0e1fdf881b11ffb4745f60ed35c03b1f6c9a1c58b40803728343f1ad37148f3e6e911cceefd7df93db6bfa80cb82a67e4945bfeeffa1d0f852a12684fc0f9ed453b0126ad6659b743b257c70d6dcbacda1401c90a4cf280bac8fa456eb48f3bec682c0b32ee951080027558802808ed5e2b085b019cabf115ebc47ba2fadd635a6af16705a8ecbf591fcd016c848502093a39b8e0e8d418dc7a12d75b9b45f11873e81bd0b6d1743b27b2af06b867134d0f5f65dc75322ede7efa630530a6f12c6a1ec60ceecdc43df6a936690397e0b26693e8e90f7fb5612b9a5174611d90a21132208b77cdb2e8299914dfab90ef5e559894d0aef0a2bdfec721aa0094e368c544d0c9dbb75264b0aaf620e28969d0d8515103;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h6a78c40501e6b194883796e22623239843b4397171442cf717b5a7260b713ead3249dc73b6ccd83829ca6b4b9fcdc7b57d398f499c3c69b5e4b5c9b936b941f7d0c96d112092589255573f7949ea30c91d90766e8734ff21fcac11d6fe2714d725c3240b01d51769d37d3b99daef484ac6b86ce96b5a40b40a67afe1863e093b201935322181ecab55f6273ccc00f85d6a1ab25a34f82099ed8b327165cb60d98766a30d1939b6258e8f99a88eb0c6b41daed6575419e280bc81f131292633bfd7c5efd737fdf062787d16a2eb9ac8d65e83c4a4f495e3f8c4d2f5711b24c0a4351278b42401458f5db41e1a6247f809b1fa693a98a1d79db5271eb0d8b30fce20b2dcfbc232fbb39e5b250bcc7e3b7d19e871379f8782dbf39af7ce70536be9ba25bef285b7554a40b196e4359f8b080b73df291660de3ad0288389aa9abcbb54ec8e1cd6b2792b5cc2d87fa850d452b9ed326e5f5b2c3c97caab9f6bb514316216d32b464a67f9be2177e0c17cb86c2586b9b2219cd13a2f8b078a9c07884ab45b9f1436d2c9712f0695ada88c50fa83f49df628c8cb5ed82ca52798f66b4d1d0b463420f934da8ce5c0762029ca025491f66593bad09991c7a3a4dd780ac3e7d6ca76a14d3776fe2a4312029d1386b778119814817c19523d890afd18d7fe8cde2e523dc877e42908e9ee2517d004b944fe0e05f2599a7e93d5b36b7c6e9625d36aaa4605fd28a26728b6eaca6ca95f41eadb9b7a248b26fe62d1a44aaa5cc557b1ae8a889db0e3b45e984765f4dd5b03e2a18856f0158650c31350b87c08f3d880b1752f2ebd4adb3f7fdec89a9c5f5fa7a96c716cd07195c294c91b0ff41e6b104a73682836e94b3536376c9f9c821ab2460dec8d64c63578e80724a24c906194d0e9567515823270388213ef3a8aa23fa422164f0440689124f9b1596fb37a4d2d5e4d56f51edead445ab1b9944faa6023ba2b3d2c1a0d9107e6b4a695b23db4797b07099ca71614c514b25fccad3492ef873038f579;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hb20cf68f11840b833d7a25f9da093ea02a0933a2c67df62054ebc0ee3179e598d408106b828a4c1f08ea0ae80d17a09c5620ed885deb912f3e07a941e7129eaee1b610496c1ac590aa631f35c1500eca1488f330d3d5d388cb6d50b6f5558959606c77fa8f42b194882d18373c5f51f0d26a74bc0f1b1516e4701ba14cfe6e1837b67f8b94edbc3e7f2205d708b5bbb05fad0028ad2efad324572601bb102882363c304c3158ded1be3184b7f5698be4820999b54373132aad4a7b4560e99d54b690ef8b0b223316841e1367377c61ebe3ca50d1542b0470d53c26603c421868fce91b0ee4e7053220af16fa30279103decd69ad4992b0c02d84d33dbc177fa38ca6a45217d1acc8c245322eff150a6b495729ce178325c703775d0adb19ea103f358cfaab5b62c9dc20ee9a82ebb3c20706a761458770ab28c9260d078d77251930b5381850ddbf8e3d96f1189a8655d65fba56400b085ebd93331358c2712a0ae5a8e2c573489cc9db3f0e7420f8515dad1cd8fef6f1f1e1eed67889dfe4c22c7996c914fd357e4a3c8545c099466253f26cd73dfabb68a153b96a28d5962ba34cb1597573d06790f7c623b883df5a587ab0163d72f4f6b37cac0e9d5a5367eab635357eccb4b170148bd9cfb92893bea372990e3305a3448a3e1252d28a4661dccca675f941019afe576df32529d3e82b801c69c63a36edfe67de9364ce7c5c2e8f94bb08e23fe4be678d853601d95356713dcffb0a60b2ef45aa3940ea47b8087dfcfe060072230346c1eb1f107e195691677fb5288b8427ba4d337306a1e0d5731a43e5960ee143fa6f4e0586bc8c713715b82514c9973ca349c9e378c50d4c143e64b824ad2d7072a299da3c82b1142c8c60e721aee6fc11170797839feb168b7dc02ff2a0b02b1b245bb3627eaec704502d08c37241b295e5ff59d93ff9019be787932f6a466dc29031351afc89b2f32e2d2209a7a7b3f76ab69ca838863680bfe560f2b309234fe576a3aed39bc7e69893b4aed59a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h6f35731f1836eb212e2aab4aad628cab88cbe9e9c6e8b4e351dbf118f54f2d14514f63921757476d8384ecd50ed01699188153471fb9dc02459b1e898212de47973cc295246f3b7343f6cea93c53de8da0209892f611a05da37551b7cf37c4513d9d580bcd345ac3d7fa78add5d7f27805056fb9c20231b342587e56d712399e45df512490825ea7f0bb3448f46c262f9f8f4e657579d457377637a6b9d5e9b814f5fa0150f14dec152917fad9c54383498e013f20e4b5492a6552abfd39e9644a1f90f2dbc4088cb9bd672f78e3d0265594215c36b0ed6423a930dfaa7e9f9a0b564d34ec4909ade68ede60c158cd0be23b373e8a4e4e760047e25ecba0177f81ada4f819b9e87aaeb766e59e5ef0bf165e43019a94b38d07ac691454333fea3bba635f8251f6d08441f12bea2f4e1785c736615e3253df70cdaa44977ac01feaa4f1440141fc9d8ef186f57b8624671dd51facb3c588972b0faee4b10b6673c52c9be9b3d8f41e7c554e9ee498b670cfd28d95255c0a495ae0dee4e27953246cdcfba05da2ce7a2d81c028bcb7b516e6fd5c67c0dc948d65047d4024ed393151bd2142b58858cb10ec3a047e4a03ee283464a63e246880d35df9dc1af3f90b48c4fe0b57bd67fd8be085f1420a10998d5091502be37df4d131d2edd38f26bbd519d7aaa4b1b9f5dbbc91ca89c87d514f6b154fb52f2ad940299f1bb5079806ce2549a0c0296ed83a2de6632bcab997d26c4a1171bb150d101a9284a50a6f6250d6b1aef724b4185b390fb3abb54b3b32ec0522650d3aa3eb5e0beb6f6b450b63bef02adeb944257d1400c37b6fb24b839bcef7dc48ae830375bb088a210131f6dc9580bbd04c7701d951004463e5db3c5546c7c7282c29c0c633afc3230bea87716acbc8669c5b1e077f9d7e1b34429bbf3be8328bb1537e8ee66606d3660984ab9a01dbee29c4708afb4c9205f8f5f169fb339d11fe251c766033d90219be7cdd13e372bd2e9e4bd5134a44c09b08eb267347b17db44f92;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h3b8bc74fa0002b0075d2124d01667f965175a83fc565c95f0f622c61540020c52f12adbe2d7629003aa674b873ec9bf5ca990059a97cab0f34068eb566601549ecaedd835bbb52b495ec9ff2bd431735088b198e4ba92f053a010c625412bb8e623b3bc3dc4bce69527a38f842c897effad56158b170c9995211401ff3651be1384e03eef2d2ea476a30d4fbd6e839150e0eda93b28831914feb91f361750a21f089851eba96bd00490b638d4ea7c0f656a98902397adebfe6ca2698d515bdfe0aa8a71235091b5dae91eab3d3f4fb9ba75f801bce2f2e0d1d9c8cbc10420e7b005783e22fdc2900efc57ae8d2b5cf0c58ed56d8733951dbded4318192e4dd01c6506a8c76607d0074d9c673eb346d54e2b2d5d99a36162b13766fe3f0946790555c9ba1604ffb35639f3e407f40869d574c0a423673dc29fe3c49c3f2d9de1cf25b8a1ed4a8d1515b8a82d002a7cc2d1c30444b34a098701011eecc29182e3feaca8f7b8e430119efd58d8ed49d6621e4b371595e149004c9677cb984439d22d4b58e7fe0b74328faad846d2ef6af04286ed351e12c924ce757c69155a48ee7add2c86af237f461083702409dbada127b641f6d71d855433212b30824ce0843aff7cc1d0118804ce249b9cfb6e7985a1ba4ea885be233bf09875725f86c965a5262d63cc625c6e045f83731be9132426537fb1ae522d3252971462526d76b56b35b8de6612936cd8629977643b5d9737cd0c7141c02aa2c73315f430575096a818e5b955bf7d6b481a8e9dd4edc73fa68f84598b793684779b7328468d65045cf33c59ceaf62a3dcc896c37fa8898c4592d52647f106fe04a11444102a435c55654bbe5be354c5f1d898592ae67d4859c78cc1f697ba82aa001241704c96304dde9c096b2f730c3ef3fb6c9d18c6e47d86c9d3ab13d159cab0afa96749326cfac308269ceba0c681a0e05cedad07af074b24ef2872d8bd496be6bfedde8d85957d48f67c423ab85f29f6eb3eae02260f094230977a669a6ce;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h98bc99a7237b7c926c50017e58e1d1ee4932974be2853955876ca851f0da87c421ef3ee923b4e54ca3177f34d88e94a9d21decb8dddf3fbbd04bc9f2135bd2a32ec77204566dfb992bca5cb6fa5bedeb03ab4d80b47dfb3ca59dc8ab3598998822254c264d907238b0fa33c92bc7b99c911e487b10acfa3d3368b8a4d632d17f93cdf0e96bbcc6a8a5ca528755f5ad92e7e939c77b51316e86781e014e0c192a641524b638874ffdf2c3a0e7e5c047589c436d511c2778a3c85850c52345d44a15296555415bb04a73197e3763d194321e7e24cfa1402af2edb1b8d6a830d1f7835a35399c226e5580ca8cbebbbd9f00983ed79b9dd3c0c2400cfb55fa2a57b6cbf44378e5db570eac4fd21783be728b749c048c728c3230220a4c85f80f45882a58b76fbd328b695a35a6ecd9cd51644cd36d19ebc3f0cd64e156c0d0a855b8c7af6589ff1593beee5707bacf29d64daa5866cf10e19bc0a200661f1a8c2e310b880ac25f143c535f4b16881e436b85fc1844d18a6012ec97020799bc1ecc00eb900cc8351ea4f7a36255e9a60b6868d358ddf4a49367df675b3ddc0315cb058e01096aad7e140505b6ebe6e7e937a3b2a6580e496a89d30dcf71d282c8bfcc554c34b315ef9f664a11162fb491b59d29541fc6f13374873c34d703e03912dd9092555e42ba9cc823400646d6f5187d80cf0340cf6d96572c06e7755bf0686bef015b5955852b5f82af5f616698a10e7dbe40431f27ff9d4f1ef030eaf48621f7fb57d574bf69aab4d62538d77794f1416c4724999061075be7f29d126cfbb9c23f6eebb0c25cfbb70694f7cedcd5e5e35a2b290ff0f90bf27fa04c5f22b0845edd5a719636f74e6f67a0311af97b76849678640200637afb0b31d9dc0615dd6b267e4ae815eaf60fe5f138feed59f05bb475dd18db25ec88c4dff36f63cf7c65af0e976fdae9e13930ce54a5782070a48a604b597096f96f1e9abfd96b04d82898a96f12c66c4467c5f34fb241e650169220ebbbbd1f7554;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hc1b7274b72660f9b112c7b1455e06c3828e6805d26eccf16450576c8c3a3063373a187a2057ad9f46f093fe320200fc9cbdb0ab773a6e966b5696508b08dd2e459f36a99d3ee36597e41a5c5789d40a8c2b88e25cdef868ee64d6951e3b84d87acdd222206ca961741736dda8de2c1879b1aa68e2bd67148bd601cb7c2c10709b87e5d044887c7e11e2f78fcb244ea2233e2056bdb791d761768a001486a9a425bb0b56cf7602367b5ab6918a64933d3614fd0751689a96606dba734bc4ada76c9d49a937f6e1ad1bd56ede4f41cffe1fa90c51fb37e505a8e78303346d9312fd35999d86d840e0f1786575e0172d74d68ec12ab7d0ede44cb038c79d5b9d059bc1817176f21ec8c6b9816b8e5a1d94f55e5446f76e08eefa7c072b48a4887ba0e011a1dd427eb14d90f223e40aadc68b3c356533e868939f452b9561d0bffffa81c796a6e2476efe4fc39eb54e51a299d73af3d9c6a20e0a2438276dd34ceb957967d6dc3678e96cf3e578a39f72a22819b149959d97daa9c68b5882cc4856a3a3a4586e6c4b67d50cede3867fee45d6ea64c789bbec7807021c2843450aafefcbe3709aefb5e988c7b58573d3f3b5e623a97da0f89fce3fd3874e2407c3e9e845eaa33727f421edac3e97b9597ab4409a32d1d37cb03c615acde611430c3a8474d6ecf90f9deb3fe8116eb807b1f83685d67f921ce307ff8c1ea49382cf7cd4e5f00034ae78485c63af95440af5ad2683e7c586a0932907c5ab614c7ee9dd30b99c65e73f2d59ad1932d408013688dc3cda6f74606f1499f08470366a6e523f66889a1af2985589f5cd56324ea88e872cb34fc0930594df38a9ba5acd98f65cc520dac55a7ec0e85c6c8b68529bf8316ea639bb5c52868a0b725074adffb3d3dd11ba9682408ca11f7ad1560c7881d68d19009906ab48dbc07acd0b45b01b4889415d7bfbe921dc385edfa952e587ad4f3941479ee9681b37fef6896a520ccddd77a9d9fcf2c330324d90e7920657084a56875a28c22737f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h920618aef5f48a438b8817fac8adbb8094baa2f5f373642b0be4a9c5bfa8e471b9283272c06ad1fcc84936e68aac7fffe2d1e7407a439937f22d68e4e9a3dd46022ac0162de31529e3016d8329c1053900bea39f1cec113df170f82c0c70fb03983f0acdbc91a733e04bd7b6a3406cfd226787d01562bbb8f37142582647e47ebd8e1305c8734240f01a67d74ca47fac16a62b349cab40fadd9407a5570bf120f83515b0c37e46bd50fadf19b88376890946b1cbdaad156dca230a25c5dffaafbe72e29d8f930f7caa4a6a8d95ebcc778ca8d620b37e20f00691263691fcdbd285a755d1c5758013cbe291836782c92c3cbb9d93a619ea9bca3c61fb636771060e005dd2db783580dddb7af00e005e60fd6a8a558d0ea2eedc58b617b756bf59dc4e90b0e43c2c273506f740552d8e45f250c3ace0f5d0ca04f113e4e15b805e26ffc1f971d4fc3cefbffb1372b93c4d8d51317c076dc570a1820b2607c50acc062cf4bc89632adb758fadf8c3192d33878d8a7b059adf1718df3924d3b4d3da6539b116c170c24a45fc4d5ac4aa5e02fde33be2bc92170f4fd8007fc47d938a4a81b9b5041a635e8af2e5b0ea11cede15f9912f79b41e9c576adf10bf0d90e3839decd906a67826c08d6c4503467f32d579302fd1f5d355765e8fc2d1acfff7ef2c914f64bc1b78ae23d1eba36c3599029cb5692cff104c68684ec77467eff747558f48158c3859e2db5180b48f5116a281b31cbf193f6b077589a278be727c7d812f9ef1db1d7aced640feb98976b8dc0212028bb32da44402bb5b5831af45317af502ef68003a4493c52c3d960bc9d337b9113773e6f85b20ae0147839b982f1bb3235f5cda02b7abf9fc9dcbca35b4da3be663b99391591e0147ab72ae11074085eff9dbc2c6d9a508873c661c1c843063da186a87b5c8c8b73064536698ef0c9f26d318b58ed4eb1cad10896f247aaf51e27a7ba50a891f93f7c8a026732a8d263d974f6a47af42e3dbffae719f8a26c7819e23594397;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hb915c0765c913e0a822b6134b59949f87a0e015cf7f365cafc3e8e220afa637e662e827e6eef72c2b502aa5a74f6dfc81777f985ef553a4574c833a49c81d006bbf3f6399c6df954d8c07f3728996f92515baed9546ac6cd07f4523a96c4f8591d6cc7485a7f47e29169b50bd57285babd8726eb5ca1e0a0bf7d34e2543da6b38f225f10e1a79283681241d6590e6bde849d0df9230073172c335743a0253e749e4196caa3a6488e38cb3ad6cdf2b34086c6f746b707949dcbc7b25b1cbc2260e797faff75283233440c0b676eeb1e497f4dfadf31b47d7243e3d7b59de8a970bffca6d311cc5015a0e8764c6ca5c3925158a55b83fe1eb5e07f91002b04ba0f340a8d7e3064534b3287c6a6c0960009631322c21a8b0291a983d97fc36b030065748265ef171d0811927882594732fc390a3754d270f41e24dab0bfed8d6e3fea584d1ab2239530f4f924fe91124e4d6f4038bad02409317dfc684ff081bb7308b7e04d57602f59d474822ff9ff28e35d3ad4dc671deda534ee61356b166e65fea653fdb44e15eec34921e5342cf43088b2984e8c6dd995ffd48218b2f24f7a69ce253b1c3bed8e29ddf5f81eb8aa9a3bdc9de09a4fe5134a2a29ff424df962abc8a327bfadec1f776fb31a9a40b73b9742f84edcfa2ee40c8809e497948e8dd0901e3f8ef24e2876acba64c4c1993bf7faf02d13184b8bc076657f47e7eb9d15ba88150097aa79ebcfcb84917030bd35185c24f19c8595013a266bd0c289ab4c242515b72518ce5a97678a85d7c6bc61dccb1e10e858a7e2434510b6a652923f316284db5bd3021b2210072440770e9b2fb2429d41867846bd2bb3cbe73900b7e469c7b5bac9b6e48ac829bfbdc30410a0b7e52525e8fd4e49dca0d5b53bcc9a18d8e05275bdeda9bb02adce6096166d6464134d20272b454479c4f0e80817b0de32111f2b22d43e83582db3d66c345d4b0d29f1f509bd6f670ea881f9d249994f72b0c3da7ef5aaef99140aa229f5ecbefb5a083d793ce;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'he9483d515a6a2ee68734f65f91ff11555bdf6f471086a5423d0eedebfd5286bb700bfd3c022ee2fb59b4f6f0cf9e9b81ebeaffd96d4edcc8ba50932260057e55e9e38db6c3368e8157888fe557a37ad65e384bad015900c31cb0c2b07c2c1476c523b3a10822e1834fee00f8011b4b8adc2cc47d4bd552759982f1d13f72a2123776cbdd0b97319bf5b54e35f950fc9889addbe4edec5587f05b7e9e876ce25006ec954f6054477024b1730a71a1bb260e8a6259f0b84f14b3fd990cfa6f40d780e7aa9eb0fc8374b2b393bb85770b39033618a80942d05535f826a35da97e589ea17cbf4fb4ebf7f9d12c373deb8753855ffdcc653e333da41519fada79f351dd96369e21cf1431f5b0d6a3192c3f5253c7067bd329e23bf54f1b27f42952e1c759ed1884d3256c2a2035ef0811cb35bd83c1618088c9bfae35ff0371f1c21020141aeeefd8481a0790d11dece04cb85be5b3dfc11f67786385789c6625005bf7ec819a9a38500ad0c52945dfcc55bcc5ef52c0f279bb2a241469d317a2c43c0f192a674572ad7e5f5466b4a1e864d92b5835322a04c47eed4f2e750716cc2d65ddb447fb7947031211e7ee1263077f9f82a6be5883d40bb26a71feb0a6925db9559abdea518418c4f4810f7b70ed7da6f83d5c3476a25001ec79778b6aefbf90bb8882fa4c51f9a74683aa45136ed9a35d7681eec887075f8c3b4a0f39a66cbbbaae06b5826a3b675e649325397f18aaa2e4dc17d5589ad7363bda3f2116bfa819d95b9990dcf6edafc7178427709f0c2a906b7f392a61b6f9349cf7677650aa346403d73b68fb19a5789d13375383644a81ec31c7841d38187b7db0806192df6d206f212caeb5e6a6ecbe2cb051e5db20c61d11393320ecf3f24c580d6374d15d0c11d74faca4e6e9b7ba3779a80bcceb26bd974a2c945ffcf5ddb83248da9bac4d964eaa2aae413d6acc8b94670f8eefb2f473391d63a8d643d1664e5a9c31d5774fcb032c3b801b88126ec810a917df2b6b6e0d38cda4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hae708aacb6ee44930206fc0647e6c5c874985e9cae138e156a82e9b0645d256d4925416a7d4fc36970738e8a153285ea68f3270731827d2043b083683c0530dc427258d474038a97772167376fcd7b3e4a97b15b1c9682e96a367b2fee988df2a0fae5c3194d72e1f6e9001062f602817bdff4ed59e14fc3c22106f01d3d4795dfc08150b256a792e152b5cff209b00d8a832f95e4e86cfaaf2800f9e7ee27e15573bd80940db26d90e60eb959cdefe5bcf4b5e978ef2f1a52c6658b5e2bcaa38f157aa58dc93c5ff5f35bd63be3af27ebeeb1d865656aa98d9a6f62bb83cd4b23b18994ecf20476615a5d2f99c92dfe2d1c2a213a50e3b03fd784b7a0535ea67edc057187b63b803f6fafcdb38899784e6efac99f787e8866c8fcdfd82f051ca48de31a8bc121f8bec562786fbf33f1a866ed843b37a7e9df5a08ecd75749b8d8154ef139783aef25681714d8da216ddee145c2da654521c582dfeadb2eea5338b2c5f9e41dc8b1f4dd199767df99483b710e52beaed3df4cc39bc2b558a79a018b4e9d592cece50a9aa8d2a73c1f4d8e784fe508177bc66bd8970a92c94bd30e2e47ced1eff23c2cee8e9000021dfc1b50361ec66b4868758ac689fb28fcd0e9f2cfecf37c5b0e415893535f0155f93e6e4400c0dfe67a826f08ec4f74f9112ce2d29983ae030d0766e93515a4812834558332f3b640e17c4a6b3b57b2251118b1906cec9485a4c3f1ab9c7b57f5984c26f4eb93b715865827f47af4dc64a2aab3995498d0e201633262909ccce33bcc67d1a933565c5852b2f828be10acfb7af852c077674b4b1dcfb1c546d90457e44bf08bda4ac1b16e61fcea346b64666842d31dc19874e2f205557b47cbfd9174966208830a5ec64c6d3819b5c517db1b2215a69164d6e29b2441a6d7b95b7334b66a5d68322fa6ff7a01394cd1ffe442f848eb24064e3cb9c69dbf56503eefec9dce3d1b5a9e5cf75d8928fbd0ae4c60e4a34b98a9591488f7fdbd463216342c53780d5d696b51a0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h230e5701f2ba088943a97743c398a09b83b42bddcaf929fa05c22320d4f7b7660d6f38d1454428c20331030e1ae1f6b510fe3ba9469d4d235852b7502b67bf1c9985ee076a06fc651287c77c9782b472d0e553727ac5fe8e414b54ead2f8bd638db74e87453fe4df16a73f2a14b317ad62bf3049a7a14139e83bc7da7bdc40cbf50f112b99bad33ffa635deafbc22f33082a03fc7d393008d2512bcb261cdc36ceb74444905fe2a4badff39f89fcf8a65acd7c817ec71332b27a0ac9debc839927ec92f22fe5580377c337b4d566ad27e6f0efe17c44d3c5aaf35af14b815e2c5dd997dd34ef3f98cad45faa7deca0f5e68a8680296789d7243c0cdb1067eb52d00c9e93a369ad4a84fa5e43a2ae4b941b12144f8b4300ad26279d22a51a42d5adb61f520d0504f5f06863f3d8408ca470cbba6a2364bd974a5f212c82ef697fecdcafb031e63d6f066a8feca6f3e3ffbc2bbb072b06dff502e54727b9f5347f8d5f69f73b8f36f5726e1af8c752767167ffc215c9d8dd5a3809090ad63dadd10b420a2f4e557090968c39ade2c01eec009d0e20a7de486193659ac10e21eaab4ac4852113220249b4459a315a32873904b2b54b9587ae8fec135fa9f762545cb6e2fefd137690efaaf4f81a2a582a1ab3b6eeb4cdc15c697b6d5a1a5f462371bac9d4afe474315eafdeeae93bff2170740fd243ae91cb0fd3fd26056e11b22fba71a8cf1b792043fadcf8002e529ff257918d9ad02bdda8dd220d067f9dff1ebd75d6c25b8a3a28662ecfda35c8ad80497ad078449a4ca1ba6969cc2b43dae8f3b1ae102fc4e8343fdf37d736afe2975bf10b9105a23be093d9955f25193cc9d9fd24a8cb1e1e9df14489ec133bf1719d4306c24a136054628938eef584e6cdf8035e4bc53d0fcd74c49edb258ada9f46e8ea607ed805dab6b049ffebfeb241483e17b87f4c13e97a17d61fc3a6f17a40db06d1ced7007f3e94ed4ca5ce72c7cef0629e539306a430863bd9b7d2393e1ea25655dca182cdc0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h5cbb80bc2886aa65e725e8fa7dfd60f99ebb775773041c0c364eb6f351976148ebbd2fda626bd8c1dd1c4a009e4ce91c521863cdf4d8a3562e581c2d793613f1399be3141d12a7a985dd3475141c09934c4b1296264f6ec8879c94e235d8e5efd6474b7e5de7e2cb49d45c293e7310e6fd3bf284824faed07cac1fa1802995dbfad62fbf3309e133610b478932c1b9affab8535458cdc4cb60f1702403a26a1b584294c64536d8f2fb1904a23b5952a93a2924f31fcdf529555858203ce79f7b81c3229362834f3408be253394a5a210fb16095c056dc4f0809c849d64c887e9de5b30e3bf12974dbeef2f333dec411a538119cfbdfb286f1c92cfcb02edf063e05baa1b02c151ae1289b18f039451a69966c55b74a62e2d9e66efa41d5b9146f1fa1cb8e922be5985c6723badece28847248e7e54bca7faeae0a7248d98e8c102ce8c046061bfa19a94b57924e4e452e6e7590bd8940489c3625490ac957ff53cf24e3261ec896b4b99427763fc7a7bfa075fa96d7d5deca39287c1077e47eee98424484fbf4068ea17f9da9b7b8c90fdb25d14be160e0245c3d2410bd19167c2e27046e3a8e2b86b8d779e031a70a18ae077c4ed02ab4fe1eed91a473879fea3bc25684650c93acb63a6615715dacef30432371527d50f5b8987cbac6f03631d61c92a0d80c196b2808d63cc917210b95856cb56bd16c9634de04398530e12c732ae282cd0997c7224268c342329beeaec0a5c2393776e278d9a21ae6ec5bb000fa5a35cf8908dcdb9944cb41b2d4b116e4d3143ebb07b6b55e9295e826a3207befd7833d37168e2fd895f9dee52e74794b7f1df6712a09384efcf3fc7f97d794e51787d905ad54090ffa8a42d643492ef500d298a1cf304b07d0e59d32739edb12c663fb0e62a991e8f66677712c557fdea32a8dbdf44118e948f3c838ff4d10a0ee15dcbca01c0abf5449f25163fbf3368a0e6fe045471393d2159827a69ab720aac0d4b55797c372aceb64ba76e5a706437998b606e32;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h373a19cea9f65923e8602c97bcba4336d825be314c33bc1c95fd4e03cd513049222a2f066d5e4eba8dc7085fb54fd2b36c9f569d21e8fec2977f94adbc3cae8703204ddacd464cae64d8b9ddc1d3c30b8d1b3555b4f1336e2e3fd7181f81b8453a5ac76257d808885f7c30fdea78d55a65c1a410629ee2cb8cb98a711f3626b673a3b6cf628d30a3f6ed9e1c21bf343aa08847021f858350f161e46e2ca2cfc339a02d5c878b4d18f976af1cf292b24b67d0f18210b9f60c97531dfbd4f149c454cccd10b1df8c4344dfd139822ad83af9a90cf21f7eea13f0a327c0e1e622e3e09781c05ed068785ce907faf75b8afaf46ba5e6f8a22994f84156c8ab73b67c27f75feafa887434b8d464918c1f022d820a3894a14d7137281c6ea6a4681d74e5a4f4442dd6928fddc225f1b3c85b8ebb251e1c2a1e644cad183245e062b234069285d9704a28cf299948bbabb6fd2bb5c000511bcefbf69c0076322fe34b48358538b079204728540dba974b75a41bb0ba6582e879ae088b6fa467daf4bdab48905d97c4cb918bc5b807102e48e23b52d95cc3f1b3ca75bd84350348697c2b2221b349992158031c06bb198bb94bc1c775dbbfb854cca3afa5d40c7191c2301c29293f5c8ecbcbfca92f06d805ee71b9f3ed62f21adbc466efa3cdf5450cc94afd60b897875c13de94ad5ce36856cf3eb4eab8398f4b9fdfb93b8dd05ebbfb423c40e2bd9866669db02ac8de767ddc108fffabd8f9c849f66dc8b65168e6da86439acaf49e02deae19ea9b2e70ab4427f9991d1964774b74e55ff3ff3a77526c56ebd98a582210ca261b97339196b2b3bf0d651d1d7d917aef67e8d918baf1f11df472c96592534abd570fd3dd533b1f3c808d861f9741f9cb20469fec2579e7b92b5b70f69fb29d2f411df00a794e9fb48fd9170e319e4d51a18bda2a3717c631bd991f4b5b3c5cd1123338a5da384e5ec6cbbda6061e697b1e30e4536ce804326b6b0f37bea4fe72b9081f0d87c5e99854dd86afe950c5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h191d7bbd185f6706bba2aea9735c90a018a8f579480ccdabaa2f8d0abceb34fcff584f5042f44546571ea94626d31d73f4c6e014dad6d151fb082f956383cdf35f478646853154f1bfcad987a9a26d0dfecef57020b1897d85bb260f409fa5e47a043d435736d374456c2d341b564695eacda7519b99d993f339cf05409ebdff02706b4a0ad6a1242d5c4dfad458f1e8743c75ce1ea47925222e0cdffd335d4bc14eb971b08f3527373eb722184c03fe1c00bc606d36f6defea6371e1103d8dd9de3fbe9119e69b1792727adbfdce044cfd1de460346d89f210a22e73d001e5824050e41e7433c030eab5e90ebdeae332127be4327e6674ece3da252092fe065a7b6442bd804256486ceb8f520e8509124a861719be2ca54c98399c1811f43a82951fdc97292e85e186c83dbb160f8355112924b7c788ed38bf731aad2ae42c62f8f484e687bdf2c3c97f5f00d8151cb0f6dfbc80455f75e34fab86ed68076feb9b821788ae39aed20fe5d9dd0656d1c886f87427b29bdc68b2450474bc8f7990081ea998daea44e01bdd323094b837cc53bf2d32974dbd960081c29f1a513a08703601c356e2773f0016a9f0f14128c0d8f3320c0023b4cb0b2195df08af36e628e191be4beb43a5df8301ea830a7c5996e001c949d644d38433a454b0f467096cf9b56e6b38cfdcbee003da5d6e065ebfa34d1600896b62cd09ee3e37ea6eccae9e04d4e8d33593d0e352823d562da132f0497f683e0e64ad25fb22e57469488bd8255b052951643d9806077c042e1f506ceb2c21cad61c0c7afd56f0ad7a7a72077b2ada7f4b945c563e1373457ed552f83cf9f11ddec394e0a68b513b0f0a570bce2b025ee47400b5e0feb69b60e6fa8522d50386709eaa21f5c1e8530d97ba093f706ab37056dc74c7d3f96be3d2b2d0bd0699d5b1680465095892ccc92c3d89a3a73e5c71878db48050a10475806d17068e138f1578ec0f7fbf3eae4b5c0d4351153b5203e760eda1a3f431606534817702c87c07a1e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hcbd5daf92998582243e0b6a90e6cf5aecc7ed443e535c2a546b0ecf7ac203188a335746d95b171f407aff94f4f390c29382066886d1af76186b32066e6df14922d5d4deb80469171dfce3151dcb210a4e29bd03264cb9570d01b4d983d60a207c839b9e33a30712c529476d72950f233eb6c69b33c124b1bce10ef39100e1e7bcdd254de1fd9bc494d8a0d557aca31a17d5e34fcfc5420e1bced2431b244cf1fcfdf15a37fc6e8721238d30441d1973fa96cc246b5d436ac8f533371e5fad3022340f385423d7ec1ee4add76a96d769a6f5e35cf7c85728b82dde8049116116ae359f5598b872b91d2218f1b0fe5d6ea747261eb6df41eeda88dc600e4197f6f08786106be2aedcbc3d71f7d873448d0b893ab04957d39b88614f3cf80fad111ac921534c2b2eded7811d3c11e12c195a5250f108a1804f906dfd7660a4865bb94a96e7475807af7bbe21052da63f84d93a6a2843c8bd7153a6f7cc66cb3549dcad233fee23f419a6b51ad65c895cbefc2660cc00aac5cd7942c7acbb1958a960bc3c2dd3f415be768af77a05f13fb1751952aa02b1d1dfc505a7ce533433ec04746f353dba909d4013e764da39294d5fab0a1eb8c8432f3c12c6236e09741efb0590c4a0dde18495f3e09ec5f834e0425d894a58cfa2e1b6dde3c6da78140184afb66256dfee9144b34f0567183abe21dbc2320fa258f340a4fd1e7391afe67335a97439142a7b7cad1998c77247327e1926a7579c68f700464c3859b80281ad28e42995308e22e9f264f1670f0f6cc1d205678b255fab16251f8e1319976ca587a62419e3541e86e184f27747d97621b3f126b44aa0306c0d81ff685fd8a6bc8c4487f56d627a1142f623dc2947629017ba0671b96bf0ad1d1a6844cb018279016c24c9431bf731aaec6dc4fb804817f0e023298019b74f9c8b2a8dff6dc3286332505de19c9d2be960718f17c5ce9f828ab57ed23937f6954b9151c3b25a8a44418ac4f7e3cb5caf3740b5b47187061b7a129ab484edb3f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h5062495b3e68d253da505efb2f54cf8e9cacd84677b5ba0b12c1054928da29e215a880f81a3654e4b3786d38d61d4718fbf60bf08b9bcbdf4de0d8b22cda4a2412425711125598df8656d0bc02aebd90928240a0fba72a045239050c9046478f3d6556e20f3111858d9f94e66ace22403853eaf6491e8deb4c0f51cbce2b57599f11b2dd4eebd93b9ae48987afa80c38669f564c587660bbee21cb46f446166f3e4f5f2ef8fe39a707d69037a090d973f0add68724de4cc20459bcc03cdc48369b30fa63564f07dbd447415e664fe782579bf16b9f83f55a09f3500685e748d7b6c423a1810dd9260b3979565eb3e3dceb9e03d877dbccac7473a9bff839b85c07a81c5529c113ea7949467cd6cee85b471b5be5eb168255822e1339f0c486891b0fc554fab276b4d7851baaf179c90a37948c996a935564ab8816e042dedf0a900884ba63231faae4a13c9e8095bf1d1333ac71900ad70ea23bfdab4c94fc606f56a2a0793db1e132d38dfaec99450143129a08f11eb56403202a5512b2cabf851baa9de80bfce1ab5bae56a62344eb33585df466f8ae34da2bed6a2937394b444559840e190ea9e0800519783101c2a8e049051bb748f7ffd8546a74668bc040901c800a4f71603ded7e1a39c720a12e99834693a12366f8e1e06fd35f4f463cca8cc14a90f0d6980d6553d4934de704f91a47dccbd4ab62a5c55f48740f5bdf4d62c0bb997192f92ba19d2a371ae843f8762c6548c7ed5c4a24f31bf6f5e31320d2124d49334cf4dddbdfc8cb3cc11e5d29e3a35a16cb760893925112509ec616cf6e3392a864544136b164e154b0b5db79c6e7c82ad957d23d5b22d83325647c860f579733f1461146245ccff43dbfe3591a178c951b237d0b6a60a2b9dc42b70e51e6f19af7bfa3325d7001fdc06b5aa215e2c418217b48232dda411ad78d9b407e771d41efdc59194702e3722302970511f6f139c756ff79bec36361bc94e66e6b0f6addf2340ad84551e8dc7378228548dcd46b2229;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hd56c6a5fa8d835accce77c3f214f73e371a8fe2ddffa4933a3d546b1ec1c15cd950c67cc8046a2364bf4de664670696ca0c44750d123fab7ea3e8f47af15c0a9e08b3bc86caeb85193bef3d0c44c610d3671518442e2e507296b56cf7fe139ca8f0df9b498f939b4686a9f9c6fffca770fabf1877693269acaa8c088014b6ec3100ab2ec8933c55051a9eb9c86f02972ce52247be72ca2769f5e084c5765ed99e3f8a52918cc82479f04ed28a6bcc4845ccb9477a8caa0851815532066d41fe6d7c2684878cb56690b14c2bfe96254c4f41402212737669b53e203132fbcf9eb63738991da4f769587a6f35083d391913c34e1251317a983366569484f6e90fcb721fbfed8670379ae7e860caa97e9e285c1350e8bab06040713f0778e425e4fbd0c4b61bc5d206f77c56f88f132dcb2b7a05e9226ce9f4f7426267d314f7d7c25cb4551a9c5d16d99f89ee974fd634e2dd1a6f3e65f7be0017cc5eaceab691b4a0271ff177ceb32a5907355141e3c3776cdb4ada41b2aaa1451d488e9fa60180dd5dfdcdb2d61a10836ebc1cd575a645a036bcf1c4ddff7a30cf7ae659c2064e9226053a8c19528aae87d2d73cb943470028f13a8a11b1dab9d2146e48cb6aa558d658311035524d826e3cc8fba046d2880efa28e27a0084a14584fc195c5b74e8a03a837277cfd1cb78d647d0eb8dd2b0fbec6e3adb16a77942889419ff38631b2d512d9a67ca9b466fba98ca189ecf512c993a6333baf05c59690f1b503feba60aca90ebc6145be1b267ec978db3797a425e32e26dc83c65474a44e0567053c4e033b4fd84c6f3fe88f4c5c960cf15e5a00aa06ef962f2a428bb5fb8cbfd66c2a8ffc4333064ce6da3bcb9bf00e5dfdfbfc79ed7594b360eef1ce0120d223afc8b82669a335b5f44ee62227eaf0cecc4d1da5301d545905d0b511c1e45fb5e9abc3a2f3fcdf528a0ac48e0be34f6a0afbede0c515dc40e889493999036e7e74580144c00fad4957329700552f88b4112ba526551b777e5e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h3ff7992e55aaf3f57f1b9e57744558cd09351c92a6af8bed43181288c3ff9053172718d5ff17ac3fc57f4d1f57a3f5232cc1cd846206cd6c50b1f672167f3bf8403636694d60faeb3c32b9d49f795b69cb4bd483c9dbac1dfcf5269a0cee25f59adc3dc3e65dd4f343384cdc1722a74f59b4c4a07f7c7ba059bca18919a51d7bf988952a8c73197887ad4907f4c0246c926ff7cb1987c1a8bf07feb03886e9dddc9b1794c3de6e2b842de0aa51340509c869aac67e6f5f45c0f3d7144801023e8137f5f58fd4ab74db82810b98d5398bcf9be73bc76dde1ae15aeae7feab57f2adefbd95e29ebf7addfb1ad9f58f80808062eaa457066231cad0c0535af30dd0e3bd9413696a2ed7d5ba51b5cf2939c0b924541bd9e66e5523bbc83a9099fe399474e2046781cf950873896b92ca2fa64ac6f0d21993de3239c9c99e947494b499f6f3a12357b93ee0be2686b76200eaecaf75194bc9f4d43d81aba586b1d252e5ac0a1e03c3f702d3249946329d1948d41b155c8574c428a72af59b9c3be1df0576b8b5c6438a0df42f171bb36451b10bb16d97ff3289f8ded09e857dd8ff17f25f3178964fa4583251c917a100e735f1bd0b3f31730b94332e267ea2f79f6785f250ff917e65223533a1f76b355ae23922f1f374e409c1a63bb702606e70b8839cd3a35f94f3fda825879d92805ded64c65690d6c68a48556902cb8a1fe7b932c5845f81cb8c0f896262719f40c0fbb7842e40d498f045ade882773d40138ef09c8f8b0ed6c1e5e3bd7ad64b099481b489c464fe59ad43f8f7fccd959b1db24ead965ebe6b5bb2636d9f53a594036b3080c922c0acc3bfaea1b4522784184475e7c3b49fd1be082a77d783069e1db739ebddcbd7bee1d2441350d07e3593af1a92ebebf3f1543cb463e0b256df78370e45028519407e6e3889102f03d38dd6627dfc27b7c79d499643cd009f9d844f1c3302491211b4142c3812631c51a7d08550bb485c470255e8aee99b0a20fce3a92580218243c23ffb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hb485736b736ec4c52171b0c61ea74716d0713a0013948bab3b2221d08a561187e9b322c39d772b1439201dc539e3e9b63a5ca7f3a42e61419fc20e455252051dad13e77f38a215ebcc40034b6e5a50d38e411103773fdb73890e2ae2f0791cdb363718db0adadb79717d2792e4ce173b54e4e9011e9c87a585000bd2fb1b4cec5b7ae34641f8ab6152de74be410fafb7f122d5e7a78bf60632562c8cff422eccedbbdd06075d03607be8a8274c216aafa65bf0d51bb4731428599bdf0493bd73cdad7daad62f92557cdd9b8720d6bc5384476d5e68e673b2ba54745e45abe2a3d0d00c72a0adc173bf10825e609cc28058542c0918002457bf871bd240ae6dddb235ecc0c86ef3b7f90dae64ac966158795b7f1c927d8ed5fe39cf4454a08ecb81882385ece0f16d4e9b3b5281fbc9f55f2f64c42250681423678446d3e679acb2758cf4dc0c4d2e8489815fdbb254bc5c5939c512edc3b00898f020cf011e8a05b0f153e57e9027aa69e9621c249b8f6022f3be51ac658c84850a30bb920415a1e7d39ae31e4123e1e51cb4940ec7fbaea81fe4ece7578e18551808d87033d0426bb41cb72fef3b59cb4542a90dccc1236215218f2bbc50e2a32ff6f5b0a37743a7dbccb71cb49332e748bb6e0548f9eed9fab6beb9fc8f33db92f051c7ce609f1d9067d927aca7f272c12b08f150752d93a6753dcb757524dc7893904f82cc50070d51001bd476d600d93869d44ebc6af4b39269ecc430579017c1e39253be11b126882afeadff7ae58aa414d5ba94d563b0f098b72c8aabd5a6a5486bd6b95bd06120d36804543132e2dea41a5e8b5519245c37854daa482ddccef4ed1739ba7b7ee4649a938c3f95ac4fbd4e54679894092eed1a900f30d1a3e9e998a899b5327901c4b61f85ddccba21f7e795808a9a6218fb0d583553dd9436e634c08a2c34e8a24604f9887d0e650510e6f3d39c7368684ae21c06416cf89a80c3694b06f1a0a97f44dec95413f54cf09dfb5ca0e33a92def11ca456;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h22562831d508e4e12dfa6d1a2296ab486f765da6a4accf4c75a62552402db46c080f0e80268642ca804ab3e53fb0b7136cd7d71de9ac9648e2d088c1ebdb6fd46dcde818aaa3ceac0cee14a06afd72b63e95a6480af689f1100847fcab6efcf81c8331bf3a2f46e5ca35fd26c36cf71fa10280ab6914b844b33c624d33cdf25cb5957beac532a3e6750f4a3d503eed97e660c07693d7c7789e94805859dac284e6512caf5fad127b02c11d6e19f8196116021e2d1136dd01f63c788d8dc5faab3b6bfc7aabbcbac783d3d1056cee21beda86054fba9670ce4845fc93dcf2dc57d4ce727d7d3a648d5773fa644ffce853b5e97a7fcad071f6c408b98d00eec8250ba990dfed14724ab9492b3bba7f01aaa2a0c2788d013a5e55d577d9ccbb620f7e21df1c565cf4c820918a5f2e5472abbfa087b0702d7b3e77c54c6cd55914705e22838acd2eb97cc1b839ef59186a8f1d5be504ef40f8aca21d997d94595b525631870aba4b4c2ddd01bd4eac8230799398f5f53d587b27cf64d97d6d627a395da2c084bb28e9a424dc5c2416d68b7b250c69b01470c15c3fb9fe9b93ae4f8c45c24c9eb597e36be16866f36bcabb925d949aefd7fa429ad2192b64f5f39f7615d4b61a9d27577bb16506fb51c81917ce3a7dc28dc7b23a3a1d0b5eaacfeb0e24bf3a8570dadbc053b3ce37fa4683e6f30b810a9d0cae57b9013e16985b3c5f53411be2414bd3e5b9cf2b9cf54202690981245c7e6073620c549d44f088bb7fdd066092b67621e6953695832a0805f7ee44883e1918c7b6bbaf6ff2e9e81dc3ba5ac5af4621e17bd50e519e24325db6276dfd9cd5da781567832c866eca3e93d7c51d28d0c6381893b7b2d47aecfcfa08de916e163681652d89f87326a2b15c8f0bae2bf0941c75bb46f1c651ac0082b9ed3ab552364673ae2093bbc77a408ffcd402b12d974a276b4e1a3e41f4e181c72e6889fa38ec0116c96be5323904eec4d137e5b25ec70256b99db89f15ebe2a1b16083c32c796835;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h40a34907119a95dd7e8673312882e05c8a5a6c2ad9c5d9430822565fa48a4124db23babf7d3bde43740bd1fd8f3c1b72d181d5dbf7eadf0f021ad09155c84fc822130b48ca4e61e73c3e91c2ef2ad61396fa69d750f75c8657fa286cd5c26aff4d282989f1754ff831a96acbd2ed1bbfb486ac4899b18e5e4ce167759279f17ce66f4f0424727a65aa8159db43bb5bdf1acf14540979bc90d0246f4c8e41cba06385c29a378c7f65857e35041f2943e43997b9319d5a25941544d5749305e35fc4c6733d754e65d97a50abfccc62004b22d74aca80e37da33ce251754d99d8d2b7610bf391e355b843b801c9b58ae782102d7ac7798002079d10cbd6fdc4b3d7365e3e57787827cab2fd4081146aece257f009a3b4231b49ae1b31f15978a7bb395f275e27d8f16155459a2800d27a03510247a46b3492499caa0b186d0c6165801b0a98ca930e18f27f9a00365056d2d687406d853b3ddcddb0441b6c41e7512663f7f528e32393a351d351c38d45202d8de1b67da2cb194444c831136e11ebe780a7e3b25daf1ed4ab84887747dae62ef3166a2cb841a96b4887a30a17991a93e1c2d264c15b63072b6cf4e8f5b360ec2548850990ee60591950f1c2c79d8f08cdd5272892a0501aadbce3cde4c4b08b87f40ad3b6260dfcfb290dd49f3ddc52ee4b0f8d9ca31053874933d5e666a93ec1cc93f766e8496c00da8f789b628113e7ad5ed5b4ea9788ea85191cb91000b04b3e24b6c1da63649d250d32635608b70888e80f7877d22f2eb6ace9885a5c42b09faadc4fb43c325464bd907a52d9cf704201c85b3b66971dd784af8318dfb72cc38ba2773d20619e6821356fd102ac43f333dbfbfd6c99fa70d0a7a3cb374ba10bc8d98f8db4deb10e0e56c00a5676d26b82341e2f626a0ebab944433b37c4ce8ec8c1c24b9bc7011e61dd17c5713967854d73fd8930f22e0fe34f44f55423807cc1312a4fd9b9d07c083d148c73aeaa2297ce37929f1020177b46eefeb37e1e3f891499b466;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hf7db54df2fd0a59a7d3fa0e4f0ac25c0cb7bcdeaaf4bcc3ca6115e5d69e623d9d076fe7894e956eaa3af43c93383d672fd8de2cfa3a519d86eebfec0743e1e0da9e78ae29da12ce68f3777f6303b64c1b8c97f5523d87a5f5a3fe1d78d4b5e555767a7c2d680301acb095132dff6cdd3b965ac5b2d3dadd5122ed3936018ddccd148233099de791f7bf87d1b616dd96d163aec13f32e00e249473235b3c2e0d178e236211fa10fb0c63bdd0de07c0137ae0b3792ba5b029b9420a4ceb2d96530d67bd103fd979b7c221aa5572ab47712d886edcc7f36128dd55a551f96f3edeb1d025761e503b6a7dff0aa07b9863ee623c6bc89bfee6bb5cbe2dfea311eb77ad8c99887989889d63bc761cb1cbc7989905d317541b3a0becb4362e57cd3673d41add444d9cadcc37f95a1d6ad1dd07b8b0dcfab8fa3fa343677ee31b47cf64829f070ffd45e4dd94520f8c0cf42ec0dd6e23beae05d3807f2a9905f6af8cf3cf909ba0d74a4787bba42e1de2a28de6ae5a8a2cf03d8aa91e1477da6066a191b90fb35e786e484471e51cc6213710f44671e595b1425571d82312f040abd999de1054abf1d20f200a7a73addc94bdfa6e6ec5b1f5b1c90052da2272acca1bb09dd01cf74862b5f6e2125ef625344162b03cf83f5eeaa36f7811efbbabeb09fd6b476e6a65fe490cf241f47052ddd682b7eff938dfa1d1dce7b3f2f05a3d3c836e4b27d7e482641e00d6c3541a937d25851d756bfb59f5f9a3f66cbfaf8e41ceb33b76ef49609def043b659b7d390cb09f6ab6323f5624069f3aa412a2c4bed6ffec43e29af1784856577c53d54e9297064844036cd61385981ec32c18a8b028a220119b98144961db5c02c233c7cf1331d3d59e6d0c73040cef229d4be59771685f73c9710904a601b8cdd06d08c98270c5a9b3ea7b832d20dffd1248658a238c2a41dad4b46882cc6b25708ef11b5c3b707a7a50e1fd4a2eddfe23d3b722fff9a188da869dde66ef6cf3d2ad9bd18f2d104fefa649099073c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hd8c09e857caadc83a779142db38c3c11e4814cb225a3da34c71250bafcaacb437aeb22feee9c4e64c120426d55622c608031317ba39fee81c8c6ff391afea5e833aacad554f770f81603ba14d496028a6edadd25a43e6f3d745a87007822b985155c9ca6d316978bdfead3fe853cf0e12fa72f7fe5cfc297ab70422499bc3cd8802dacc4c9d4f1a337139517d4350fc2e2277c0c1194827a582ec5ba43955dda7d15e1e627bfbb7f068d27fa15c99a53ed99096c0440f82df7cd21d0d6794ba342d6c2b7a5241f62245c7eba14a86ad143d24b8ed25756c5d378fa0fe81d8bd2850d294646ef0a085383fce4b7849f1713f99e485312866b0b6c28e894c44caeeb15ef49a915e26de9277357a0bf1e0f41fcc7c02a5369a15c54c0a6affa21df200be391b0b8f749c8c102aabed8775eb6fbf41d76f17e3c7d3e6954fa38b51a6f8b9fbca3a9c51e1a9fa756e7136fbf1d6146bba39f1b11f4b57c92f8a3c71ae61a533ff23699b29c9e0acb8a5a8cf4de65f9ad9d08d84024c937bd0fe612dbf9263e598d1d6d7cbc258902f28881ed323994dead88d9c973eac5ed872a7ad613249bcae1dd89b128d1281f645a6dfdfad4c9ecf0bbfae13525ae6388843e00ee66b19b228bd88de6736ccd24b26991bd06321810bc34e1343987ec75c589c504e8e7aae868b3c6126dc4e9f1109e4783ec95913119f4ec58ee24f78f036afa31fc3783117e30089fe7ec8a385a9b60f607cab5d4625890876d5cc0a4ca689cec805a39c682b49ba0d4fb37ee42a5f08682eee94b41c35865cd74edf80f0d1d17b5122f36fe44593e1c94ed43ceb81479ee457285d7651af9cb86594a48ac9116909cebce9606ac41c1f5517a47655a6660fd7fd0b90b25cc973542f30da398d8c106cf2c21ad4bc389f6b05ebe8e6844a78b8b1db5d222cfc3aeee8641ef622519a2eb96eec3e4ae2be11572d2834d6fed3b10b703a51f1390533ce6edcfcec331e06780fe71ebb4d4b3df219213cf1e564ff44578aabf6d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h3975c8ff96586f086d36c6d2185e934199407960a5416ec0bb194ebabca594d59e9929e43277a46f50921ec5e61cbd22df26b037a75d95951119705450048a374431376cf9930d4f80fd0e03c19bd1ba29aec23d8704a3acb2a18bea7b961b17dfadae220987e2e425f011d4139bf08db699e601517a7aa1e8e9c31b204ee07b9e4a1fbf860b25fca39fd5dff3897ac211a982d10f47f4f98fb46a2e67512d2076da2368ee4d44eca987447cf17ff0d724ec849cc75e97845ffb3d23fdb6f4b4c0e6ef3126356748597b1b4d0be534a7e78abc3ad0da5b9cb399554427a5b657f18bad76715d1e4ad9dfccbdf578d0b104ca91850f7ebafdfe9dabc4ebada861586841eaf9eabbc7ce3c135d78555e74c776a43279bcba8ab5c7c1c45f12250da5cc6e66dce2648f7ee81d53f45e6492d8913de85d3ae8be752294a24f606379f4d7412ed6460190bcf15cb05bdea2b542248b996d9c37847233aa2acf15367159da5a9ccae55cbbd30b8b6d51cddbc34040f4d8d4fc17abfdccd4e2c3787d6ccbf19eae6359c21c41dd66224fc054ed04d7092211446037362d2ff3c1d3b87e3e110351161021d56ad08883ad2da45d59abdc3dfec69c7d3038f46b27b28875559a9cfc3f5416c19c57a9c9cd2be85be8760f022445c3a9237e55d939f4cb542303ad6643b04e9fb5945942082c90e1f8d9b70f07f8ecc48a19ccb80aeb88c84280affc377acdca746ddeab18d7536f64adfa2e8173101004afa7e43f42f740378532161876c6514b72eae643ac8f89dd0b8d4a572b045ff401fdb1d88b18b5f1899170fc42db29f0148d16760e12f2807955961632d98d8acb2186a3519eca030dd178980feb216ede8e9fe93d0494eb8a64b681ab6f71db3763a0c0c827d6e7a72e21d3e94affe5c4edaf37686adaf8a44a4021024803add01f74b8aaa0d2e82f69010925d92a465ba30be11cccd53f52457e7a7635f4534a346ed26539dd862f40814a3b255346c85f242891de33ea00b9f3c4a9729c56;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h9c62c3b00202969f7ce7c520581509d997985789838cf0c74150ca27d30a3869540396a3334ca7a59d1c981022585b185099ac083af31ebe5195c0d9aa3e1240fb41bb8fbf9481bd6412799fd9f6a2c06615314b0b828b7a91b1d19d3ee0f135cff173dcd7598c56297832ece6f22c9dbfcb0c8665320627b72aa92ae97dd11239066755873eb382745c68a83ac63746af6fcd975370524ecb36dfc0e6bc16bf39049c05844efd0ff7ecf6c8776f64e3f2c08224ab432612ee06f47894dd751b332a3e6347b757b239ea1f3172470610b88d1fa77d5518315fc3888ef27167340fb588faadf0f9e4630f5fb9d28078265ddaf434b36b62f325e1e805890f29721a3f10091eb50c80a088263fbaf2b6e9b26c9dcca049e3ac5b5b6dfe069e65396f2ca5cfce05155d3ecc302fd41cb49a17d01e94de633301593ed9b5da047a26eb471dc44ebecb519f47a66c9d78680b713c5831ebe8f798338963c590318b2e14302eed92aad7a23ad1698887789e51303b4f414b9a37e5cb77533384ba6554bcf54b6802d816072551dd95680676df44e8d854815fa6809bc53d1cb50ac34599fa4a6f97a7ce07f169999c73e866b6f167e68205557d5087c31856b72a90c0db3d29c6d467c04ed15c090efdd097b3937d11e2b4784a40115fd713ddc072e83c8b031d5d849302a6cab6f639fd8f4b822138cd6337472d96edae750b00b60ffd73f931f8accac87a09dcdf904f9521c3f50870f9895ee9600529337b7cb1ce5208f2643ad3d3ef11926087bc641e968733922f58b4c87d1936fca1a753fb4d589b05d9deb811ef2ebba64f13d9a7d17617dc4ea95419f8cbdf4521686d7b3a3db5ef1c2d99ed8ac51ef3285c2816719484e41e7f54f767d9e873256802255aaa3404cdbd06004df6a478afde94f600993e5613869ad8ac6eb03e41d6fb1bf1c494466c9e280356e8f27dca6440715b7e06e0f7d758579ed2614ad1a43c08773e91265ada666b90f705f58691a25d51e0e020a46f40670d01;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h85784622e406d3a79f25a1f3194b8fd3cfaeeaafd09e775ceaf963e8a71930ebd477d653cc22d87891eccd1b45a5af31ccb90f96c911957ec2763ff30ff56bb02805e9da41cea083f3438ca05cdbf99c003275dfda98e16fa011d7285cbfee91ac6c73540d196af88703b4c685d5c840c7bf0d9825f10d359eb668f2b19e2d1198fd5c05dbce192d1d9391d690d955e6a078d99c9bf0f03b78d3843fa13ca5fb5d41e6f05257bdc82366ba781efe788828d824ba6b9c359c08dd5b617308d5f56d74ee923508f8d26d49f917868ffe46805fa1246179417e33ec444d77dcb3acb68e040951ec27795267cae77eacd6875c77627cde99100b33d5635621dde908c13539db444653202206f0bcc80b358f3702026c35f92fbef8eb7fcfc2cac3ba0d10a2dac7f10f2872f35f40af8b745bd4dce8f75f3da5f94290bebaed86998abaf90ced5087dd6abd369e926ca75c8002002d529dc7206d36eb67a1d6c826a1d2f2fb9e1892cff906fb755abbc4af4b09c02d6a27f847e162ef7fd6ae5dc01665d7b6e1181a2feb161f6d51285e33f1c49094fe3f1e4ad0249bf1944ffcdc4a0931de651617c73ccfa51aad9c48adefd616b3d9f10185411906bfd6e29293f218c5b3d89b1f0ce5cf8d684b7994336f7c1bb39f11dc7faf734f03a8004140fe6549bda5779c872703e26868299369cdf894e1fd49bd8269f7fa59682de3fa024acbcc3b737589b02ad9c1bc9600663fa318909681677345018e759a3e8ed2a02a0ed22189fffd254670d0f8e5cc6fcdf7a4ad82aca3c05394c664acbd8e2cd96bd53c1e09297dab46064e51691da7138c1a2c32b7c41ae327e7f423126c95db69f7243cf0a46c1fcaab5a23b030df25bc95a9ee5838d8a9c4fcc74073eebcece4f2387b81891845661126968c0d086e4c572fffcd758c0071b81ba3ab03f04f6c6d3c6267b64aab4b67549a8d317b5df256592ebc7de75214be8ae2eacfc1fc7ed4ea17ece6582ac8075eb5218ee0a85ea0ad610d8a8b9313;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'ha011b11d21d84b8736f2ef76b8eb17d8af419bcfa8166059321b40cc3f799c03a88fb0ca5e2a8ead438b589ec6d3b49da2dba996f6a52357931ce0cc410483f631efda687b802e58af1227919379bde33af79073c532e8d94a0fa976b0da1406d4ad0af946959fcb31ed4cfe9b0814ba2ce2bc3e1d4fb241487cf888f0425b549510579c96cf7cb37211d9d661a53dbc7550a0f941c900d3577aafc818fc4c0cba41ab22a472d6916758ca5f0ac55f7278036d9f9443fd57f019242b5a8e2c2e2e9cde7fd4b457f4f9ef20e1a73b7e24422cff18f1e7e1efdd615d4bfd8a407dd251c83c121349436e53e05ae16a8e5c6cb07e5d3bc1c12e91400e30b39a868600cbd8a9961fbcf11a21984e0c3b4e06aa81e4eed4a86c11be9213c7951d079d114fb64822c630c6cfafaf93e156d61eaf6ea248658765d1fb76323c5edcdfb0409855b48149e8fad8816e3be40250bc1ac33b89005ad07bbcb9c455dcee66387c0181455f5b65d9c1c41056f88f451fac429e42042bfebd11fad40962c48beee440bd4b218e35a42101d7ee4553d81d5609e423238f903b2cc7afcb17b10c284181004997d4cb3f409308677cf79a1b36ef13dafbccb7a7c524d9a687c7aa269d40772d5d6b5cc677ee6a72ed819bb58a51f72713950a029bbd430c3808cad0aef336628474862a43923b1a9366e99ee816f97b35e6d0194d9a4a413b9833239c0d15a17168ea8755c350d6683e6cebd8a594889e159f38da00cd57e22fb4e8ec71f7639005d5600d0e03410c0ccec47633108e34979979bec89c666d49625adaee9aa31c04ed8112ac78e129061583180e0270cd53ac3172ea0f8fd04edb38de19c58193235429ffa6daab0222e5a41fd3015be63f2ad8ebae5d09a0c692aac94a9753850ebd0e4b3503aed2201e2657315c7bfaefe12f2c1cce68813bad711cede28672f5d5c87649eb0ea52869db8ff6bd3cf34b3924324858512b9d7763f8f204f7a1bf42f4bd157c99a545d05696a973aac36896e741;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hb9b94b8b711456954ea1a74156f48d2c459599b9b3ea587889e8b64ac6d4075c83c32c95f66485bd713f565e4158454c9d64f1b2b80d41c857e763434dbe26acc19ecd9db949414efa169033916a640a1b23ff10b7b0129bea8f3e4e44fec567585d777cbf76c95d3bf900e7cadd30ba25da56872764d125a33603fc48dffb2b65e4cc59fd42534b8b14c1c1554a4d4308554a5df704cfb16e7bb5841d15b0fa32abc797497dd1096e6042e145691ec32a02751afffeee94b347a979d1cf6b2baf9edfe7175281017e21fee1370ef17d99946f946cf0d0c870836019eb1c9afa6b33591abfe513b11fe1c27dd82dd3d2643517048351eeab36e5379d3967e88b9822952441cc2a80223a3208aade86200342277fc50fddcf4d1e8fd49baeeb164392578ecff9ab5ab59bf275bbbe4a8fe1202f0417f6e3e2ab019e26189fdf8e3304a5451be0fab406ae7b0214a3e9ad18c2a34026f9b226d2e3c0465b5aa41c1879b0ccf7f05d7a7875afb53a54595232f2c9f4ba753d0e7f31db2bfd10655528a4ed993fd8f397550a8d141e6d8a86435f6f43537c697b64168a2155330ce6e126e1c003dc5206bfd76cf77b1f6ee63f548f75c1f135022fbb30958ad33c40fe9f0fc8706ad93f02da29d23f86317c4372cae5ce334e5f9aba6558345d19481afcef8e6a7faaab04aef600c5c21cadb6bd09a4d53e62f9ba5ef56b50f0c05b34e5311d07e2b8a4bae1cb44ac95a08d49e41fe4d93d491fa29852cce132d1da8a8c56f87b3b4b02ba3e0a72548b51f443472a67b5ce25e6633989a0c9b0f1d45f26df08f36e6e90cc6330570c802cd197c55b7600f20f35ba09c573ce4b66cd726d0fb5cef8a2a1cfab71bb56f9dc6b7e2749ccc6244da18af144217f8e5e70f334bb09088638ca67c1ab0339166aa9b776c58c670a93874233bec9181b1ecfd213c45bba005db8732069954ba27e8793eeb128e3dd2aa5f1430bc66cd8877385e0830b8494666ec0c2b4cd863afd6849924e88cc2ce7b0e0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'he6a4176e9739b40d1ce70bd408e125113379736d4a8675dedcd9076c31fddcd7d8452a660f2e2a28708afd384728cf8a055e992b8dc5dee71231b4f14567ade3a94f5ab6f9e7c49ee8bfc765bab3659c1be873237256fc7a42b35224b81e97d4efa3bf79a08284f63c224b7eb53d9b074541de744ba8a452c8b46c55e82a70e37f9650c757807ccd79f939d9104a8098918a3fa7c1fa3c6fd1e216c36d623cb1e2a99274e172d33711489b10172b14abf0324e7d69bd4b15ebc356dd12cb1b06ef6770e92e728a7fc1451601c6d0527c1bb4bc3e482393f4c19e6a164bd7de4be016b1f36ca2cf67f895c88a47b33d6afdef0469b9f47b5301477f3ef80cef56e3626b77ef5a7ee06f54cfe76741a9719843f2d6c55ea49d1a67b9c84d888be813b1d58cdeb64a27447ca3a83f51315c156553b682529a5e3b89ce4a70fdc35486b42ce5a5ab952fa0cf97ce1e4119f34fce6f478645c731e1b8c9462171bbb57fb5be62c4830b7648d502dbdbc140a6f5549d30b9e248967cda1f0802ad4c5d2391a57fb38622c8d476e412892be66dea07e6e05c5485ee885635a747a904a49bc218256d79a5c7cf1268b571724e17a445b4056c3269609e054bc572bebbf384cf59a7ab976cca2262e4889bd24b33854626032451ce779f0226759602ba818dde983e16a5362b0a76d6b9c3901be0831d0ae2c8c63d822fa9f19fbcef0f9e79a9bcf35ac0d344b17a8ddadf1ea294cc0e57c5bb66cd3a651e80d39ba43adcdc68b25c769e4180fbbfd8b5d24f1738dfd2fb364287b26f7092fed3d45e25440329ac22753833edee5ba205a4b4be5e986bf20b6ee662545e1fbae5624c8bc625c4126b63d8a9dc685653f29089b97cae5679127e31c81b4dbc3a47a791b9482b417ce07af9e258412c9dda50403aa6272362de6322fe5f708f360647c818552d88ad4859406630abc55b9805e13ecb85d33c07de386d7b92e47848e7f7d57a5a58542118216ef5a939f4ca8da41ecbc3e101ce7b6d61245b;
        #1
        $finish();
    end
endmodule
