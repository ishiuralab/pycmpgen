module testbench();
    reg [20:0] src0;
    reg [20:0] src1;
    reg [20:0] src2;
    reg [20:0] src3;
    reg [20:0] src4;
    reg [20:0] src5;
    reg [20:0] src6;
    reg [20:0] src7;
    reg [20:0] src8;
    reg [20:0] src9;
    reg [20:0] src10;
    reg [20:0] src11;
    reg [20:0] src12;
    reg [20:0] src13;
    reg [20:0] src14;
    reg [20:0] src15;
    reg [20:0] src16;
    reg [20:0] src17;
    reg [20:0] src18;
    reg [20:0] src19;
    reg [20:0] src20;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [25:0] srcsum;
    wire [25:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17bacd25876b3b55a57e9bf9cf87ef1d9a9278f92df5da81d7926198d0e4b07cd09245007d4938893d2d40850fca558a2df056fd4ef1af3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf5c89458b90ccda54d260b99aeac3288cb7a50d320e326ef5154eeedc666bbb912e249afc11df09770b0f7724c189409e6fdf6c55e6464;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f061baa36cb5a4aac377f556e506660f60f3678a1b0b8c1358931612015a5a819cb0a36df5818339289ff4d9e17ed8586dc68ea67d6d26;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1133a09479cc1f43728ae2add52b48fc301793ee307cde73244970d9594492ec462d15fb79053b549b343a3311626e1738784f4efe2986b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5414fa04a9ba66f2ebfb58f2d200c285820e91bc26c9c65ac2a9563c9b520c140454b9acab01a579978daa98e5df2310582ce32b4e83e8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5297035d42364c52aa007ded2366b75b64765435cddd6aeeea74608c81caf10cca3b85e821065f131bbe579a7b3a12f08b8e50177e1251;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc6d7d71117129fb04bce42eddf7a999c5ab9c62175b93bd2accc424d03502cbd91c684d47ca7c2a7271c4db706fcfe64de5a3fe61a8de1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h71d788b4413934862b8a96a9505c6a68fc9dea5d335ece46ea75f4a77ae65a0773b9a474f528a2a036c79967b0f3c6765471776fa02297;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1de7845f4163b490077daca8f5dea01d02b6339e4ff35a83ec6a2fde5470633b0cf028561ac01fd8d75691c3b84094c297ba77e599e2149;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h647e994e89396c5f4d1ae712d2e596b05c20d7682ae44cd9c91f575137e17405b21a94a184811351dc8a66ba87086960f6cd31ec5887ea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16d3d8a5845c44241d4cf8182ca05f865a5f8992d5bd0cbc21b1cfacad26f8f2a3292585659f6bdbc74acdd60e6c2364f17023c02f2dcb9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11bdc2f1da40b5c8220e80ad4c511a4604cd76b905e7fe1a1e91189c8b2fe4381e56b28fb3739c806214bc2a037d8ca2d698456d80842bd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h81259e799723939e614183444d81cee1bd05abbc3620e21690e2a69ea75e9b4d211dbd1a4f93c83caee5fbd00279ee7d6ee686edba89ec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17c70afa2ca8fc388e80116c70bdd13e784c7f00db97c77970dbf3e892d8d5c9ed6f0931f43275692104778192a56f0bc89fb7e221895eb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19e5849a104ab656f9f56ec1afc0f5fa123a4a981cd45f224b27c8b5305c25b15e1f352d5f9379bd149b87e288f624c25420858fc8396d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dc208c1e0b9da6565fedaf1d169d877191b8eda52a9c37512a19e985240722fab3f57a5794d0fe6cbab061f651d85dc9b5015a2fd9ba7a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f511f9d12c6c0ee379e85591a6022512548746d8fdadda2e92f2c883ec9742e06717cce0e0c9ff097e68aae07b9398ed53c9034c0938b5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h140914401eee9665f79edff942e4a29f8a1111896affa8f1aee38ff85a6e7c63fda223cd58092e074fd04a3468d68eefc8eb46355b6dce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15d10b371cb434384fc1e95b23a77947aa3026de2f90e8d590f17f9e136794b22af28ebad31f6987b2eb0aaa1425178fa828b337c04d7e2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6b6e607d24f610ac57b37a0c7871ac728900230e522b0af8cee8a9fe375d375b897c8c78507d5d9417c54ff2bc828321a8399a668c9edb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a6bd5561e802db9b2694353748b5f04b8a94725f6a3681eedf2a0d61b4935aeb5a0cca2636d17a6b034ace298393367a002a009ef7506f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h61e01c12d10c16a210b84f4274ed2804697e68fb07cd54ec09854c608cb3427bf8bbcf2215e81eeeb0fb4c2a5eb89039feaff49980bcd1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18643e0736630be8d96633184e6147ecdb68a2de95f04189d5c401ceb09c7265efdb93d758b37db0f5061bd674487eee85889735e2a8f02;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha5ff7e844af1dcadad7d93b8dea51648856114d03d647136b0177e2ccfcfdc0d83c69fa0a9443936108379fdea95d1be174f5369e1c101;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18a2eded008136af82d48125d3ac4eb4b4338b59f5458b0e61669babbbe13152c8889596e7550581ff564de1c5c1d73f7698aeb22024246;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h716dbe536e0890cf432d19c8a2a9ef30381ab84b539c058708c99a07690095ed68f175bde252cf87ca48bfce1e93a15cd425e810fb05b8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e46e596f4704c8acac2aa24a0f55a0ef5be9642848cdb35218fbbef64a65505858dbcbd34dbf4aad31a510640b721be143967c38ff1418;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12e60dd6dd24255d58b1d92179a83c5a30e643dc2b46b2317713f9fc49a358ce97fe04939de34b6baefc3115f7b1557cafd11a3cc24228b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h199f4ff00b3bea4a80ffc0ed4d53fd2ce1bafcc48ea8c02d3f19e5b6f0cd7fa4fbcef8f0bece4d2364a03c21e7a8803401d3306637b7d58;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h64d4893e6dacb3b298751561ccc5b62ecf194465f8363b639acb49bd7a458734fd67c5d57c270e6ae083562546f4abd5b3d6ce67b8e86d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2846dc5e8e64b08cf362e90ce9958915d42d593696f95bbe5e1ec927adcbbe7263684d0d8d5881f228d86776f5447f3f93dc2e280490a7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hae6d489c722bfe6fbfca8c65a1f13161030a5a4209df9e7fdbd8025e6cc0ca79fde88933e4c0381dcfe5a9b89da2bd8fbc493dc697ae6c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11f65309e8b24933966c555d042f14f34844654a5291e504df23d914a3783f1cbc3a9ee3a1c7f207f19b76aedfcf5f7924bf5db9e71d02;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfd319588e724213d4365909f2ba864ed8b098d26df783ade584d069fa998f56fd7f06e5c461018ea2c62855ed5d7ae488f77af4939b458;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he9519059d5ab944bc21b34b8892985b8cb3a753a6a269e10fa19184367f207e228b816740435b20b677a92cf35f1676e93a22cca457ce9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14a32ae7c066bb675dc31265d8b8b3ccadd7f03998e07f596416fab32c11e6084ccc4f1ed12b93fa814a040f0e61783ad037802d68be1ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19fcb65d1b099b61fe5cada51d5bd68689572d61b2aca27d0edb3b964d2d57620431fd70bffc178ae432aa14f13b44845dbd4d98f293e09;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4f3e5b18a5d2c3ffda14ccdb44fa781b7297fb085aaecbcf37c9e75589055b67cc511700ab92be5be6ab535d6ec01c5e3297cb5411a12e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17f1ce14b3bc1f7bf390f9b0920e987a9eeb935469cc4691f764d7cbf8bab10e5c984d9478f1cc470cffb52cf689d8689f6b4370bd8fadc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h129066ba68f85d9a2d989292d61e7342c9a4f281c7db5c0270240857274dfb02838919fdde05e324f2de0349227779733565ce7592b3f02;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1979a48874ff76fa9182f3e424e84c03fd48761feea14c55815a2dbc7b3988466ced1184715690d39d1d20cce60974e3f69c32b45b0ccb5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1427f703a4ae64120bd5f2829c0e282dce18feea5ce20bd81304a330166cc040b891d51820a22357a9c455d7e8c4c35a982246b6ddcf152;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h90a489053826f071c78d8b79eeb35989b28a97ddc4bf9c0af5515d190c5b719840e730cdc3e403d85901466aed6cf7d0d596d691988513;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f62294062597ee91e266ac5d60bb4c311364e8e27d86a3c3b44e4f14d679e23aacfa4e3412c17ad5fb490524153ad25a020d11627943f9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e4777f6f5a6100872b679820cdcc4ffaaa8544249057f978b1e33775f6d559e1f96e7016cfe4b69de55aa0eb8cf34e98040a35ebc582d8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h164a2552e24aa575745a47e4490e3472ce9f22c8a1d938dea4801c802742e83cbf099a946c69f17317c730c58440f1511d316e08807cd7a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f64c58fbcfec4180a66da9d1f4fa58965b478e803808135176939661e5b4b7c511db8cfa658d5a3bf33c8f468f5f3099ec0e1e44b5fa80;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h193c0185888704e64648e9c50203828df25bb084ad758d81d99b1897b9fe9612366da93c3b57eb82e453afbb7bc45731fd86e9823d6b5f1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9a5196ef9adef2f078993be77d740dab3730b321c2f41eff2d3c856045415e336c364a9670322f996db88cbaae153c18d08bb0baa384ca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h89bc77fdb0beb87c95d352d2954de9369b6c514acaeb536ca23a82355b38addbbe78dcd3d896d99d935f37e8699d41a13c2c9ec69feb15;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6ed57df4617f1c926d4af1ced42dbfe3caf04485b775378c3fde660cdb0b171588b46b4e06851525457c7e9d9c1f80a89a9efaacf3dd80;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha451ef36fec0cf7d5e45a52ef10d5a1ec9997844ca49c097efa5be62667afb2f122f3664a4727b1199aaa794035abba407432b36c60b46;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h598815c190e56f488483b914012febc4ce6a8602d62472e35e544986cc7544bcb01f405c306aac7055f26276088c41b2a406d1c83340ce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h102cebc4709bbe12c6f1a052fc86f25e6b38f01d866787b190d671501f38a6fc06996e3be6cdd09517c42fa2553e4b73dec299eeeef120e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haeb83507831b3449cbb74c445e2c08cc0486a987e27d5e082338c8b013fd3c8d314c6c1efb37cd5d6ec44bc0d318033b659f4500586d4a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h39abf6d11cb4057c6bddbd848797bcd6c4b73211c0249a37ffbfc50b0849226a1d3c56d51f10dc8e37ac8ddc1bbe5e716f0a42cdc9df67;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c0219f68497fbd04f05d4bab969a7c868e22a8b05e17bc962aed1d56118514d03650b381e378fb0b81ac5f5341958a7b2a1d6387e6f5c5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1746eae6f89f292ed4d5149ff4f45e043e309af71728dfe32c32bb9bf119a4b196665dfb7861aa91c51f9adf3d603c15e998f2cee31be77;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6dca1894f4ada7972271a103cfd1cb80d2db547f091cf560f6fa746fec23efaecf515ffcb417f65aeb47b7c3f5484b3324a2ff0f608c60;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h952e414ba6e646fa8aca8ce73fce3d5a5359c5a22cc5214e7761b77af76f3af3ffd66d2c2e39770af2b03ca44203f17d5101ad81796d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h100496d391fa4fc7f1f2f103dec0dbf0bd5471a47113e4a5306cbf69ac2ad85f7659f68e39297a3d1966905e822a2219007146bcb657fbb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h108666b58835e518fe7e82668943a04fbeb90ad5c8464f90e9dcb67a1b47f0f7f5c0137638d71059a5f0cd4a4932809ce82531417fd6a88;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1765c0e887c40eff2b959f15431e03a6db67bcbfc7ee71ec184b8d96f32bc3375076410bf2f33f43d70abd8052e9b2fa26a6f78f59949a8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h162f00b90612c6abc4cfd750c06184daeabace8432a52d68542f423fe4fd0a0f74eff51a47e33b460ac71dd95a6450ae69affd19295e328;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7bca8e7a9c6987ceefa8cb379021fed529332826498309e0fa96d868c886793994f23e51d57b85d0148095eb7fdf8f19d20118dc1d3c38;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd234d399b342b35d52799c787cbf7b47e204f58fb5df0a04d3309e19e247d196d11eb1a57f54724a98b4b1b53f7426a25bef7326901b21;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c704dbad74f6b62eba7743bd9e39698f8868ad8c945dbb55cc1add6f202d409acf0bbe68499686937cff726087c80445ca5daeab67e007;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e94c51cf76c1074ce0ce81b3244dcca04fbac46bfce092bf0dcb29b25b5f5afd3be825b8ba7dafcb014bcb2c6f74c0feaa8bbd3029002f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13588ed6873ad43cb47d3594c640172bc93f504a8b8c645c7a140f6acd89ffc3bdb329ce3c9012c43cc7c72b813b900b2f96d563bb67ccf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1807b87820411e586c48a8280f787ffa297604628509027faf7ede298e5e36f03bfafecac1e7e432fe8f8a89fd2e8aa71cc0f2658c85e02;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8a3e1586f665af6f584003b356144b85090399edcff340cc1a09b42c5817368eda0a3d23dddbe34a51127120f0dc6b3c4ded9de83fcf82;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f924559279db56dd875e03e797a0afe3064606f1def72c0ba2934118137cc6144f57951a74c17ee92c6873b289e438ed2583e15462f025;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h32417a17993a2d1ef9f7e804ab8891485ce7277d6cf0eeedddfdfe53b597a2918d030d2f09173d9abd2a26564a1c394d90291b69edfacc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h63e116dcb32317488fb81482090e9a9aa67f21f41ada76f9111fc1caad193140f673ecbe852cf4fb91969247f199c81b7a606f0b4c4ec5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12c2a0eadd36082cb65066e1dc4c934b3193dcd9d1fa9d247d6d1bf7b0d37209c6f32469956ea06bb85c87225d51d867a6abdc8b858aaf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h158ae9c889d43b1933dfea82250fffba8097018a768a919087aed24621c85fbce791e6adba7627396611da4ca256716335bf00d8bc97792;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h195a6b4d7d5ed1040a2d72afff2eb64e3a5edec31f25c5849cd2d850e47ee8382916ecb909677baeb03c626e4e2c80bfc6cea531d4e248;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h79c6b3810a67c2bd568277bab82a672e8fa8d1a9edfddcd4fa68dc0ef8e1002cf82e972a625f89525a76c69d2cdf614c894417dd341eac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1489e87865caa81080bd1ea076ed3b5c46eb2efa2caa7930fc9d13c6a7cf490c6e298f312e515a155b4b4199965baa91e22a3e6ce3b0991;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14b0b6826c17b85f49d0948f59edaa67c992b58ed1770209d42410ab48396196c10fa04c264e57e158f115f7d4b7691619a82a7a172c916;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15e5ed9b0535e8c548496b65824dfa76b3c547575ccd83d698157492e3e9b018b9597c4731b255461418760917119c570f4088dbd2e23d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h114547ca4c4c5b334d9b305f9e114dd37d1fc22937a2585662aee4eaad8864bc5dff36fc92e24508d43856a043ea0d15e9773e68ba98afb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b56a2f3607a98eeecf01e22521060796bfe272feef9707b630cfe6f007c9cbb0487bfbc77c3b7f1c21b9e68508bbf63f79377693200785;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbca3659942d5cb699d7ad07a94c410beba58b55acca4d5296fca0b73a3be00e0836d7dfddd80297cd423a180bea51f3864f72a1e71099b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11630b0b7c7c8a4f06dd7289cc5a6b3fc5bb64aef5e2f54853172ec0d4a6aa34e1c75efd1c4bb4f7335745aab9e51237a3c97465f0e0e66;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b30ecc11376207248b2d7138445d9db78501ad3f9b4e079b3f92927eb63d199f3bc8ae01fb35a82522f493503f8fd4884f2ce867a6a0f4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1201fac7906be4632e766c3a8d6fced50831408977d7ad831f5d75a01705936d54e1ec27e22da2fa1a4576bf3b952ace20869391ddd7ff7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e6955030bf0e6add8a8d7865fb241ae13db45e4484c5d0dbf541acc75c1713a0ed9df271c96c683efef76d517d71df99d2f80cdb4878b4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9dc47b62d0ce4ea1f2c1021e11859b61fede4d3f7d98ed2af304621cd9ca6101132e354ee2fd7b8469dba0e0d176ba61a686587ebf22c2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h130d676a555c4abfe87a02013c688d17222404dde200ad3d238145a8a197d564b7ec62a2430ad74eef2661969575cb7d4fa88f5c2998e53;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f8b3ab62743fcb760ec442f755407d7643f3d857a79456db32762d9286f7aa905f2b9c36f81363892166dae974696673788c23b4bd6400;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ca5eb124d18411e561392639e18e5fd458bc6295b496532affc41db821f212457a3a01214761a6201b37f4fab68aaaa734df1be8488aad;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd0a70b45b9fe2c0e218f30d95e62ef89cfe44ffd773db88df93c68a14268fabfb66abc1c93de820cea86bfcc251daade6a26d357503b0c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfef100d5967a036a235b5519e256def0ec44363fe7498bc02ea1f918c1ae221d6b98d369df2b1baa980fabb86601a64d675d1d39cbafdc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17991aa5dc25d82e7645c6a8545b633addb4ba6942af76c99c569305da0b58d7c66fdfc9c7df7f602a769ba3bca32694a34b464ee1253ad;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h77ae03d1dce92e6312758454a70af25557234f8e7b9531494a26eae0f854dc8f9519933bb76b347aa5a46d3391acdf0e1bc203a56431b1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3712b3f858799b965718a7ba39857e29e24ee59049c3d8d7c63d6440e6ca9aed7a09f0dbe2b0ebe315efda1664bd7afd59c7934f96c90f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14f8a9c7c0cd51ca6013071d516bd2f4eb706d235d906182b1ee7b2ef09b756575bb44170a1e004d86086ab25494d0870b7b9df93bdbe7f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8156ace6914a6515ff5a917c45bee19022961607d2df66a1b849ba34ffc347df9336656511d0865e164dfa26d3f24ada1941af0f5892a6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2fdf4873e9cfe26f9d6874051ed1f2216af656e3a0ff8e861f1c06107a4d0d821d746b2bee68416bfe56ee4365a02be697255e47e1dcb9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7657e0299629a9adc5a3bfc5b94dc71fec25622558d05579997048f77ef17671ced9c113398a22f2c167bb7c9e1c883c6d95bf158f19da;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fedc507f055aefecaf06e9e015b9ee516310d55174e39dd46b0113168b4d7786ff6d04bc27a16153f6c9040041da7573cefa92da40a8f6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h107beb9428dc38607f178cd8d4f8edb5b47e8f20ae0c03cac3524b5990af13f5556e57d33c68541164dbef420bc9636eb596a15203e89d5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h164831559f89f5f3c0e50b40bd19ebc20fa871d519bc058c41db8a416b26d5d951065890ccdc5e4f2e1150b6786d8d7d845d29710ecb4ae;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c6e8eba3eb78aaf6de09ab138fccbcd0ff72fb6bbe706393ab016f0d19edeb48832eb05b2ef49f9dc3eaa776166ea88bde97083486941b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a7dae48332714f8c086de4cecc84930466b77730db10184a50a18b861efcc22efc3fde8893951fbc3314442565f3e115ca9372148e9274;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b54bee312678910c951e6b76141fc48cb309a9a9664f5f1300729bb2526e07d7e110572056f4dbc0cfe78e2f13878b3fdc34c0a1d08be0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h31bb891a8d64fb75f6d96dc3692e01b1daf8c3ce334df42dde40fe26f2cae05b8b89ad1353a6e8a4b1118026612b65883111ec7f54fd4c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d50b28533ca74d2cc2f847755d16d5789af2e8784ade98a6bf602c7045e8d548e78aff55e4f6381d026ceb9bf810da1799a7c76960e42a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h173fbdc75251f8e2614019ae35bb584e18337b236d3843c9196db7985a8a48331fbd003ca059cce54dc0f898b2b7e82514da36ca4ba3eb6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17c1cc043280f0639c2f4f808e3ee3e4b8f3bdf581a436358c01c8751a88997146137e2d78cf1da30a03d2b4ad592763abf61c4410977b3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h541bb0667d362608f9ffe11919568da7e72dceba7ca3c99b943856eae48628312589e617e57552ff320211dc347a69a4e6f4f4053efe80;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1afd391153d86a54ddd73b7f730a2d3e1c9037122f00b889c83f71caf5f0ade18f21fcf479e0d344f0c32587d35851633d596137480347b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5e81c22042fdcab39b17b34ccd65f43ff42b689ad9fdc6d6a1cab14a9c0fdf27572f71f336509780df194f292c3f4344ff4d3c832f3688;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18ff891bf33a49407141679daf0e095f5642cc559d4fa06b3a4b066d40e9a13c3d8cb656a68d9987cc3c60a5f29be093c1275edc3bf53a4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha85b5081dabd63333cecaa7fd20dc5c69eba96ca0d20f9cc117d084c5db39549ef855faefe235780f461b8f8ce3d20b7db3996390005b8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h76bab022e8b2740382658813d62913c5f1c775e327357dde4a5f26a10964947ae9bf05aa9ee03a389d973f6c22f3e9c88406074fd0923b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha78692a2e76b96a4ed0b61ea245eaf8a8203bba71ad7255980d612ca71bd292f535588dc56fe7420ed0e504e2f58ff54e5fa948dd90f59;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hff855abe31945a0bece5e2e638505a36b6858e3f9464bbf2a3003fe61dd10d0f1f9d7b59207a3badd2d1cdc9f5cbd9959a33be1d3615ca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16f94a925b8afd6e4eb78a01802aa38a47ceefdfe49bb4aa6b054c2787d497825e4fbd229b98f597d0a7eef9be6176be8c835ebae26cf60;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ec0a4fd41512bd332052b5b31e4214bf3bbe41c463b904d26d80b55ecc7603bc0ac3ddf07ef401bd20f9f910edebf46f986eda1e9e1c1f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha622f58f547f8051b6abcf0d5cee484cfb436d0b11001b2fabd28c4dc86e095aca4bf54bf63b2046bb8ad077898e9346c7c3e2a6fc394;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e67eddc853cf5d9fd5282a7f3a2c620276db1b34dd802699f5341212d8e99006a55e409592b59ddaa1055ddfe94e8d4161d6265e8d2f9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14b116c97df9dba8987c1f60631460739f6d9ef50a159dab75e3e5212f5dac798a6a4eef11ab25c292db5f052271876ea593a19e49958ec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c824427d49558d76123f2f2907ef56b4795799dc03ee2116b26b445af2288ae1654dee24b9f0ae34f7228a4885b06d2cda60db78697f50;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd4f697dcd7c370c0de8b01f79d625dedd80af643d19c2460fc979937ea8d330992f0ca82d968b65060f535345a6fb94ea446152e1528eb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h107ab8d18655d600f0a87f16e4932340e11cbb770f3e95fc9e2aba62a31368a4f627c07d5c8eb7f2adc0e9ab1effc92694e634fe1df11e4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c7911c2c41b763c41e326675b1ed323d1ecdb27b73744b744309be088cf07b7b43bbb2ff7c9934154d5c980fde6a8d880770708381acc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15ac5b91a296d6c8a324cf347f22b0d3a5f7fa2d944c6bdb3ac312e9ee4246cbe97e433db79004ac7393c942ad516389253f2c65d4640e4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1aa993cc066c53a324a29393da89cfa7fb9921219b2f8ee3315d30a45fccdb48ffaf93dcf0592e814bfe6a2f493789f788a407baea0b2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h190bdc52331668a731a5f2b2802b44f6edc91b34f120a12a01ff18825150511d39f7ca540df437fe6fc0c43202bf5f9dcc7f9096cda9d25;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h121255cc7150672a7a843dd3172766c147aeeba194142a11da7f5ec7c1146f9c25876d46e830da0d0db4d138cd990de37037b4ff30f6fb4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19ba97e3d774dfd6691f822b9a5b8eb8fde1ff707faae60c5a8247c5ed188ceaa729ad36c9831508df3a94627af7229912457f9379d7219;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h615aed92e2f7475fe22b4c9096fd7fa3dd2650eb0809cbcf21ab1ceb11b01f9a3d19caa4ef330024de6b658a2ef55678458cc457a68e9b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h190e3d48f32b21f9bee34a53b997582f0ba2a20a93ec984652b0a045af114bc1d31010022c04c0117532b1c25a066c7ed3528293a5d4610;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15d13f4715cc1aab48da39abcb47b6acae4236e8653522606932ae1ea52049eb8383f693e75956008ac565daedfd192ad3fcf10e34dde6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19b5bc1ea74db85396dd6d98c22d910ded5ed67306179831b1fa7511e0d02212b8cf96ef9f530f0ee7727a221d649c2ce7bc865bf9e1f45;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h184531c682ed03a3103954ae5aaf9bd2855fc95f4df64e24db734e2b425e394f0e429412bb656014738c026bfc6a165c9c62c7372eb6cb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h133c7d56aba7d95abef3fd5c786ebc296f4b47c6d61c40e3fb1a0c35bffe06fa6cda168f98eadf9c376c20cd1ec75f26bfe0decdaac0d92;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6a73dd5cba31ebfd819826dbcd6052d88c2ab099c85044518ead4b6339ac9f855e3d9f767bf58873d5b29afa547133f657e2e2609d59;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18b019f2942551cb617fc1edc068f41a74ec1af146c6401c8b6f4970632734d65aed472030e9fec262faf8a972e7f79dd1c8fd2fc4e46b8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8092e9dd35f411ec276ec909dedfbc7d3744d36b938592538bee917f091256971a81604fc4981ddee2f49678028f2b7e1dd9bed3d7176d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcba068e6d14d69bc387e724905dc73b62587c6778050fba15e4dd6e1d5a9cd7428133758c07efa76d2c49561be95c523c871e77a22e704;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7b7450822f77d29290cc31ae5ec99d7f0fb78d686d3c08fed1a3177647c3910099406f5919198f84afff425673d6b8c4cb232ea9071c60;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14d6965e7cab3fac10cc42c3dec987865706b099a5eed6909de1b4444872d35f3b73c7af8ea4cb363b9d21f2c495e9f87fdf24fcdd9ff7f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a9faa2ef38f01c1564a9a550042c5f58a5c2049cb8f6f8fba7d6927406f10249ca8c2e6d7b6df4e42318f17e32fb0d399298496881dde6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17caf7de9903fc7b6f1d3bdfe774b740bd9f419d7afa16ccfe5964f0ba33959b201560f7719ffa7c136359b13692afaa2ae3005b40ab4ee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5f6937b44734c56a04c868da24ef391bce83512eeee6ff67a11744be4b477788149bf83237acc6a8117cf6d0d1ce8ea5ba15c78f437047;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14d43fea40a03df10a6796345e6a9f1429b1102b132eecbe3eff21448714fc4b7d57d2ac263d9bbe5b36a1c46c87dbb4c0e620850f65f23;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1830dd48519da0ebdc3f472eb9fca62c534f3e2656f5fa747c8bc546f7749648c5d4d0f16c88b0a171234796689110464600802759af501;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4c7f19588422bb350b1dbc5a1b764856de314367e99c080a412371698aa41e03fd46384b30d92825249fed81a26c623d3ac189262cb7be;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14085f76d1e4134da909a1e7c187db4a6b24c2806518dc1afdb9f05cdc374ba1bcf2d12c1e706470231516aab3b725627f6c6153f577787;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19803bf66ed107a196282c2774693585d17f10c14e5be0bce43b28190d9219c60cd7e810ecf36b861c357555ac4b9cf0a4adeb7fe7aee6f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h146d156c590f0c481dfe2e9e877c560f5a0c43da691f4288b2d80fd39c6306257810deb247469411d1783b265404191b02ef838c2068f2a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c5363ecd8af5e1bd249867ca2b601e2253100055d19b6766bf7f1f554b2d35a4736bad181b7de6b1a1a52adf9d30ae5d28c8fa37716dfb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7b17846611a4a0573f7e8dbdd2574e61cac8c59fff3f3f8c9766f6055f842be093acf89dd9ae23b93d9a7afa3915d993378abe375081dd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15a1f775670d65b7855dbdde438ae407ca9d159b4386dea189ad3fca102570523518518ba65461a70cefb685e615320af94197524c9bbd9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1279003891456ee79a4b6d09ae79c79db2afcdf23c9aa61cf41d7063ca701e78d21ef63da337e715c05e22aa32213857b89a28d6cc195b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1244fe638ab35d417d23ac234f13be55d619ab3943c9ce29691f82567f4b5721af51bba3f5a7f6541fe7eeb1b25dd6f89a8957448e2e681;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h209ec1be75acb0c9b032f7141473f4a6b175e7acd89f673695926533fb53ee3855d8e54e78c9fe3a1e7380b68e01ac3cf4ddb882c0bb47;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he457803d71c7ce593c081ba789ebb16da4c8416161a2271e4dd7c550cce8d04b7c573c85c1b2e7db279b1ecff461d6cc0dd1749fb5a677;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14fc8fcd8a0928beb10c90bfb68d6e2cba4ab9c0d5c991abc981613c832f6178edf8546d191503f066bac8c2ea6a686e3d563fdb7da7b5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a18b6301cf4421f146b1aac8fc77b2027352f3e1e087eac2ca683a15bd03488d503b2ea03a86843cd9b8fa56245dba9cc21f4dae4ca9eb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hba0dfcd16254b14656b8ce2a852225c26cbac2f0e4abe0fd3aa201183676e5a45b1308d043aa8d76f7363f8addad21fee423d98d3fd299;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he289e75d5c4ac191b0eee3da5c71cff2305751acaa52f1796aa2a83f30ed383e9db0bdf094bc4aaff9393349fb126ef6c1b9054076142c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1981e2e6162bfed12a96ceb72c510a962f99a64de89a626a8c0474583e2e8a5c02237b4ed0aac47f3328a76166c28c573f3d9cd8f5a5091;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h146e1f31391656f25f4a87bd935c2b9e19bd1f373be50403fc608d9313441a22236ac218650c32ad05b97a26f77297c94255c841cf8ba3c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16e24fbb9475a3e26959ed218f0bef907b1a5b5498606dc6bb51ce325d86d40578aff6d032da01ef14f775800237aa02be93c504eeffb21;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8d873984409bf6745abb503fbc7d9b447272ef8dd84342a55f8f36b5a8f1ed5526560b793f420fcc676e650fbae9aeb94536c6e8a1fe2b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h509998fd2b496ebc8ac2311e34e0a61e8868e579f05355ae4b465d74bd346f7524804007527b1721e0f6d0513fcde5436f13ca939385eb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h268f92af8374fe7300c2391c32dca3c9487a75c6307fe399a0a4f4b2f71318fbd1e6d35fd59ec2b9e201356d0a91ddf9776c3fa4898323;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1909b2fa38ada7973305b7d1be5f8f45ab49b3fc1064f6a023f4339013e53b87adf9102af2bdd16c88b0a45df491138044837492969e150;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1196fb78dc930c0d3b2a33e96b3516f8d941622bbed3a4269b1231c321835d017449c398b779395fbec437044b0fc881867fc32e8d1aa36;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h134e465cf91836c2169c872bd729b53889bb03918e28b7840c75e20e5f0842c45b43cb169df22d3d2780e18087557dd84b1ad188d4e22c3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h107116ba8358570d382a9ccb3bc5a2e4df7213be6157043381a01ce644baeff8a2ef91b3a4011ee3c7bd0e5e6b3bd84517622f14334dc44;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h190e64977bd88b510e5eb038ba4d8f9b39ab8f19569beb89e8d63cbee75b126d7f13a3e80307e5fa2ce35861b50f60dc2e55d1c784893a7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1637a18bea95688ac396987990dceb76f8898d12f286045e1b710e41e0b28ea920c24872d22bc48ecad71f40e37808f39b1c19f5a0710e6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf098ea2587fa7bab290f218932fde598024baa5093423fe002193c27e68176bfde2f806284a7361cfcaae891072a8321b3edea1e2f5a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17da5c8fda43d9c83c74fc5180e7fa664ea097d348c405e54d2f23e462519602c1a06dd2c41a320cd12f92346f35d7321e1ed023db6d7c4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h43bd5dab2597098075208a8e2d540e30994a5b7d98794f24b1993fd8206e0c7e0f87fa078a6d7f83aa9fe7523c0fd0fc1f5cdcecbecb7c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h190b9572d8cdf1945bb6168a8950a95baff0186f12edddb6fa5ddad1074d4437dcd188f4e97258022d5612c4ad67b79e3b7b720e1e270a5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f3e564fc58fba97ba969e82d19fedd65e73829302e947a7883cba3018aa01e65155cb91f3389948e009d3c67a135d53629b2015f477e97;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1908072357c5e077c3404952fc358bceb71ebd36547b7df459c9f1d3c472aaf20f6101250f7f1fa7662a2f4f96db4911b43c14da59500be;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a56649fdca71583193f911aa9d8987df3f954b1c42d60b02757fc1a0b2103f917fcda94b6dffce5f4e98d88809fcb73bd59dd2ff5730f2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h305673dc4fbc969917f71fb871baa11ebc576ee22cdc1cf8c1ebe21c0df845e5bcece21e27eac1e36334a3e184abb4a0192811f85fbe42;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c1cfecc329d826713687b3b763e2b1dc127475c26d1810a7a7d066c337c7a160509f08bbbf4ff553da4e537d4f52aa5b55a5bfd4b7f1de;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1396be019e106f4a73f397e8054b77e9a2cc6b73c6faccd9b82b59e3de3d43eafe6c29058c16b9a14516f831797bea71dac965b1ef47bb2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h187ae4a0fe282deaf4b969d2d1d71d9d0f8a039667b36adbd890746d844b8307c0efb4b3c6280340d9d1797e1889562ed0acfcc64066460;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18bd7c4c79aef848ed215669dafe52cd20b30e30923843f5c507364c558ac6e5657c66a92c4b1963eeed1ae83eb08d8af3705691647eb4a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h107f73ac1e7592b29bbdb9523f55f7217fed5ade6f85f749b674ff800f31d800acbdbde7b23db006ed2b3b976294d1c449941fb14c94140;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1346cd528552f8129382442938030bf851d2ef4b6cd51c177d85aa720ed1942f02235a5de299265d83654d08eb6d2a51b48a04a227e3be3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7d5d19bd8da29b74a28cef7baef26678e70ac2dd1eaee229389bb3fc63c2d4bfe0339d0f9eded71056ba5b0a286bc0f5d202a2bf6483f0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4d0c98c252228ffcdaa81ef4cfb5837d0d947fa6698c8d1bcffac4f1f4d758780367a3bc8393711e07ebb05a2c2c7b7f704cef6ae07f7a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b2fef0f1daee3d13178790a2265089fab1edc3759bcf97fe867750041a1233882a374c5a7037b4eaccd9b755d2eed495986522312ba75c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1673ff79bef76b4ff566783f1b6b8cd353e1b83187b59d7705740f4ed0eabef0a32dd8e9b1aab2eb6377885a3269f8871d4ed4afd528d01;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8dbc9c311d68c0c30cf8660986522239fff3fac6b2c42ca5d2e4d7409a3f83cfaf3e0f77b40504c5b2d24005d11d670b9f734d42f1261b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h115fd5afa9c33194d852fea7fd36fef9d5291ffe2f56f95e939af740ef9616baa4ffdc6032166c6cd32a4526eefb2636ff2f653217be980;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11af6fa29c521472aea9dce6aa6c22ac3865ef835c651c29a6239c6f3a2410e9b4db700badd574e0592abf223b7171d091c7c2d9036ec4d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he8e8694e5ef71068f365de045eae2cfe2aba296113e10c54ba51be16386240f4081d8116f62ad7c2211b0cbb2dcc19ddea4f6eab136b7b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h144fee9795700f84c47c59a3434bfd986feaebf65b2a58dc938c0e04177d0857da48b7946b0125dc0c7af71a281220da4d66ad0dc119f43;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8e923dfe85fa0847135eed8d68ed990469b12e6a59bcd05106ed9dbf8088b0356cc11ae64cbd9fe068bd11802e9608940fae3b8fe9ab6c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h67708c2463389eff07c9d96f751b6efb9521b877c6d1e87c2b77826ada59a1941e94d3256708d000dadf4d1357b2316173ba6f098e2b37;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dd945a620e4c2202d0b08d27b22005fce1b2f5a2c227374e396650f34d7e06986269141afdc6c347266ee878f15079f59803c072f4248;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11cb510a30ad77b8c95a686bbbd58b56866178c2ab22c2d276f3504a90df47c2b7313d6eb2260f06fb5ce0218fa6396427315ab834f1c92;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10d9162b45f319985a755c98d20bd5b2e48d02edfe55a9660303145dba1d24ea2a295109aea34370bca59376f0214af544e29e1273e3960;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16e42bfa2f55da49e3aa15a05a931caa73768a6c4a9fea779f2fb7d0eefdb14cfee0866ca06744973409d93704b92a7c942253fae4d338d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16c325a8ddd96c7aa9ff26f974fb9657aa449214010079fa17f026229c1c3a44628c30c4a585c83dbb2b411b935fbdebb35329fbf54e3f1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10c70f1684807c03c3ccf98c8eaf387108a5e9921129dd4eaaac32241d806aa51cbaed785074c0d96efbc9474f5a3cdaed5a263b4e8eec1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4d83a083054b10b2fbd361c67453c92c9bc021656951d7c16d67a25dc464a4a890176cda46c8d52f91cdee25e4f00a303c4e5ee30ee3c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6f8b2a2f00da829242a185b6494b4de3bf032e38447c027eb1780d24d9ad938fa949b309cef365520804db8399a9715569f8cc7d4f8559;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbae2291918981ddbc9a7a1b69aaab436fd614bc44eec088f89b2db6f4e90091760a7d3205e0360b5e8d594452a09f38d0032b389baf34b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h60399b976848939447cf80c0a3044cd6ebaacc5ff1f242c5b160bb3b061afbc8c519383324b574c648fbb7132948263f16f20482e68294;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1853761c4cb551f13a45f9c7c26b2494eb03425bc7ea8081803aecd567b5eafffecb07a53358dbe0038fd892bd42f9ec06f6810aa4b2a97;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1439590b8562f8d09bd1a224a620edb682ccc4e8116abc24aea3ab4e73659fc10b33221eec44533500289b49a045bf049fb32672ea9b654;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16e9e53a096af9e15a5a53f44ca7dcff164ce63bf114d4ea205db5465bef54ca189dd5d75a329707792574a025c9af811dcd26d3c345e13;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17d33864c77e103588f79bf0cfd9c098338deb11a4a9b8e05268f517d77d80456ddbe8d520abd2ae82e2686599ddcde5cbbd13f2d1e4c9b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8c516804d999a9ba3747d179868c92dfeea8bda6ed5ad4914c37ed037cfee6c68c8ef16bc9d9dca72349ec974622c7f2e5943f4a3105c2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1213e23f9939dbef2b413d79ffae35d8305f00b792100b45abc81c763b8d0451150a6754c5ffc03c52fa525e6c8d31c565c8eadce42c9eb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bb30876ad42dbd00cfc81140284c057436469c9e8e9128a7415dbc4a585cdd8771dcac57288e326755a0181da525c0ba17bd6c6f553ef6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h136a8d09977ad8ba02a8d53813bef028f71e50b1d9f1f0ffbadfed91096786fdde4e9eaa804f6a08117e458ae90e1bab86f33dbc3c2b884;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4019eb31f2b6bf6763c3a9d241aa25f79d81a26992f2ede06e71b00b47d1199952b5f8d572a0550ba0c9f950b344249ce84ea7955827cf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h47009e2321f7027bff053104314a983f229f3f29efff685a272e037ff86b601fa9a9486697bbf1f515e2d74ad436cbba3e429ad7dc7e24;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11d870873c0178d8a79c369abd5cd2515c0534429d02d7a2f28fe790e2526065a0983128cfe7b3e2f0ae89b6557f5efa2ad358d7d51f934;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h146b9a57e16d61ce173ce915f0f52e72a5ff90b438fc6263895a6355aacd28791ade9857b0305b32c81a5499f4879c347ba741acb2f826d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h34717ae04b0a6883d249bd9ead1a840ca29ea5073945af7da0cde9f3e969e7022b6b8ada457fc6661935186d80b25641c54f8397ab60a9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbaa2785515ee10f244ef5f05c77840a976a654109630fc1020c3606dc88c6dd4cad4f103ef226c05b3b98fc9d8878dc186d17f4cdff704;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cdd1f67297bf17b7da24e0d1bf6470dbf5e8c8886340b8f43ab7bb0041c7089639217d9008fed7a78a2abf95fb6a04cfbd8a0be2b67333;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h162f6dcddcea6a5012a3997c11242ba2556323d2f2d494cce69b1c5f98b5100a1a5a5c80d74373cc371a5c4a2cf6b1d1cbc9737f3fdc24;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hafc5a253589b559709a1a6a5522d260ca37b5200d39966c89741a978740aedb657b9e4a6da663b9eb2341d1bb3b145fa542d3a49a3eaf1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2915492a9fe5d353665a430bdb5ef4a0dbff3ed3ce3532078f0ed3b9ebd4b28b5d47e9672461822abd7a0c1ce8c980b45ee19e5918c2a0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d5ab68d00645c3e20f5df754a8b06225fe0236aa5355db12ce5de0694b1eb1179673f3166f3bf1dceabdf13b471cbd94c4c6a3e7ce85d5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h78f8618be5fafddec81b4212f74523810de62b521045e5900c85e20ec64f4812d32bdd3c29aa3319b3c451ee2200a03247ee922a9feaf9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bef9bfd070a619fba18dc4d6ac8dcba6e4de5231c699532c07bab36e52c2c489ed6097d7569e9a39555a7399e3075077e888b49bf1d794;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13cec40c3001731b9bfa4535908734f4681e17a62edd912041d8d9dd8b203284f0ccafcdd1b1a8f558bc4514cad5d0dca0dedb7638e7ec7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc9c30066fd2223d9e6851c4e41cba6a0f3ca571872b6bca40fc5376986ff9487c7cd8ff3d1a81ef1c55de0d4278977cd53c84dea533bb8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c76b4431f41b08d34c670913095494037856d64f3e33f245d1fd860da32addc63428e8c9c005cc053a06ead8731fd2d96569c4859e7652;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a7cbf07cb8439fffcc19716121c00dac9d8025421fb94c25e3cb093001187de67f93e939937f8b1d643817bc59c25c998f78aa6cbf8acc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd23980eeeb16a00a2b7b005efb49dc735537e85fbd36a4366edac199cc922c444607f00d080d0f1f3023e307f54da6dcf2dab1c609064;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h181c24348c6adff47390aa28bf71f4bf63ecdcbfca828341c4a80c1aeebf8e0eaf1507f38ec6dbf237890e376fdeb82127385c27735bd07;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h199c462eca6c485aa1fa7251dc0bdcb293af85294e5f2b1e5307e804a541a263a317449456103fa9cff656975e549d803f795187025856b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h345fc6d6895c653772f0a11f3e511a0dfd0a2ecb6af9e49da6890782a757e405e38be3dea9aaa49e0016eac1cd427e49628f3a33a2ad9a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10bce09eb7ffc2e87590f85c0b66812181b31e40797d0aa779d1ebef857283f73b4227ce303910adb6d0372fe85210560bc4b6f29d5cee9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5827a86ef4446f1c2a8eb990f22a4f9e03928c95fe05882029388ae69d57a46b38bb97496e7d7f0da14284191fbe942d8e5290aa09935e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf03c078d4479a6170ccd3ccb4acabf5a0f97fe955a7d2ee07e5e50a439424467f3549dccb828648d6ad501ff1b2feaaf04a75763538c3c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc2138a53b19f29c0cafe2584f4764b7f19c308a37350457eeb42471bdd6d164ccf8c3f844463f23d8d280f089c30b2da2cc07137c0e27f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h49c71c2e0a0c2acbb16f3fca8b2e3e479c72b227856828e805e4d601619d52057f258f85333610e7525b145465126c3ffe2c8904578081;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a827e7f50db6cedd4961d129c97244c99abf8991b27607c8b7dd8b08d13ed98c90b813e89c7629cb7900bc53b1912331e653d85454a615;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19fd0875e9454d1f0287a7b1ddc726f52c4e926cce4073e1bb6448ce4044d3f22416cc4fc0a787f7c52529f1d06503701078d5da6049864;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h85b2a44e46cd875bd0ebc78672ea929aa5db7e0db3fb1881c50261de46ef5f34af153450c4fe543ad38adc158b8fb0d7e1c645eb00814b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16f414dee8a908c3f8df93636089b460bfe69dbb4f32cf003fdfb6d156dd991259f84af7b5c83a9a70dfcc29fbcb21d91ddbeca33957e19;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf03bd20f99e239a0286045d6d074b9df42857cd43d0fddb889b641096d77fcd2c21a39c97dd59cc576967b4979248e4217da285f043c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18b0356df8c6ef45cb7a061e5d0b7a934734ea6369f005ec1243f5a848cf69f2956672cad554d9602366fe4287ec3b794614c2b46951d3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b3bfecda3ac1555585277e043244526c2a9af401e4c81b135e0fe0e63fcbbae9cb530c2a67a0da90195e2f301e50f8387124d94f9557ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10537541cf927665144d927f12090b8e4af136e7be3912707986a636407a1114035c7b5b4df64117cedc0be6fa3eb3e05eac7c199baa1d7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf8cf607141b4c38bec7226ec0936c85afd0b85a603893cba40fda2867916a9a55adf15126ddf6c87bfa049fb07f39f777eb1b6f1a77c2c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h30fa783f835a9f5a8f2989fe9dee84ba0f1db62ddacba693f8140a436db1a5ffefb7f00b19abaff8e0674ddc7f1370d09a821f9196787;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h184399cd2d55e4edda2e1d3cf71c12264fbdff6e8427c8d48355901cfb2bd744d3c0af6388e1b7f4e5822a6b17600d6f793d8c5e7fb0d4b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16b87ae90ceca245534b4bc8ce2fe2bfb5049a8192c1993140b92a952f05e769ab7e1d2efc91b5d57b8071ec25b19c3aebade207264ec13;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h974ea886af4ef628944ad41595b3ffd50c26e611ce2286f5abf1ad5e89d42cfe2b69dba4a036f8006c263bd36a6a9a2c9795a5b93ff860;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f09433f8510dc732296abeffd1c93f50af3da1f26d6b9b8ca12e501487826bb7e39f95f4d75802dbc57b438d0ff2e7497dd20540914d16;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h86a6f5ea7a1a58c4f7039f8f7562ed3f8d38cc8c0f2dbfc12943323cfd897820aa7ea4d01c686238094bd7465d0a7a93b3efc615b52663;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d10e3cd86e45fea1a947128073f84b339a6184f61c01231704ed9233c1a2c2b13d9fa64c279c35f9d32768f2ab186ad1a37f4e12ef9a02;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9209307ac5813401586c5cd8c274e1141bfbd9ea3d929dfb787ce010bcbea41f431a7535193917d186824f255e219ac012e4ced9e5e18f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h104e3646d44f3db925418f4286edef91c3a740f9a2ba9c1f88056c29e3c35b014f6920b5a52ef33a5bc844df2d7cd7fe38632a3f4c7fc84;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h75868b6118f0a22ddcd2edb3d6b527d0395f8d94b75a35751af266024ad592c94de1a6b264c536f8405b017de69e2c01cb25190356cdc0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h104d6c975fa996cce1912d014c66755d3054332f615a2a2b53c6b7042ddfdcb24392bce0fb4fb5da6df9e5b3d95373a60f1f442b8e39f66;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7880ad47ad01d81a60cf2b6978fdc65a6b0d839b976f182bd2e9e94b962a0e7b500ce9608523b010de788c179d537e0b2613e112bf9a02;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15de1a067039d49078ab44c906a9ee8e4f000320dfaf5769b7a8c7d63c3702b2e86e68e6456127a0db339af00069c07aa12c8fd874c2160;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dbc8b0c56a131912d2e44c87ef5f0eeb9a6dbb0e143f4c1f3a85561c3268f8770811129d5a251f29243c532b24a1c487cebed0a32c8b80;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h188634c9e30f38231b2b06dd063eda6f0a593a9d4fc379c923793cc4053a04efdbcfa8321b6370701d3910a16694320ff60a79f7616fd87;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h764564c081574c22dbb89ebb8fa30f04644f19ef6424ed70ab3e2331c105834067f18a1cc93dd2a46751c456128e456fa1ed3a727430bb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd794298aa066bec2299a9bf90c62fb55f5c9393a80467aa538aa75cf74fa0277a8743f2c3aa6a8b98c50b8dd869fb51c3b2ef7f6c8887f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he7e102275c4ca54ae04289daa07a63572d4faea7054b3cb9ab2f66ddab9097b45302b19413136b801dedd2b1a6baa7f1f51c236e964ca8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dc36e6061027887325e82ecbef9c6e1a04d59128ec3fe83c8f0f58946344764d558ee526987aa606e6828cfa078ab74f8f72cb51a1a8a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15c95cf295464e230aedd7c244cc28b3fdea9872ad31361b9db644595f7cf3ba1edac5b9bc6d0541ae0d2dc4b6f44b7f3588ebe187a07ac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e6090cfc6ffed21b55ddc06f79ff3565954a6481bff46b2089a33378ac7b34686079b37180a8a243d0159f9383b81d853106ae28ba53be;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ec211cebce4976a476337fad7b1f355d79f557c5c349924098b4965700fd2c930121af0fd0b8781684f53beaa137a09295f642b8a798f1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e358483ab9c09125ddf53e03008d3e7938b921f7a3987efb0895924a168d21e93cbb584be5eff341ad31571f8b9b6bb01b95a34b2d762f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f0ada68260f119b561078cb5d631009be6b68418b6406482b079984ce7db7fedc002a12af2898296947daef46986377fbf3f795e6e1834;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12b23f0ed43e08559a656f35114b79d249816503f99a1ecdd0e4ff094ee0ab6f3fbc13d56268a5c1f33cd6865b89b0b2096f98c60714fe3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b67bdefd881122e27859128453571f49b94ec3039b7c0c3f415c4dc35e59e463a016243910ac7c84922e0f8cbe6afa28f7e77a8380c8c4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10d637e03a51bef6e1e6ddef12799def17fa4d988cf5bc022eecc07c380c235ca90845036c3bee0fd4dddf1f10a68d98a8d23efecd483b5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1689205faa601b9fde083cde46927446d69326c2404a79a22888c0cdeaf0819f5b7f1ac6f66fd736c1af3ca9bb9d345d5e68bd1264ebd1d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h844f991c61bc49b1c00a23a0bd49f76e6a5f6d5baa05533d26045b47f3879706eaba3524a2a4ae3218ddb49ad7bc6a55b4d47ec8a36f8c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19a9a198e45862b5cc23d780ba7d03942f031d3a77cd22b9f02dc555d07008f4bf46d39f71b523d64277a09292da259806a988d9aebb7dc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19328245148339653f852fcb5b5aed08485bc4e4470ac6617373074255d4e24f8a349a758d3158d004b3871d63564a5aaa768d97480413f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h131214f43618a593af1eafa8fb9119b66a988edd29874caa3c3c4fc05bf4e89aa7caa952f1e324d7c86f44605a5dc25c8696bffe942abee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ea9854566e0ebe642ade7d34d94aabc570ca07d95f3d10f28949c3882c0bded4e9970923cce0eee95144dfc3fbd66ccc02799da41b09b2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1edf5012996680829631cd4775b6ce9345b8040601c10d02efd350413229b32e95ff75ad2091af125d2fd55c5d267844b3aed8a0cc1c33d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hab8c7a2400ad8f822ebf10b7711a05e157f6bbe7a9aa64d18dd6ee0c03e0b7f53e2cea27d73d7797148f4186dee91974b81cb6c9314780;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14688aca207020947146288666757fc2a2e78331783e445c32d6dc27ad78ab56fdccfbdcd0bc196350e1bf7049c1df7723858375c3d2cf1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hef6c31ddfea8540b722a78bbb116898b52c9119146046225d022f2ec5873abe15d292ed2ac681c58b6b1d344ef102ffe0f0fc2aa121af5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11dbcf47a1d4d85959cf769f6d63d98b2b5a810d0c23ac10914a648c840d3da7cecf6512af0b16fa2382478c83f445b8ebf31a0293e7c24;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h23abc584ec2dcfaf88a692ef2f34a30aaf50db3a8123397c98874c8d92cfe769afa8e738833dc57d4e5c467623c1cdfffe232c91b104a9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he9483bb998f30f5b31b42b60e0907736000fe2eb059130aa2d680c80d0ae725f929af1df610305407264be476455865ec2f4d3762e3ca9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1126d6b2a8d341ef55976bace2287cfa81eef32566fee5666ea940b9bda196903b7fd6dac46d00dd37c173e9b49511caf75766d018bbaba;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ad1dd8c236ff0db11b5c116dd0d3f3ac96f3e6920fcab8ebb118f45d59af9e2a1f6b6178e32ec5f0d11a9a9eeafbdcd2bc37267384d16e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7ee3bb7e38505f630609ed688e53c1dd14e346f30be0fa05832f4b052c1b0bf355d0f109dad2f66274be54366f9e0bd2eacfaed4af1317;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4f6e83e8d483a8549bec97b684f2941815eaaaf220489615f0c28a12c030f805d1bfadd921a3d28139439575aaf59cc217254430489dd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1899b8cf96577f7c99db42baf4e8137246df8de6e7172f5c6fba5da303c8e3141caa584ef9393a9ebe1865a26f3f43c73811e5ad55b4c49;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h194e16989b589bbbdd877e0a093bc3c15c5f6c8f67b61b9c5d8bc228d5c15e04ad3ab227dd289340cc5c4200203b62e24b26d3381667099;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b8b773c51fb4f4e196123c5ba667f53d90a10c8f25a5b96d6567c6de6de945ed0773c472d3efbbc2ebff769643158149e3db6d1d8ca8d1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e8ae9f13850b3fdea9aa74327232ef190e8f012c26edf7af820c7f9c8252b82bc5c7ce23f8c69b3527a176834278fc364f9db4df3700c2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d07f5c3de7d172fde242bfda0e4d163c807f0fde60193d719ddc967aefcb18f0d8899d2e0e4d32191df4c16314397e9ceb2537bb0ac00d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h61fdfd90a615de1d2c7f0d8343e12284fc0a60d5783c4e275876e76b27db53d7167b9bf0414eadafb4c2784141e24a9973f911774798e1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15f52ca7c5ebe219c29d0d4db99e9e2b1110d8ba0626a65fe9b68a065a2c2a723a7a700f806b231d0171e3bd34dd7f8a18ac64154007309;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dd8751da41789a9ae364aad206133c377935719e8b2f533c4c5024bf6b87fc76d9cb3e151230463281ee0201f16dc7709e6bfcc932c1dd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16d5e419ee3f8251b0f0dcc9ce8aa7e40aafc88c980f681fffc88c7ec8958ec92c3df993a7fb4be714aac3c4e95085732d7763c6e813c46;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8565f1a6a12e11b0347b17278951b67edc356d9e9320c231835b7fec9204e57f9272172fa105da3ed3316599669074f0ef99f44519d922;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1071944a6c0179eee7ad93a817a41123af6e911459302be2be884d13efe9876b9cf799787afd3fb5791e9c79a1fc57f1060bd72a09aa375;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h175e6e45fc414579f90c359d84101eb9e62d1d7f6961e239ee04a6004d052cf33e0db838ea398c1e91046424f1e5d446dee1167365633c1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10adf39a14aed06f018a1bc3b7ed58ac0d56a0c83a5ca0f187cdec8decadbe6c15754d03c3df42d12862d9ac44568c060e60dc1ed6cecd7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ade5c81178aed67824a290975b109835756f2a6644dddf312f9a3f02893975414ec0afd5ef26dcdf5915f61b4b458f396ee90d3a744c95;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c911bb6c545e4b7ed910cc393a2c4de4287cd8a0b749d85f48598fffe3b0c881faa7f579c95d68a0e17851eb639a032c9e5808ccc60e6c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2267ef316d2f126ace24dec28485bbc258178ab96628820df7c53fb572c6a3b00cbb65a35b4e5d38bf7b8e0ee17e4ee2fa352e48daef70;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ab75232790bdc54cb91ca06d1a86d6c8a9c5de71c9502df63946f7bb8e2cc16ccbeacb8331588d5afe22ce3722658c6696c8eba40120d0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbd480bd491a10c89e986b3b1096e879811b1448b8648b9f316681fb762cdd8cd655f979e368c267dd868036827582d594a6651b71302d0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e05aeeefacb2d402c0101263a0448a56fef24d8e3557d97fcae89a00f7d40063db454709a9b0dd44d30e4580b3db4dfa92aa78a22e7edd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1df85e90052eaa61584f160967e2392f82fbd643ff600418c58e4c60a8ffa47fbd6fba1abd123792da851bb221927d6d6e24b83338748b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h38106077513fe42a62df84a535466de2e07da99814b6fc0e1b3169157d1c8de56d3d2fb48a1f459fcd0dd0531fdb20c3290dbe74e1da65;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8c9ef5a5ac7a241e4d6991cd5497556bc0ddd61c3b79f7056ab7a57676efb33a997e81ccc23100da53ef0d5fa79b5531df245a2ec222d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h981ffc47541fa0b8926403d46924a6a0c6367872450eeb4af4197ac42b3414720ff4e67c1532f5eb3dab1911611e9f78eb964f81a5fa50;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1092a6dfce582e2e22ba4cd57a8f196ea341a841ec4855d4b35e1ee7210cac5de617c91f82884ddd2bc41be5183143d719cdd467e7b6ca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e133ab04a6a05fc41e5827901793a6f6b3d013b12a68de871c2522ba85caadc570fc7905c5bd897d09e89409db72a21b88beae1ecb2ed7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14eab3a82a3bd4e87165f1a8d0fef300869ae3df0eb9f51c0d8f807edbc02bcba75ff2ee24e6fe53f632c53748fc974b05bb7be388e1a3b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b812b58f222973b35b8f1553f9046c796e388ae957074404f377757a557a1426d4271f77f092cc9ae69c157023c202b52fa7814aa3ae1c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc450f7dd00ee833fbd0ce29ea638e0d50f92d35f01cee4f26d21801a787300afc9b9ceed4dae55b74ce2a52e0a4280177ba542663c3a7f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1955053f9e43eeee7b98973e6bb9754d4b499f35580c95c738de903159c863b6269fec791cbd4503547790fed9cac04f0d1ac1b84b63eb5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h112ec707d35db9cf836930c9e0f97b1f3e40a0df3b1951c0840025ac56216eaaa36a93b3d16d2e2ecd97db042636f3c31a98ccd96dd5feb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha2e607f29c63df815253bd539c1404683715589a6e8d2eee519a2645940bb570a0d3caad0376d25f3e7a2c97c151134200794a05706155;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he11faaacf2303bfe542457d977ff6dd44709d52db3eecb0f5f1ebead3e10999e4fac3d8354f93f08f457cd4c403eec007515e20df560d3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcbf3d1b8086ab6f07fb134d5af737a01e59c323b28b97e3582e69d4194691b2ad7554918b176b3b8c868728a0fcfb8e7f72bdbad78ebdf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e987a52832ccb000c13045cab0ae258e345089f58c94b4d5574d0aa82027ec0bace1896d4446664145b58a1ff4cc3109c90b6bd35886fd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12d640c62057fe2d0aacd40e947fef8113ac780a0c696af2a43606e289b2e9e84007e891f9ebbc6b61d29a66e94ad16f854e4af27ba1ffd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e10c6ea63a4fc214451819d120d6ffe761ac2024059aaf085eb21d6d86f5cb19597fd9041dfb0d1b05e4eb467d5e4c28dfdaa007e8e837;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h71a9ea20caca9dc801ae5857c403c9618a6f29c02422cf9ab75921d4796917934875efb768dee911b70c5cd2d7f3b64bc98e6cb764c907;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1663018c57010d5d45239109904ccc19a80f3dac94eb1eb32badb2321b21e0ac9405b639a1dfe720f66cd6a42ae07e7dc4e1fa018a80c2b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf519b26bba73f04095dbc8cec4ea5e5b88f49a6a6fa385abb47db9a575a5b571ba9be3cd9cf6815a22c186b09c923de4c38e9f2aba23a2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h470f44ec6d52a19e32d771466440a94d16fc7d999a5eaaa0e9059d1aa67d3c4ecfdcac882715ab0072ae11f142e381f505aeca573b1f8c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc0fcdf68c40ce911fa038defcd5996a0cd41747ad9287d1966a5a0466fb8453fae40a3533b630c0907574e934edf861d6b25161711bc81;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bc31708b2594caf126ac6e350a3cd2b69bb5c2a6554624d1888294ca9cabf4270a9752bbf0bf89bfe0292feff0d41b6148dcbbe398a1cb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b99322b5c515f599ac58532b926c8a843a58b2b581d62d73b65ff5a8058f27e6f4768e31dd9abb4f0d581d828576ae680e3ae9df5feb23;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc12cd05ff7703d8b97968f0a3c01c86d165f5c9890fdeb5ee146172b0f271a9563b12be7e2439a0b11a2ddc4d143d8b6cd4036eecb5117;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h936508cf6862837e83efc58ddb989d39068204e4a26e0d7501459363ac8e91e69abecbe6b48897a06f003de0ad0754f59c1429932b8014;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1aada2f5fc9a42e41b21192bb38d615102f20bf88def51017524aad298dd33f891ebbbc027cde7892c0245f6b39cf1cec0053cf960b7a49;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h74693672afb67c6a62c43f49f5bd5607f92b2d7bd38da07a464a2879578d97b290f88570b8ad61a7dd1f90c8d45f6c02a01fde2cf3060a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1669ba855299175188238610d3eabe07e1c96c6bac82702af39aca8c55635f00184245753e53ab444d75e58587200d715b716b999e5859b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h495a19e902e2efa8694f6a0dca73768d97e4780a03bb86327e400fbafb7c696759559a243a138eeff4ffc93b28d10e2535b54bfe98e8d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h977c419e6ba734f546344617bbc4354e00b53d2e698d3a3da4318b6046e4cbc78db72e00dffdd33adc39bef022b4c15c67454352c65cc6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d3209cfe0c64ebeff72a7b6f1bf1118e0879a35001c416ac5241324085346703d56aac4931e6ef71b347938d25d95790d615568f835f90;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h194cf63adf8348caed9635026e81c1be1fb89643e21ed82c9599d71208436a09c675ffa99db6b330a722f1eeec7f145fc4f404950e31c0b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1de11aa9212275cc336fd897c2990a7123c27c14b42708e6082ef1d77921367279a96330e3381b4110a0d598d7f5765afa40160be9a1bc9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e6dfbe0926e2c812b75a0ef3382c598f4c9ecd45a01bb4661f4d047f5da95e2eeee201c921cb746f7367d9b84987d62c2ed02da18a3d9d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc3f3f3f726ea1d9a389d16adb486416617796e0fb5ef0e415784bc6c41dd8770096f636298f6acb0571e7e12e66d67c54977e07b698faf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1767f9312bdc8304d100fad677c36e149d5959158a00c989a1a4f24fadac78b02a78e5c14b8bae6da919b2c8d25b9eb10ed4d86db49aa04;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e25776a68b3649e15a216da371e632c23778899d7277c2572208b1e1186369cc862f6d21c851bf89a33341e63c5bdd50dd7da27a7afe19;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h440b09247ce9d62434c259aa81229ba3ea0e7dbcbfcbef3b6e5e1f7baa1b11e9e7309bf3aa1827594a7aa811374ba173a49551092fe431;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h120b34f415c48f0e519276ab6ba6d8f693ab0cc26e224bf4c786772447e60f80deeeb98761c537b6f322daddab2fc013d839fab9ed90a11;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e66e9859ecf067fd55fb47ab4426f921b30d45d4a5c4cf431b1d6b1afe9fd0dd5259e6c98924c74ad22fb08a38759d34dccf5007306ee0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h88d1827fbb9de8b1a82d87def1a3624e84c001387d48b17bb8b41d738513c508348541efdb544aff2483b7d0fbc5f34811493288fb4950;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h342484f93b9c33433c4b3ed152fb1cdc7a0f1b6ee9933fa52700b47033ceaa81af3434712411280b529b52d4700143f5820ff7d066b5e9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd05dce23cc0d14eece3617e370c87d585e06db8158adf6ba6db869c27083c10cb6edfb40ac43145af43b90cedb8fc4ddbf75e3acbf035b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h203328a67b0ab9a63700ee6c3d5b39cf53c6715fb9a2d8539a568ab3ba437c52c0400ad5e111d8520b72e666306efd2834aa7c556db2a6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17452a4e4aaeb11276d7e54c2e33c6e05b9b433c20b3802200742e1e65db5fec8bc1120ad3231ab900aa92df488d452cff54bf35570b3c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17ea924684caff5c6a8e76a97d7db2984dd4b8a8aba771799dfec383301588fe763cb717bbab1069d519135f4200ee406f18f205b26ec13;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha7f184d340dbd1e5551a4bbe25684251eb37ea75c66a0919c76f31fa8f29fcf64bfd5b28767acd9f7752de605292afa0fc80601c42d14;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b911759d4478c2cc597014fc15318473e4084d9841b9ad6fbba76957cf30ef064671cb3fc5533e3a5cd122b41d7ecee1183dbf68f55395;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f3749611bb28937321502164b88d4b463f31de45deb548825419deb6277ea2a4e37dddb3e33588a4cb9f6ac68e4e83b95423b456ea2ce8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13608fbfd7b7be71fcfbd73ff0f37c30e7e9b1e1cbc07114c65b7beceac65ad687dd24859c4eeaf0e881d1184be1a7091925ce262267e55;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1305d0364ac228eb5e12f69bb93efdb12927642dac309ea007f5d7474b26442877700609560715cb571c6b0a0a6c1910460cafde0a0ca90;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17fc1278ae20e5ef5cfaa61477e4aa1e9af34f95c5cc0f9c3aefdbc57b0c57ef14e71b463e797e8b4a6020ae523732c2709b1b4113b93d9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3831a333e8a0e5e31dfeb8e770b377838bfd608abef543418e0d707a75672592c410de7318eff6db97a1d0a283095120011d69ecb3cfe3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h26c1a6dea5bd80045cf1cb18ca82bfcda9c416944302875b9fc4ac05fe830c3ec4d58ab41a17983d2741bebfdc3a191d6e5128dcd6c3bc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1080abd6a2a95f6c113291b27a7c940fea532751fb04eaff0f521fef1a5083346693aed255f1d039e979417ded5621e01794bdfc93064ad;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd11d23df3d831c04aeb164d73902a7865e80a83845b5971f55ddba3a85bd66c7a42b64a869933b856c13ee0e3f660debc8b50fde9582de;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hde094755e4cece12a2f32fccd1b8502c4547d078d8d062594b8d976f00df007e4d51c2a6e66ca97130529486ab9282801d0ae0d255fe68;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4b73bf493939fcad8a2ac262ce5e448d175a2dc2ce2ad7f0ad8d8461aac8246fccb8c3baaa82f8aa8025c6769c3ca879161048f29fb2ec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15f4fd791fac8c149c2289b11850005905a8deee1e1ee482cd07c9dd3b16ec51670580ea9385d1b859ea442db062628092c68c56e48eafa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h611cc3bb6ac058c469edb5a896e4e1e5f013aee9edb0c171d1ffa873e9d43f197a6bb54798849421ec9a67197e92eeb64ff2050d69a11b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h187948efaedb283cd1591b7809625778aa7e089d8b571a31c4d4a370650ef7954aca2a3859d75c6f44733fd0c216ad5ad7dac86035f6be6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h852773831595ffa0c2fcfac15af2f1dd4d901d1a081a31657b05d3fb03f4ebf5bb1ee31aeda6c6d9d7c90450ef3a4695be044670c8f9dc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10600e310c6ef22cf6d74fd0026dd3f253a91de849929bb077f2af9bd90db625eb13e727a13d0fb2a5bcc5adfe534af7946f0e13029115d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h62966e9ffc0bf0092d32a148455bff8c62796cf6cbe968f5b4f3e8f14c300d1f661d125f0472cc5e5e108f734dc5978edb349059a0db7a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10880b1bfb4cade4cbb9c7cc664b904de262a324bffeab9c41d2cfa2126476aa3c5b97fdcb45c85a61cef2dfde06f6c7cd366ad7035f894;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h118284e456719478b8d06182d43a0899ff9d5baa27b842ff947d29eb1a5fb90c1fb7dc00a28dd9c9bf8f518ee3eb4f71f3eb3be255b4c9c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4702f537aaf581806f05af9c68f2c98f4cf603524279d6e097303587320e3da0699f61bf7c8ff9473aac373f1eee031894127bc69ad899;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18d2fef58948e525556c20c47479df44f17eef19d50015b7a3a47154b3bad49132b9b2a98861a4fbc65d13aba708b56c06b0a12d5be38a6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h206f5649adbef9671b7663834e6d5f73701a3be4efaeffb509724c53b0dfd03deab1bddc15ff4679eea19aa1e465845c86d7476eea612e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he17ed2e55c1a937d633868a47c505302a5795bee851c2782069ef3b2018517f55bed3094cf60907724ce747ba6e2a4bf286abde8f7815f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2b87b48f9d1067b1e1cb697b7dc9665d3762516e5fab048366173f9118beb86159b08454fcf33bfca56174eb566841aad0783cfa73837d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6af1fc1dbda891065c5426499e8fe6223179ca2b3968afe0bbbec353d70edb3ab3cffae90e2bca2f39630c84ee9248cff797796b7ff164;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h59ef85c239b9f78705379e624bd308cdb090108cb7a60f4e84030f20dd92ff339c06231196d1ee7667b3b17ff53657c61cb58cd2ae8440;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6157ff4f46e4a7ffde7e072921c35dd84131e27683c09e1920d1e63403f2f29cc9d4fba059517f813d1a71aa3af6318c6d70e358e1d921;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h651b580836274a8f11819fc535809926d16c91f71a33ffe55cd2517fc9665e986dd87d7c0ca3ebf79acf123e3280d7ffc04a19d38eca2b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h93d94921b8e08c65ff3e5a6e9773a566b7010093e7760213dc97e1d8473b01977e294f8cbf7a1ff3e1438855e3b1e25f341c91443d3958;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c6af39d46662a0478bfe62b48e47e5d62ac0f02a314adf0956c86e4841cd20d8bee9e8541efce1af573bd244aeec9ca505c79072be5ad4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1329bde7fdeb9a6384c2ede4462faed5698be81980d562744e24b23c8519558c5e6e8c3887e43dcf7b0d613ecf79b388c704edf13edd129;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1290feb1ffe136c31fa3dc36c8845b93792d47e4eb6cfc051a35ade9e9b98aaddf79422617883b91650f804a98969051e689d65793e688;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha030bbf5d30aeced7d221d2eef71dc6aabd68a4b62022d1d8515f94d372745ae07e50c17a3040c44be81382ba53f6390836d53b6710870;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16e5ed545bf4272bb09758fdde6e1c70bc499f7592d1178c66a19345e9b64d40476952ecde31d6dd4f48f10085bc4259b0ae4f3dbaa00d5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h763aab8d3075c6e57b30209e0dbd8a9b4ba512897b4edd820d359c2039d997c9c916cc2554713c804978d358bfcc49a5e8c0e678595cce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2da96f3c23133a2f84a366e68c6582e75f40aee13bc7ea983af11f1bb72b97b3d33d25c9a724a6f20803f5a6d48d28bd17169ba013c05e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2772cc32d8a98bdd83d205ebcb170921588426fe5abd9f86ee27de6b828473a87ffc407b62a345069ba6079f228e3db648c819f7afdbe4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd24613795bd0e877f8f6fc65cd025a0534d42f9ea1307946fec8b97462b871f092a6141614f40ede05a66b5c3b67002300e6bcc2e7dbf1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15ca63e932030f48df7f034202eae25f87c004d62e45dd607267737add73469528a5494699eb8921fe002c671476ccc8a0498804c4b36c3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13569b17e9ac354b29e4dc29e6d9809802ca32f8ca02c4082b1f8fa0e3226feb358de0be377f88c2d3e91c0490a1cc0555606f143493082;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h137f424e466f1c0ecfb99a073027de1288b2f16f0b8d97ea4403a7b4704ae0063ec1d4b893dcfac5eb75e949daca1fef19b574ccea11ec4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ac02f245a685bc5aa9d2d1613997bc015d2b2c336315cd086f4becc4d11462d0b19b748de871516c6d78b2d95e2fdf6b60f758040dffe6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h97ecc65cbddf8171e62abce815da6efe39d1731489da71f7eb79d5667fbeb50564839f308831c99555f80a85cad713299b9eb111900259;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he3137d29443e61be6491e4eec22c371851f5e8757ea4e5ceb6c829675a4c1d35f662760b346f622c001ba75b5be8fb1ce52c6a4db3f4c2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7f286786129c2d35b1f93c247e030327a5a5ac66959f8dbeaed366b00b17d44e9c45cbb1008f62b94d8a4ba2de5cddec953ff4407a53b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fc410bae3d925f218a2d20a5b3b567cb84a0386a3fc594e3d103d92fb18c500eb5caba0ae2ede200828b8946a06fac108955a5547a52b7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf01f75d2f9d584b9a7a3fedaf7afd40beb9c4d5584409982ad0ae8d28d6dfb71fa84fd0c5215476638269e7b0b8d65f4426b81397b1572;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h124b0ad9774203c7fe7cf194a569b72b3d0aa37e37816d9486ce87189c3bc92608643f56d0c4b2b37f87bf0ba8c427cb84d812d7fd3425a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h133bd61c34b0645021d5444a86cbbe0e5f137b9e1e400e8f266e3c12305f40896905b36ed745fbc64b3be0839b8e12a9c078ac6f26b7a16;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1600a3980d789ba521812ea35b891bedb3f25708e886c6e26d5aebb4db528167af564fc82ca745c25ea0009b75304a9dd0db74105c9a540;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ac7ea557c969f391cdb9b49508409d9ab675f0f37d05f36b78f200c1eca81ed30400dbf66307adb8176ed8b4c55ba68a7a9a76e0be0433;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fe714a34c3d14a3b3522091289aeede5fceae42eb321136fa9e82a2ceedecbb14b32b2934d1eec5475126f9d7a4c0b3e2dc15e41f8f324;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fad604dac12ab0d92572448cfdfc20228f32f973051dcb8520a429e8f9975ed05c8e87e2f556b8c4de5643336ffafeac36df2cdeb52a94;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb752fd624a00043fb2bb250ec451f61745b6481bfd5f951630a29710a8fa08b727352e3cf24e990b409031bed517d92143c58b4688d2b7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb766305dd094a48f39fec43afa280440ca4acdf7a38eafc9a28a337d7add0e5c356e9e1686f62c5caba7f3e225cff7588f63b3c5b61384;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb290af76d78c6737d3b62088b9e5369fe03695a320bd78d7ca7c6dd1d34600e410d6454d776a896a5daf447aa89e9bf0583552a3a48e36;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h42d8c0a4b22bb5fe39699f67f822386aeacbc3adb677aeb774dd03e1f557590e8309dce1181b1900a97c3ffe3bec6a01511aaf2b506879;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1406c53d14fb86460ea764f2eafa66dd560f578c79e4cc35393e054fdd7ab0df07a90f725e3dcbb01055a79a4bed09b5de0c9fa6a82c8f5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19782040775c4ba4393efc52bc4ad67d8c21752e12402407c5462208f3aa754cb90d89d4dfb97384d0ec3cf6646a576521a3009318a09a6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1154f3f9927be89cf71f077fd8b8fac9132d5e4b3e10c41b5a2edfe68f736ca6cf1de52b7d0b36344033f8601b9d70b747369ed7be9b022;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h601b6691e1015af73347ed2658f2a41223cad31b9728688b2b9ef1f8787b502c1f1fc2bb4ae04253a7ff9f8a4f4d9aa2cc044e93f85240;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc0caf0fb2e2dcdd1fff7d9d733f1d635dc8dafe65c13b766dbb0e9c71336c72a1aadbabb6ebdd473c60d89d34e262d05ab4f10f057aac2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11d503d22ca2ca8e0017798cc8123ee043ecaa0c9c61e03f31c2aabfcbf4870bbb7b1f27ab3ba8646e71f44224f282309b036f73c447718;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he6ad7077bea13b6de611fd86c1d308958bec242eccd05ee646bb63c717f9b4f7e121a6022e1762fd04e8159b667815f88c5d2e0576016a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18addf79d45d789ad3055bd3508bc14d3ffdabee1759d7dfc1fbc5ec41ecbd6dd05d4c64ed2512b319c4225cceee747dab5acaf14585438;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ed9b32dcba5f08c2551396605df5984f809f46cd46aa94b5aeed49a3879b02543f7942c0590f7397e8b5406bab06193aac615391571f4e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2a7f51ab1ca81d4162013c2dae3991733cd992b81dc083d57c3f5965e40676bf5eb345d535e0a7f84beb96cb37c8b0e25382d2987cda80;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19c109616526e34ac8fd46a21ed7431c86b5cf52269a234dfe6618e7024ec293d6ad30c578e2d25478201f5531a8363dfe9375457017a7b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17c8e227cf0cfd1e6e5ac1a049dcab37c0cf6ada88dac21be7f70d73e3abecb8379515076a880af06901fb1bfb342164081c67a5614b528;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1516e03d126eecb5a36c379546f4e050813edd423ea902d1f2d8313574f154fa0a4e8d519a3b788eb74c5121aed63cae17160dd7882f69;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha87b4a62f6bdb1cf8889d99f16510783756f3e2cc2640a0f946ae56e1e8bbddb925dc075fd053ed3ff0b157fce31d4417d496f042e267e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h91297758da779e15a341084f3924eb7670bb3e236e996450d2623de4770e41ce7b80a0cdf43e5d67b6d9f28b9ae0d1ba00ae0df9c4075b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16127ea1d43478ef271cebf1b4c99a68dd61de6af503088664e05cb7a78cabddd807174a6b2ee492d1450564d8fb0c905a99add5947545d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1db537d6ca5bd871c9837f6ba93a096cc3d557e397b0d9575de4db1ef6a4270f32b35800c9736c2914ad83bb513ac78b199e51db155d00d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc04ace1ffa7f98be8489791524d7c90eba468642417d2e44580b9071f57eca1cdeb4d12e2b770b97f16b1d7b5abdcb678f24088aad6d36;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f69e2b51607966abccba0f95e0e663957733baa19861ee3bbcf1a3cf78caccddcb156b36a5128461c1da5849fb9ea3171d719dacb5fabe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14298215f847f105f7ee74b8fa2ff8e5057b12968505ea15a45bf1a68dc4b462e4a6041988a2bcfd12aeeeb4e8cf3852e6351e7578f6acf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b9c7b9607939c78f5e078b6a75c12fd1ea6143e5c5ce3d369428ca3f7b3afe37e12c87676ed5bbfa7c28f357e876b85232b12ca57fcf76;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17211eb81eccbbb5f73c03b33f69d4eb9ae2c69b45992ba3e064db22d26e7f9926b5e3f336508d3efcf7d9dec5534e7bbe50938aac5d5a0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1de3e595b493ef4f6ae04bba4087bb2a0ad53339b4e1445467df215180c112db25f489ca046d3e2e6edf5a46e704f18639b755635b25b29;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19a0ac3f7761dd0061e329cdbb6ab40db22d6143b1c2627e9cbf6752d8f5f86c5e29d4c6d179b686231115815fcf5f3d3679a04e5371b5a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h94ffd8b52b1b65ba43927d4b02028dd69c6826e7487e0c9250a0618963dc6d3da7141d77f159646e5cea5ad6adff53202a41884d635d11;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h22598e94ddaac29d7adb6ff1b61f2bd6e3e561b74f080e56bbbd1a48a82f4af35938724fc2ebe6ea5f8bac2585c1d9fa53c80cf8bad1d8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f81b05597cc178f06a0fa8a17283cea70d55ad0b945aebdf4324e860ab8aa9033a6e79b7fb2be4ee840889572b092023a9ecae4cfa326f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h728c06c8c8abae0e34305f9b144008b5b35d80e70dfa1a4a57d39d80b5045a47d774d9f5dcd36e1c2a27ea05640f066a893d8a335a9ce7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15915fb7ba4d2d6c406a13199dcc5d5b31ba50974bd0f826764a676fcc1b6cb367c6e400163bcf70150a2dd6ae9f80808e8caa30a31bcd7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14b53d46cec62924f65819667cda3c3322ae2a8bce6fc4b8e0409dfa4b5f812e59920d61d38b758195eba0b5317f5bd5a3964eb944dc6a6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f24ab74de7f14763623d712fc7a97727ce71311bb2f7c43dfb99885174ff30a464f5040476e349a016d0e5ec4af84b6214dadb7b4ddfcf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h183a0ea924e0ebad552269220c9eae3a04834cee2d509ec133aed5e77338777ef54f634b889f15fbaaa641d9473f88cfb888159fea9f7ad;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fdd16744aa52bd741779e7ca594884b2cd5ab3773b9d2d7023b9ab3875883bad01c9ee9288677cb3cfcdc766e2c3ac82e0febcdb872e17;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d247765452d6322423050e557df88e608512c59c11dcb7071f7d6eee9171428752147fe6735cbb7e5caed7e809c215076364dcd3b8ae7b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h75ec3ffa73c0a9e9d3af9524b655f33b589ebb546af025cb7298760b24f754535eb724b43e41e2eedf9df819b715c81802517fb65400e0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16c359d52e118e173482b4ba74bb39fd8c04d36ad7c5d338fcfb2649afe8d6a345c5e24b6e5a80dd1134baeaca216ecafe3789fce26b39b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h799d5c5cc6a561ab15174ed0c11d053990f4f26fc5d1bba314d7a4b1c83e4da4853043fe34ef9fb342c644e6198f8ee52a6215842fb37a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h711900817731e4602d03a85d29e5cff16b2fbb9c087b3e05caac6652ab2232d4a163a33ac093a84040a7bae4c422e79861e37141babe59;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h170852ab4ffda419725335f17084f0b4636d9334f6c7a4c4b8a874dd77a285ecd57183313234919838cc14c584066fb1003909168af9037;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b12637c546cb2eab2edd2ef398f9b0c89ac336dc883524e1ede08d6660e809a709d23410ace1a8be1d96febe0c1a2cc897b7cb6825ee2a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h29961a4d3b39d9bc29bff053d5d76c2e89758ab9e008afb88d7cc3b8266a1af5a63753d0215b629fab79773f58a9513f22902beac1ace1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he91bc6da1c00e14940a06807db2fb54d74a3b4675c77d7ce9fb1605376679edbb03651051947a5bde90d7fc2549a8c778ad0d279ebebf6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e43cce0e4194fb232afd08b0abb48634aa766d00d09cac1739144fb005bc2fef345237fbc1ae4e7d3a647224b646538c9599d4bfa941e4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcc3f3c24941e8620d0f2bd14082ea40adf83c50b21b6cd2e49514f03a80abfe9ec8e074b2618d2296d1b610ff884b07e2e46c2f136ef9e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbdfda3543d59cbd029d0d41edb63e9c2f8a08319fb7083516c8f680961fb397e63cd0cafbd9810e5295356c9987db481f783426dbc5073;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcd9af1628c99877af563b8494ca9c1b7b210360eca8fe1000752320969fa8768afd1543196ae7681125f2381707159d666e4565f45f2ca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12c42d68094196ac2cc83bc4829141e2dbceb8d71143d0d85a80ef91472cd4dfb627f75c7470d448e607b5bb6031cd4467a922b44ec2bae;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h175bde1339013f82acb152f2dbab849943b8854ef9ecc3ae68d6d3b88851a463443474684daef054e49762e081275ffb483dafd3cdb767f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h74935d1feb9c2447fddec1b9bbe94911a3e4843a8ecaf031e7e767258c5b70045ce96148b263305cd8508ad1a452214c5ef618ea51bf11;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h62b6d421e855382c749471e169460fe5f1354f5ee8820a178355bff14336a817e27b055ae39fe599cb6e3e5def3a99e7a33ad0563c9ab;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h71d2adf5a0a43f8dd478a40e7401a2be0529342cf482f195a8abd51dd748d5f87683a94e78d91d997802b4b5325685f722f726aa2ac01a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h133f7bd172c2490d581940aa65b36e8e2591c2e6a01a818eadb62a4c21e2505f5748e08cd0e285ca407403b7598869ba2bb2e68a114a0d7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he0573ad2f9e869a2397a8ea6e7fc042f4cc619cc1cc1d10733e12734aa3249e2c31cbb8abdb81b3be9fa96ad37a22abd76ffdeeb26fb55;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf109b41e38a453f5d30044d08e226092e0c98907d8be26969af772e9b7a852883c079eefad12c3b4851922b0a4f59ce40697f5627a50fe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2884b93bdfb8f6d59b466e381c14b4310bd961d388853baac56b51a4d81ef15908545e27a3ab47636962ffcefc5a8516e5b409e8ddb1c9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h191ba8796ee8a0a4d0677a5b4915763150a6245ca72e95876561aaae58e5bc115fa22b50987b44c9665ffdca5f9e076e3c1d90ec01d1919;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8c8a1dc590a5966dc658cbe2b77d52279b5840431cd164aad15cc2fb57f5482fe5db9a66cae7684e3cccb12c68752d9d90b7d7c6f6d6aa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h560c372c41a4fda646a815e9c13da55fa549f12d6451b1c1c9c8ed0688a58178921dd7605f29453b2dd47b7fe593aeb5afc65a8bf75013;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf8bf602a51c69be3fcfa78eef5874f1bd0090b723a220b64f16aae02d8c34b2d232876317f0e56b7a3a80f5318b033a7ee063e221ed620;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10829e2532db9fb45ba922e58d0abde7d5dfdd51b662199a552990c41e2bdd0b062cfb02755c877c1c2f673d40db6ecfc8e5f52a36f46dd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17138f52f874ab591261829d935f62b84d8443bd9d4f9512e8c78430eed28c66d10916c1a5810080391707430fea4bb552c7a4b769e55fc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h61dcb16b7652c96f3ebd92bc75eb1714bd8760964e6c0a70a25206f8c18d2725bc2fb61a7da86026c639a28e0ac00c324ab6607f594d74;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11746e21080bff3eea7da1181ab5812cefcd6d7093ee7fc24d340710bb4e7221b21db03c8f8a59acd47cfa7226b28126e09f5ad0c59130c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf8c86fca6b89fd862ce4866bb9bbf6b80f3773562b0aaa919648cf75aa69cec310efc264511c6d5da71de3fb0f2435b82c8df9d148a74b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a698cb3e903d7723a20f970d76fdda9b085f273f9ba62539aa6e8a7e7bde55b432cae8a99478a4956187acd59774935d7f96b9ab55137f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c3f8c6dca3a8a32851afe1b6622f86484bfc0af65ba8ceb5b1124857f619a42091a9327cca7ab9c2f994e5a92d281c7329165a2cead8ea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bb1404ca2b7996757226796ed668616af427a1bfc8bd31b15e6cceed53a8298e5285fce6ffa4e3e20b6fe6dde23bb3bd4b2c902244c440;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1da07594e4cecd8b8a16f52de30b8844038133ed720ec235cbf546d9240456cd5a4f1f4588611efde288c0093bd7b3174cd39044267c18;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hee024a0977546b5293c1ee095169e139506caa5c5e4eac3d52c687696273b33dd642dbaa806e901af249bcedb00d025142dfe4183a105c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h33babc0644c989271ce9ace382a776d092714ed9a2e0cc99b8643b497c5615093f0047c5dac1c448717c5391a672f9fd0f74bfaa8c7101;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hca6544bc93b914f7def4e6e7351a8329b9deb2083d8bb3e24ccd583ce0fe16a08c0b920c87521b913488f70311df56833d9f312ab1af9d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3768c1164be9a132e895eefc58976626e2b5c5da542f6e210ac4e2658b99e2947d044e8295d45bf7d6be44dac5f42672269d8db72266ec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbd650ee855209c2719e4f52ce28a7e4ee9a5978e4e631953166cebcd754b34a3477ba5c6beb31cb877f297c97cfbbdc8576de5d4a6cba1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hebc24fb5dae7603e4b425d7191625b9fd653b1c0f725f31d6c0fe6d75989db973c23367246c499b3ea118254b28e79ac80af7c49991c85;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13ba61880e9332eaa37defdb1df2453faf3051ce3b020cb6e0c98babfa67850c5ac2876146bb0b12376bed4e40443ae466b82bd861b5c83;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1596b31e99b36c201256ccde4b58ea81be67525fda3a5e4bf41305dc4c8118f677a11f6130ed69af0707d31f34835efebf531dc153ae1d0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbad420a206a99672e89096d6571a1452d5c19d0c2e4fa3693004b9f46991ff8b13d065446829089ac9781562a5e32b330aae2723ea2b9f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19d91beafc6b28457856201f8a0e74eb2f527cd78635ab22899494e574bde5ea18df0450fbd69d14ade4af6bfdbcdcafc70a917a82806cf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18cb5788031c8859f06e94203bacf69dc259d7fc7df814855e2d46e73834d9eeac27eb2e9bab25a90f3585bed61cd62dc6d34486d082660;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd0a7a152445d5b5ba10a03d67739ff3cf14636a900fbc3d4ab50023b67f52d424b2fb8c24ffb7f26d81e4400f8cfd0fab5f04d3db1dc21;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h126a82df76572fa58a1a20910664098ac7e9a966c66bd50d082815bae890bf69c1f173296cf030099a0e4bca122284b6f38e4fd11e8241;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d17152b2db9d36a4f9bf5404fb8223fc70f4d1aea5dc41dfc20950480b2f8d1aaeefdbf713fe18f30b5757ea460f4eb59724faf66768be;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7c3399a2bcfc66eb66ee30deb301fb9ada9bd34bfae6c94e7731877e543234612224003ed1833d274d0ee8e1d2af4d548d284a6fb32454;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h122ed89cf91124a3d41626df29a55881fadcf6f10978c590dba924020616baafc2b6383b3fa1dea00c0ba52e42ea294b3c375cc2e4140b5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1805f8dbccb7c00766cbc86543bff7a0507b12b6ea8c748ad91a0eaa3f567eb3f1b866922d06a8b2db32070f03428b576cc8da5983b95c8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d70aa43c09338e69c1c8e860bba7deedfda9c863c8b55fbda71b1337c2abbc9c03edd0e59ce1031a94818c2b4527be23f30839beceb4f9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h104da13c6bb291ebfce97adb5b22453da4da66acc15e5faf8f1b5a19042111c406c382c2240b09671efcf297459ad18fe704c04fe2a3024;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb268ef070fca6e5afd90f4e21461c458b723fe4a3445c624dc6a649668e0f2aeb551cd2acf5f5bbf9539872c6adbee67928beb68f3b854;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h131a6abd15a008c2f03f65315ea47d2d81d059e4f919caa693ba6d04e5057174af498057caa6b40bb12992ddaef2ad5589ce03a9ab33bb0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf81b3c267f448eb8894418708daa71d7f3640dd16069bdce9abc52ba4d4883fd82efdd0feb4f21a6899a9e7c164087edfe1d346d04bbf1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10b6ab2b4faf9f52799746ca634869feafaf900a6eb48ef49fa595ce1ba36302ddbe3f4c0e772e0ba37f32431ad5de9f63dc803d5f44f5b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1714e25cc50739adfc17bc49fa1c872f93b19755a5430004c7181d34268518dba93e023074f964a4191f888dc5a5c10257cf12b5218ef34;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12805da425d4e5151a744cdebcae2bf2b5f56faf60475b95be2c8cce89bcad18003b5e1436c2aa4b998fddd2e5895e2880ab493db32f7b9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h486cbf107a5f45327310e182f138441b08ef0d777e2e40752934efb1dd705743d6dd80da3f51155dd8f90858c7acbbccc5c95429b59fdc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a3514bb16a41f05443ee64c703d18619364cd12c37455e7244fd318335b48a1e465119a226ea4c2496f206506a9b09e333e381ea24f686;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdaf3061b29a2bbc6a7780915768cc5637d29ac035c9b0b07b8775e589888911a9ec7ccbdcec16ec6aef069422db0a8edd7211cf339bc8c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h164bd236f1935d162785fd2a20551bdc5e668cacf464b1f6dec0b6c3f0601aaeb77905dbdb6da3ee66c6ce2d10b51025512148238e13c8a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fbad27314545cbd411bd97acca2894deca2640dacda782f909b4ee505fe72b045819be9e4e86cd7808c9a2ac628bf995f8faa404e85162;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cfc5e7cdd23993c949cab5541af91ba3d31f4fa3dddd536091bf8bccbe1bf130bb61934bf78be72067bbcf6fa09e17a34d6b103e9b2c24;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1390b4ed8d3d3a0e48f4dc1b62fafd31590f96c20d1f098db9ed5f2ff2b99de9672707754699d823dcf9bc688f3ba61596a6ef71ab18edb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h171f2c7f77753dcbf064492b8f7e87e6e9ed46dfe35174aff51202fd51ae45e6955eec4abda8e0c86720e6e2a2b46fed2a023ac23d61674;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a91e67e8d98f2fecf8746d2e625cbd3aed59692138d9715976e35da721a8aa60f380a64820e1c27ed77f22e92f89a9665b849290ea26c5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h36f465347fb230c3a8669a705b93252360804de62a432621f9c7d336a7c1609110cc42984d1e34462c9ca29e56026051cbb018ce127656;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h60b68dc189d9979eeec58a18d17b05cb2b30ce2e04f7b34243064773d08fc4a805c5f29e1e88771b2ea0b36a35df35d65d574d0255e329;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h66f17033b0d2b5d9f61cb7ea3ab907598567939935c75549c8489b66c6b50665e8cce22ce3d9d5745605a339273037b915dc9161223d3b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fe79829ec1a7b1a81c5ec4be2a7d6bf43b80f0961248a2e4b18174bf87d22503dddaf6ad1b26044f3214a2b8e4b46a88d78794d8366fb7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdb44ad26f72e3a459b4b27f5e04d18cfa69678d05ec5ae3c6e0f3d5beb01b22f6e0fb0361c4a7b165493ca7520732f93dfca7f849747f5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13c8e0ca223a039c0fee74f20004df86ad9d7da4ba47b7914b365807ad2917a63c16d0d0a120e51b912da468d2602e272f05b7241395fae;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18be33c3f7dd528f66a695093175359e9db11aff147a543db283875a579dc6f651c07659553ff62fa31c92af36324ab3024381c9dbbf20;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1856f27abe47901f94082f8400330f075f2f669584418e31522ceb370f6011eafa3b6dd6648bb04f9d2df680af785d6b64fce25acd10cb2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h104f1bbfaa4aeea8143fe40829c55e7c064be2915a8e22d63abd49c9160997eb902f9f61c7c3e64d189a90914699a0dc8cbe01cfcc214ed;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12bd75c75b471fb8478ec43715c5a92a7e1ee02601a866c8f9633820ad281adf8ca94318fd4b39a1f0b630b60a12adf02fb155e2a0e8af8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h168187cbaf19372f9099ea36da9b28d8a5541e91589cb44519253d135bea037a7698d931528cd0993c6785c8b680bbe125eb4a05ffc5107;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b5ce13f679e8763b992dab6ee4882e515b566425c9b0976b5a4157fdc0419dcefa7cd094a378717f6abe23d3d4864d7728ab69ec333123;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2987bde654b75e7b624093ebdf13d9073ac325d9e62e8866ae6138aa6f3af3b57add78c471a094677f5d32a0f19934b3a8d3e99c2cca81;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7128c457e53a4dde4fca39afa51bdb33b5c07311c66d94c464d996922c6d74520ca2e8c8a4832d0e384898172eda439a422fa803e0f893;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4059c307cb9b5bd16f68fc97c35e2349a2b6283fb9dcc88a3c019ed5fae0aad6cac5c3cb6a9c185581cbdcaf2afab5ce8fabc62ea25063;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12c17ae9a1d1a7f2664698157b0cd1e5a01deed38bc04c7ca0d8bda2a6e550856368fca751aa0737d1063944f9d0956d626f0dae1e0e960;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3f1de0cd32b9a728cdba0a014116aae023a568f8411d6a21908a04be9d56d4919840c9e05eb6d475196ec7b0130dc98029fab480689469;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14b357803d2aecd84081d65789184ae8f757c5b51e567e50a788e3ca13f03e2e55e9d7189323cb2ab78f4864284aa080d9be47e71bdb7a5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6a45e58603e5808534da6e746748ffd3efb584916fb504550724f979f9659fa66a1c4de1a16deca9563fe3a0d00cd9dc0860926673b019;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14acf95a7f40fb3af5e592bb7c94feb249b0f23eeb3fa86e31cde1eddaedb4d4138353cf818df1dfb88e1e1306baeffcc0d8ed297f4449f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1286bd0f58e9f3ada7fe5afcd801de95468ecfca13e11621ec564d8f12ca71f7243d7df50cfb3abc466aac40ed7fd9231e330df53f37590;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3e45d46beebbd81b838812433d66648608fdf8f3acd36c5d092c885ffd95a66adbe194d72c53c15f764be16d20519ee4a80144b40e38a2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h633e2d0f44ea3893a0ba03ff891baf24dbac9aff8739791201876f6e4e9ac3bd6c709211152b5f1b91de13d1c2f46e731f09f967feccbc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h103e4fa5683380630a5834fc9c64c487f55ec759859a50eea5fcd67060612c0b356bad7372ff8d220579f088703cc8756e48caf65ac15b9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12a0b80fd5dfbabd320752554e8b4254f8db347730c92c8a5946e96b6a12a9c2d5a306b1562de1ca14d1162a5f5f2c4e5a420caeb751a05;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h149ce03041264771a59febddd2fc506cce41667cda49542724a504d11ba610791d9dc84d8e49ec2d91db9fba6c0dead4d8e9b460a340708;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6a2c02946e7026ac7336271b093726864155fcad3b49dc65126b74dc9ed40f697cea53eb11c4614a856bdd728a81676bc21d2eeca671b3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8e0c65b9ba5490143eced2b8f1e214f166e2625690ffea877bab1141d96e54ff540fb46ed7535af8656789f81583bb4a6e1415dafc76;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h130c3d42a5c36a9f0c5d788c20031e3147f681f37c652aa86fabd61a611eff89fb6fa0b16847cfcb862e818186580642a637337ba72b99;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13f93cbb3b6f2a999801370774d39ac8fcbbe67bb878ff5358d395c6760aebdc07b7a1e2c7e953c96c5571083de248b978708c5d9af34dc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haab3dcac21b25ddfda7a73d06a9dc9281511bdd76841d9997e530ee6732721e20100bcc5f67f75b9521c6be69ffd57a8dc9b38531a5aa4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4197a923fa2ae7aa59799f432b33f5b260f639a284366e3eab1b0a40fe163b64802f74dce87e6136c1fb482e4dba4896fb8ae444287ad6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha270f0e45bee7c2268a81428ebae45e7f1520490fcf4b38cf5e46d36a981868ea6ed60e9b4402e99c91f8d0695ed12b1fdccbe1a4e9338;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha5d8cf66a1b37c649f0535d15a6fab8f09b629e9a3f3a8281cee6e5c8cbdcc65041050d28f9e5e7fe56866251ac9a30a6aedf07620e70c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h866afaa862e084efe31456d847c2cfe88d6b5a6189130d41560e664b45525cf4aa2544d53036968d444ec88016e5f3ae3e1300171a6d7a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17a28ffa9fee439f39ece7b9039dfd803e5679abd64e692be64fd0fc717678b289e8f9cbcbe5e6e6df8402f9eab3831e28376dff88c712a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bfa543d0afb218244e633c57c99e57131648f3e79bb7181a3394dc39fec9bb80e99d49fce2bf3105b0dd35f3b09778dfffb1cb06c29fa5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h131d3cd6066855137acd4b79679f5b1aedf004b050bd45923d306bff35a7ab4fd5a79ab5714a3bdd0c1184533e8dfcc47c1ff475934c41a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15342d345fc355412e041027f4f93d0adb6ebffe476aacad72fb86cb3365ce5980f3fac4ec7c482f4f7b387f458a939f7fe71ee31f33e0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5b1850a0f87cb8b4ee2923f523152d1a804b5deba0ea9ecf612077e198a36f811aacc69fddfe8f567ba0d43d8485651e95d5fa4b5d3325;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10f26c33dcc9a110d0645bdc6f43fc0a0a4b6c9d978b9eece72d8f16db098dfe35be6494b401a1fe6fae573f3aaccec9043bb6c81ab7c61;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11335e28cac09fdd40f52438741fe2e83beaf595bbc4fb5d94370ecd448acdc3fb934b736f7e902c8a632ce9db7841d83ebd3868ee13853;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a40b918b357aee6ce3baca2df6da5f89731f33e5fd51af65e0278ca8fadea261f668bdf87ea1a4765d255e4f7cf5f8db5f946bcb025bba;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3d98b8e6f593e8b2ad0664673645dee630e5c48571cadbceaf6f5a6b793b22a9a690324d3e1005df7145ad1213a50bac0750673b4ac43;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1783096681443f8651d9252b830620b7e9b211546620b060b898d00dfe240539363d38ba08631a1bd305839ea0a74a33f7407c9ad12686e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h170f89f7b33abe4bdf0f8942c79de284d4113cf8f890b07b206b1a354b0af00d7c9d632ee2c8c7c653521ec3961cfe4698f0b43f1d868c5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f5142871057090f622f4497b8c41fd9112fcbc5edfc1df9ed782fc19948f51659913fd1834cf55cfbad3b340f2f1d572e9f2d587a97046;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h101f5b29e0b92b61eaf993587458154c130f14da64f6665f9bcbafe5159b81e8103fe6c65dbbf06d3d6e226e8c8b087cb3c91ad13ccddc6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h29db91ce25dbe38eaacf7e5946206f84741b883d351295285b7702983d65adcee1d25c526013ce1e59797a1f7900e3c114949f2f6ff01b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h104fa0643919bb4b044eb1cd5eb74c997fdb882812f9386fb73759130e45468d7091abad6e2d37252a27dec9686181ede0404c20f5878f7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he318c55cef3c4e592a1439b7a32c9c585322b78f8d851ec58fed525f73a06ff00131a391f00d2fcf61ab14c2da25fe1db4633de2562e2d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ba1ce2124d8d1ffdc87b5253282df388690c488612cdb488e9b63a08014ecfb63e1226151d29e6525bfa9fe20247bcb2beb3b4ecd13603;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d9fcbd279f5bbbcfe7c270dff5fe679a81824b1c8f58119330cf76ff71e8dee575c3dc0013de69caa5497f454a529a1c5c648f0a4f7bed;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bbb93103202f3073ec8eb4e24152a982721e2781fca5ef842e3614aa626fca16c47e8b36a067f81d675d85fdd89285e2654efad19cb322;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14b30e0781e2692a3e142ec58575a8ecbea40a2b25379c37ed1c08c174c3e35effa4f0c677f7ec8629724c63c957023e0debac1e27863bf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c43d59f780da47237f86a2148ad2b97096768025f5a4b0d8c85c68630639a7bb71bd435e39a2fe51400f14203d5c2b3e9df17a527a0359;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1384b3a1482998f39beff03dda3a6fe1fc085f58d8610bd12fc271f0660f911b90564c3922d946c2a52f4c7be18f5de4db80308b26f8818;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4e26c4ed01b56716938aada59bba29f32a7edf906ccd2791eaef2f7e44f750a1776d2da9565226fc9b3e68f327227b2839e48a253530c5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9935298b310778d6a9a287e61be57b1d7dfe9e12ba70c0501b5d3c6f9a73ae571827b7753870501bb8d4381fd03bd062c6cb99a977d5b6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19035c42aae68c65bb47523f701d0fb60d2508bd74cacb8b58c749bc4528ae483b959784b20a1375e1890dc8b9ec0dbdf82c1792bc68839;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14a13e86b3775966fc1a2ca3ff375ebff1bf3df58c95ee8145f964c941498ca7ad5ac6263bf8cb2485db0180b01b65a5fed31da40d2dc2f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5fc0ace2e3a3af7bba8f69ac5309b224ae165d97e699232e53be272f4fbc548645bec778a8def1b8cb53bb440abc5681bc9ffa279b94a8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1da625e810fea84538e9e7d283ca0bcafb99b2e43663cb9dcb9ea18567145ccb9bae7c0a8444d150467b4160dbdfee01aff79e21aefa4fe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fe7066a14a48dda113cbfc13401130802e14feb7838e6a8b84ee44e3e9d09605f9398a45f84c032d7243f65b4b6b866c55510508dbc0d8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10238005018885c17148c8d16f61ac963685c4081d867192396663d684598da781c23a2cfe2b0093ea4c481407f1933ea2e1af2ec02e990;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e1c928011d0b0c1ad7c2e9ebd66e6ee3bfa339a3fba8e5a0c9e7d55e6dcac8456022842648b4b5dde35f66865a8be665b77b5346bb397d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ed5c3a5f341bc13f063753ee930d0d3e465072e4d084f96cd8931dffab8fc41d87820c2e72530bd3a90df298b9820dd503321314b47aa0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h31cf64e1049110d0656589fbefcd487fdc55cc01c3cff1d7755314f33f593633373f83dffcd01073c1b7495cdda6bf35362f911827e4d9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c6e4f42d93543a1f84a726fed91137b6b2ead2402ca208ca56241fe5bab28dccf78e64544eecada89864f6828a9c4d2978b215188f05a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcd9e93a23cee6e083723861befffce817a094682a2afc2ac1983e54400ecc01dd921b01d8603775c1ae48e258ccd850720c3f796c512d5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdbdf5fdd5a50b2883067cc7371413c7f46fe1356dd1ff3e7b45da82a23d9c591da0df3531107282e0f6395f8c49485d480346a00824c99;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf9b9236ec29947bd44d9410e5c696b31d372ec090a60f01f8fdb70dcb2e8d69d3ec798c7c3e614dfff54a40670c4913de9ea781d1cabe7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b57a147a79cc04620388db59721bf75e209622018868c8c131f47b6524b0c96c1f427fc846ed8653bcb169b775a1bb481f365a53631beb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12e92191dcab26731d0a9c55fab9a164a5c7725d2b6ccc953ffba525fb49c501968ad7feeb9208c3db72b20a00e168f4e6c2c8c8106cd20;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h161e479aa997f1013c44ca1cfb630fd013f88c18318fe481251e124dfe1ad74b50f2c4d4b9f7a74450778be60c64ea20d323bb8e2650879;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h179609b8aacacafcc7150b14715f7c9eaa4e44b7d7c02c15fb022a6d1e274e5b1248947f9101dc7d2523cee3926004c9f3f04daa241bf67;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17d98b31ebd2da0bc6710f2d06dc721d21ac663ec4fd615d9c7a219d8e5aaa3b3419a9b357d14603ac16c2d2fd838eecb504b7ebeadc0af;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haf3affa68a1524ae3efd1ef1651feec106b9eee8743cf7916ed715fe73ba2bf223d21959bc7697642d0888d761cfe00ca4e305cfe0142c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ed63439f4c83fe7845b8e33e6c8212b90eb4c11555f1249eb22e6084f9a99770c0e2c8356916f4d501fefca1097fc08af7e08f4967e893;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h162c26f177cb2e4dd692eadd6409b322a3a3e93453577cf3b0c0813ab4b5978c87ff318355dd0d2ddada56751f0261fb8e2929cc9f19198;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7a557765464154b47b56150192e5a099aad1936dabbe5da4e6ca8496f0254dcd1895530075459d5b256ac1450aaa27af4e62b219432583;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heef220fb6f966af508bb6c73007e1a635619fe91eeadef86523b2f27d53f0d8962e310b50754ec433b1062b8b8958a03d6e0dc56628f15;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h694f7cd398ce42a29485dc3299f9d4ab66c234a1f12e3968f89dda902ceefb15740d5b9a539aa8ffc3c12c3c34d146a33283f59e29264;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17bec8ec455a83fbf4efc7b59319782015723132c856c77808e2715fb5ad0a14d5f86fee4fa8a0121e4b444ba9b0a07cedbd2b3b88e427f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fd562315aadc7e84b5199bc843775f778022a3e85e5a1e18d5e3ce4073e432261e6b4453bda71439ace61fd3f2b0839ddfaceb824b6551;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1caef9547be81a2298126ad6b3119451830a83fc0cd65f281acd717c868b65ae8281d0dbf805ae28c069e88f76785e17e12614786d2ea91;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h129196e3308479bbf5f96d01372a33d8c26990b9a597796b64456bb0280928b72e820d0d3e4b44be3e8a4b080ed57496c1f62255aed7d47;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15d7ab2246747f2d76184c39214da28e97a973351d1d00afa519c2edd397da83020863590b94abeb6d9ac16a8c741780b06e7f0a36c354;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc15413a4f6aaf79dc704f1da2a0cabd8cadd69b924295459d98b019f99ce2cf1c9a6fd53563d7bad848462e1375b3cc1060098b4cf6275;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10a642ab8c4c25ab13cbc92720be2dad3004e63a99ddc38e3246b6e0e7efbac232970ed11f8650ebd84a4b1227b9e15a8d14e00e85e62b1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1752abb20cd0d6fbf5f668807874bdf8b6171438439ba5f5bfb2adb8745e7465982d5b5ea8fc6edb1dd4886d93692c8087fa2ea6e5467d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5b917aba09a1c9750f73446f12c44a768359014b4872eed0e9a1aafde17bc3a26e83ded2e41451cd720dba257d322aa49cccfabc446eaa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf1de6f69654ba52a9843242190e05a3ac8d5049cd467d68c4b3b263e9f1d94f82e4f116496b0deddcb897571474c701383d2a0e57ac083;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12f7aaff4eca2058d088d3fa3451b25ecfe36e685892e626a0a677b1a3a86605ce72f62fac115e88d4b4a0edc84d70a05c9d7c01c348627;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcabada043c07317eec420bd12306e3188b3e857b18cd67f44e3c1b64a5b0b043e83ec5bf10434463307beabac9cd40b60e8fb2813ffb83;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15707c4cae86e231f396902ffe909b0f7ba4480fbf8a73b48781900b646848ce5dba1a6630caac83c66a46cd97890b2157b62421b001921;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4bd03668e93719ad5c98566de35400b62fb2f661f23055a76ae22d396f1551a15b2bd5b959b2768132c657f0fefe9d732688423c1159f3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hde85ebbb9981c5a1e91236c3b5e4cc6c02681d9d0f7dc77bfba207e35536366fbffca9edb1df7ee4a025c65216bcc64ea4e7b142017281;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f983e1d7d2373493a533ac790cf51b1625d205d63f0002257f2e018181d8530f4fad6f476408a4be942ef627aa1f572ae06a83e3143146;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1006c51b731755d9713ee64a2efadd877b1868f0e1e09db0d9d1d1ff634de666dc59fe82f2d5fd7ec01262efd9b25a441b5879fc4212387;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hda8c573bf7a6dc5b5c7e46568f5a9e97243d495a2187f3a2529d7a70fd331a64ba8cc35286c77246f644974d324a90378b990d54cf53d9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bbe9a6c301ea00d9790f8b1ecf20e7193fe3beae424b47bfc0d3b0c574d70dfcd46fbddbbb453cf43feecefb3a5376c08ffe7f3ae7ff80;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha5caf2a0e5b4f3e350c1a57a0b81c0239f0cc0c550654224e026602a8ea2ae41c96336f1345dd5d4bbf37a74cd4a56271bfc94b49d8e7d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ab0feb27d48e836676970d14e15eb25caa9b5ae8619fdcf8360f124a566ec43bf9611cc708888aca3ac2014f9bcd153d18cb92cccee308;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd5ffde2ae150fefbe79bc8589b485c2eb0b6f51482f21cb27849017b494292bcbb5aff4aed2b6451f0b12df44d923b63e540981a639eb0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h98e84dcd01fffe019e3e64b8cf965c33d9750de4092c59586ab46113edeb096155b5c25cd4346c44caa1d68f6ebef7edc9adbb4298bbe2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h127fef439e0191c9e72ea3ff6a4a2fd6a83ad6ee6f86eb40a6ecd82315eeea61a7adb575aa483923f912d208fee32d1d6268b337499989d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h132669aaa66f0a90eb5119797bf465362d0a5fee504fe0fd2ee93629e9ba0b73f9ecf24ea91ce1d6c876cb5a29e7d992ae8e1b5040f57d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14cfeeff353af1476f08b633e35ce1779a5a12e6064931e22aeadfce9696f8ec9d52e5fcfb218db47b00160a07403b8c0043cf652bd09c3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ea201ac74d92fee0c81625e7fedd6a4e936bb503ad8947ef6183dbdc865049795bd934453231d8e12a349b6a70fe9dacb2910bbbf77a3a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a93bd67394962044c7d82c95a84ad055e35b5949b35cd667cebd0c2b6687b35a626444c764a762487603a2ac1ce61d872492ea93b3fb23;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e1ff6ad36dd1c0597cd968766d1c966ecbb5ca652569a0d0983aa0bb3de31736380baf7e80130095a9540186ca69b2aacfb18daf027959;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11a745e9a90dad59f8d77558fc489f3cd818b0ce100e6c3637feadf5a056cf5d55c0676362f5653f5350c3f3fb034922cca09b50b9e6c48;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h112853ceff664b35cd5e4eb37007df1da10c3e0eb1383d257233fbc3f66fe25f7075dde987decfcefd74e7dd750db751b4cefa346faff86;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc16f4191079046d008ab51b3dfa8052dfa30bbfb99c8d144abd0a9ac3f90c1b8988869326224e161d39388dbcb8633192f22a28ff6b336;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdeec7ba013e943981e3c3d9f6fab8867b01eadecef00d8aebbf6b9011fa88c9606b226417018b971826df676cf6f5b0373969a6f800d22;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h141b9e43c97cdc6ef0a7169049445dc67d4c1bd1b7ddd2ce7c81ad05517fba56eebe5e1762a553c209db99dde25570a41e327b0191f9567;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h145af35985b4bfec8ad5eae6335cd92a755022e26fd2784e02178cf9e7c04c29f56c0c34a9327e1039881c54d11bb11d7ba8b6130bb6236;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17d0ffb020de8d4b08d3f13a05aa842c6aa5492b2c2efb997243f5a2b95eb204778a47ff3f1f80fe89e86d8e4912b039b576c28e077e735;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h183484973d3ac0422697894dea54bb6476da9aae87e505ff44125686ed49fc2a3d0b366aff2084233bbf905e50d1eadb569b2f61ca35868;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1436cb6c977e42a38e94f3573b9b14beda8a024e5e2fb4ff6034427cac97308db17da35a275dcd47063247ceed54a74e37218a0682b9348;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h248044ece79f387dd28def7ef5b167c66f36cd7651dd1bb7d021411d7d7b4cc26622fe9d5215db575eb1a65c33930b0e04e3a1753919b6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7a9b906791cbe1a2a0bab11b9a254bb85ddd320728f0ebb5f3ce633f17d6c9a22b70d56a046c036edb3fbb9289e102433bdb835c11d3d5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb48feb139002ca53b0635ef6430a39b958476a19e90e1c0840af4424a86f9d314961f3d6bcd8ec4b8391c882d74db655896dd0539147eb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10f38d7566b59c7d13b4ad71a9aa5e489b2b6793eecb9de3975573cbd0c114ebed5bbcbec61f8ce48a51371c1d1d1c263bc871e8098207d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbaa00e0ff753c0e04c3700e19f97af9d2ba1cae9b336398d1838d2f9d68841313e07517b02102c374b00291a50929e7d2f8cbf25c182b3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18158e38aee765b9dcf33ff8d856c62ad8854de8734c08b553980ed4f4754e760ee2945c817c97bf1763a1669e4b37133f526c11c6f9e8d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10874155c0fb2e910533537036d0c574569c5bc2fda94db6b756089864fd596c81a8818ef6f2466dd208eb406bdc9aa077597c41f67b5c3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1be6f1ed270436b0c053592d2a1339e3cef143703eed39210a8880e388dd1ed865d226bf2e7f2881cd3cc2fe8d47c8e25cc614826e79e33;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11529db2da650d03db18652f3bb49dac544d7ec48075671be21e034ebb2ada8c5b84d2e4b99524d5bd0832187ca7c0f74d07bddcd433a79;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha96f351d63a0fae6a3d663cf4bb98d5e3d5bc165c3f145f89b7e16030bab16645048e0f068b7766510b53c4e14aa46c3c363ed7b36ea73;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8d8dcb539af3640b63232abdaf91304f06f257794c7d9a138af86a0896dcf24e1ed6301d5126b76657cd57f880e23da200742a9301a67a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hda76f8b708fb058e0b734c3783a058ac07d7d2a7e22cbdb0d79289d09aec93774e60bdbdf8a906d76c971334c0cdda45658b15d58bff5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1203ca1f83e3063b785154b48ef43a1c847e0518ef5c7097abc0e0ff240df3859a5efa2a6ef04c9683e0b1e8207f312b3121d18c071aefb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h92a6a7e4cb5a7a9ce24520cd94248651bdfd03d02504235cc385614309516a0e769bb0c4908523f00476bb0bb3482d0ede89d9cc6adea1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heb946dd91412999f7459856719a451efcac3a43c94ef2604508662b3870b71d8556f4bd14a76a027606e068ac4584302edb27d2cb7b6f5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18266821e42fce8fe4abc65a9dcfff61b519fc14cc482f3209dc72551a63b15ac58713b64ac3d0aeef82b5cac55614e866e8884e6ffece5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha59dfd84e982f7d07a60156508f49c6561afedf544a518548383ae648aeecd7042cb7b1bbb15281c5be11f74706d9824145377a368d352;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17cba4e6e5cf309d6f271593e3b6562567d8bd3c0f3985954ae7a43369fa4ff22acc2ec68256e26a002e25c4e7efd9439dd863b78ce2f03;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h90c0bca335144574285f1903977ad2e8a4534d53d46ecec9d01bf3665927079fad7f4e2a95584700a4e0c8ec6f0598ef46779c85400b5e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ca200a30adee98712a353082a75e71e637ecafc19fb1bcf9d878312ff4c36669591f3e082ff290fe39ebb299645c0d03c472d23cc45197;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cb45fd8855c77eeeb23452212161c05b0ce50dd53a25005647497e5d27cdbe17e9c7238611576899ec281ae862030a28d830942d4238e0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11a747a62bbeb500f1294f19e891e5fdbf788fbd4aaff7bbc14d32c56d09aa2cfe9c146cbb7e07a29c33db27f0dcd003818a717617329c9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9aaeb293b2011a3037698332136ba28b5cca5f16fcd6edc1e082886ba11bc6d6d4a70728aed2dea3e2c5b2e98af52c764d4248951ffb4d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he675bad5d261b7d01f66b7a868b9dd3820d12b2c3c786a7ede7e790ffbbef9c3cf054c870ca34736b53a7f1a62041b960dbc8970659e57;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10ea81e4755d0b19959317e8040b553b3ae3bacae0cc8f5dccb39b2330bd59ffebe76a01c65a8c40bae4df25e745f3066e32cbabae943c6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7605e27deedf72a5a2fe95c2c2f5499162d4d217510aa10288554f2b89c518aaaf485fee4acaa655e829b3b06cee27b3061807b695f459;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12466cc38d1ea9645cca9d655571d2c732ce718c82b85e3c7556bf3a1b551f8787f48ccf8df7a8d9f7c5f721c398b0f8102d276eb516eda;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h140466508812dddcb789863e1c803d7cd2e6f4f858ea12959975d3634c7d9bd8db8a90ef7b698c6e057c5be5974c4c15ffae4b9c2ca8393;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18ebdf57b1c73fc11d2093025a0a7143b6659e34025d8f76289ae382443ef7c01c9c99cf34b3076dacaa31686b585f71b2c4b0db00d31e8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3f8891905cf8c76f3cb5f6d9b484deb4199851f3e113ac7fba981b5d878bd0d556be8201ed66bb728bb003c90c1c80b89ce9e20d0dbc9c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dfb28dc0d82fd34f923470bd9c357b550bae9959c729647f685de7301bc6cd72e9c09e278cec9692afe212edca40bf4bd36f0b26903ccc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7302cd8dd9be4a8d48a2f67fc00094ffca26efdf2ecb4f7b4fc30773a2c49b71467047091a6ac0e6125e8ee96c0fd1cf3dcf14d2ec8a71;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a8e760af4221d1adb76ab2b243f801be834669ac4d4f7ee4eae72f53586a8a27f0cd77b74058a36d4c72f08c9808e3d0c81b3c01fe5b92;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h189d1b81cb9751d5a2ab5dd9ab868a3077748176766fd968bd50732fc02a93495f7d5cc8ea5ab16def433e624e498b646237f40a8cac137;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19a23446b97f850bb52ba2b1df9b7653dc60a3a81ddbaf3516742bd3fbbbb37839a0966898ad5ad79a146d000401a9a908e332d8f692b4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a15a6ddfb62877b1a7228270436556ee34e87baf5b637f47426dc64ffe7b47bb6f279871b69c7e60060db016a63e88992a3874cda0d159;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1521cd807c0be7b26443c21df97124b4a7df0d37654453fe8d76000483b890850e2e0db10c5956473cb41d298586509ee97b54cab3e4a08;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bd90381f334c001e8d1ec0fa316d7757410c2ce6fb33dae03446aa9e63a4c8d969882ed97a56591d37cd6b2417436844451a11fc311e50;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h54d98500e3aa2fa2ed9d6e193bc0a0e9eb35de5f90ddb0b42d7a2103c2e4ec37afccc747863eb3da278f816e63c21218837217b7116809;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd0a2a92918e08183894e79f103fcc91ab4067d1ecde1acb2b882da30de5353e5687cda58c6a37798e1dc4ce40bddc3f13496384faa7225;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15e258c5d35c534f7bbb405c28f0b3840ca873586b44ee0f960dc94fff10505c4556b6424a4bda439f1c4dd89e279489d6ec3ea7397c094;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf852d20312a2f968126b4b2639d0c798b6dc3cad9f4dc37aa8e032b26b4c2193d40797b7a0e097da7e4a2f1df3184d5f298fcc8beddd12;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8f5ff9ef4a416ee7f670bae16f350ab3494bcc953b0535a06995e4ef4477ca5bd03bcabfd3f44ce691f0c4bab323a0c61d8814df1799fb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h89bfe7a57fe723234f54f3d2777b6b25c3254e0f794de68711ff988cb60d4d9d2c6cfc799f414b38bf758ce813fbdc7045bf3deeb845ff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc5ef6f64e7629022de0592db37a8bd5f56b0b2f493926dd80652e709ce3c610aa4bd453dcf168303fa34ac1eaac9db0082b687d3a1c2bc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he409d348c3b31925a90b7dac687e5bae54c1e65d0dd5fb646b407b8cfb67a7a1ad7ece539cdd8978c91e09f067ba7b8e2280587779881;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17063f7e8ac822ca2200c8ea1f08e5808e3170557b3eba894e087318034f53b05262b803e968c2b85dc57d21013226937850f46e56532ba;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h185940f75fa88668b4c06b6dd1c3980cb7ed1c94ae26163e68bef9778e7361f4c0f3314a123ca15c92fa4b5a981e78ccb9ac089b3c4500;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heea335dad37f2b516400f8556e25d4e5ff6ed90b7869d4d3c3f085be4a0b94d775c504081dca10890f10c0faf34f0f02b5476f7a3dd603;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc4176b25fdf15b403f37a30efd51961cd89d1edf6fd1a453f6acb7d5198d9c104c858fc909a7d0c8d2a790b4a6834aa36a7dd509833891;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha2bc8bbacb2ba7819cad88ce1799d95ebd48bca9c1b4af7d0a3c4fef71c4a315f646ec93517af718b8ebe0a20b8e7d4a64b1af41e0de87;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he2852aaadfa3c93b7a95446d29d59cd4681c22e129d6194e4a23e739654e52d46c3396174e37940c987e09be2661cf84cc9e42d18bc472;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd3d38bad56d53236732f6d9e7d2899b3be80fa51863a411521dc11231f1bc04b0ac068e01202ecd2a88632597314aa60abbdcc224eb902;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14fd37eba5da477667d9c135a7b4f3e66af26817c63483cf4932d1c7f43ccd6465f902d3e9bbd4b0d1ff08ac77a51a2a178367963f95dbb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha1a40e74b903532b33e4973b9482a60ecc77a4ab11f25e0b029c0eac68219a64f7d79f1dc70ec44bb28057ae4aa09096e5ccf91cd9629f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3a1d0d04c1deb1047fa3975807d9f3f7a2832534c47298b3554e526c3d0b86bd19b6b036e6e4b34a61d3ea553ce8c249ab582e1230e1f6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11c13258741c9bd91b8dae09e01aee180b035c1f0916a161ade16a40088e8b120dff5b406844ff5b046dd4835e548faf57dc238b93571d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15201996a4b81c901f66c979048a65188380519a512096ae2b6534946e2247a5c814dc96a20b7f58eb8795aee64b1b463a04058ca27a36c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f38f0fde292a59c8dc7282f24dffa49be43ba6ed5b10bd577d2adb59b46b789dd63bdf934905fdcbc6b79085eba4449c572e5cb484fdc5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9f7f9b1fdc83e09f7dd03a7f7f22c0388aa6ee333ff61275722066c2cf9524a056a2c803c17fad38f3dec68430bd40af2d9b3df07b3527;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6fd52e260bffa2c252be4389872c2069ae37eed8a6ebac49925a9e6a56e10420932f752474e4c5eebbfff63ec710bfe621eaa46545023b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b6f007c9c2f9ea5478545471fccdc83c9ef0cf24288d7875038a8cc6eeda64374a7cee01d04f24b39a467dd9d266bdbbf70f010355aa3e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1089b1303e398c33c0a551adef38edbb8c665c06191d3018f0b24e2b10233b9cb87c2add11c66f1041fca0f8ba9e2fd9764076b74b2b16b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1275afbac6532c21061babbd76be7971d732adfa40e5902089dbe75cfe8624317b3a162a2ae9b0c0df68017d185123ae2a59bda261e0489;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1912a143ec0daa4c17214201517b20dcd180fc83a344605715f52d9d89963005a0458c47810f5e8cf1fd1330532032748258c8561107fb4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf2885a6873a590f63cde58953862c35b65dca79f3b53c54f9b9e19d76b6750923a41d368f213e8f18ab09864c9e9ddc812610a0d65ea7d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1456c360a864a0c90f57d2403ff6f522eb267f38fb2bcf6206ff9d96f87a55733caf011d823273494e129205069714b3fb3cfa967d233a2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16f01771baf8a1f916f31353ca149e58e6a5cbb2d2a27fd025302a67e4a2937d76c5c28910ee7baf57acf4951ad1d2fd93018b44c6b702c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h142b84a928c02cd045db5a5f00e3f9bd5adac022a4307aebc50fed22a4c8f81011fa59c99c6281286230a37bc73e9d11d8b4be577b135b2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b2b648c69efa4d4e54d1391139a0427a2a2afc921172841b5b0e7c3add9551916f64c0bb2ed3d6a6900126fecd17f5d219a14a550f5344;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17f9cb726c4275c93dd0df168ac02d505b54315e6d9fe054817cd836bf9a611abb2b1b88dd141fc5acba3a959e4e2774d9fc955a3d9b32f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf2960921382b1f513daa0b2619f35f64f9a5b6d5adb23ffda84311bb896cd5e4d79ff15197cbd94caeeb6466c72908feb5b991bdb88d58;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15111673a899f7b172874543da18602498d583e33ce5c89f0ac87796b77363cf2d42a7f733cc88dd1f84f4a1588bd1707e638bc48b701f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he8d46652c98df1b2b64fd0300f496ba1fafced4c389180c4d716ea5b8f82948681d681eb037c32de624bf6a4c87e77eb1d12a6d678eff2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eb16cd4dffe8aa1bbfadb1420eba69d245061d07549dcb7bfd9fca6945aa1f0536b293927b138b359ca5d0823cc226c69efee086af46c1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9db78be3a400fda768c2c1263c96575fc52078f84d1bb8424cc6ce20155ed7e3ad32493bcd4030a228f2b6496d752424382a8f372ffd64;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h168cfe3307a25b40bf70a84e0a949e625e6aff216c8b91a282810cab4cbf8ebb8aa95e38d2f9fe1c24aab86efa956a4645c79ce8672de6f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc4eca432b2324f7c537ce4c57abbcb0ac8861ba53fc14c1f28e19c6c47ecccf5c0ef4124bb2c22fc9be88a95a3bd3868ec32459a711fb3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc39b7f16371a7da6b1f1e78cb11095345c73c00d1a280bc773a0cd93b636053e1d9989fabb718d7e5e7d8bcde0dbcaa9a64735d66ea05c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h196091710d8b7ee91d446316d0060a4c3934fa928d37010c304a2d68e024cc435bc522987c34243142bb715f4f16ac02c220409d2dce339;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h706d3b67443d3f9d57b7bd2160905e5a9b4a54763f4017f84893b6e53e3678fd6805de03e4182f20b3b720f14120a1004024b275c10dcb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7821a7644461f06483c8d1036d60fd1f373276459abeaab443c41f25a441552c1ebc7d400c8fa3d045e073c8939d897de1263fbb07cfdd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbbc82d005250439838a307ecd87307fa0d911420dbe5b3afdf0b7c24fc5457dfe6cc4b002736b8b28634abe673cc52139f3ece32b70d1e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h63a86fd20fcca073b3d68fe83a7e09dfa9aaeac45a428cac4c3b626ed50add0106f1d0ea48b5ba04366652110f9379e57229e646db563;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11290f382bd255f1c999e2e00f909390e5724f4f1414e25e07d172cd5865b8e7520ec51a8fd109fd343d5df915816179edb1f002b0b3a4c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10d37d1414c40747d84133fbf2375c0ecf65da1d43df7b6c2272f262a7fbcae5f3f07d61b0595d374b4b83ef14e4d39fcb73d4227dbc014;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h117054369d35f265eb7ec4dd73be24399c7ae015319138d3a3e9698419f3e7a90f324ff8a196869b597545c59078f26523cecb0c4fa02e6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10ae1227bb7af2616b2aac0a755deca3f34307b6085672379a8534437fbbfe4675905835b002a50930fb3eee823041bbfadb20c677a0d47;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h67ab80bb6161f31e3377f0785bdc4d7256e39f21a0966e6f50af89abf1c662152688a9c4f68ce90c829902a5a174c109d6b3eb41ce45dc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2e570c2e08543067011427fd7883bea5b5312e2b6f9fdc9e15f3ec97eec11db1dac67b683e380776abdd4bca94ddbb70298dec7922f26d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9c11ecc828637710eeda3878440ea0d0e411de12b4e366d902c0695ce5bc485f4f953308f921e340861cca457f9bacbadb7b9ee9a90431;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5e7e364b072cf4a469fffb966cbef3fd05bd17e93804d982918a35cc185d40e740ebd37e992b5c8d90e56e0b59b9e86b1442f5f4af98d6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c0d35e616c472a07eb6d692460695966ef92c0cb093bfb45bd92ee4355db82499211fbe32c3572b45d34bc5818b8fffc2063c4e8c5dcea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd4a150750d40d69a20800fbf455103796e220144c81efbd21f47fa88a019d6f69e98abae0775b0f722ca9fa9471eb470a5bccf5b498e3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h351873ac450f1e4d766b70c09b36d76008720ce176eb64e0957a6a4c8f79781756344415ed32935dbda7d79b4b4a0302feee45d160fe1f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h157f594429526cf2b25af84aecd71abc351d6241a71d04e993c3738ac21c6256f9eb0090b1b2bf34ccb54e858beacb648ccf9bef3fdb8a9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb98759b48bdeb73b391ab566fe25d03194478515a0d3ab09df86b4703cee4dfcb802c8faac62b55e10bbab3020b9b15ac0f38bbbf6a849;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he661c42662414965afe8adcfbc78390931e19afa935a40c2f8ca2ea2db799f5742f4c1bc98efaf2937e659785132b3599553c1d1f15959;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha7fed0b51c74fa90944892da2d5076ef198c259283fc0042ba6db3649a28cabc599ddf0f9cebff72ea7a4e1fcea5146f114117f76447f0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c953b54b1d6b187fff73c819543b276796347e1166983625e0422f4ab976afe9cfad581b2f1e25f40fc2a0c4bb84dff68aadb836043fea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8055e2b2a06f146ecdcb8be99fdc5ac803851a391684000d383336ee0b485a0067f8aa61f5f62d67d82535909f7d4eb9d5bbc8ac4bad1a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h112bed5bed9c74a3cfda39a120eafd0a4b663852eb3131dd8271d58a561b28f8513d984ab2ec564fd98e51e231fbcc839ca24557e49adc1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2758942b3ff1609a29750f7a9cbbb7df67a6c1cdad6cc5ea3d4d08294179565a74f63465625a4fcbf66b6e3d569281710d176f333d0a0e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1039778344ebb50d5f2507416d36ddf4b941bc3fd6c940360325d34f39086cc618e75835599073584572cf313949ef3a67e0d3f73a90d71;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h78abfe0f4f1c46cdc9e9368f3820df1d6cc1c7e5edae865e70541bd12bf95d09ea8bba4ee627058db8cd25b03d9c7db8eee2393eb63406;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f762500780194527960d7fd7bc1a0e42fa8bde3f8fab2c598706b7ad8dfb44ef221ec050fc4627a0361219502d47d2ff8fecdd20fff7cb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19bb3803337aaf34d7b1e4427bd23a3a6a3cdf22333b8023951a331c021fc546524d7fb842cfb2b722b92d93f4efb37832f3a12e530f9e2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h828d98b935f78da235ca65d31b3e4419558c70a35bd865411223199ae57505ff64be5e20c8d711bd68fff5add58c189e214975be4fb79e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ffa8d2d1484442e1aabba2d77ab05045938cc3984883cb7549151fa3881ecbe7903c749165a536fd50739c4ae1571183a4fe98b640abee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d1077333775e7a71d5232f8d9ff6cee3ebe153759e9a87f64d50ed60b5baace0aa34f08a5b82d55c2a5e16a95f54edb16693facdcb299f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haf9d4580109887624d4347d763fd08c0d78fbcbbc2bef1d766d1076a0365752bcb68143f5c82218239468648460c46d29f5cc59325647;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c17a7c27f5d262b6579168e264b4dd90d1a5fb5c1099fa698d2f6bf74bd3f69b2124e08e55c9eeceaa1db5b10a36e2a12251c9b1234d01;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h581f7f2bb0284418267df2b6f56c570ae69c35db387cd69aab85ac23e86a92de257023ca57e7ab4cea61388bcbe428379a02fa3404bb7d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18b99c955d6ca1ac7a80af060c3ccf3ed1075169f191da84c5d73ebfc5365f32f1d0378bb35d3d9de9b458f7bb56db843c7d38971a9985b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10cba5c524aa6d607518556c9abbe84e463c9caf4ad4d629cdc1e1acb2510f967d7b1415ca84c6b03930b007eb55bcdc0984e79517698fb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h149dce26c8a27ff298cae361b8693e9b17dc01afcb104044dea65cc96755e70083925cf3cca6df36c45a14ea16cb589fd0699ff4fca7141;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdeb61efcaeaf5bbf0b99606e20bcf8cb84f30f818f9b00cfa2f091c2da513f7f50877f1cdabc716136e5e70f7899448d5a195ad75d7cc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd75fcab783e7d5c19d2b1371d1ecdd1ae95021d6846c2644ba436fdd55291263379c7cc09cc3cb44e279fb01e50ed0220385ce6e8984ca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf483b9028db13b8a45723a02c99e876a3162973792d835ab3b32340838a22cbb9315d94027a05ad674b514bb934e553640abc2d0c72a79;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1743cbe716281fa7c7734a6425d2be5c7fa4220db48581a867a0bf8a1694cafbd8505e90cab2681be9a1e848551ebf73f23111429265ea4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dcd86c4cf92ee7095cfdb874e9dc647131f89ca28c2384eb9a1b64337d496bceed41b6cd38d280df2f2f8975921d526f3e0400ad85cc52;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e5540da49543bdd4f41240695e03ff68c3ab9edea7efb0c5720b6a12b57a6cc7db7ec58868aff0cf45f5d924bd540e0067800f1f06f918;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ebdcb4bd232b2f90840fa97437212c9ffa7c919d1907c4e63e879255c1017a233e97e0f3c37a84f8dbce8beadf504a82f0b2f46834b661;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd95065616824e87276878a44b98c766cc4178f987e6731f5f88bd6e4627b7cfc57e2e2c9557d5f458396d1db85b5ac4c1e9fd020541e0b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1226f32730a4c05b7bcb847a2c397cb6db3ff5cf811fe125b7e3332cebf4ede12908541af735270223b4b54d2dfbe37ec22dc1d8dd4461f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfe2be4adf56332fcde67ff1c53b89c6f05189bc2638f25b75c38d1896690d6ad3f45ea825fac4a974f03c2276a6fee3abf214e99fd0848;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a309ac10df100ac64a8e459f75243508e589890ef086ef3733848ad294c4efb76098d8fcc6a1b3d246ff69578e229533ef8e84b4e10c2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4f9ca12b80038472f4c34db5da05a488b059747704372bed73194cf6ba2f95ccbf647f2bb56f853892cf9b808f0e6217279cc7d8e97b0a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hac01b765a9fee83fe8f12dc60d429d082128fb63fd97aeaa32879d5bf10804bc7b74962ca5ef7559ffacd447b10d9b2e6ad5bd4545f606;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e7c653b4280795e767144d4d38c6f74a1a4f0870a1830a5a40f17068c7f59698a6bf544df7c6aeaca4d047c7aa545e452c0426c238fee4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha5225e8c9bbd6d8b10db849e08c6ae33107e3dcea7a0cb0e07578a2221af8188e31ce9140d97ef39dee26123fffc744f8361df01e43870;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f40b83679ebe73d2d98866b108b2fac5b2ff6f883d77f03ca8128e8c7ddfb8902730356d50c785c36c355945c211b4f3813eb1f4ddbf39;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11a012392d873070ed27ad5476bf71a22684a364d64c1c4d3a9c6b07bdc24bfb43c1f88c4e83f9563b4b64fbbf6cf8e006dfd5acf22bd3c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcb8ca2fedf145c614083a9715738164aac71d24a5d123738e84c6461ff8e46fb45b1a44f6dd89791912914250e85ac60b59b0fe99ccfe0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc296643c25715fc332fc78576ea5881ef7262dcf0f1382e78ae43cf2b72b033d6a9e9e55d606faea22a4c91e1c9d7e9890d89ad128c288;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb42de98d41977e94538274f55eaec39488a3c8e0df4cee63bd2bd43a651c5b942fd18d67dbc58b07c8ce0f05e382d178c531cb741575c7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hde978e691e68235b50602a2a8376813717a3c6c1a4bd222b633b0872009cfd7ba284308f3e3456dc07fb37b73feac98f120bf61c54d805;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bb89eaf06c3d436b93eb05d41296f9da87c0a52b66fb514d80fda27b0431ddb3dda55e1056a50c632a0ed50d87863fa1c3c90a8d3f40f1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8d3afebba5d07a5e8811a1a051f8b1ffa46b86e3d19710e0de799f1857cfa21e68302f3c86f15ad1ca23936ab876e107707abd536cb431;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16658578059c206df6b3fc582d2c1e2ac376d9ae224265a7daf7920d5522ef6b9dd8ae0cdb8e5e71d70a942286ed02df42e3a59e8efaf72;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h334464ae6c17d4dad3546aafa884b6d38f58dd5fc320b0c53dda6d716fbd0a3a12920fc5746fee3bf263179bf715b8f357c66c9d3b3b01;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a52cb5403f81dae9dcaf2f68885d21a6b7838a79a09de89646aff9a439b6c47dfa3d8eddca696670e5c69f6e0654fcdb4f7d572f24bef4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e0aeb48bac758605197b263c0691ad684ffd0b3fc7d42f01116b7afbfd2c5bc7132c1afe29b385f6ebca399c85f2ed9c33ea0a923cf967;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h789e25f042067e79db39a08096ea51a00149d85c5df2c7268a7b9b498789c6f25b0b8fe8137eb105e1ac7abbfe48638d8142606f9d8c0f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfcc3df309744d7d80f976590363397bdb5b2bb1752b33cc02aae8aa859fd1483d92c30f4cef41dc41ef5451f78e1cbd241c3e89c0ae7ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cfe5efc1786b2643d928533fe6801e0577e1b376e834368542da672e42d1903325f0b12642b2f2aae77558d9c28ab7ae712dd94114e4d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8bdcb0c4416fcd9ad4925e7ac6ba2c677d25ba88712a24fcdfb78a6d7cbb75feb68f9a50f53b5cfd4c8ef3e22957dacb003fef0dfad364;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8adb15a19b04ef710b7033006d6c26aa94e0b628770f8a0e3923f5c91c860745edce37752f16dca48b31c9defb411bda437a5c123bc28d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h156983ac76b38760eca4210bb4e8691c2665784f922a4b21e7a077288a48ec110e1c0acae9b3f76f6e448dd720abb5bcbaeb32cd39fc6d0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h97b743a03bc01a799f04d3908dfcacdf58de1a5e9c8ecc20dc174b87512c7a89d56d87963ee2c2a0a92bf2f8d2a3cc7efec6ed38baa0c5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10394706ccbee9e27dcf0216fe2f22b6a3e6482f9821c153340019f8dfe712a02b1b420c55643c3da6615803ce7396f15ce9e68662865c7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf1e58aa4c65cbd0a46354e475bfad0e405a85948394d06df59d619156ea6db98aaf2ffc40c36b8ebd6695fd414c83316205bc66e8760ea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h406a4a9615720381c11680043b7c6947a5001cb3501219c8cca00a841841db8d307de3dc4e4f694bd0858e26b4ed930011d9c06d52e775;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h36d6d41705c33df3054104a9b6ddc4e8b08b088e7f00a9f9512211334cdb4f281c19c61db32ef500e2f05ef4e089c9216ba44ea07e7e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2b0bb44fe0054bcf78f30b987afd08258b3d0485ec83aa576ce29b3d86b54a0ba2c8c44332a1620c344f2bc65e7e62248ef64d2d006a6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6fa566e4382cba5c5d4a5ebcc2a0ec3baf0dff6a553641c40b98b312fb222fddf517e905220ae336c6665693cacb3738fb3ff2ffb67745;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h111417c2f3cf4bdb4ce0e5a19669bfa683a5817e98905545724a87d0f969e497e2ec4843f8cede5f5df685ed12dba79afad561a3e7c6898;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6d31ffb83432fb7e14ad4f2b6717cc708b9d73cd52603041d39de364ee7a8986cf65e91b43b8365b0587aafc1d43caffc922961d5c7611;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h176f81075c238d2aa0ba57238570034240f180d6bb012da21647458254b59d919d19091ec100995e243187a4fd12e27e36ef7ec1e2333d7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he44c59f5171d672b9db5e1c064bc8999945937df2e89b9102db79ea0fb5cc8eda6c400b339af5f5bf5b263e39e6646b0b8721e4effd8d6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h91e24c7caf616dbbdda49c9395b92df1c3d6539e02f03e81d9630faf5c1cd7a1737eb3d86d7e669c6f185a7c647aebe8fef6f4f0eee649;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bf148ebf11b2088d8bff781c8ddae9a83e3170c3390a583a5bb16d1afccd6208b7b5300656ad39ea9b645d64ca587b4e9f564860f9096c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c5add79f0d5a2bde215fbd7044a28d3aa0c6b6ccbf7d8e82e2cabcb00c906ebfa75c38fd1ec5ab3d48b5312d278b1e98ba4c209beaa6e3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb23876763dc5bc9861e7d0bb851a579891e02ba809bae5cbc412ce4858ce9fb652710e088b2ce59d64008f0965b56b081b62bbbabbae96;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha4cdfb23199583dd5abead4eaf51b0a5ef44ceaed9d18e7f242ad780b171b6f4d4f2c2863616be377dd327762612d1b5efe48b4ea5c3b1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f99c2308c9c6559915559d96b0e90b3dac4922414cbb20ba94bbcacb77f754a3c4040c13d23a155e23be49102dd53912f248874a30e7f2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc6f8653d1af92a0e135dc240fdd301afa07383271fa299aaa4087609da1bbd5311d2f578ab551a20f10f9a9bd6eafb872f1b4b823048f0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h106752ada9b38b2271337e7faa388eea9ebdd3ede0eea1c7896d8da3560a9217323dbb519e24da01347e76997cb32209bca24ed9a6ffc09;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7b65aa4a2234bc13034e725804fece75f6a9ceec7a2441681252d6548042ebbc0cec0884edb4ee766c40fa6a2dd0935aae5bca7c540c80;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h493a9cd83e4fdad8a521a847acdcb1dd6daaccf83cfbe701cad5e8409849ba0c2846f49687862582929c853e279ec52dee35c00e4d23eb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbf12cad2a8523788fe88619e723773b6c5c7d931893faf371d9ac42d950319b736dead0d5fc6aff5a9b2ad3f061187bbbbe503bff8c59b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15427145444516b0bb0b0a722e3dfb1c48f46277d8940362b517c19a0d717392fbd763ce1179df41033ae2eea170ffb6a509593e785c9ae;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7c28a23d189f7762addd8da68150e43fed2da3dd232aa5d6f282808a0222629129a9b40c52709039f7a8f2a01a5ab10d5d7d2eb5551f8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h27d102200de1e4330a61850ca84304a9b333e9c4f0373687940b738ceb72f4d62fd8f22e2498dc4ed559d75d95ceaaa8e9f395f915d4a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1263f34cf7e45bb5c59a083b90379537cfb5d1754972f10dfbc73b9366fe08048b13e7775eb4071ba95abe6b32226a7cfeb82492e5ee5b2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2fff425c4ce3693498f77d9c066755940beea22146bf33febd9b28cda1c853f99193954990f434da49be8e5d2a1c2effd930a9157ff937;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e64a34559711ff75f7e05fd88532aabe4ff47598287c95dc76ffdccacfdb907f0153d40093995d56317b1df84a1b436b4e3a839bfc226c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c602ffcbc479dadc3224179b0e2db993ed8a8f1b65cba98f567ec08b6ae53ba9409ce2ae571be34a4d873d3ea399b19ddcd6a8ec23adc4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d1e9f0b6c7e9fe1ae0e414eed84e66e0c558b4241266a2114d2de29abe6ba38aad13cf347ceebacc5385b39903862ad73982e51a92b7e5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1522b75547ddae9304d5ececd56718bb392a4e2015b6028a573aaa7ead273f846c053c44cf602254b563734351615b023bb4f80e21514ce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd7d39f13999536f88b8b495da5002714f74271855f535866f8e87919bfbc7a8291037b105d31010024c7d6059f908bb29769a89e8f9864;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h91ff9425cc9ad210a9af6d718cb902da602c0d11077e9a8b9ad9a97ea50faed43f4044dbd7a1b9d47d80540d4870d57b2a604d09202613;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h83c8a84411f0b286d94b76a28b7474c5dfb30a26374682920a90c4ec736d2f9a72dfbf419b27359822d6f6854c05aed8d04b830d56b9e2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4fede836daac778f372da9260253cf8d0a7923e9f57d1055ad9e3961cd874dd3ef45194930baa74817b27c8a4c744aabfc71edb1299a99;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a403def4e51bdaf66304f01aa8f4f63a407da5e4a508ec96b11e3fe150217033bc7e88fd433666c42245256b9ed995d3761025b5046e18;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f64f3e7f825a3df90781fc3c13bc9d7f8500a37f64c5d3c5a924dcf13f32a91fd77c270db31dcff2caa381c350eefbf07916b9d80ba3fe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha0787255cd21147732a4abb81709331965ddb288baffeae104d51a87570083a869b9efb8e36a2d09cc491a0f8462d5de98d732ab4a01cd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h32f225c9988e7e818636c95c4ce57b4191b73e14a43f98f412d5c49a1ab386c1350531fea872f595fbeb62df456e0f6deca0f654b4549f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1342bca0d5c24a000027da20e7f6c1664be090e0aff1b1e6f72d308233f2b9272a41abadfc6bcf5e8279e7781c2f5872abdb4b9922ab224;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5bd579f5af8f56130bc6ac1954839b84d0ee9d182e09cefb90c3f07133c2aade66efb5568bc228de3d79563328503a6a71a49268324b6d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h78e3540ead1200994c5bb86f9eb14143c7a4efe717931a4dbaa31de5f1bbc878cbb127326246d3a66ba45173f9921a9866f3be2748a60c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15788dd8fe1daea2c89420cfce34aebf157138bfd9ae6a3fd7a14c10f451924cf323ca523c110422ec1e8e4b60fca72b80870996cb0e9ea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12a304906e499d553636706e00b6617a46318acc5577536ee03f0a4581e034c7802031204c92e9fb148495d2572a78d55f0e7a15f89b300;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2d7d4eb9803e376a69b4fb2bfa2f657384032c0cc097ec660338734fd688efe004e240325bb10b1cafb05527d39bd146a2c90d06fd4668;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18eab1fa075092d8b898c99bc05a0eb4449a1c5cadeb0f3453265862dbab687221077aad6f75cf0fc8ca4d2b6337eb449f7f88606e8aeee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3865c6c5692c69aabb02a0d60b7ac41e3d53b33439352ac452858187b04b0d65f1ca0277ffd8a49b8dfd3de3b94e88d64e080e173943c2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbcb4a00e95323432d48be8d47abea0c8e8da8d7d7d70b33b861cdebf0428d06b6ef6df26ccdef5436e7b41874bd7f1c65b520a8d09825f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbe671f8ecac94141293fe09c4510cccd8e8418c7ececffa9c86bece4597e8827a8e231ab59ea489ae7fcd369379ffe7ecaca2a16524eae;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b09a902a0d8d382f8226fbfaca184b8bd38d1a6cbf6d4b747739e522ba04bafbaeb49fae6230a05e042e32fe6ea5654a24bd0479ba55b5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14233ed5649859c457bf70ac2944352b8aa3d51906ebe061d05d5478abc5c5f3cc506e960fb2e784da81dad2f18e36957309693f29ee438;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h63a1013920f49db583a36f3bd7382c3bc5824fc2c4e669ed2383e3cdc695bbe17bd9ff14ab6b9ebed7eae78a57ff8fb41fe8435accd7f3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb6c1ce31744127b47b58ceeb541ee2932703525b8582efaf5809ef529f0bbae7cc3a8256fff76519b705bae2730e78e9cfc8491f93d59f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf178c8221e79e2d7665a46554d6643e6d34ce8dc6b2e2847918500c1864a968a04e9a53ca55dd69e3604ad62fa1a3888f853c835330326;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdd3c7a26a2162f9a2758fc3bb4e9bbc62b1112a0c83cf37e87527018ef9fad083220f66d74dca2ae60753c80bf667f609b2cbb3319ccd5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfd85b23bd374a067d9a6897578ffb968812b0d16a9a1a230739781474286453d144052b9a3ca9ef4706a207f88b1b3507827597fc1f39a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14f5705c8271869a4a0bdab97cf7b82d785e81dec077ab4e1bd627a1ae277eaa505d7485fab780b4665c860075212adbea5d175cdc95e0f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bce58afe3deb4a177dccadd74f05db66e66b6fa7303c9291528b02f288cc6c12a74ff58952847843581652b3e2df1903b4bc5a55fdd528;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h145d32be131662305b2627316b30b0a495385661690eec357ca0be0487457a7da2264d71af335e5cc45462cd3285cb0b8aa7a75fef89d8a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7d5686e60e92cd646bd6ad67f7cc005c8fa483b20012509d1dea3b06576817818fe56d69ef40dc13e494d85f4feb05588aa15398b65fd0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16af472f566d6a33147ea3c888991521cd6b7740e7958d23591b40896937f4337d27e27d8282f6ccf2b1388eb4a8db846faca4605f236c6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7efde4ed35f6ddabcc8d9a2ac313e049700586993eb8ee06fd272c23f4563a4835b5ed7bc8ba40c423c91e5cfe6e13c9447cbf0a7bc08a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1255346e066ecb599ea621eaaf1775df6f8e0c8e9ac154f035b8a8233a195309d07ca659bd81e2f0ec38602df56fb99a7e7adf3c44afdb6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf2e0004fcf709289c29e2fccdc8d9cf96f9f97bfd22bcf3ff012ff1ce2cc8375819b25db476479980d9ac34b62db3386f038a47b65ac56;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h63632af41eca093babac85831ed8247d5468a80fa91fedb097ba34127a779febe8d09b526d973ff4c7c8172cd57bb4a0bac2c041aff80b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19b202973dea10d51c7695df0d3e95deaf9099e315abf862d6e5df42a3642780d9266153046eccaab47c492903461d33aa9e23841478eae;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11e3434a17f61cca5cb295046ec726b23fe1e35930a9cc0588c632afc6172123ab7e3afc1a016e81683c24e23ef9db8f1158295491a2ae0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1243e7f84415fb2d86067021d6a99be766f8955542002bca9f84735187f16b8dc97107bd7e19b1065aacb99b4ffff18a703464d3ebd9a85;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9b31f6eb9f7e1f7bfa6ce6f9095ee72291eb6a18f95eb8cfa24ce3beedd6792043f2200406564bb0a5530b4d2bde3c887e8d147b4655fe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6628af3b9ddc31211ba0fbbb9c7bf4a1d2e345850fbfc3b162d4f9f6cf0bcc0811a522923d66754453e9af3c7f5e1d0f7f16f00f8ba531;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10de9b377c874fd0ea01805fd0bc70f52a7478549326f1d797fd9cf547a1b5af2a40cc437b167da2c0d04b2c45e30738986c974705859e2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h67c0a5ff8ad215489fbe7b837dc3f5af169701d2a8c4911fedf7c8145f1c6311246fabe5a5d47ff78ff74f6e91129b98841eedc3c4a9cd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a62b15046de2a5ddd76c1b0274d3bb22abd874c0dc991b103fc9a09b143a3159c4ef94a4e227f705b86f4707c3d150d72434eab5421504;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19a65c5f488119d9a6d633c500b8c5150957a285307514bb5f3dbb0e5f4306db9228a72feed7226743f1b4e2f28dbce88a1ff3a8ded33f5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12e2dce1639b5eac48b70b8aae3c40254a8f3a81bfe71d59c7184202b4e877048f81737fa2782e58f826527cb31e4d5ed878ee9cf7e2e57;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a0214e2058b66ddf8b4a326e2e9b9a91c1e196af56827608bbfd8f33e0df3a2d3af37c1d0ae8ee6220043854c1c7a3d90adf03a4c410bc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he5181ac351862c921d5a09fa4910a5d29f29e84cd2d1781a7ba2fe3b03c21c06b81b32b655994f056ce811461328d1e4b3685870fd3c0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14ca0877798dd1b70c8eec58f4f4fc26efe1fde5a462bd0d6fac145ee86e61851324d81d832eb08c06353f6a1649f321fb2b957992e516a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14b86fad5f637e60d8e8b1e43b28cb5467dac128bc08a9473e092b36cae318542f813373c024ccd1a6da3712f950ef3e33eff26922e5097;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13bc5d30db4e17e226c42ba6832e55e22605c3c14255fd7a204b185270a49bc4ab9aa4afcbe81c0699967060779bef509d3ee1a96c03b1c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc69b9db1772471a551c53b15b8f887440391d53031094625557dff2f37cd88f0b4ae5883189a702d63b44f3ab767e6914bad662a4b5b2f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3f6836c81a8b574b637fa874dce592b411cb09445f8fb89767ccc2aeafa5ea2c3e841be16f3592b5bc6fdd0fa64a42c6a02e7617e3629d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h88bd937a92fed97423ed7a9102187379a6a0eb63353154b57784dab901d5207963c243d30582a4a33f8716055f4d20b0fcd284e2d3f59d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b39356b9727094efd77433c3d4b5a221127d05239d678e1db68b945538a9cffe00b05e90fc43bde12358bf50838f83ccec88f8b68e625e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h164f8f01572c56fa15aab2d2632b188304efc27e5610e2388fea4992cb176724c677cf5de5b4c00baf19a8eaccdf15e37e65e187d52eace;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb94040a519c19a0b517df5b1aca165c91039e1415762e45673ab5f77704609deac97399d179711c585b8f83dee63aef7a0d47960692433;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha10190a3280b3104f3ebd08817977c20ec25cdbe71aefacfde903f7713adc1689070e7a3c5f7a2446f6239bd4ff9a5b9148f0cb1704f55;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4ab6fc47765f3d87e4c674592966622f8ff44ef1678ba8ede8b4ab8ef8bcf68640ffb6e5397e13e5cff9441ba57631039db235ed4ac742;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdb93f32c522f3cfd3212734e2ac50ceba60d5484c7f951b74cd49d20ea150394135d25e44b5f2bb05a74116da096744ab48602e501df89;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdaae26980d0ac3884b464647c3249a4e3bc55532b73a690c55eb76a65e68979b337c8072773cc4a3e6d106d8fa6267aff64235fe6ea590;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c016e04a4a0a7e781eb39f485000e498fa8d32a02af6888deaa0b5116cdd0b78d8be8dfbc20962c76737f19d476ccdc459a849c34520e2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4f9c403ccb728e70373346b8b1d59f364f01f4382453d44e0bccf4eb4ac6624708d17dbf1ad3fa8d60a05598771caf8b7a023abaef744b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1063bf35181c512cbaa86bf12c1a87eba72746c29d43a5b57c4bf6ca76fd1956da5ba5500e00d30e90456453ac58a0ee41cf307fdad37e4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h187580ec35b50c7241201655d7793ffeaa1273ddcb2b9be464a590bee2a1c845635616ec5238069d2912dc71f833395417d5b17c1843170;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ce47f7ebd93bda99ba6a30966981644f4c00ff893dafafbaaccc2329ed198fcd10abb1c01ddaa246eb471bcef2f12abadb8787d38f3495;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h67661883a6a5686c6694f3c4f44fbcfe4845e24126815afcfe9d0752615629a0fe0f499a16a280c2da6c67d3a04b8b36fa95073c41d32e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf686b0e330e1050661ed2c95619841d62a097416fc7fb6e5ccb9daf71939261553da000981af7e616de0522180cf7cb70c2a5fce7a38af;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h58b3b9c41727668379d2ea5ebea56261ba283d5ab230f37e029502c9e1cd4df49dcdf18a710191876c10adf582b3e5b63f449c0dc06e54;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf22820c55e4b9b32fdb29d4908275a73f5e89b4f62469fb28e4b043fc2171931fa42457d3125cd8a9146180c6a07ea7264965619280a88;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h184b226f5b347e61d3cd9dfddc35aaaa40ced7068227e323212083183fd8758e567ef2ba0ad50323f052c5b77fc83c762f5bd017ba0e70e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcddd41f468f97bcf6fa778745af9ba1fb007c9082012cf0f8b5a0fd5e1fcd698ab30da556df8990a9240dccf42805baa8d4a432c92a08;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h524e54c26b3b2d81560e3f54f02f7b5dcff1bf4a1690f4e1a7659295a22c6e328c3532a83cd7e0cbbc5ea7361c76d15f6f1721de314ab0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6c079043bbb9599a2a6581682de7252be1ce88dc2ff3540653a02e583870a9914adfd2b2441d71c9cf6617d8d8a3ffb85de8fb44da7de2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13ab35aaf083a0c486ffa38964dd862491de084d927c57d47df1bcd45f454a13c6b4251bfafd4d805cf92777c2deeb6d65db3b5939f075d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h199d1847c28b0097c8c88f1284a218efc161cca5abc47f6ab7d4800522a6076357c352a6859071e137a18f86c43c8d4c3e499552d242d0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dd34c3fa5926c7c75d43fe6ee91a1b03d4b36d97bebba82341e45be5f015a182a4798ccb3ad7b09c3fff559970eeb28dfaa61c3ce69843;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h74e61fa46df09741fff9889c85947170407aec9349143138455010ebb9e3ec33001b18ba74507f67156898102bb07df5b2e1e8e7afa142;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heb0897a140b727513b89877efedc868cfcc14e9e326d8204f4545738db013852ab1aafd994876fb2b8bfeaf8b09e25244d48358fdf1788;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b3af4fa2d9f60faf6b605d7be42c29a2b35dbbfc790c461b34a8ca10b7640a1c374af44910c8d8ca9714cfe2f7fca044e23858c871f008;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10778ff57ddbcda021e5946a277565cf810129777cd9cc53d8fd5e77604f2140f4f30033a871e1792b4770517f4ebd8fa929598e2301acf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h167c69ddc90e387bd08fe72d5cbc532b2be75f134b0399c625b4a8ef0e62b89606ffb7af78ad9a1996e69beb8dd5274a29d1ca052514ecd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15603caa9be864e9117b2abcb2143b465243f72d8282ee9f9257e55c11e7b10b49fd21a06957d251eaf88f73c11e600101af4d6e37d6799;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1402f28e75cc26baa8d0a9c85e4ba918f62a7bd49062c07f63ce742c69afe0ee74208a6e4a304a4b82a6d0c038ba9ec934422a4d90c691c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h951893cc79706e54a5c54e1431cddf2692f3820489adaafe828b1aa934be910ffb0a7e5bcf9108fdcc7a476b5bc480024afa333f3b2d12;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c9bde1c718f626e7a30a194c09a2706c62c713526a555097ccef9cfaf310d2def826dbcb836faaee08743c7ae82e4e1259eda433fa687d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2e69d6d05f7489de84eca77f5fdf5c6f158d0be27e17b5a90cf945f896f9ba082113275abd1adaa157bae6c9bbef980370c0ff9d32adf8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha542fe8662391001dc9578acb5a5ec2ce50f8e9d3343c7f656a338d726ea43cf296b8f9a167da40c6d83945ea3d9fd79fefae3e5d966f7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h60ac590b0d58db1300db66520ce972840dd8222c17f8e47896a36f22abf4da5e3003cab6d576b71eb1edb077f876c47c18cff9964e9bff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11e1c306c49dfd2c0ca4206b45d9d44d75638b3bec47c99a0a09ca5e4ff4e25ae378897132ebcdce00d058d06ef0214280def3988e161d8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dbaa602634abc58ea21210f67f0bda30aa03b668db889ae49fd81c04a7d25611387902cd81ffc0ca1687128b3aab49ff523b831f9672b9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6d0a8eccce31ac894f2bd0e13eb837f67a2d88aa816f621c656cb2431c5a99afac7da7e14ff03288240eacdebcfb54df6f926f394d7614;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb5fe12e8cd8e0ded2e8c2db66dde99d64eb110d5469ba0062e088d5897ca08002004d1006c17a952bac096307b5e11ce60af1bd31d7d25;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1522d560b143ed0084bd3d43b547bc9f757a1527e2361f9244a62104f5e201a8a719383b0fefd0d4aa50eaeaa9f200a8f867034d2cab375;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h109941cc4eecf9332238d4ff52bd3b8b0712a2879788df47db9cef9d3e783a414b912f9b2129f8b1247f9d3fe9ed8b00a1d8b0d7212fac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12b4ee24a65e8940f2e6173f14fdcd2b4a864c49ee92d243b797dc827d48538f4f2651ca5c755af938496cccd4fcdfaf819c9b95910647f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h121088e51b6e1e939988b19dbf56f5edd2cb28f1a3b7241a5589542922d80f53311ddcafdf0f1b688abfc087670a065833b77c4a23294ee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hec31050ea0ccdad1843f908e321f50a81e9d7c1e40436a942fdee221df4b97d70cf202e7a34b85612888833d0c110dd5e43e8969b90ae;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haacbe5e7c7af36b5e7cf160de3b757105d1d3a0a7b91ce2a6454695e0c87164bf4393475eff32220967dbecc8d982fbefc395ce01f9308;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c400d6c4f620e084efc582de174a070965b2ff77328068360f44c3ffa38b406ce3439482169e810019c4f6faf381f5053dfd098888ee43;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1537a1fd74444be4e0a1d6133aff3743010b4d2e5004588bb210b526347fdecebedd34a6bc0ad266e04b12e408870c60247efd0f18fdfea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19b871b7024ff5d397e85a97b28cf6511360f7af8cc55761055022e80afd0f1d7abbf04d383459150a8a16e4d7a9406f9005a0752070905;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1264d9e3e439c4c172a949acb1a5fdbcd3f611dea5d3b716e3f10a08f63c9bde0c4ae797e5edd131bb539ddd6425559754454201f1241af;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a7b7a743fca4b26387265a023c0648e87f64ca69a6be778d479cbcf740283bc24e48fd66b72631774d410cb4aa11250cf179b3d10266ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h89acab0b474f39edce72290dacbb517c202c4f0f07b0fbde58da33b19befff8e648c3649ec3af2bf0cc28978678e4c8de020b8239a2e0d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h189db1fcb81c30c3b018cef3a0c34ab5796d1583c4b426b06dbcdef1acc011a0f124bef7ef8924b017b809adb4146e269e9ad71b68ca571;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10c69267049e3fa094dee1693712af79d9ad5f88b9f49d5bab7e14059920ef7d7690821186e3bdc1e109ccbd45829b2548883403dc85e1e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'had8fc475e1c9c30f467a27316a5d546a24e572242aaca5bc4808a61a6b7b2c4306046d5346d9aa559e068af21277ff4d4f3cd6ede5edde;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c46bb2077006648f5aa6667111c90ab50549bd6239f3a6254bfac5e243d29e7418704c5cec5898fece9478ea9f9d98033763383db2804f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15739ef46f2d8f41f49639bfad0c9751059d8660fae76fcf0f0484999ec57d36a681f1908107bc6ebe7bb1cf28857d93285e4379db47ac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h130ffec6779afb5ceafbf776de3d4ea76bd443f176930411f692966188218c635937bbaa9a2c83376d2d15c5ec55c2ac3b77209dc40678a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13ff09363bb0feed0eb12ecf5a333dff0d6010f25107f3b5a5e8c45fe0a02c83e6ebd32a72b81e85640bf129038a23d26e0acf128a74853;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf6d75c546bdc664d1a058280a0f78c8e66333527c6b8b5e439cb8c00211910df63f7e13bebe5ded17ac0fd092592b9891f0d82131c7b6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h78a6d5d73572176889cdbd996d9579c5488c968d33e615d3a57e48776ec38896b4cbc2c190e4e56ccdec9f1f116df4845318bd168c6e7b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18b708fe9a3387b5e32c82399e337883cf24b99e2c4da34b494b1b90fc1ed974e7b5e17b8f16c087c7c7384b785d7bedddd4d0f00b3c938;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h194df8e60f10a476291dfcbe1548e9d14daf4c5fc92a875c6dc732316c616c7021f44dd03ffc7d8fc825f99467afafa2cf396fba9bcd1e1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h74f959892a5af67b10ee1a185fcb676843d82a50150878341a46df789a0ca0daebfee5ac60fb01124d9d45b41d56a442914cb77fd65632;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h94e23237c08f2de6fe4e41ce7775adb6a4bbb787c3e9c71a95d7c3eddb4176f9ad463afce51573eb5e7711bc296e22fb9081cc31150ff4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9511f4aae6876e5969b7ad706b8e42e4ab2d2467f723ba5dd2f47ce2ec6353e0f853ae443aaf3163ab526f9bcffaa5b7521900d770d7dd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eb637eda2fa2b67935ea9ef76e95d1a734163bca2b6b268947198b058f205641056ac92926a2e0af770198025c0698c255c65586985bcc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h985fdfef39788850f787839e597e080a358c4140afed33136d0b4e9da0d121eeb07f396bc08fd97ec19ed499abea3b89cff1e40dea9ff5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bc996eaced799d849ec8656216beaa977c51a75e6554fe143764a6d2ba72015e6c62d5a07a229dcf04ee3b214a9262155cb06a636bd6bd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h160705047222a9f290e9db1255ada427c56bda95d6a51f32e3d850b700f030527e0f3274e9f62b676fbf3df52f3a7a29b080f36f95ee7a7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10227e9f00eae26e12aaf7c008d40cb0dc66b5a3699ff13310e822a2188b40c32a878e31e8b9346a4de93278710d4995f4a281d75499559;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc44e3c61a33e46df00cbe14bb00a1f8ec4deb7ff387f191a00b4cd75ae94825511a0891a5537f21b0d7e6094d585f583287fa4e412e833;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2e3ffac01d254eca25412778b6e91cac0f937cbb76e321e9fef2daa28f92b01df40fd7c868e2301d0df88f781e0a6b056b7b92e49fbc3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha8342a018f430fcdd6c18b78aa78e8c786066489f07eedcf4c9ff492207d6e7191cbd89ca691417c2de90923b7f2c2117545e854f0ac5a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8a55c19d1bfba14ecafd1baa5a0d20ec2f8d94607bb6149a743a9300971150c4cdeb883567ac510ce9575ca3c98c8cbfb5998bb92851a1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ca10377f77c0dbc0e3be77fe80c3beaab99b9fdd4e05a431a362ffe0fd70f09b3265fc33332eeadd265d6624959dff310ae47cbef50540;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h87237b1bc87c1a049bcf9b0946ab1bb43f3f7ae5d6ab1ffb02566e2a2ea4fb4a9def61daa19528681f4a786ece0c1e06b0dbcdba10b42f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19ff83611be4c5dc9b5406aed1552cf090e675e90d00e7fec86d2af5abf5f80b1bde9fe2114376ae9e52eee68844d9eaedc5ff45e1d8448;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16cc4e605c01b31c4c7925329968a10d7012b32dd06f14e005e8829f96c5b82d7b9dc1a0c506e55148d993eb866502cc5bf3e0bca5146b1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8ba81937846d60f1b635e70b46b032e78fd4fe87cc889d01fdd59116f12d68ecaddc8a7b660ab3d5c52cdc8053782cb9d4c512bf6e9c68;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbb62ce5b351aa56698d19b78e740391f401b0ae934c21d16f71cfdce15a2aa645b4057708037e1922ee312e38bb34582a437aea159d45b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h491e73d0933e5e8a31c8994c3bf37492cdcf75cc70fba05412ef50ba819df1950597db516fa12f69b85118912bfd02161a4b7509ef9718;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1efa03ecd94de5c5dd929d8c500a673dc83c7589028b38a4a23bf4d1a0214099e432ea438f93f3380f3936900534058eccba6ff751fd093;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he4ef7e14214e1c1309ebeaf93741e4a754222207b109b67f39360893e11a0eb6519f68d29ac89749b6222cc634b3d6802a27d934e4bc4b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5e2a78028ef8d5fbfc81a3e3168276b7c980c4f84176d8c12929c8b31b89f843076cd096a684c2031030b93bd1647c9a5ca7c9e79d6efe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1194f02e01568c6a78971d5666f12f8b3c0b36bac990ee8c270d6a8faf5e0799cc22c92914c14bf7858988b6966cb74d7248ac3cf9afbca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d1089abf6cbb9ded4e2bb383cfe9622282c6df30102f03592e38b876123d3582356c2b6daa9ed96cff1a9ca629435c9b0ab0837188dfbf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h116ed58ef6e315e0c6ab414716f608f02e2d4eac21961229c4c5cad7189d976b93744868ae609239b42e483e381cb847cf6ba9cf9e312fc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h322ebc97f5620a59846521ae09e6bf755465da705d30d57cddb22111857696c6b973e6bdc03a3a2d64815ce4afcaa7b4f77e456a2adedc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a1e46d5c0bb5ed03fbc4970cad0612ba1cec21736cd59c813b159080856cb45ed401a70c3054632c586b7fb9429619600f36364c2c9f1a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he74dcb5561605fc0ec659045c1e030867b3e5dca05a4c1fdeddc51ed4bc429afde53f8d1982399f15ff9cd0a3fddbd4c1c7227180bfb9e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h68e4234d1b167f817acf59e8b0c0fec794dd29aa4d792daa0aba861fb24f533a05d9aae9af3f22be05b860954dd31301c9d93418692097;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3dbc0eda5e5a4b46fdb01da708b413a141ac0ef7e37320174d62c884ef6f3fcacabd1832b643b4c952c9c5505412f4271b143555bc224a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h403474de3cbc73a04a653ca8cbe035b041f5cf74b00ce7ae09aa883e6a2edd491f1510edfe6c763e1ce77ec970e483ec0a2deabe0274a6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f078944b0366f2af38b03f62340e282d3d8c522efd21cb0fccf1b4ac9a639777ef5e9c98a5e3966c11deb53f0dd78bf25bf5dcf9d4a7ae;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e12a84859a6893a86e7a0ff4d61db476c7365bc6f73a032e34e9a0cb7a026aa61c58f439e3ec613dd8791c3a3d0b86c22fc031266c0e90;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7a0d6d33040afb7f6d5396d7d3750372a7945c804f65b61ae82a5baa5e2f45fac6d4ea9076542b22f0f03b8c06018e505a8771f7ea2ac7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10d044b467da2d4ac53efec638cd8390feb3bde6795bc6aff2dea1c09364aa20da9ff254730094089d88ab52fefd570622db9150f4eb39;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h186caf16329549ec4f6e4495e8b0f09617b33f2ecc67bed0e8b116e140dc3615397b734bc0ce077ed9dd6cb3c4a2a65cab8fea7477e0173;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he7e750f0a43178b2c93ac11cb8f1d063a44aa0a0b63db5a9de9d42aa4a34e0a91b24b035e790c09c4bd73725b12f5e84a77e2681aedf5a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12034e9dc44ded760b3ce6766156249f06659b9362f2ef768e3dd1fde7b41ec6b953efe9ce445de2a6443e7b6e3fd4c23c4da4d5b0bf642;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc15c2d098b7d354d6974c62509d28a68555d4d1f390a78beb9e080bcfc888eac292de8d6471c2e4f434cd35e592bdfec89dc70142a55c4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcb3477b44e178681fc3f717e7c37cdcc0876a70ec32ad39d73907e0b986bfedd58da76ad3b878cc58d9e5b8e7d76eabb5fd6429f3486db;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h143c19c2ca66e1c5f787d81049385fe3dcae6abbb9cfb4a213e382efe3476a69595a3206aa9b55412be8ef564ef369dfbeda643a0cc455a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd382144fb83ffcb99d8bc3243b39c50224f41b64cc57cd989ff3ff2879181cf68c354610d6c8570d9e9c0a3907701a113485995cf17fc0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h126bd3c763256d8ab277b51acd2f1d9252fb03d1f85496f0a9dda32a2dfbe2106974d74f3b81cf133bcbe3ac09848453f3b4514c26cdb1b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10aa26912e80ac1be769ae3e82c0c7ee9035af27c36d3232daac17e5283367b9859dfc480f93401a85c67cc9c5bcf696a8938f0495add7c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h867fd9902bd9301dbec28991a3d99196d7c4677fd8cafe7ef37a8737214de70575a5783e2d1b5ecc4359d91c2aff48bccf8566cdf17ac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7d4a60cbdc705a76a6f7c56ca2102f4c9469ab3844e92a6b6b9f89061799dcc1e2658ef1717d6ea4d24e2e8332b401846ebc0526e87a38;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8e68aedb0ccb7e845429001ac522d45b8a7e2c273f2ea3e0d22ca9881c4451e552d8d3358eff584ee6367f1495c36b5a2cb6ff7a20dd2f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hda8e0b28285e3e9fefedf02008ee717cde6f3335bd2106bb2c3dd31fcae06f45bda9393f6737c54a9bd9bc4b6b08826fec1740d66681c4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb0d9df5e0754ebb5582014d3a2d5f5bb42763f566b5e3b0ce084bc34fe04173f164c336ef2926cb3728eb5514884ed31ba9937e73398b8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eb9ee00ba71e5518ddbe68ea0e3a038914c21fdc1594f01de9ad46cec065596e61f9058f34fbe57a3fcdd872d032924c5e9e4e9e7914d5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc488414dc36e88251158d3e1c50a0d16f58023e19f67a3715fc787da59e0993a37552a7484d2fc8a6f72221c6445ac0eea24182faf1449;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb076d45237ca09a6aabe9406fa8afdda4599bcf294c19593824b3c635d73a10e3a0292cfd268c9cb7c6ffe789fe192c4464f21c2428e6c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10fc9a8e77e6bf32abec707778fed386e76a476f6e5957237cfc14a778657424d5bda85100ee65833aba7bf00199388c0dd4c417ef8fbe2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e398fdb0d30567125a2e87b3f3722236db651ca8a960b3881e7861f60e0384447a6895654267452959e14d4a351ab5d3b3b934b2002b7b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15af4e5fa21b1481141339d265d8e44d24c54bff70044c7c6988725788b4f608b67fdb0b07bc552b46983a99d0d1ee0369c3d081ecaebdf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c72c7f48633cdd63af12e615e9cbb9002e4d0e46e61cadabb92bcf4c5f0daee6666095e4f3b16e11675aaf12e4cc8eed6272c548e5f7ba;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbf72247dc29f235bb9c222ff764d014e887fb8abf156fa44a2255283917cdd9c03a885fcdc3ceadce47d0a2bad2cd4a39da73367c89ee3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ffdd01df88db1756baf14a7720fea9841ce9291cab04661d9c932b1ee5d3bd7c7ee91a58be5ce9faea66737a6f7a9576be1c3e7412ed69;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h163e05117b138e0e229e6526fc8df5ccede7e433a675459f024fa50a93c5a18e71ca587bd3c066514309d57191d99ef23e2ac109537b886;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h552963b8dbbfcca46dd4b823403bd7d8c8252ce313ba02bde0b6e04da735c4c8193b37e621f38360ade5f97212451db22dce30b2706a43;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ef1772d414505c95e5be7aa9418410ee8441bbd3000679ba9030d4cba9fea76a5cd1d185873b9faa8a018b136b338ddb84705a849796b4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h129ba97e86eb80406bece25d4bbe2efd32700b67c7c4f3d44d917fd0819a5b802d42b4eaf29fa4d4a6847ef426db0393d941b199609bad1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b27bd7e40cbb873c32336adf327f2efc6fb07420d7774d11f6a40e57cd597bc94f8d10f49fb0a107abb1290e52740eb6e1b139193a6abb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1511fceae5ffd44a18f68295a4c44a72c247f5ffbdc7cadfe3a3ff4a7ef133aade592cc1025a1dc8951c8b145130e93a57b79f3a62dea52;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12048e51a68ef3a4cf0c9d1467b2ae237b9115ad57d3c1d492c297fabf69220c74e7bd11d57eb089d2fa03cd4b97ed13fa741c67336f32;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ab103fb86273ae37f7de73546f00569db435aeb632398a2349449007a8ba6b064d95bf244515d24c1f90c8abc3b67121a27f3ded9efd35;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13e2c2db30684d4621204ebe6539ebd9bde6c368bb08f63f87846645ae05893eefe656be067a43cffbdcdf4f74055f6c01ab74c6946970a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d90473c7ccb459520f2f636dfadb12392e1e8f74240eeb30df7a4c04f0c84ac13b37bd2362a14db697ed2b2234b206d80d943f6c48da4f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hab9d7035f7c74ef1749e4002fabe248463905b4e6d7b66855189cd84e9ed24d249a919613685425da63dd90ef07a82dcf5d545f24bfe8e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h98dac934297514e73e497733db9097e1b2b9fab9d741eda2a311f32caebc2a2e8f01036fb605265f8bb457b776d3394693e7fee2f516cd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc3ef88e71822f0d375f08759c46bd6b45de031019c093e854f04ab04edb1f416a90f43cbad19dce19801d8f603cfa2f6c2687ac2848a7c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10638d756506c0dcc68565781407ea939339ec42aa6ccacea5ed4a572134eb7a4f45bd0b8dd12d7d014ff8acbe73834aa9ca1379a8b3d69;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h28b85eaced919edfed1998b367f53779b4f7af4bbc5f864308a09453c72dc76cd939aba1befccbb29dadf844a4c17da8473e0785309564;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e09098a3effd8bade6dac0eb3f811b29fc48a958546e9943eb3e866954faede7cca56c29672ad68cb2d9f9ee26f2642b5c650b77ba17a4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h170e85b8120e5c35c30a51ada6bc0435c5b1625a117fc32c5d4e47448208abb09cd585aed00d5c85b54f627253d095a57a5bf21ad619f99;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6e30d07c2d8e1d1266bccd86e32da1a1d61cf4bcaaff2ec9343367aa2f2cae4bdefa9f7be867804680db9c2901c1f24c55ea4e8d5b92ea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19c865bfa3de0eae6493578b9383a1df01ebf2383248ad11d8993917d08ec4993f42067438be322c0a841a60264433873000f39e99f1ce5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h33f5c1c15fca24865fc5c7856dbc3997a5d7e455ced114b8aa7fc15af3e5bbe09a6bc09f013373d22e0ead11ef2a8e19d1d0d8aedf0fb9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf7795b1323d8a5441f9fc4e3b6e2ed42df404ce8e6cfa4b7241db6532670d06910edfb56b0aebf4b1c441720d17a40f6cba42fcaaf087d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17c1d74a1c4e011846b94ca22043a513bb3ee83dc2edbe4b67f16eb4dbb3f8c3bfeb3ab88849512ca79545c6c4e6d3d2200126f4ae67b63;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13810e59f4a2df0a8740c4ab179a07401610d0546576a8bbaca0d8ca77990a5c3c7d4fec3bf02f0567fc7fea5376d4919d1a6cb214c46e6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heee0f97788fcf513021cb68cd83fa32c892ede2f65a120c58d498ded49ef2c01414fa664f51a3584269cf126ec3b4d8450239f48b4f606;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd757a711992595373a3a0acae05b237033a8ad81bf18270abfa7fd91d34df0a15dc0b95e3195c927a609730b5e1d16e3d4bb4411179e1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbc612043cb879623281570e48020fccd94e564185a48775e92a8acdfa87d0cb9627b139f92f9191965aa596307873ec3228fccdb3de198;
        #1
        $finish();
    end
endmodule
