module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [6:0] src8;
    reg [5:0] src9;
    reg [4:0] src10;
    reg [3:0] src11;
    reg [2:0] src12;
    reg [1:0] src13;
    reg [0:0] src14;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [15:0] srcsum;
    wire [15:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3])<<11) + ((src12[0] + src12[1] + src12[2])<<12) + ((src13[0] + src13[1])<<13) + ((src14[0])<<14);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hffffffffffffffff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h846fb6c0dbe21f1f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h942499f6d57d91d0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha33e99dd836f9aa5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb376b5c1ab61489a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7e15ea3f68cf8e6a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3a0a03fbd86ea1b4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf31a27358a742a3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haf0f46690b45446f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h14a63e63003dae71;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb984ba753c6ad5a0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4ad596f1a800f4ed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hacfc1e945502d7d4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3e1b6314fb64078;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdde130e32f4c193b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4a418087a1b6d213;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha3dc9b9f085f1198;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7fd026a5ada4d48d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5ca54ad2fbae594d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9c144f8c23bdb5ca;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h714a4fa85ff63a31;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdecc40500aeed68f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd994a2833a0ae711;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73f338deb74192b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hce1f0dfacfcda46a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he0050d345b467f33;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h79b3b2cb989a89e5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h964407f8f843423c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfcb2ece78bcfa1f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h40b01c8b89faa87;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h42375d55e24e9352;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4e0a9f9cd42fc78c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he9d3d1d215216469;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hddc39a9b25377ba9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3ed779079607509c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6a5898ab0b1cc4c5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f898c9c99094998;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h614ff917bb81d6f6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfc7e4732e386ba2b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h186b32d9c31ebf1d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha716d135f5a773ea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5178c9392d49740d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf07fae06cd835671;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha9c6f62b912b16d5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73f273e1059ba3c9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8992a4d1dc0004e8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8199745762de74fa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he857623cb8621836;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hecf10c3a514f3398;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h44a17bb33a1e2c22;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd78e05b5a52cd7b7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf08f50799fb8d999;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hefccc34c9e46619b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc62e90972ebcea2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heedfe65a64954eb0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c6acdb05a6cfcba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf94165ac2073f2c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he6e84241d77ee53a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h57732cf7407a382a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb3757b3c65269367;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf7821ade653664e0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h698cd95a5ef9da62;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8ed80e9bb00ade9b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h874fe1b90f579a7c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h68a45337477a7e46;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb1a39a78d04e5aa0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd37e7b76778c353e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h46e62b8cea270768;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72d306b072970ea6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5e1844bc6cc72460;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha6e016ec16799ac;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h65c163f682d2faed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc583c8eb77f23086;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb1b2a087a95f410;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h50e59090f9b399c7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf7a416b6d7b7495;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd9349069f1f8751;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h414dbef934bf748f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc775a311f989b15;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5af382db5656faf6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb5cf8ecea7a9154;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcfc7aab1e9b1f504;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8cbbaf4958618e77;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f1a17426b534664;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h854b7fbbcc479335;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd8e08553040c2317;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9583ef8d74bc1068;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdec283086f29ed94;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8017a3d4a7c7ee81;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hff1c917e70f85dea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h817fa5705546f272;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2644c896f7db6566;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h17cf7fb70d835459;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a137f8701f1e2f1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf33153a0a9db4504;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h456e334a9b35b72b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h82a87fbacf8705d2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd171f08393b3193c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d779fedf7925b60;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h614de4544de2d44a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4b8e62fc7e17fa8c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc414a97070a7f035;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4feb973030c61a94;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hca62a6b527c7f585;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4ced72705ad84a31;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h21f649694ca81527;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdac3c882cceb9e59;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha514db9f6484e911;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h56e8215fd51c2ce2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec7343161dd2408c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd385dce3dc6c819a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h68901d62dc47fc49;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcc37ef6a76be7fa0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2a7b163d9d61f4d8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5097ff98b23f6a0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h508d74614936e63f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc2f1f6ac2303f77d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbf23da13729441b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f42cd60f19f6ebd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9c469b26c5443840;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7fff8bfc2be6e773;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7e3a15936f78c61b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he2269a9e6cb63b8e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h720564d7710043ea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdae7cdad128671c5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hffb60882600efbeb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4f119e83a5df553;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h68b753a974f396ac;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf9bc587c593faf93;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h963e4364e867826a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h22686bfa168bf1ba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd9ebf6898e05d6d9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb3eaf01fe31adf15;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae56da3f1eb6cfc8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3e950a55969ec421;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h161ebc6640eeee66;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2f0cb2d75c643065;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1890b1630c1d8efb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h822088d16e27a158;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h245720b864c494f4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc9c3efc3db51d59a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3c21359b69970624;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4186168db2ae9ccb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2df8169ba799cac0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfebe92c2263f2719;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf119308e1e9a149;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hebcfa528eeea8719;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haa5c4046881a36ee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcbe69ae5916c125c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4b9d9776ff9a3fee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb3f5a2ed438dfe9e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h60aa1d7d8863229a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb42ce188718d6188;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h226ef8b765de4297;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6368f49d0f383d07;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf6c5670db56725e5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h89df595e5465868b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7c0a8019af287e0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heeb3a3f2ecea01f9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c64fed479d6ed76;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e9a7a59db97287a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h42230a59c32be1f4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h97361cdc036819d3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h949340727d737a2e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7eab22388ceb8631;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc5e7475403c3ef0a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hedfb8e4c70ce2ffb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hacac0d47dbef45d6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h86da923b2a82d400;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h418a1c567e68ed54;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb66cbbdeebf908;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc6f1145cf9d5c787;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h15a74a26259610f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc8c34916a3972b08;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h66e5ad562161af33;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hac48278a093e4eb6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd37ad551e197ef58;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h29d6d8dad7938c52;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hea13417c6de22498;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd04ca2f2bc95e311;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h74321cb47a99a643;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdd76399ce35498a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h79e1a6ed9dc0de58;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9ab495f6ebcc2f82;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4fc6422587fba018;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h902cd4c7a60d3aa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbf2092222d155761;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee306deff0cee568;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf16ff33d8c756ea8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h58ca72b6344ef471;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h246ee61b7da36fe7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha7da796b2ff4df80;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2c4e8e767c5988a8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he7e8629833372de3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5ddefe0f4915be08;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc9bfc9b83b61a103;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h247b2e97331e5f77;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5c8927194080a927;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h558119a3cafbb647;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haf8cbab87e02154c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73d708b7066fa8c7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7bf5591fa520235e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h23044e4a0c0f7d7c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h12b077a7fb79b4cd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9aa801d8991679a1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h23df0e2c9dffd32d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h11cb8cb30e3ceab;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h794bb6d66816c2e5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb51d7ed91f75dc5f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb02abe03d2fc56c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb256f27b5c798c71;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb068330b84626e1e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4efe2f2663475ca9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h56a6a93aa9e91983;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcc7a8f61890368e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5fe53e61320433cb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h29712d0f668d2899;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h40ecea7eb801a16d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4b2d8bd9151a7f8f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb08da7ab99395a12;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h29b2ab0609736cd2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hac145ec40fade2b6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9d443716259fffb7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc613d10f621db1f7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha4461ab580bf836a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he9d6974333da0f5f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf5f3798940aa805a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2466d8bb89e84083;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb1dc2b754f7daa43;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h437f7ee4f588e3dc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha054766bd20f39be;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6017a30ce2d1ecf2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb1dd489fe7557e30;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd09c6e26c3889613;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h903c720842bebe75;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h698bb46842d465f7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfaa4abc9062211d8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he4d9e3eb2b3188b0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf7cd6a6ca024f217;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h670d0f6572bd06de;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd07860d12f9be5a0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h76e68c9712d62541;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3807345764f9026d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6e781a078290e6c0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf97d922e4fea50bc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha749ce5d4104a552;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6aeb9cc0f1bfe6ce;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h987ad0623503376e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7c90d033ddd8cb41;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a8cb942eb3847d8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc08600405ce6d636;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he0b1ec061d3dac15;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h55d5f980fddd4121;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h773618a25fbe2e2f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h591291dd50580ce3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1f44bd839492a84a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5214828276adda42;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd07f947682f16ce5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbd624743369bbee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h23fbb60b426ef70c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbdffc2f53c575808;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hecf6083a86c5e56;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha5c22aa540d358ae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ac79ccc760c86f9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3066ea67eb38f138;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ebd58002ad0e468;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5d367722995e6e1a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he8c3c58e2951a8e8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf0498d8d1ff15a42;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h178263720a8bbb92;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb140830d59ef6f09;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc9aa7908faf0e092;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd603796c1393b961;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb523f8e3ed36277c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5f87df9259138b02;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf06361cfffc1f9f7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc50daa040b74a810;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2fb93742d2e1ace5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2764287fd6ffe0a2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h510f2d4850174fa3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd113c8a73dc9f6cf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec33143badf5e394;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hedac5116c5db61bc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c57717073de180c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7aa4d313d2df3104;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha1ae02c545f4c83f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h486282fd084c11e9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae459a003a4b33a1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h832fd96332422fb3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h27eb95414f66255a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he5c3082d09f9ff56;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f6bcbd08b36e8c5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc291c8318f59979f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h70d2137ecabad198;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9af2d426703172b2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf4aace16965cfc53;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5d62cf4df7496631;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he2c0b389f21d93da;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5fe67e88b38c51f9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72b31b77a748ca3b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hce9523a4c17588ca;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6214d98bd5a3a8c8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h57af2df56b301243;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h419d1dd55c3aefbb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h717dfff376544161;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h953c7487b118b52c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfe18c811758bb06e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h68a12a41e1bbaa74;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc454b1c1e8b727d8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hac221860375eccd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3e6bc1fc1e94fd39;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h78a8b747104ba507;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdd094d509e8ce743;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6f62a0b4e392e7ac;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73f7ca7536846434;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6d4460b8a5d6ca23;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc498df4d29dc8b3c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h25f3e709958007f9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2f2203a57919db63;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h89b32bfb44124bd7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9c0afe6e84b649d0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7e155dfd505d3844;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha67ff059af40f2b6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcabf360090c3130d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hca83a9648d9de6e8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h792cb4964ef8ff25;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc5909a67ee15c503;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h412990eb90a53764;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc9f51c3b10e57a66;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h77305bc69df6c895;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9d9aa7365c6f2020;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc4aa68b4efad4f9e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb6114148fed93ef;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h97a13df31bfde32e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h55aed1456f1b553e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h53ee361e3cd28a5e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5220b32d7c3c2950;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd480c2428385a46b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h53d35270ce934bcd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha524be55d5da0679;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he673792f0ef70926;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h833a2c082d55c4de;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcdd675991fe2c56c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h392c7f529db1ccca;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h83fcbe6fe11db182;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5170abe77d47b6b7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h794a90293ee610d8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h155d95621b773906;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b84476ea290a53b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3a82f37388763be;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he65a6356a95854ff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1e788774b294c31a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h730532aab247c116;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h76972f7b82281406;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4229d3ad7c3041cd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h217e6481aac121b5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h61ed5804c17bfce5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha5e4c5a6117b4958;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haaa11656df9eb4a2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h89b3702e598cbcc2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b2306d08112e3e3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1d355e214cd2ca78;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hca49ea330c3197f1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec3445c5d006b522;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdba48baaa2fbcad6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h87bb0d7e6c86864b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h205fe11819acf819;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd963f33990d4ebe5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2cd4f119673c9fb8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2bfcf666f8543e89;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h589eed1f31a53a39;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4c5d41f99b77706d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9650bb87aed76659;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h41c65881279766ce;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7261b7f0f7303f64;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1447ecaae698aa16;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hecf11e2f69fd95e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd71aae66fc844a71;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd221797e9fa80bbc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6872eae2b154844e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he9cfadb088c18ff9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1809f2817f98e099;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h61147e97c7ac8bc8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b793f53888115aa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h88a13e4d0a2a6a63;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hed5d6f3fdba505d3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b365355b64d83d0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h47696c95623af31c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf4c5d7de425d16fb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf666295e7ad8705f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5d0eddb4b44c0ad5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h31be05d70af429eb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6e515d3c1bfb73bd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h480bea1394662819;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha4d22ba23fa34af8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5650efe3e1cc66c6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb3a7e61021871587;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf658a71e09773372;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h983ad44683395df8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd74cf9dd3ed0aa7d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ee08416baa5ec3b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72efa3dde5621edc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h99a958419d8fd738;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdbc85bf71dd0c64c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6afb93ef20a75df2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4b54b4e702aa4f55;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h45452eacec9ac13a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h12a5d52edc9c094;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he3d734556dc08398;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha9597231d3a6ee97;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2e5d872a5081f554;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6ba9c5ce816ca635;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hed19431c32696df8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h65b30ef896229dc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfde1755c9bf09b5d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h542d7af2e6ed4ef4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h371442b9c6412ece;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd9538e5c06d71d6e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haa8c954d31fe7a62;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha6759c5e81000927;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h991cbbd4f07f9fbf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd54db642fe309ef9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1883aceebe0baa6f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haf74a3fe56d469d2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'habfb4d6a20effcc2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1809ad69174ad682;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef18ea2e8f3d9632;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3837b3dd2f02e898;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf80efd36d4c8ca25;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h231cf7324f41565b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6a87862ceb627b69;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he0828881c12134ed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he0bb9011a62c1c91;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc94f6fce6cbe397b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf86c47cb55baaf01;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha469c97c856d5774;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f75a93ef67b319c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha269f1557d65a65;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2d481f234042262d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f273477d33f4851;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h70d5891acf16b98;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h58ad0faef754ad78;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3ec0463a0bd84cba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf9b63bb6678bcc36;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h67dddf39f8b11035;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h83325a1481dc3ee2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h906e63fb33890fa7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c4eacbaf0d1a98a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha45325250867658f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8680661e55924f7f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha8a539a64ad30b20;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b64ad675cf5d5b2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h403b0ae2e8bc21da;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5490397a8574b3db;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2c9c21c827e0fa7d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfd24a1e18ba5e444;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hab394f13b4e0da55;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2a25fcd796efbe20;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb742936e87564dd8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf743595db062fe7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hed7158849b06805a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc151f39d96b4965f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd3a7c878a04f0c99;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h194e530047aaaf8e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb8cd6596f7c83822;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb3c5a0584a47495d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7f1716bd1e2f171;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb35a76444b2512;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h31866debf7f7735d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h15584e17d1ad3dee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6c95a80820db3f30;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h10b5c0e2c71d417d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h80f1cb619b683508;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h293d397c2c9a8db3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h89f1a945b8aca3c4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b2999f481771a48;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1d374f405804f93d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he448830103b4d6e3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf17234ce8af078a5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9905c126e81108b8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h70bc2079148e3fcd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2653eb72d47c3844;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h81613a7165a4c031;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he7c360e6b9f9a418;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4729c5dad91f97e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hebb6c3f0b52086b5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hccb1797486d663c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h25ff90f29120f873;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc6f472332c57dd9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb1c1da6826e0d4dd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h206baa95cb5fa3f8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb3bae87aef5249e4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha4b7062d720315d2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd3e087ac7090bb2e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6091be69d2fcfd84;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b79d9f9ffad7efd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb89a05cff8f55dd1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4d21992d199894ad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha224adeb9add9cf2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd81e22c158fcbcd2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he059fa638eceebeb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h589edaecb5931fb0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6c95fb2667474501;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73e6d8cc8d7b6901;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h489a5b78253beff3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hefb9287c65400ea4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3c891356601e1167;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8001a0822ea382d8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9654a742535347f0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2d8dced2086d5683;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2fbd6d15fbc1a4f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8444cc0773c6e8ba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h85b9cdc2ee60b3b6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h418f30ec72ce8a9b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h29e8a5342d24b0c6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf04d98b8d81cb518;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9ba05216e6bfe969;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6f7c06e01ec23b77;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3c9fc89ad484b5c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h49ef041325ffa4f9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h39108ff9d47c52fc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h15236f57ec1c9e55;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb3e758c9d84cede;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h105925d3e7367ba9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h81f21a790a71bdc1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc9c4fb47436155e2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha2290786c4a8cd4c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hffa34fb18849bb2e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h679d40288f7a746d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6c1b1cb125b329ba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha7a02aa7611377bb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'had3ebd3709eb3458;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcabbdb2b61573f45;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a9d522a8c823925;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcb665eae17903edc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb6d77cad06174845;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c9b249bc4dcd411;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5dc71acccc56b48e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcf5ad1b920418f6c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb28cf6948df537dd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h77f196da0ba021fb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hebdf14c72a05a01a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6506f5a63cddb036;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h64ed48a035e72a0c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hce8cd7096003d6db;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcc4940e9eb6b26b7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2ae6dea639649c5e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb6d4b825118c881e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h695ab041593dadd6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee1611e150f8abba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcb9e54e6b6de8344;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h719a2d03a6f764e7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h314130883a732b19;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8252b30e2fc1044d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha09159ac27cdef;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd15f68cf333ce2d1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h761cf25d77614fdc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd79bee78750f3505;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h68b9e4f90bc5c0d6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h274af7045c943783;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hda05bbefeea7acf6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h232844a36f35f431;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf45410852bf55db1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb1816312cd745db8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3a384f2a89094d37;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hacd5f26eab3014c7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h60b0f3ba17fee9e5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd6b8734a15826c4c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3b451d3200c29f2e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1471addfc855d811;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha142b889e2564b94;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7d3c01fd388e23ae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6acba54241b26e19;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8541deb30bede440;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he4dc2237695cd6e2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7df1ea273621732e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1803f205868e4a3f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3119be5dd810ecef;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h82820e598a68943e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4a3306e4b2d3d48b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2426f75764947ef9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6593b8e03e72a53c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcd2af5c36fdd9c8c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h723ef601593a1173;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h104d66bda692e475;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2783d0808b08236f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haf9198e5c663008b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf2348c29b5873c69;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha8cda2bd03220f32;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2716cd9df8eb27a8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc6076f6aa4b336b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8bc0fac553944992;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h17263f327e845c8b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h534d31cd91283ddb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbcd890888327e4ac;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1365b3509fbf3447;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h34aa0eb0ede1fad7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h29ebd13f27d8198b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1182283f80e9524;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b9d6a477762a8b5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h93455286ae79138b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3c25c95c1404ce75;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb66cc17bdaf96f2d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h503e3f7a284c16d7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h12a76de313ff4855;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd9ef6e44a98f5487;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hddd3f4eb9582030b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc2c8f10daa890383;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc91177f3e856c972;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9238d38e329c414f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h911b25d740c87c0d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h384435f9beb4eb63;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7c537cf466c95dd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h77ff625ccb83151;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2d57a490c3b2e934;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h27e5047d90e2da09;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h448063519ef2ad3b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h602ab2665d74b511;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdcd5273268213cbb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h74376aab1b42ff7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6749f27cfefca750;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h61221075eb045b3e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h16016a3adb33df26;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd1772675d1dc796f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heaeb05cf75cd2c38;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hecfa68da76ee7ac;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc359bc0ade2a2a34;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f34451f421ff689;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4c27bbf00e9640f1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h548ed08f76a98415;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb6606b7b48a49c4a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4970f19dea8d24ca;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h477d6bfba0fcd643;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcf57807a28b49980;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1f178d21c587dd72;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha4a3c255155d1a31;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcbdd3dfc2334df8f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb001618a175d5ab;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb69aa516ee67ba5a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd5c005bbd9aa1a4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb12f6d1b54a551cb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heaffa1ac838ca8b9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'had8d4d5cb13e7658;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb19d144a66a5a160;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h42d9c29d4ebd8544;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h665431d7f7a4d42d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a70afa1fb4d92e8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a69c02f0dae8300;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4af567b65e3cf2d6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb4be1897edc8829c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc29e0ea78d7aa4da;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4a4fd210c615da44;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd55895d787d6deb8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4638425d6cadd56f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1a48f149504cdec3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h527808cd7a507f0a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7493d1e889001b3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1567c9031337931d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5051129a5df9801;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6f0d445f27251cd9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9627693ff9de1593;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha59f1b1a42ac2b16;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he8d82b30417ff1ea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h61dc44e976410f53;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9cf166c5c1e18cfe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h28d116e94083e14;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7a0825023cdb2b01;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb0a82a5866135047;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6957be21b108c6e5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc7be1f9a10236a01;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h207ece8c9cec846c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f9a78bd287885cc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h32d7f7523bd16ee3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he42b23ec6f77ba73;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha630353a2dc87d25;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd6f77b0c1e32235d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heee77e90cad42995;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha62f764a8a1c3a3f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7088244d48fd3d0b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb0faadca78699bfd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'habe610656dddc8c5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c5833f865bc16fe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h43957e08ea372ce4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h21eac7700579f4f9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h464886fb6620e082;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h348d6bb9bf96862;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd56d9bb380f983a8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2a70abae67f02a7e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he64401c8d5a6ba1a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc65998865e371c59;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h700ff26d169cf3c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h678a7fe7857768c3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h30ddf2b96f4def6a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h50ae5bdd712467fc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he9b7f55dbf96159c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h89e6e1f43f4be3e7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h43af210dcc5bc18;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbce7b3c5a506b0e4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h303e6a86800d49db;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h587229b6b195446e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6b7a720b5cc1c672;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf5ab568a37af0f0f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a1335eb65423cf6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2638b9356340d9c9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcc166f31d5d07eec;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h947b26c62862390d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4f2cfd744cb3fb81;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a52842fd273dde0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha2117aa28fd62dcf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c4f340502f8328b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbf16f3b1aceb0188;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haf5d6bfd0ee82dc9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1f7e1e550b5eb738;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h197b4d01d4060452;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha00f3559b47ac7a7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4d86afc3e0af4b56;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb2f1aeeda7b7a6d5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hada648ebe6d52197;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hea017f828178245;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd9768d835488b049;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3efd43883b3c0517;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h61c6edb260cbca53;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf04ac17adb2bd7b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h718d99955aebf992;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h20f4efedd27a3b4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h492b5214b3ae4f5f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9951116a28a1d2be;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h11860dd4fb80a968;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha88f023b736624a3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h601ce79766163010;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h34fe07f09c500084;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7c33e1098b0fb958;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3db4af2efc200a79;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc7c1f765ee50dd34;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9ab133ebf0e006de;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h81148e613bdff019;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha38a363a781a7bd5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4add9f14f4f0dc9a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4acd69e6ee882372;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1fb5d0918a4b73a8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hedc8dd35dad3f32e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d6f1f264733113f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h67a6b80032b62d1b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd4e9615eab6f48d6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8b389253f7d3fff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2d45e08949131081;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae390f6938fa51c3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcf31947b0162b49b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf487deb936d3a02c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he42cb2f38950963d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5854f1a18442feed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6ec40c0908242d5f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h54c1cbc38d598f8e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h40d9ff28295c7094;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d66c45017b2936;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4de951bb02607c9f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b71053451105143;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfef9927ac8e13599;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h182b5b3edc0d178;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h365c8fd19f41d833;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h555f983e87ca15e4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b79b2e1a6030d5b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb25703286dac9e77;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ab6ade89129d7d7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2794777d042ae061;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2cbdd064d9616c90;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4624da09d3049a62;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdd7ad9b5020a4bd7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h31ef9b581d1482fa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haeaee6f5397e02f7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf7ca236f7c04a5d6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf3f8cc214de90e00;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7d6438e3d04bc590;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc1557c35903ba17d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha8a4f04155b57187;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h55d90aec49e48bcc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hda77b39032af6da;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf662b1aa7454e44a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2726c8d07e94dffb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha22c571bc7069597;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d71f37480d55165;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h91b1a84f5278ba70;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h21f2769faa5b1e48;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc32f6787db8b9c5e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h19da58697bd8e708;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h69ee93f15e8e395a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he3440dc1c198b9fc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd678e16b0661b761;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb94837073e9e45c1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h903a8b65ebd2fe15;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3de7ce8e4d87ca1c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc262211b71b0ce08;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hea037a8dd4be2842;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h355754bc8aecf48d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5db102a855415a9f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf39a76704878039c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3e9455386ab4c0e3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf45b1600d3b13149;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h36b5043e6e7f819b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h422bba2bd8250036;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h585d04b65fe5bc23;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4737dbfd6749b366;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b32892498c9dcb9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfb6cb956c808c77f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc2d33e82a39f52a7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h422a56f84b0ef464;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h183c0c842767b1a2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf4bed013029c449e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hba279cda2ddba58b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha62633197aa0f394;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc47a1d732a535243;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfbb344bf3b3c0433;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb46c6f66b940f60d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h689f16ba9d662710;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef0071380ef689dc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h78aac6cf0bdf5489;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb17e3ad488d91c79;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h765accc4b392c518;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h50ed954741103a03;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc8953f5159fdb80;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h35fbd4178bb317d3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h659ed049c0c30c43;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h182d7ab5b0c5178b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcd9cd6a4cf5e89e4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd8cdcae0f252c4d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3e929d1948fecafc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3801e01af91fa937;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5d6b4370d88d5149;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4b5b1a11cf45319d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6c65bcf0b8460589;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf1413ca053852dc6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbcd4a1462a71c30f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h236180a5f2b47023;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde8ccd463d2db76;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha7f82381f5279c38;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h560f05f53a04e2bc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c5e4ddebdfffe52;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf985066d9c4c3583;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he75f4b0c02b6910d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h987666c170f78831;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hca37efddf183859f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ee455a0884081d6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h999948cba4b55ec;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec67b076a9ee9b45;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h75c0a27e2c3d98e2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h44353590ae082a85;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf14229c179f3540b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h172522023c64c5b4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8b18d85ff6cc974d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4bdd332e6a84df0c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1e4de12b807a69f0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3b7aa1cfe12ac1d1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6af0cdf6bada09ff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7e97cc02ad4c0280;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2615f1944f8de2eb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3bd7eb8a21a1a10b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he3ff570046654ace;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h31818cf03d8e5997;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf3cc3530b3491624;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf7f63bda2f4ae80f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae98de6df6eb26a4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h52d8660ee7769f7f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb7ed4102d455b66;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hac820399bf8cd3c7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h75326b730f5c5b97;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h85fa37d50bd02857;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6f36a308d31ed74;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h93965340de1ee81e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h53d244dd61dbff84;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h31878d77b1d49bfa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h92c7896acbcaa363;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbdf83db5757fe353;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcefebddfcba0969e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb4139d91a4e23f76;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h31e277321129ea78;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3e0bb401696875b1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7112379e42e23139;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3ce39f51e4775d4c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf581c3bdbd783c6a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h54a3ff55ccffbb5d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdbba2ee4089867f1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4decf888dfc21754;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h32bff162225abd25;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f4a9a101df5e6a4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4672b4abb177aa60;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf6407e30be6d77dc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c3d110efb73b847;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6cf6472a5d1ed915;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6ba28ccd97339c8b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h587bd2aeafae2536;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbeaabb23f884d787;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc2657f20aa6a3373;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc865bcde56282b9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h826d1d5bdf9fc9af;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb6fdd60abcf4b3c3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d45d3060b2c74a9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h29c22c464d66e3df;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h83c089cdbace411f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7dc1f31ea85186ee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc7fd7c47eba5b85e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h715569fc38c8fd2b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h482cd3570920272e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7a3f7d347b6e9b80;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha1b18904386ee909;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'had326856aaa84423;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h59177d775fd6273c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h81804023882d72da;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5b29d1a5b5a6a973;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h46a57d119d55f3f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h91ffbe6c184b78cb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5d6055bedc7a769e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd02c199da1eab742;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h11572ae3d807422f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h77e8f8f68da5a2b4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h574eebcd6b56b9f4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h15c6a4da89147c2e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb68acdd69d2b944f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he5851aa80e4b1bb1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5fbf2a584a3dc288;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h300a02baef14a954;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f6da1f0ff3baf6f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc5b7ad073011ab6e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1fd2f9931e235ded;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc69f4a732930980;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9be30cccb5e54791;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he3030246840ce93d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b4f5453bf91a5bf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf2535f5103049236;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h550a38433ff4338e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h189815d658625c5d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee1f02872923ac91;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha1c6ec02604a0809;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h12050a7e5a4bd5fb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd53af42840b8c085;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfb9d4589e9e04bc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb456311978b0619d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9cbdd8c2426b7f03;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2aab80b0218407dd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7eb58f91e1b4bd08;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h670e1970b9991fd1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb79a0538f64e5178;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h20b845e63fb18303;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h606ff570d1c48b82;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4ecbb92695b1c8c6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc2d19efaf58c347d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf4fe5ac756f7bbb6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h404ed61d233fa17f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9ff2fc8e032247c5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd35d4676f4246587;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he46eae5128547429;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b6424ba37edea72;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7068891885fd5e36;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbb43e525e411ae24;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4e1423d44ee50941;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c7bf98875711950;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8577eeec9db293ab;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h86d4d761ab73488e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hce887d4727e1351d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he79a3fb8bc6489ba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde1f398b5c134b1b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h27690c88d0957713;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd57f8b5633f670ce;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc77c78fac6fd1483;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9eb9c237278e9832;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc862759741799a79;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hceb2d1b663796892;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'habf5f8f6089b584e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h57c3d9cf7d7b5a4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h45af5ba2f05bb5ec;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h33534e13186aedf4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf2b5d7e639936345;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9bba404589e4ccd9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5ab694b8c1ffe82d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h17c57653e5704f05;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8de81eae8abca8ed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3cb43922287d32f6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4dafa257a848524a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4db5744fd599c19a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h41ab1f3ed18a2fcf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb6e21337febcbab2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72755e2e217c79bf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he5efe82435ed22e4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb77c6813b8f2fb69;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h32ed8d6d3b0f5332;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h667e3ff89557362;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf890dfc071f4b8b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc1dc7809da1d46b7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1166897e08ecd994;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd734b5aba4bb6162;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h54313b963888439c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h608aa3b85c80d76e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3fe280582b8573cd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2d06670d9456e101;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcc47c4d9e90a4573;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb4101b99d6dc6996;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha159e6aea31caaa9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h315783f30e887b08;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h20852aae656958ad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h627f53f8a75dee11;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2480f53b694f5609;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf405681cbf96c280;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h84aa852059ad34a9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5450a0b8a5a22888;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b36450cee3423bc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h66a9a80cb4f18504;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h47b0bd3b24fdf4b0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h96b4ab589a9a32d9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc11d9a8136e5ff5e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7f8df57a093c1b7b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h119a3dafe680aade;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd1cd765bfee92cfb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h610bfcf71f8a2aaa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b44ae38392858c9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he4273b2f96c418a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4481eaa1b1868bb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h768344a5468ff36c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae9406e3dc6f2b64;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h76d6d10e8ffd5760;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hce1decaef686e708;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h68b4760041f6a539;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdde5a655fd7ca1e6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbe63ce5e369b1ca0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he92af53488077887;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfeb3ef65a272ffc2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heddd5336ed3bcb37;
        #1
        $finish();
    end
endmodule
