module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39);
    reg [161:0] src0;
    reg [161:0] src1;
    reg [161:0] src2;
    reg [161:0] src3;
    reg [161:0] src4;
    reg [161:0] src5;
    reg [161:0] src6;
    reg [161:0] src7;
    reg [161:0] src8;
    reg [161:0] src9;
    reg [161:0] src10;
    reg [161:0] src11;
    reg [161:0] src12;
    reg [161:0] src13;
    reg [161:0] src14;
    reg [161:0] src15;
    reg [161:0] src16;
    reg [161:0] src17;
    reg [161:0] src18;
    reg [161:0] src19;
    reg [161:0] src20;
    reg [161:0] src21;
    reg [161:0] src22;
    reg [161:0] src23;
    reg [161:0] src24;
    reg [161:0] src25;
    reg [161:0] src26;
    reg [161:0] src27;
    reg [161:0] src28;
    reg [161:0] src29;
    reg [161:0] src30;
    reg [161:0] src31;
    compressor_CLA162_32 compressor_CLA162_32(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39));
    initial begin
        src0 <= 162'h0;
        src1 <= 162'h0;
        src2 <= 162'h0;
        src3 <= 162'h0;
        src4 <= 162'h0;
        src5 <= 162'h0;
        src6 <= 162'h0;
        src7 <= 162'h0;
        src8 <= 162'h0;
        src9 <= 162'h0;
        src10 <= 162'h0;
        src11 <= 162'h0;
        src12 <= 162'h0;
        src13 <= 162'h0;
        src14 <= 162'h0;
        src15 <= 162'h0;
        src16 <= 162'h0;
        src17 <= 162'h0;
        src18 <= 162'h0;
        src19 <= 162'h0;
        src20 <= 162'h0;
        src21 <= 162'h0;
        src22 <= 162'h0;
        src23 <= 162'h0;
        src24 <= 162'h0;
        src25 <= 162'h0;
        src26 <= 162'h0;
        src27 <= 162'h0;
        src28 <= 162'h0;
        src29 <= 162'h0;
        src30 <= 162'h0;
        src31 <= 162'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
    end
endmodule
module compressor_CLA162_32(
    input [161:0]src0,
    input [161:0]src1,
    input [161:0]src2,
    input [161:0]src3,
    input [161:0]src4,
    input [161:0]src5,
    input [161:0]src6,
    input [161:0]src7,
    input [161:0]src8,
    input [161:0]src9,
    input [161:0]src10,
    input [161:0]src11,
    input [161:0]src12,
    input [161:0]src13,
    input [161:0]src14,
    input [161:0]src15,
    input [161:0]src16,
    input [161:0]src17,
    input [161:0]src18,
    input [161:0]src19,
    input [161:0]src20,
    input [161:0]src21,
    input [161:0]src22,
    input [161:0]src23,
    input [161:0]src24,
    input [161:0]src25,
    input [161:0]src26,
    input [161:0]src27,
    input [161:0]src28,
    input [161:0]src29,
    input [161:0]src30,
    input [161:0]src31,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [161:0] src0,
      input wire [161:0] src1,
      input wire [161:0] src2,
      input wire [161:0] src3,
      input wire [161:0] src4,
      input wire [161:0] src5,
      input wire [161:0] src6,
      input wire [161:0] src7,
      input wire [161:0] src8,
      input wire [161:0] src9,
      input wire [161:0] src10,
      input wire [161:0] src11,
      input wire [161:0] src12,
      input wire [161:0] src13,
      input wire [161:0] src14,
      input wire [161:0] src15,
      input wire [161:0] src16,
      input wire [161:0] src17,
      input wire [161:0] src18,
      input wire [161:0] src19,
      input wire [161:0] src20,
      input wire [161:0] src21,
      input wire [161:0] src22,
      input wire [161:0] src23,
      input wire [161:0] src24,
      input wire [161:0] src25,
      input wire [161:0] src26,
      input wire [161:0] src27,
      input wire [161:0] src28,
      input wire [161:0] src29,
      input wire [161:0] src30,
      input wire [161:0] src31,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38);

   wire [161:0] stage0_0;
   wire [161:0] stage0_1;
   wire [161:0] stage0_2;
   wire [161:0] stage0_3;
   wire [161:0] stage0_4;
   wire [161:0] stage0_5;
   wire [161:0] stage0_6;
   wire [161:0] stage0_7;
   wire [161:0] stage0_8;
   wire [161:0] stage0_9;
   wire [161:0] stage0_10;
   wire [161:0] stage0_11;
   wire [161:0] stage0_12;
   wire [161:0] stage0_13;
   wire [161:0] stage0_14;
   wire [161:0] stage0_15;
   wire [161:0] stage0_16;
   wire [161:0] stage0_17;
   wire [161:0] stage0_18;
   wire [161:0] stage0_19;
   wire [161:0] stage0_20;
   wire [161:0] stage0_21;
   wire [161:0] stage0_22;
   wire [161:0] stage0_23;
   wire [161:0] stage0_24;
   wire [161:0] stage0_25;
   wire [161:0] stage0_26;
   wire [161:0] stage0_27;
   wire [161:0] stage0_28;
   wire [161:0] stage0_29;
   wire [161:0] stage0_30;
   wire [161:0] stage0_31;
   wire [49:0] stage1_0;
   wire [55:0] stage1_1;
   wire [55:0] stage1_2;
   wire [75:0] stage1_3;
   wire [94:0] stage1_4;
   wire [53:0] stage1_5;
   wire [105:0] stage1_6;
   wire [65:0] stage1_7;
   wire [53:0] stage1_8;
   wire [76:0] stage1_9;
   wire [92:0] stage1_10;
   wire [66:0] stage1_11;
   wire [55:0] stage1_12;
   wire [85:0] stage1_13;
   wire [68:0] stage1_14;
   wire [59:0] stage1_15;
   wire [106:0] stage1_16;
   wire [63:0] stage1_17;
   wire [81:0] stage1_18;
   wire [66:0] stage1_19;
   wire [60:0] stage1_20;
   wire [79:0] stage1_21;
   wire [81:0] stage1_22;
   wire [90:0] stage1_23;
   wire [66:0] stage1_24;
   wire [77:0] stage1_25;
   wire [54:0] stage1_26;
   wire [66:0] stage1_27;
   wire [77:0] stage1_28;
   wire [74:0] stage1_29;
   wire [62:0] stage1_30;
   wire [97:0] stage1_31;
   wire [44:0] stage1_32;
   wire [18:0] stage1_33;
   wire [10:0] stage2_0;
   wire [16:0] stage2_1;
   wire [16:0] stage2_2;
   wire [34:0] stage2_3;
   wire [40:0] stage2_4;
   wire [27:0] stage2_5;
   wire [30:0] stage2_6;
   wire [33:0] stage2_7;
   wire [32:0] stage2_8;
   wire [31:0] stage2_9;
   wire [45:0] stage2_10;
   wire [38:0] stage2_11;
   wire [23:0] stage2_12;
   wire [44:0] stage2_13;
   wire [36:0] stage2_14;
   wire [33:0] stage2_15;
   wire [43:0] stage2_16;
   wire [36:0] stage2_17;
   wire [28:0] stage2_18;
   wire [27:0] stage2_19;
   wire [37:0] stage2_20;
   wire [27:0] stage2_21;
   wire [33:0] stage2_22;
   wire [43:0] stage2_23;
   wire [34:0] stage2_24;
   wire [30:0] stage2_25;
   wire [30:0] stage2_26;
   wire [32:0] stage2_27;
   wire [29:0] stage2_28;
   wire [32:0] stage2_29;
   wire [36:0] stage2_30;
   wire [35:0] stage2_31;
   wire [40:0] stage2_32;
   wire [23:0] stage2_33;
   wire [6:0] stage2_34;
   wire [1:0] stage2_35;
   wire [6:0] stage3_0;
   wire [9:0] stage3_1;
   wire [9:0] stage3_2;
   wire [22:0] stage3_3;
   wire [8:0] stage3_4;
   wire [11:0] stage3_5;
   wire [16:0] stage3_6;
   wire [18:0] stage3_7;
   wire [17:0] stage3_8;
   wire [18:0] stage3_9;
   wire [14:0] stage3_10;
   wire [14:0] stage3_11;
   wire [14:0] stage3_12;
   wire [17:0] stage3_13;
   wire [16:0] stage3_14;
   wire [15:0] stage3_15;
   wire [12:0] stage3_16;
   wire [16:0] stage3_17;
   wire [16:0] stage3_18;
   wire [11:0] stage3_19;
   wire [17:0] stage3_20;
   wire [14:0] stage3_21;
   wire [22:0] stage3_22;
   wire [12:0] stage3_23;
   wire [16:0] stage3_24;
   wire [16:0] stage3_25;
   wire [11:0] stage3_26;
   wire [12:0] stage3_27;
   wire [22:0] stage3_28;
   wire [10:0] stage3_29;
   wire [13:0] stage3_30;
   wire [16:0] stage3_31;
   wire [15:0] stage3_32;
   wire [16:0] stage3_33;
   wire [15:0] stage3_34;
   wire [4:0] stage3_35;
   wire [1:0] stage4_0;
   wire [5:0] stage4_1;
   wire [5:0] stage4_2;
   wire [10:0] stage4_3;
   wire [5:0] stage4_4;
   wire [3:0] stage4_5;
   wire [5:0] stage4_6;
   wire [7:0] stage4_7;
   wire [6:0] stage4_8;
   wire [7:0] stage4_9;
   wire [7:0] stage4_10;
   wire [9:0] stage4_11;
   wire [8:0] stage4_12;
   wire [4:0] stage4_13;
   wire [5:0] stage4_14;
   wire [9:0] stage4_15;
   wire [6:0] stage4_16;
   wire [12:0] stage4_17;
   wire [8:0] stage4_18;
   wire [11:0] stage4_19;
   wire [5:0] stage4_20;
   wire [5:0] stage4_21;
   wire [8:0] stage4_22;
   wire [6:0] stage4_23;
   wire [7:0] stage4_24;
   wire [8:0] stage4_25;
   wire [8:0] stage4_26;
   wire [4:0] stage4_27;
   wire [8:0] stage4_28;
   wire [5:0] stage4_29;
   wire [5:0] stage4_30;
   wire [5:0] stage4_31;
   wire [10:0] stage4_32;
   wire [7:0] stage4_33;
   wire [8:0] stage4_34;
   wire [3:0] stage4_35;
   wire [2:0] stage4_36;
   wire [1:0] stage4_37;
   wire [1:0] stage5_0;
   wire [3:0] stage5_1;
   wire [4:0] stage5_2;
   wire [3:0] stage5_3;
   wire [1:0] stage5_4;
   wire [4:0] stage5_5;
   wire [1:0] stage5_6;
   wire [6:0] stage5_7;
   wire [2:0] stage5_8;
   wire [2:0] stage5_9;
   wire [3:0] stage5_10;
   wire [5:0] stage5_11;
   wire [2:0] stage5_12;
   wire [2:0] stage5_13;
   wire [5:0] stage5_14;
   wire [5:0] stage5_15;
   wire [1:0] stage5_16;
   wire [5:0] stage5_17;
   wire [4:0] stage5_18;
   wire [2:0] stage5_19;
   wire [3:0] stage5_20;
   wire [4:0] stage5_21;
   wire [1:0] stage5_22;
   wire [3:0] stage5_23;
   wire [5:0] stage5_24;
   wire [1:0] stage5_25;
   wire [3:0] stage5_26;
   wire [3:0] stage5_27;
   wire [3:0] stage5_28;
   wire [5:0] stage5_29;
   wire [2:0] stage5_30;
   wire [1:0] stage5_31;
   wire [2:0] stage5_32;
   wire [4:0] stage5_33;
   wire [3:0] stage5_34;
   wire [5:0] stage5_35;
   wire [3:0] stage5_36;
   wire [0:0] stage5_37;
   wire [0:0] stage5_38;
   wire [1:0] stage6_0;
   wire [1:0] stage6_1;
   wire [1:0] stage6_2;
   wire [1:0] stage6_3;
   wire [1:0] stage6_4;
   wire [1:0] stage6_5;
   wire [1:0] stage6_6;
   wire [1:0] stage6_7;
   wire [1:0] stage6_8;
   wire [1:0] stage6_9;
   wire [1:0] stage6_10;
   wire [1:0] stage6_11;
   wire [1:0] stage6_12;
   wire [1:0] stage6_13;
   wire [1:0] stage6_14;
   wire [1:0] stage6_15;
   wire [1:0] stage6_16;
   wire [1:0] stage6_17;
   wire [1:0] stage6_18;
   wire [1:0] stage6_19;
   wire [1:0] stage6_20;
   wire [1:0] stage6_21;
   wire [1:0] stage6_22;
   wire [1:0] stage6_23;
   wire [1:0] stage6_24;
   wire [1:0] stage6_25;
   wire [1:0] stage6_26;
   wire [1:0] stage6_27;
   wire [1:0] stage6_28;
   wire [1:0] stage6_29;
   wire [1:0] stage6_30;
   wire [1:0] stage6_31;
   wire [1:0] stage6_32;
   wire [1:0] stage6_33;
   wire [1:0] stage6_34;
   wire [1:0] stage6_35;
   wire [1:0] stage6_36;
   wire [1:0] stage6_37;
   wire [1:0] stage6_38;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign dst0 = stage6_0;
   assign dst1 = stage6_1;
   assign dst2 = stage6_2;
   assign dst3 = stage6_3;
   assign dst4 = stage6_4;
   assign dst5 = stage6_5;
   assign dst6 = stage6_6;
   assign dst7 = stage6_7;
   assign dst8 = stage6_8;
   assign dst9 = stage6_9;
   assign dst10 = stage6_10;
   assign dst11 = stage6_11;
   assign dst12 = stage6_12;
   assign dst13 = stage6_13;
   assign dst14 = stage6_14;
   assign dst15 = stage6_15;
   assign dst16 = stage6_16;
   assign dst17 = stage6_17;
   assign dst18 = stage6_18;
   assign dst19 = stage6_19;
   assign dst20 = stage6_20;
   assign dst21 = stage6_21;
   assign dst22 = stage6_22;
   assign dst23 = stage6_23;
   assign dst24 = stage6_24;
   assign dst25 = stage6_25;
   assign dst26 = stage6_26;
   assign dst27 = stage6_27;
   assign dst28 = stage6_28;
   assign dst29 = stage6_29;
   assign dst30 = stage6_30;
   assign dst31 = stage6_31;
   assign dst32 = stage6_32;
   assign dst33 = stage6_33;
   assign dst34 = stage6_34;
   assign dst35 = stage6_35;
   assign dst36 = stage6_36;
   assign dst37 = stage6_37;
   assign dst38 = stage6_38;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc2135_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage0_3[4], stage0_3[5]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc2135_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[3]},
      {stage0_3[6], stage0_3[7]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc2135_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24]},
      {stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[4]},
      {stage0_3[8], stage0_3[9]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc2135_5 gpc5 (
      {stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[5]},
      {stage0_3[10], stage0_3[11]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc2135_5 gpc6 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_2[6]},
      {stage0_3[12], stage0_3[13]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc2135_5 gpc7 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39]},
      {stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[7]},
      {stage0_3[14], stage0_3[15]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc2135_5 gpc8 (
      {stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_1[24], stage0_1[25], stage0_1[26]},
      {stage0_2[8]},
      {stage0_3[16], stage0_3[17]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc2135_5 gpc9 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49]},
      {stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_2[9]},
      {stage0_3[18], stage0_3[19]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc2135_5 gpc10 (
      {stage0_0[50], stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54]},
      {stage0_1[30], stage0_1[31], stage0_1[32]},
      {stage0_2[10]},
      {stage0_3[20], stage0_3[21]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc2135_5 gpc11 (
      {stage0_0[55], stage0_0[56], stage0_0[57], stage0_0[58], stage0_0[59]},
      {stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_2[11]},
      {stage0_3[22], stage0_3[23]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc1163_5 gpc12 (
      {stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_2[12]},
      {stage0_3[24]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc1163_5 gpc13 (
      {stage0_0[63], stage0_0[64], stage0_0[65]},
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_2[13]},
      {stage0_3[25]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc1163_5 gpc14 (
      {stage0_0[66], stage0_0[67], stage0_0[68]},
      {stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_2[14]},
      {stage0_3[26]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc1163_5 gpc15 (
      {stage0_0[69], stage0_0[70], stage0_0[71]},
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59]},
      {stage0_2[15]},
      {stage0_3[27]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc1163_5 gpc16 (
      {stage0_0[72], stage0_0[73], stage0_0[74]},
      {stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65]},
      {stage0_2[16]},
      {stage0_3[28]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc1163_5 gpc17 (
      {stage0_0[75], stage0_0[76], stage0_0[77]},
      {stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71]},
      {stage0_2[17]},
      {stage0_3[29]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc1163_5 gpc18 (
      {stage0_0[78], stage0_0[79], stage0_0[80]},
      {stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77]},
      {stage0_2[18]},
      {stage0_3[30]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc1163_5 gpc19 (
      {stage0_0[81], stage0_0[82], stage0_0[83]},
      {stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83]},
      {stage0_2[19]},
      {stage0_3[31]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc1163_5 gpc20 (
      {stage0_0[84], stage0_0[85], stage0_0[86]},
      {stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89]},
      {stage0_2[20]},
      {stage0_3[32]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc1163_5 gpc21 (
      {stage0_0[87], stage0_0[88], stage0_0[89]},
      {stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95]},
      {stage0_2[21]},
      {stage0_3[33]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc1163_5 gpc22 (
      {stage0_0[90], stage0_0[91], stage0_0[92]},
      {stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101]},
      {stage0_2[22]},
      {stage0_3[34]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc1163_5 gpc23 (
      {stage0_0[93], stage0_0[94], stage0_0[95]},
      {stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107]},
      {stage0_2[23]},
      {stage0_3[35]},
      {stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc606_5 gpc24 (
      {stage0_0[96], stage0_0[97], stage0_0[98], stage0_0[99], stage0_0[100], stage0_0[101]},
      {stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29]},
      {stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc606_5 gpc25 (
      {stage0_0[102], stage0_0[103], stage0_0[104], stage0_0[105], stage0_0[106], stage0_0[107]},
      {stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35]},
      {stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc606_5 gpc26 (
      {stage0_0[108], stage0_0[109], stage0_0[110], stage0_0[111], stage0_0[112], stage0_0[113]},
      {stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41]},
      {stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc606_5 gpc27 (
      {stage0_0[114], stage0_0[115], stage0_0[116], stage0_0[117], stage0_0[118], stage0_0[119]},
      {stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47]},
      {stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc606_5 gpc28 (
      {stage0_0[120], stage0_0[121], stage0_0[122], stage0_0[123], stage0_0[124], stage0_0[125]},
      {stage0_2[48], stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53]},
      {stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc606_5 gpc29 (
      {stage0_0[126], stage0_0[127], stage0_0[128], stage0_0[129], stage0_0[130], stage0_0[131]},
      {stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59]},
      {stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc606_5 gpc30 (
      {stage0_0[132], stage0_0[133], stage0_0[134], stage0_0[135], stage0_0[136], stage0_0[137]},
      {stage0_2[60], stage0_2[61], stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65]},
      {stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc606_5 gpc31 (
      {stage0_0[138], stage0_0[139], stage0_0[140], stage0_0[141], stage0_0[142], stage0_0[143]},
      {stage0_2[66], stage0_2[67], stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71]},
      {stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc606_5 gpc32 (
      {stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113]},
      {stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41]},
      {stage1_5[0],stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32]}
   );
   gpc606_5 gpc33 (
      {stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119]},
      {stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47]},
      {stage1_5[1],stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33]}
   );
   gpc606_5 gpc34 (
      {stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125]},
      {stage0_3[48], stage0_3[49], stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53]},
      {stage1_5[2],stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34]}
   );
   gpc606_5 gpc35 (
      {stage0_1[126], stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131]},
      {stage0_3[54], stage0_3[55], stage0_3[56], stage0_3[57], stage0_3[58], stage0_3[59]},
      {stage1_5[3],stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35]}
   );
   gpc606_5 gpc36 (
      {stage0_1[132], stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137]},
      {stage0_3[60], stage0_3[61], stage0_3[62], stage0_3[63], stage0_3[64], stage0_3[65]},
      {stage1_5[4],stage1_4[36],stage1_3[36],stage1_2[36],stage1_1[36]}
   );
   gpc606_5 gpc37 (
      {stage0_1[138], stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143]},
      {stage0_3[66], stage0_3[67], stage0_3[68], stage0_3[69], stage0_3[70], stage0_3[71]},
      {stage1_5[5],stage1_4[37],stage1_3[37],stage1_2[37],stage1_1[37]}
   );
   gpc615_5 gpc38 (
      {stage0_2[72], stage0_2[73], stage0_2[74], stage0_2[75], stage0_2[76]},
      {stage0_3[72]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[6],stage1_4[38],stage1_3[38],stage1_2[38]}
   );
   gpc615_5 gpc39 (
      {stage0_2[77], stage0_2[78], stage0_2[79], stage0_2[80], stage0_2[81]},
      {stage0_3[73]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[7],stage1_4[39],stage1_3[39],stage1_2[39]}
   );
   gpc615_5 gpc40 (
      {stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85], stage0_2[86]},
      {stage0_3[74]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[8],stage1_4[40],stage1_3[40],stage1_2[40]}
   );
   gpc615_5 gpc41 (
      {stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91]},
      {stage0_3[75]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[9],stage1_4[41],stage1_3[41],stage1_2[41]}
   );
   gpc615_5 gpc42 (
      {stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96]},
      {stage0_3[76]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[10],stage1_4[42],stage1_3[42],stage1_2[42]}
   );
   gpc615_5 gpc43 (
      {stage0_2[97], stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101]},
      {stage0_3[77]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[11],stage1_4[43],stage1_3[43],stage1_2[43]}
   );
   gpc615_5 gpc44 (
      {stage0_2[102], stage0_2[103], stage0_2[104], stage0_2[105], stage0_2[106]},
      {stage0_3[78]},
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage1_6[6],stage1_5[12],stage1_4[44],stage1_3[44],stage1_2[44]}
   );
   gpc615_5 gpc45 (
      {stage0_2[107], stage0_2[108], stage0_2[109], stage0_2[110], stage0_2[111]},
      {stage0_3[79]},
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage1_6[7],stage1_5[13],stage1_4[45],stage1_3[45],stage1_2[45]}
   );
   gpc615_5 gpc46 (
      {stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115], stage0_2[116]},
      {stage0_3[80]},
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage1_6[8],stage1_5[14],stage1_4[46],stage1_3[46],stage1_2[46]}
   );
   gpc615_5 gpc47 (
      {stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121]},
      {stage0_3[81]},
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage1_6[9],stage1_5[15],stage1_4[47],stage1_3[47],stage1_2[47]}
   );
   gpc615_5 gpc48 (
      {stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126]},
      {stage0_3[82]},
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage1_6[10],stage1_5[16],stage1_4[48],stage1_3[48],stage1_2[48]}
   );
   gpc615_5 gpc49 (
      {stage0_2[127], stage0_2[128], stage0_2[129], stage0_2[130], stage0_2[131]},
      {stage0_3[83]},
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage1_6[11],stage1_5[17],stage1_4[49],stage1_3[49],stage1_2[49]}
   );
   gpc615_5 gpc50 (
      {stage0_2[132], stage0_2[133], stage0_2[134], stage0_2[135], stage0_2[136]},
      {stage0_3[84]},
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage1_6[12],stage1_5[18],stage1_4[50],stage1_3[50],stage1_2[50]}
   );
   gpc615_5 gpc51 (
      {stage0_2[137], stage0_2[138], stage0_2[139], stage0_2[140], stage0_2[141]},
      {stage0_3[85]},
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage1_6[13],stage1_5[19],stage1_4[51],stage1_3[51],stage1_2[51]}
   );
   gpc615_5 gpc52 (
      {stage0_2[142], stage0_2[143], stage0_2[144], stage0_2[145], stage0_2[146]},
      {stage0_3[86]},
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage1_6[14],stage1_5[20],stage1_4[52],stage1_3[52],stage1_2[52]}
   );
   gpc615_5 gpc53 (
      {stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150], stage0_2[151]},
      {stage0_3[87]},
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage1_6[15],stage1_5[21],stage1_4[53],stage1_3[53],stage1_2[53]}
   );
   gpc615_5 gpc54 (
      {stage0_2[152], stage0_2[153], stage0_2[154], stage0_2[155], stage0_2[156]},
      {stage0_3[88]},
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage1_6[16],stage1_5[22],stage1_4[54],stage1_3[54],stage1_2[54]}
   );
   gpc615_5 gpc55 (
      {stage0_2[157], stage0_2[158], stage0_2[159], stage0_2[160], stage0_2[161]},
      {stage0_3[89]},
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage1_6[17],stage1_5[23],stage1_4[55],stage1_3[55],stage1_2[55]}
   );
   gpc615_5 gpc56 (
      {stage0_3[90], stage0_3[91], stage0_3[92], stage0_3[93], stage0_3[94]},
      {stage0_4[108]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[18],stage1_5[24],stage1_4[56],stage1_3[56]}
   );
   gpc615_5 gpc57 (
      {stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98], stage0_3[99]},
      {stage0_4[109]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[19],stage1_5[25],stage1_4[57],stage1_3[57]}
   );
   gpc615_5 gpc58 (
      {stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104]},
      {stage0_4[110]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[20],stage1_5[26],stage1_4[58],stage1_3[58]}
   );
   gpc615_5 gpc59 (
      {stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109]},
      {stage0_4[111]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[21],stage1_5[27],stage1_4[59],stage1_3[59]}
   );
   gpc615_5 gpc60 (
      {stage0_3[110], stage0_3[111], stage0_3[112], stage0_3[113], stage0_3[114]},
      {stage0_4[112]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[22],stage1_5[28],stage1_4[60],stage1_3[60]}
   );
   gpc615_5 gpc61 (
      {stage0_3[115], stage0_3[116], stage0_3[117], stage0_3[118], stage0_3[119]},
      {stage0_4[113]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[23],stage1_5[29],stage1_4[61],stage1_3[61]}
   );
   gpc615_5 gpc62 (
      {stage0_3[120], stage0_3[121], stage0_3[122], stage0_3[123], stage0_3[124]},
      {stage0_4[114]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[24],stage1_5[30],stage1_4[62],stage1_3[62]}
   );
   gpc615_5 gpc63 (
      {stage0_3[125], stage0_3[126], stage0_3[127], stage0_3[128], stage0_3[129]},
      {stage0_4[115]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage1_7[7],stage1_6[25],stage1_5[31],stage1_4[63],stage1_3[63]}
   );
   gpc615_5 gpc64 (
      {stage0_3[130], stage0_3[131], stage0_3[132], stage0_3[133], stage0_3[134]},
      {stage0_4[116]},
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage1_7[8],stage1_6[26],stage1_5[32],stage1_4[64],stage1_3[64]}
   );
   gpc615_5 gpc65 (
      {stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138], stage0_3[139]},
      {stage0_4[117]},
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage1_7[9],stage1_6[27],stage1_5[33],stage1_4[65],stage1_3[65]}
   );
   gpc615_5 gpc66 (
      {stage0_3[140], stage0_3[141], stage0_3[142], stage0_3[143], stage0_3[144]},
      {stage0_4[118]},
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage1_7[10],stage1_6[28],stage1_5[34],stage1_4[66],stage1_3[66]}
   );
   gpc615_5 gpc67 (
      {stage0_3[145], stage0_3[146], stage0_3[147], stage0_3[148], stage0_3[149]},
      {stage0_4[119]},
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage1_7[11],stage1_6[29],stage1_5[35],stage1_4[67],stage1_3[67]}
   );
   gpc615_5 gpc68 (
      {stage0_3[150], stage0_3[151], stage0_3[152], stage0_3[153], stage0_3[154]},
      {stage0_4[120]},
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage1_7[12],stage1_6[30],stage1_5[36],stage1_4[68],stage1_3[68]}
   );
   gpc606_5 gpc69 (
      {stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125], stage0_4[126]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[13],stage1_6[31],stage1_5[37],stage1_4[69]}
   );
   gpc606_5 gpc70 (
      {stage0_4[127], stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131], stage0_4[132]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[14],stage1_6[32],stage1_5[38],stage1_4[70]}
   );
   gpc606_5 gpc71 (
      {stage0_4[133], stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137], stage0_4[138]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[15],stage1_6[33],stage1_5[39],stage1_4[71]}
   );
   gpc606_5 gpc72 (
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[3],stage1_7[16],stage1_6[34],stage1_5[40]}
   );
   gpc606_5 gpc73 (
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[4],stage1_7[17],stage1_6[35],stage1_5[41]}
   );
   gpc606_5 gpc74 (
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[5],stage1_7[18],stage1_6[36],stage1_5[42]}
   );
   gpc606_5 gpc75 (
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[6],stage1_7[19],stage1_6[37],stage1_5[43]}
   );
   gpc606_5 gpc76 (
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[7],stage1_7[20],stage1_6[38],stage1_5[44]}
   );
   gpc606_5 gpc77 (
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[8],stage1_7[21],stage1_6[39],stage1_5[45]}
   );
   gpc606_5 gpc78 (
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[9],stage1_7[22],stage1_6[40],stage1_5[46]}
   );
   gpc606_5 gpc79 (
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[10],stage1_7[23],stage1_6[41],stage1_5[47]}
   );
   gpc606_5 gpc80 (
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[11],stage1_7[24],stage1_6[42],stage1_5[48]}
   );
   gpc606_5 gpc81 (
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[12],stage1_7[25],stage1_6[43],stage1_5[49]}
   );
   gpc606_5 gpc82 (
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[13],stage1_7[26],stage1_6[44],stage1_5[50]}
   );
   gpc606_5 gpc83 (
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[14],stage1_7[27],stage1_6[45],stage1_5[51]}
   );
   gpc606_5 gpc84 (
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[15],stage1_7[28],stage1_6[46],stage1_5[52]}
   );
   gpc606_5 gpc85 (
      {stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[16],stage1_7[29],stage1_6[47],stage1_5[53]}
   );
   gpc606_5 gpc86 (
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[14],stage1_8[17],stage1_7[30],stage1_6[48]}
   );
   gpc606_5 gpc87 (
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[15],stage1_8[18],stage1_7[31],stage1_6[49]}
   );
   gpc606_5 gpc88 (
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[16],stage1_8[19],stage1_7[32],stage1_6[50]}
   );
   gpc606_5 gpc89 (
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[17],stage1_8[20],stage1_7[33],stage1_6[51]}
   );
   gpc606_5 gpc90 (
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[18],stage1_8[21],stage1_7[34],stage1_6[52]}
   );
   gpc606_5 gpc91 (
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[19],stage1_8[22],stage1_7[35],stage1_6[53]}
   );
   gpc615_5 gpc92 (
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58]},
      {stage0_7[84]},
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage1_10[6],stage1_9[20],stage1_8[23],stage1_7[36],stage1_6[54]}
   );
   gpc615_5 gpc93 (
      {stage0_6[59], stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63]},
      {stage0_7[85]},
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage1_10[7],stage1_9[21],stage1_8[24],stage1_7[37],stage1_6[55]}
   );
   gpc615_5 gpc94 (
      {stage0_6[64], stage0_6[65], stage0_6[66], stage0_6[67], stage0_6[68]},
      {stage0_7[86]},
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage1_10[8],stage1_9[22],stage1_8[25],stage1_7[38],stage1_6[56]}
   );
   gpc615_5 gpc95 (
      {stage0_6[69], stage0_6[70], stage0_6[71], stage0_6[72], stage0_6[73]},
      {stage0_7[87]},
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage1_10[9],stage1_9[23],stage1_8[26],stage1_7[39],stage1_6[57]}
   );
   gpc615_5 gpc96 (
      {stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77], stage0_6[78]},
      {stage0_7[88]},
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage1_10[10],stage1_9[24],stage1_8[27],stage1_7[40],stage1_6[58]}
   );
   gpc615_5 gpc97 (
      {stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage0_7[89]},
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage1_10[11],stage1_9[25],stage1_8[28],stage1_7[41],stage1_6[59]}
   );
   gpc615_5 gpc98 (
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88]},
      {stage0_7[90]},
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77]},
      {stage1_10[12],stage1_9[26],stage1_8[29],stage1_7[42],stage1_6[60]}
   );
   gpc615_5 gpc99 (
      {stage0_6[89], stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93]},
      {stage0_7[91]},
      {stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83]},
      {stage1_10[13],stage1_9[27],stage1_8[30],stage1_7[43],stage1_6[61]}
   );
   gpc615_5 gpc100 (
      {stage0_6[94], stage0_6[95], stage0_6[96], stage0_6[97], stage0_6[98]},
      {stage0_7[92]},
      {stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89]},
      {stage1_10[14],stage1_9[28],stage1_8[31],stage1_7[44],stage1_6[62]}
   );
   gpc615_5 gpc101 (
      {stage0_6[99], stage0_6[100], stage0_6[101], stage0_6[102], stage0_6[103]},
      {stage0_7[93]},
      {stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95]},
      {stage1_10[15],stage1_9[29],stage1_8[32],stage1_7[45],stage1_6[63]}
   );
   gpc615_5 gpc102 (
      {stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107], stage0_6[108]},
      {stage0_7[94]},
      {stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101]},
      {stage1_10[16],stage1_9[30],stage1_8[33],stage1_7[46],stage1_6[64]}
   );
   gpc615_5 gpc103 (
      {stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage0_7[95]},
      {stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107]},
      {stage1_10[17],stage1_9[31],stage1_8[34],stage1_7[47],stage1_6[65]}
   );
   gpc615_5 gpc104 (
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118]},
      {stage0_7[96]},
      {stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113]},
      {stage1_10[18],stage1_9[32],stage1_8[35],stage1_7[48],stage1_6[66]}
   );
   gpc615_5 gpc105 (
      {stage0_6[119], stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123]},
      {stage0_7[97]},
      {stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119]},
      {stage1_10[19],stage1_9[33],stage1_8[36],stage1_7[49],stage1_6[67]}
   );
   gpc615_5 gpc106 (
      {stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101], stage0_7[102]},
      {stage0_8[120]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[20],stage1_9[34],stage1_8[37],stage1_7[50]}
   );
   gpc615_5 gpc107 (
      {stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage0_8[121]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[21],stage1_9[35],stage1_8[38],stage1_7[51]}
   );
   gpc615_5 gpc108 (
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112]},
      {stage0_8[122]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[22],stage1_9[36],stage1_8[39],stage1_7[52]}
   );
   gpc615_5 gpc109 (
      {stage0_7[113], stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117]},
      {stage0_8[123]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[23],stage1_9[37],stage1_8[40],stage1_7[53]}
   );
   gpc615_5 gpc110 (
      {stage0_7[118], stage0_7[119], stage0_7[120], stage0_7[121], stage0_7[122]},
      {stage0_8[124]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[24],stage1_9[38],stage1_8[41],stage1_7[54]}
   );
   gpc615_5 gpc111 (
      {stage0_7[123], stage0_7[124], stage0_7[125], stage0_7[126], stage0_7[127]},
      {stage0_8[125]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[25],stage1_9[39],stage1_8[42],stage1_7[55]}
   );
   gpc615_5 gpc112 (
      {stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131], stage0_7[132]},
      {stage0_8[126]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[26],stage1_9[40],stage1_8[43],stage1_7[56]}
   );
   gpc615_5 gpc113 (
      {stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage0_8[127]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[27],stage1_9[41],stage1_8[44],stage1_7[57]}
   );
   gpc615_5 gpc114 (
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142]},
      {stage0_8[128]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[28],stage1_9[42],stage1_8[45],stage1_7[58]}
   );
   gpc615_5 gpc115 (
      {stage0_7[143], stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147]},
      {stage0_8[129]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[29],stage1_9[43],stage1_8[46],stage1_7[59]}
   );
   gpc615_5 gpc116 (
      {stage0_7[148], stage0_7[149], stage0_7[150], stage0_7[151], stage0_7[152]},
      {stage0_8[130]},
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage1_11[10],stage1_10[30],stage1_9[44],stage1_8[47],stage1_7[60]}
   );
   gpc615_5 gpc117 (
      {stage0_7[153], stage0_7[154], stage0_7[155], stage0_7[156], stage0_7[157]},
      {stage0_8[131]},
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage1_11[11],stage1_10[31],stage1_9[45],stage1_8[48],stage1_7[61]}
   );
   gpc606_5 gpc118 (
      {stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[12],stage1_10[32],stage1_9[46],stage1_8[49]}
   );
   gpc606_5 gpc119 (
      {stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[13],stage1_10[33],stage1_9[47],stage1_8[50]}
   );
   gpc606_5 gpc120 (
      {stage0_8[144], stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[14],stage1_10[34],stage1_9[48],stage1_8[51]}
   );
   gpc606_5 gpc121 (
      {stage0_8[150], stage0_8[151], stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[15],stage1_10[35],stage1_9[49],stage1_8[52]}
   );
   gpc606_5 gpc122 (
      {stage0_8[156], stage0_8[157], stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[16],stage1_10[36],stage1_9[50],stage1_8[53]}
   );
   gpc615_5 gpc123 (
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76]},
      {stage0_10[30]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[5],stage1_11[17],stage1_10[37],stage1_9[51]}
   );
   gpc615_5 gpc124 (
      {stage0_9[77], stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81]},
      {stage0_10[31]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[6],stage1_11[18],stage1_10[38],stage1_9[52]}
   );
   gpc615_5 gpc125 (
      {stage0_9[82], stage0_9[83], stage0_9[84], stage0_9[85], stage0_9[86]},
      {stage0_10[32]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[7],stage1_11[19],stage1_10[39],stage1_9[53]}
   );
   gpc615_5 gpc126 (
      {stage0_9[87], stage0_9[88], stage0_9[89], stage0_9[90], stage0_9[91]},
      {stage0_10[33]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[8],stage1_11[20],stage1_10[40],stage1_9[54]}
   );
   gpc615_5 gpc127 (
      {stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95], stage0_9[96]},
      {stage0_10[34]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[9],stage1_11[21],stage1_10[41],stage1_9[55]}
   );
   gpc615_5 gpc128 (
      {stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage0_10[35]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[10],stage1_11[22],stage1_10[42],stage1_9[56]}
   );
   gpc615_5 gpc129 (
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106]},
      {stage0_10[36]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[11],stage1_11[23],stage1_10[43],stage1_9[57]}
   );
   gpc615_5 gpc130 (
      {stage0_9[107], stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111]},
      {stage0_10[37]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[12],stage1_11[24],stage1_10[44],stage1_9[58]}
   );
   gpc615_5 gpc131 (
      {stage0_9[112], stage0_9[113], stage0_9[114], stage0_9[115], stage0_9[116]},
      {stage0_10[38]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[13],stage1_11[25],stage1_10[45],stage1_9[59]}
   );
   gpc615_5 gpc132 (
      {stage0_9[117], stage0_9[118], stage0_9[119], stage0_9[120], stage0_9[121]},
      {stage0_10[39]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[14],stage1_11[26],stage1_10[46],stage1_9[60]}
   );
   gpc615_5 gpc133 (
      {stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125], stage0_9[126]},
      {stage0_10[40]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[15],stage1_11[27],stage1_10[47],stage1_9[61]}
   );
   gpc615_5 gpc134 (
      {stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage0_10[41]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[16],stage1_11[28],stage1_10[48],stage1_9[62]}
   );
   gpc615_5 gpc135 (
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136]},
      {stage0_10[42]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[17],stage1_11[29],stage1_10[49],stage1_9[63]}
   );
   gpc615_5 gpc136 (
      {stage0_9[137], stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141]},
      {stage0_10[43]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[18],stage1_11[30],stage1_10[50],stage1_9[64]}
   );
   gpc615_5 gpc137 (
      {stage0_9[142], stage0_9[143], stage0_9[144], stage0_9[145], stage0_9[146]},
      {stage0_10[44]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[19],stage1_11[31],stage1_10[51],stage1_9[65]}
   );
   gpc615_5 gpc138 (
      {stage0_9[147], stage0_9[148], stage0_9[149], stage0_9[150], stage0_9[151]},
      {stage0_10[45]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[20],stage1_11[32],stage1_10[52],stage1_9[66]}
   );
   gpc615_5 gpc139 (
      {stage0_10[46], stage0_10[47], stage0_10[48], stage0_10[49], stage0_10[50]},
      {stage0_11[96]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[16],stage1_12[21],stage1_11[33],stage1_10[53]}
   );
   gpc615_5 gpc140 (
      {stage0_10[51], stage0_10[52], stage0_10[53], stage0_10[54], stage0_10[55]},
      {stage0_11[97]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[17],stage1_12[22],stage1_11[34],stage1_10[54]}
   );
   gpc615_5 gpc141 (
      {stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59], stage0_10[60]},
      {stage0_11[98]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[18],stage1_12[23],stage1_11[35],stage1_10[55]}
   );
   gpc615_5 gpc142 (
      {stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage0_11[99]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[19],stage1_12[24],stage1_11[36],stage1_10[56]}
   );
   gpc615_5 gpc143 (
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70]},
      {stage0_11[100]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[20],stage1_12[25],stage1_11[37],stage1_10[57]}
   );
   gpc615_5 gpc144 (
      {stage0_10[71], stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75]},
      {stage0_11[101]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[21],stage1_12[26],stage1_11[38],stage1_10[58]}
   );
   gpc615_5 gpc145 (
      {stage0_10[76], stage0_10[77], stage0_10[78], stage0_10[79], stage0_10[80]},
      {stage0_11[102]},
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage1_14[6],stage1_13[22],stage1_12[27],stage1_11[39],stage1_10[59]}
   );
   gpc615_5 gpc146 (
      {stage0_10[81], stage0_10[82], stage0_10[83], stage0_10[84], stage0_10[85]},
      {stage0_11[103]},
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage1_14[7],stage1_13[23],stage1_12[28],stage1_11[40],stage1_10[60]}
   );
   gpc615_5 gpc147 (
      {stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89], stage0_10[90]},
      {stage0_11[104]},
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage1_14[8],stage1_13[24],stage1_12[29],stage1_11[41],stage1_10[61]}
   );
   gpc615_5 gpc148 (
      {stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage0_11[105]},
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage1_14[9],stage1_13[25],stage1_12[30],stage1_11[42],stage1_10[62]}
   );
   gpc615_5 gpc149 (
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100]},
      {stage0_11[106]},
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage1_14[10],stage1_13[26],stage1_12[31],stage1_11[43],stage1_10[63]}
   );
   gpc615_5 gpc150 (
      {stage0_10[101], stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105]},
      {stage0_11[107]},
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage1_14[11],stage1_13[27],stage1_12[32],stage1_11[44],stage1_10[64]}
   );
   gpc615_5 gpc151 (
      {stage0_10[106], stage0_10[107], stage0_10[108], stage0_10[109], stage0_10[110]},
      {stage0_11[108]},
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage1_14[12],stage1_13[28],stage1_12[33],stage1_11[45],stage1_10[65]}
   );
   gpc615_5 gpc152 (
      {stage0_10[111], stage0_10[112], stage0_10[113], stage0_10[114], stage0_10[115]},
      {stage0_11[109]},
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage1_14[13],stage1_13[29],stage1_12[34],stage1_11[46],stage1_10[66]}
   );
   gpc615_5 gpc153 (
      {stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119], stage0_10[120]},
      {stage0_11[110]},
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89]},
      {stage1_14[14],stage1_13[30],stage1_12[35],stage1_11[47],stage1_10[67]}
   );
   gpc615_5 gpc154 (
      {stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage0_11[111]},
      {stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95]},
      {stage1_14[15],stage1_13[31],stage1_12[36],stage1_11[48],stage1_10[68]}
   );
   gpc615_5 gpc155 (
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130]},
      {stage0_11[112]},
      {stage0_12[96], stage0_12[97], stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101]},
      {stage1_14[16],stage1_13[32],stage1_12[37],stage1_11[49],stage1_10[69]}
   );
   gpc615_5 gpc156 (
      {stage0_10[131], stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135]},
      {stage0_11[113]},
      {stage0_12[102], stage0_12[103], stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107]},
      {stage1_14[17],stage1_13[33],stage1_12[38],stage1_11[50],stage1_10[70]}
   );
   gpc615_5 gpc157 (
      {stage0_10[136], stage0_10[137], stage0_10[138], stage0_10[139], stage0_10[140]},
      {stage0_11[114]},
      {stage0_12[108], stage0_12[109], stage0_12[110], stage0_12[111], stage0_12[112], stage0_12[113]},
      {stage1_14[18],stage1_13[34],stage1_12[39],stage1_11[51],stage1_10[71]}
   );
   gpc615_5 gpc158 (
      {stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage0_12[114]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[19],stage1_13[35],stage1_12[40],stage1_11[52]}
   );
   gpc615_5 gpc159 (
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124]},
      {stage0_12[115]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[20],stage1_13[36],stage1_12[41],stage1_11[53]}
   );
   gpc615_5 gpc160 (
      {stage0_11[125], stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129]},
      {stage0_12[116]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[21],stage1_13[37],stage1_12[42],stage1_11[54]}
   );
   gpc615_5 gpc161 (
      {stage0_11[130], stage0_11[131], stage0_11[132], stage0_11[133], stage0_11[134]},
      {stage0_12[117]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[22],stage1_13[38],stage1_12[43],stage1_11[55]}
   );
   gpc615_5 gpc162 (
      {stage0_11[135], stage0_11[136], stage0_11[137], stage0_11[138], stage0_11[139]},
      {stage0_12[118]},
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage1_15[4],stage1_14[23],stage1_13[39],stage1_12[44],stage1_11[56]}
   );
   gpc615_5 gpc163 (
      {stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143], stage0_11[144]},
      {stage0_12[119]},
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage1_15[5],stage1_14[24],stage1_13[40],stage1_12[45],stage1_11[57]}
   );
   gpc615_5 gpc164 (
      {stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage0_12[120]},
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage1_15[6],stage1_14[25],stage1_13[41],stage1_12[46],stage1_11[58]}
   );
   gpc615_5 gpc165 (
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154]},
      {stage0_12[121]},
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage1_15[7],stage1_14[26],stage1_13[42],stage1_12[47],stage1_11[59]}
   );
   gpc615_5 gpc166 (
      {stage0_12[122], stage0_12[123], stage0_12[124], stage0_12[125], stage0_12[126]},
      {stage0_13[48]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[8],stage1_14[27],stage1_13[43],stage1_12[48]}
   );
   gpc615_5 gpc167 (
      {stage0_12[127], stage0_12[128], stage0_12[129], stage0_12[130], stage0_12[131]},
      {stage0_13[49]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[9],stage1_14[28],stage1_13[44],stage1_12[49]}
   );
   gpc615_5 gpc168 (
      {stage0_12[132], stage0_12[133], stage0_12[134], stage0_12[135], stage0_12[136]},
      {stage0_13[50]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[10],stage1_14[29],stage1_13[45],stage1_12[50]}
   );
   gpc615_5 gpc169 (
      {stage0_12[137], stage0_12[138], stage0_12[139], stage0_12[140], stage0_12[141]},
      {stage0_13[51]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[11],stage1_14[30],stage1_13[46],stage1_12[51]}
   );
   gpc615_5 gpc170 (
      {stage0_12[142], stage0_12[143], stage0_12[144], stage0_12[145], stage0_12[146]},
      {stage0_13[52]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[12],stage1_14[31],stage1_13[47],stage1_12[52]}
   );
   gpc615_5 gpc171 (
      {stage0_12[147], stage0_12[148], stage0_12[149], stage0_12[150], stage0_12[151]},
      {stage0_13[53]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[13],stage1_14[32],stage1_13[48],stage1_12[53]}
   );
   gpc615_5 gpc172 (
      {stage0_12[152], stage0_12[153], stage0_12[154], stage0_12[155], stage0_12[156]},
      {stage0_13[54]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[14],stage1_14[33],stage1_13[49],stage1_12[54]}
   );
   gpc615_5 gpc173 (
      {stage0_12[157], stage0_12[158], stage0_12[159], stage0_12[160], stage0_12[161]},
      {stage0_13[55]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[15],stage1_14[34],stage1_13[50],stage1_12[55]}
   );
   gpc606_5 gpc174 (
      {stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59], stage0_13[60], stage0_13[61]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[8],stage1_15[16],stage1_14[35],stage1_13[51]}
   );
   gpc606_5 gpc175 (
      {stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65], stage0_13[66], stage0_13[67]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[9],stage1_15[17],stage1_14[36],stage1_13[52]}
   );
   gpc606_5 gpc176 (
      {stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71], stage0_13[72], stage0_13[73]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[10],stage1_15[18],stage1_14[37],stage1_13[53]}
   );
   gpc615_5 gpc177 (
      {stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77], stage0_13[78]},
      {stage0_14[48]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[11],stage1_15[19],stage1_14[38],stage1_13[54]}
   );
   gpc615_5 gpc178 (
      {stage0_13[79], stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83]},
      {stage0_14[49]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[12],stage1_15[20],stage1_14[39],stage1_13[55]}
   );
   gpc615_5 gpc179 (
      {stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87], stage0_13[88]},
      {stage0_14[50]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[13],stage1_15[21],stage1_14[40],stage1_13[56]}
   );
   gpc615_5 gpc180 (
      {stage0_13[89], stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93]},
      {stage0_14[51]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[14],stage1_15[22],stage1_14[41],stage1_13[57]}
   );
   gpc615_5 gpc181 (
      {stage0_13[94], stage0_13[95], stage0_13[96], stage0_13[97], stage0_13[98]},
      {stage0_14[52]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[15],stage1_15[23],stage1_14[42],stage1_13[58]}
   );
   gpc615_5 gpc182 (
      {stage0_13[99], stage0_13[100], stage0_13[101], stage0_13[102], stage0_13[103]},
      {stage0_14[53]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[16],stage1_15[24],stage1_14[43],stage1_13[59]}
   );
   gpc615_5 gpc183 (
      {stage0_13[104], stage0_13[105], stage0_13[106], stage0_13[107], stage0_13[108]},
      {stage0_14[54]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[17],stage1_15[25],stage1_14[44],stage1_13[60]}
   );
   gpc615_5 gpc184 (
      {stage0_13[109], stage0_13[110], stage0_13[111], stage0_13[112], stage0_13[113]},
      {stage0_14[55]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[18],stage1_15[26],stage1_14[45],stage1_13[61]}
   );
   gpc615_5 gpc185 (
      {stage0_13[114], stage0_13[115], stage0_13[116], stage0_13[117], stage0_13[118]},
      {stage0_14[56]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[19],stage1_15[27],stage1_14[46],stage1_13[62]}
   );
   gpc615_5 gpc186 (
      {stage0_13[119], stage0_13[120], stage0_13[121], stage0_13[122], stage0_13[123]},
      {stage0_14[57]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[20],stage1_15[28],stage1_14[47],stage1_13[63]}
   );
   gpc615_5 gpc187 (
      {stage0_13[124], stage0_13[125], stage0_13[126], stage0_13[127], stage0_13[128]},
      {stage0_14[58]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[21],stage1_15[29],stage1_14[48],stage1_13[64]}
   );
   gpc615_5 gpc188 (
      {stage0_13[129], stage0_13[130], stage0_13[131], stage0_13[132], stage0_13[133]},
      {stage0_14[59]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[22],stage1_15[30],stage1_14[49],stage1_13[65]}
   );
   gpc615_5 gpc189 (
      {stage0_13[134], stage0_13[135], stage0_13[136], stage0_13[137], stage0_13[138]},
      {stage0_14[60]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[23],stage1_15[31],stage1_14[50],stage1_13[66]}
   );
   gpc615_5 gpc190 (
      {stage0_13[139], stage0_13[140], stage0_13[141], stage0_13[142], stage0_13[143]},
      {stage0_14[61]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[24],stage1_15[32],stage1_14[51],stage1_13[67]}
   );
   gpc117_4 gpc191 (
      {stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65], stage0_14[66], stage0_14[67], stage0_14[68]},
      {stage0_15[102]},
      {stage0_16[0]},
      {stage1_17[17],stage1_16[25],stage1_15[33],stage1_14[52]}
   );
   gpc117_4 gpc192 (
      {stage0_14[69], stage0_14[70], stage0_14[71], stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75]},
      {stage0_15[103]},
      {stage0_16[1]},
      {stage1_17[18],stage1_16[26],stage1_15[34],stage1_14[53]}
   );
   gpc117_4 gpc193 (
      {stage0_14[76], stage0_14[77], stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82]},
      {stage0_15[104]},
      {stage0_16[2]},
      {stage1_17[19],stage1_16[27],stage1_15[35],stage1_14[54]}
   );
   gpc117_4 gpc194 (
      {stage0_14[83], stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage0_15[105]},
      {stage0_16[3]},
      {stage1_17[20],stage1_16[28],stage1_15[36],stage1_14[55]}
   );
   gpc606_5 gpc195 (
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage0_16[4], stage0_16[5], stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9]},
      {stage1_18[0],stage1_17[21],stage1_16[29],stage1_15[37],stage1_14[56]}
   );
   gpc606_5 gpc196 (
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage0_16[10], stage0_16[11], stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15]},
      {stage1_18[1],stage1_17[22],stage1_16[30],stage1_15[38],stage1_14[57]}
   );
   gpc606_5 gpc197 (
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage0_16[16], stage0_16[17], stage0_16[18], stage0_16[19], stage0_16[20], stage0_16[21]},
      {stage1_18[2],stage1_17[23],stage1_16[31],stage1_15[39],stage1_14[58]}
   );
   gpc606_5 gpc198 (
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113]},
      {stage0_16[22], stage0_16[23], stage0_16[24], stage0_16[25], stage0_16[26], stage0_16[27]},
      {stage1_18[3],stage1_17[24],stage1_16[32],stage1_15[40],stage1_14[59]}
   );
   gpc606_5 gpc199 (
      {stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119]},
      {stage0_16[28], stage0_16[29], stage0_16[30], stage0_16[31], stage0_16[32], stage0_16[33]},
      {stage1_18[4],stage1_17[25],stage1_16[33],stage1_15[41],stage1_14[60]}
   );
   gpc606_5 gpc200 (
      {stage0_14[120], stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125]},
      {stage0_16[34], stage0_16[35], stage0_16[36], stage0_16[37], stage0_16[38], stage0_16[39]},
      {stage1_18[5],stage1_17[26],stage1_16[34],stage1_15[42],stage1_14[61]}
   );
   gpc606_5 gpc201 (
      {stage0_14[126], stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131]},
      {stage0_16[40], stage0_16[41], stage0_16[42], stage0_16[43], stage0_16[44], stage0_16[45]},
      {stage1_18[6],stage1_17[27],stage1_16[35],stage1_15[43],stage1_14[62]}
   );
   gpc606_5 gpc202 (
      {stage0_14[132], stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137]},
      {stage0_16[46], stage0_16[47], stage0_16[48], stage0_16[49], stage0_16[50], stage0_16[51]},
      {stage1_18[7],stage1_17[28],stage1_16[36],stage1_15[44],stage1_14[63]}
   );
   gpc606_5 gpc203 (
      {stage0_14[138], stage0_14[139], stage0_14[140], stage0_14[141], stage0_14[142], stage0_14[143]},
      {stage0_16[52], stage0_16[53], stage0_16[54], stage0_16[55], stage0_16[56], stage0_16[57]},
      {stage1_18[8],stage1_17[29],stage1_16[37],stage1_15[45],stage1_14[64]}
   );
   gpc606_5 gpc204 (
      {stage0_14[144], stage0_14[145], stage0_14[146], stage0_14[147], stage0_14[148], stage0_14[149]},
      {stage0_16[58], stage0_16[59], stage0_16[60], stage0_16[61], stage0_16[62], stage0_16[63]},
      {stage1_18[9],stage1_17[30],stage1_16[38],stage1_15[46],stage1_14[65]}
   );
   gpc606_5 gpc205 (
      {stage0_14[150], stage0_14[151], stage0_14[152], stage0_14[153], stage0_14[154], stage0_14[155]},
      {stage0_16[64], stage0_16[65], stage0_16[66], stage0_16[67], stage0_16[68], stage0_16[69]},
      {stage1_18[10],stage1_17[31],stage1_16[39],stage1_15[47],stage1_14[66]}
   );
   gpc615_5 gpc206 (
      {stage0_14[156], stage0_14[157], stage0_14[158], stage0_14[159], stage0_14[160]},
      {stage0_15[106]},
      {stage0_16[70], stage0_16[71], stage0_16[72], stage0_16[73], stage0_16[74], stage0_16[75]},
      {stage1_18[11],stage1_17[32],stage1_16[40],stage1_15[48],stage1_14[67]}
   );
   gpc615_5 gpc207 (
      {stage0_15[107], stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111]},
      {stage0_16[76]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[12],stage1_17[33],stage1_16[41],stage1_15[49]}
   );
   gpc615_5 gpc208 (
      {stage0_15[112], stage0_15[113], stage0_15[114], stage0_15[115], stage0_15[116]},
      {stage0_16[77]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[13],stage1_17[34],stage1_16[42],stage1_15[50]}
   );
   gpc615_5 gpc209 (
      {stage0_15[117], stage0_15[118], stage0_15[119], stage0_15[120], stage0_15[121]},
      {stage0_16[78]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[14],stage1_17[35],stage1_16[43],stage1_15[51]}
   );
   gpc615_5 gpc210 (
      {stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125], stage0_15[126]},
      {stage0_16[79]},
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage1_19[3],stage1_18[15],stage1_17[36],stage1_16[44],stage1_15[52]}
   );
   gpc615_5 gpc211 (
      {stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage0_16[80]},
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage1_19[4],stage1_18[16],stage1_17[37],stage1_16[45],stage1_15[53]}
   );
   gpc615_5 gpc212 (
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136]},
      {stage0_16[81]},
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage1_19[5],stage1_18[17],stage1_17[38],stage1_16[46],stage1_15[54]}
   );
   gpc615_5 gpc213 (
      {stage0_15[137], stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141]},
      {stage0_16[82]},
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage1_19[6],stage1_18[18],stage1_17[39],stage1_16[47],stage1_15[55]}
   );
   gpc615_5 gpc214 (
      {stage0_15[142], stage0_15[143], stage0_15[144], stage0_15[145], stage0_15[146]},
      {stage0_16[83]},
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage1_19[7],stage1_18[19],stage1_17[40],stage1_16[48],stage1_15[56]}
   );
   gpc615_5 gpc215 (
      {stage0_15[147], stage0_15[148], stage0_15[149], stage0_15[150], stage0_15[151]},
      {stage0_16[84]},
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage1_19[8],stage1_18[20],stage1_17[41],stage1_16[49],stage1_15[57]}
   );
   gpc615_5 gpc216 (
      {stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155], stage0_15[156]},
      {stage0_16[85]},
      {stage0_17[54], stage0_17[55], stage0_17[56], stage0_17[57], stage0_17[58], stage0_17[59]},
      {stage1_19[9],stage1_18[21],stage1_17[42],stage1_16[50],stage1_15[58]}
   );
   gpc615_5 gpc217 (
      {stage0_15[157], stage0_15[158], stage0_15[159], stage0_15[160], stage0_15[161]},
      {stage0_16[86]},
      {stage0_17[60], stage0_17[61], stage0_17[62], stage0_17[63], stage0_17[64], stage0_17[65]},
      {stage1_19[10],stage1_18[22],stage1_17[43],stage1_16[51],stage1_15[59]}
   );
   gpc606_5 gpc218 (
      {stage0_16[87], stage0_16[88], stage0_16[89], stage0_16[90], stage0_16[91], stage0_16[92]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[11],stage1_18[23],stage1_17[44],stage1_16[52]}
   );
   gpc606_5 gpc219 (
      {stage0_16[93], stage0_16[94], stage0_16[95], stage0_16[96], stage0_16[97], stage0_16[98]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[12],stage1_18[24],stage1_17[45],stage1_16[53]}
   );
   gpc606_5 gpc220 (
      {stage0_16[99], stage0_16[100], stage0_16[101], stage0_16[102], stage0_16[103], stage0_16[104]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[13],stage1_18[25],stage1_17[46],stage1_16[54]}
   );
   gpc606_5 gpc221 (
      {stage0_16[105], stage0_16[106], stage0_16[107], stage0_16[108], stage0_16[109], stage0_16[110]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[14],stage1_18[26],stage1_17[47],stage1_16[55]}
   );
   gpc606_5 gpc222 (
      {stage0_17[66], stage0_17[67], stage0_17[68], stage0_17[69], stage0_17[70], stage0_17[71]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[4],stage1_19[15],stage1_18[27],stage1_17[48]}
   );
   gpc606_5 gpc223 (
      {stage0_17[72], stage0_17[73], stage0_17[74], stage0_17[75], stage0_17[76], stage0_17[77]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[5],stage1_19[16],stage1_18[28],stage1_17[49]}
   );
   gpc606_5 gpc224 (
      {stage0_17[78], stage0_17[79], stage0_17[80], stage0_17[81], stage0_17[82], stage0_17[83]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[6],stage1_19[17],stage1_18[29],stage1_17[50]}
   );
   gpc606_5 gpc225 (
      {stage0_17[84], stage0_17[85], stage0_17[86], stage0_17[87], stage0_17[88], stage0_17[89]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[7],stage1_19[18],stage1_18[30],stage1_17[51]}
   );
   gpc606_5 gpc226 (
      {stage0_17[90], stage0_17[91], stage0_17[92], stage0_17[93], stage0_17[94], stage0_17[95]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[8],stage1_19[19],stage1_18[31],stage1_17[52]}
   );
   gpc606_5 gpc227 (
      {stage0_17[96], stage0_17[97], stage0_17[98], stage0_17[99], stage0_17[100], stage0_17[101]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[9],stage1_19[20],stage1_18[32],stage1_17[53]}
   );
   gpc606_5 gpc228 (
      {stage0_17[102], stage0_17[103], stage0_17[104], stage0_17[105], stage0_17[106], stage0_17[107]},
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage1_21[6],stage1_20[10],stage1_19[21],stage1_18[33],stage1_17[54]}
   );
   gpc606_5 gpc229 (
      {stage0_17[108], stage0_17[109], stage0_17[110], stage0_17[111], stage0_17[112], stage0_17[113]},
      {stage0_19[42], stage0_19[43], stage0_19[44], stage0_19[45], stage0_19[46], stage0_19[47]},
      {stage1_21[7],stage1_20[11],stage1_19[22],stage1_18[34],stage1_17[55]}
   );
   gpc606_5 gpc230 (
      {stage0_17[114], stage0_17[115], stage0_17[116], stage0_17[117], stage0_17[118], stage0_17[119]},
      {stage0_19[48], stage0_19[49], stage0_19[50], stage0_19[51], stage0_19[52], stage0_19[53]},
      {stage1_21[8],stage1_20[12],stage1_19[23],stage1_18[35],stage1_17[56]}
   );
   gpc606_5 gpc231 (
      {stage0_17[120], stage0_17[121], stage0_17[122], stage0_17[123], stage0_17[124], stage0_17[125]},
      {stage0_19[54], stage0_19[55], stage0_19[56], stage0_19[57], stage0_19[58], stage0_19[59]},
      {stage1_21[9],stage1_20[13],stage1_19[24],stage1_18[36],stage1_17[57]}
   );
   gpc606_5 gpc232 (
      {stage0_17[126], stage0_17[127], stage0_17[128], stage0_17[129], stage0_17[130], stage0_17[131]},
      {stage0_19[60], stage0_19[61], stage0_19[62], stage0_19[63], stage0_19[64], stage0_19[65]},
      {stage1_21[10],stage1_20[14],stage1_19[25],stage1_18[37],stage1_17[58]}
   );
   gpc606_5 gpc233 (
      {stage0_17[132], stage0_17[133], stage0_17[134], stage0_17[135], stage0_17[136], stage0_17[137]},
      {stage0_19[66], stage0_19[67], stage0_19[68], stage0_19[69], stage0_19[70], stage0_19[71]},
      {stage1_21[11],stage1_20[15],stage1_19[26],stage1_18[38],stage1_17[59]}
   );
   gpc606_5 gpc234 (
      {stage0_17[138], stage0_17[139], stage0_17[140], stage0_17[141], stage0_17[142], stage0_17[143]},
      {stage0_19[72], stage0_19[73], stage0_19[74], stage0_19[75], stage0_19[76], stage0_19[77]},
      {stage1_21[12],stage1_20[16],stage1_19[27],stage1_18[39],stage1_17[60]}
   );
   gpc606_5 gpc235 (
      {stage0_17[144], stage0_17[145], stage0_17[146], stage0_17[147], stage0_17[148], stage0_17[149]},
      {stage0_19[78], stage0_19[79], stage0_19[80], stage0_19[81], stage0_19[82], stage0_19[83]},
      {stage1_21[13],stage1_20[17],stage1_19[28],stage1_18[40],stage1_17[61]}
   );
   gpc606_5 gpc236 (
      {stage0_17[150], stage0_17[151], stage0_17[152], stage0_17[153], stage0_17[154], stage0_17[155]},
      {stage0_19[84], stage0_19[85], stage0_19[86], stage0_19[87], stage0_19[88], stage0_19[89]},
      {stage1_21[14],stage1_20[18],stage1_19[29],stage1_18[41],stage1_17[62]}
   );
   gpc606_5 gpc237 (
      {stage0_17[156], stage0_17[157], stage0_17[158], stage0_17[159], stage0_17[160], stage0_17[161]},
      {stage0_19[90], stage0_19[91], stage0_19[92], stage0_19[93], stage0_19[94], stage0_19[95]},
      {stage1_21[15],stage1_20[19],stage1_19[30],stage1_18[42],stage1_17[63]}
   );
   gpc117_4 gpc238 (
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29], stage0_18[30]},
      {stage0_19[96]},
      {stage0_20[0]},
      {stage1_21[16],stage1_20[20],stage1_19[31],stage1_18[43]}
   );
   gpc117_4 gpc239 (
      {stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35], stage0_18[36], stage0_18[37]},
      {stage0_19[97]},
      {stage0_20[1]},
      {stage1_21[17],stage1_20[21],stage1_19[32],stage1_18[44]}
   );
   gpc117_4 gpc240 (
      {stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41], stage0_18[42], stage0_18[43], stage0_18[44]},
      {stage0_19[98]},
      {stage0_20[2]},
      {stage1_21[18],stage1_20[22],stage1_19[33],stage1_18[45]}
   );
   gpc117_4 gpc241 (
      {stage0_18[45], stage0_18[46], stage0_18[47], stage0_18[48], stage0_18[49], stage0_18[50], stage0_18[51]},
      {stage0_19[99]},
      {stage0_20[3]},
      {stage1_21[19],stage1_20[23],stage1_19[34],stage1_18[46]}
   );
   gpc606_5 gpc242 (
      {stage0_18[52], stage0_18[53], stage0_18[54], stage0_18[55], stage0_18[56], stage0_18[57]},
      {stage0_20[4], stage0_20[5], stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9]},
      {stage1_22[0],stage1_21[20],stage1_20[24],stage1_19[35],stage1_18[47]}
   );
   gpc606_5 gpc243 (
      {stage0_18[58], stage0_18[59], stage0_18[60], stage0_18[61], stage0_18[62], stage0_18[63]},
      {stage0_20[10], stage0_20[11], stage0_20[12], stage0_20[13], stage0_20[14], stage0_20[15]},
      {stage1_22[1],stage1_21[21],stage1_20[25],stage1_19[36],stage1_18[48]}
   );
   gpc606_5 gpc244 (
      {stage0_18[64], stage0_18[65], stage0_18[66], stage0_18[67], stage0_18[68], stage0_18[69]},
      {stage0_20[16], stage0_20[17], stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21]},
      {stage1_22[2],stage1_21[22],stage1_20[26],stage1_19[37],stage1_18[49]}
   );
   gpc606_5 gpc245 (
      {stage0_18[70], stage0_18[71], stage0_18[72], stage0_18[73], stage0_18[74], stage0_18[75]},
      {stage0_20[22], stage0_20[23], stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27]},
      {stage1_22[3],stage1_21[23],stage1_20[27],stage1_19[38],stage1_18[50]}
   );
   gpc606_5 gpc246 (
      {stage0_18[76], stage0_18[77], stage0_18[78], stage0_18[79], stage0_18[80], stage0_18[81]},
      {stage0_20[28], stage0_20[29], stage0_20[30], stage0_20[31], stage0_20[32], stage0_20[33]},
      {stage1_22[4],stage1_21[24],stage1_20[28],stage1_19[39],stage1_18[51]}
   );
   gpc606_5 gpc247 (
      {stage0_18[82], stage0_18[83], stage0_18[84], stage0_18[85], stage0_18[86], stage0_18[87]},
      {stage0_20[34], stage0_20[35], stage0_20[36], stage0_20[37], stage0_20[38], stage0_20[39]},
      {stage1_22[5],stage1_21[25],stage1_20[29],stage1_19[40],stage1_18[52]}
   );
   gpc606_5 gpc248 (
      {stage0_18[88], stage0_18[89], stage0_18[90], stage0_18[91], stage0_18[92], stage0_18[93]},
      {stage0_20[40], stage0_20[41], stage0_20[42], stage0_20[43], stage0_20[44], stage0_20[45]},
      {stage1_22[6],stage1_21[26],stage1_20[30],stage1_19[41],stage1_18[53]}
   );
   gpc606_5 gpc249 (
      {stage0_18[94], stage0_18[95], stage0_18[96], stage0_18[97], stage0_18[98], stage0_18[99]},
      {stage0_20[46], stage0_20[47], stage0_20[48], stage0_20[49], stage0_20[50], stage0_20[51]},
      {stage1_22[7],stage1_21[27],stage1_20[31],stage1_19[42],stage1_18[54]}
   );
   gpc606_5 gpc250 (
      {stage0_18[100], stage0_18[101], stage0_18[102], stage0_18[103], stage0_18[104], stage0_18[105]},
      {stage0_20[52], stage0_20[53], stage0_20[54], stage0_20[55], stage0_20[56], stage0_20[57]},
      {stage1_22[8],stage1_21[28],stage1_20[32],stage1_19[43],stage1_18[55]}
   );
   gpc606_5 gpc251 (
      {stage0_18[106], stage0_18[107], stage0_18[108], stage0_18[109], stage0_18[110], stage0_18[111]},
      {stage0_20[58], stage0_20[59], stage0_20[60], stage0_20[61], stage0_20[62], stage0_20[63]},
      {stage1_22[9],stage1_21[29],stage1_20[33],stage1_19[44],stage1_18[56]}
   );
   gpc606_5 gpc252 (
      {stage0_18[112], stage0_18[113], stage0_18[114], stage0_18[115], stage0_18[116], stage0_18[117]},
      {stage0_20[64], stage0_20[65], stage0_20[66], stage0_20[67], stage0_20[68], stage0_20[69]},
      {stage1_22[10],stage1_21[30],stage1_20[34],stage1_19[45],stage1_18[57]}
   );
   gpc606_5 gpc253 (
      {stage0_18[118], stage0_18[119], stage0_18[120], stage0_18[121], stage0_18[122], stage0_18[123]},
      {stage0_20[70], stage0_20[71], stage0_20[72], stage0_20[73], stage0_20[74], stage0_20[75]},
      {stage1_22[11],stage1_21[31],stage1_20[35],stage1_19[46],stage1_18[58]}
   );
   gpc606_5 gpc254 (
      {stage0_18[124], stage0_18[125], stage0_18[126], stage0_18[127], stage0_18[128], stage0_18[129]},
      {stage0_20[76], stage0_20[77], stage0_20[78], stage0_20[79], stage0_20[80], stage0_20[81]},
      {stage1_22[12],stage1_21[32],stage1_20[36],stage1_19[47],stage1_18[59]}
   );
   gpc606_5 gpc255 (
      {stage0_18[130], stage0_18[131], stage0_18[132], stage0_18[133], stage0_18[134], stage0_18[135]},
      {stage0_20[82], stage0_20[83], stage0_20[84], stage0_20[85], stage0_20[86], stage0_20[87]},
      {stage1_22[13],stage1_21[33],stage1_20[37],stage1_19[48],stage1_18[60]}
   );
   gpc606_5 gpc256 (
      {stage0_18[136], stage0_18[137], stage0_18[138], stage0_18[139], stage0_18[140], stage0_18[141]},
      {stage0_20[88], stage0_20[89], stage0_20[90], stage0_20[91], stage0_20[92], stage0_20[93]},
      {stage1_22[14],stage1_21[34],stage1_20[38],stage1_19[49],stage1_18[61]}
   );
   gpc606_5 gpc257 (
      {stage0_19[100], stage0_19[101], stage0_19[102], stage0_19[103], stage0_19[104], stage0_19[105]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[15],stage1_21[35],stage1_20[39],stage1_19[50]}
   );
   gpc606_5 gpc258 (
      {stage0_19[106], stage0_19[107], stage0_19[108], stage0_19[109], stage0_19[110], stage0_19[111]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[16],stage1_21[36],stage1_20[40],stage1_19[51]}
   );
   gpc606_5 gpc259 (
      {stage0_19[112], stage0_19[113], stage0_19[114], stage0_19[115], stage0_19[116], stage0_19[117]},
      {stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17]},
      {stage1_23[2],stage1_22[17],stage1_21[37],stage1_20[41],stage1_19[52]}
   );
   gpc606_5 gpc260 (
      {stage0_19[118], stage0_19[119], stage0_19[120], stage0_19[121], stage0_19[122], stage0_19[123]},
      {stage0_21[18], stage0_21[19], stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23]},
      {stage1_23[3],stage1_22[18],stage1_21[38],stage1_20[42],stage1_19[53]}
   );
   gpc606_5 gpc261 (
      {stage0_19[124], stage0_19[125], stage0_19[126], stage0_19[127], stage0_19[128], stage0_19[129]},
      {stage0_21[24], stage0_21[25], stage0_21[26], stage0_21[27], stage0_21[28], stage0_21[29]},
      {stage1_23[4],stage1_22[19],stage1_21[39],stage1_20[43],stage1_19[54]}
   );
   gpc606_5 gpc262 (
      {stage0_19[130], stage0_19[131], stage0_19[132], stage0_19[133], stage0_19[134], stage0_19[135]},
      {stage0_21[30], stage0_21[31], stage0_21[32], stage0_21[33], stage0_21[34], stage0_21[35]},
      {stage1_23[5],stage1_22[20],stage1_21[40],stage1_20[44],stage1_19[55]}
   );
   gpc606_5 gpc263 (
      {stage0_19[136], stage0_19[137], stage0_19[138], stage0_19[139], stage0_19[140], stage0_19[141]},
      {stage0_21[36], stage0_21[37], stage0_21[38], stage0_21[39], stage0_21[40], stage0_21[41]},
      {stage1_23[6],stage1_22[21],stage1_21[41],stage1_20[45],stage1_19[56]}
   );
   gpc606_5 gpc264 (
      {stage0_19[142], stage0_19[143], stage0_19[144], stage0_19[145], stage0_19[146], stage0_19[147]},
      {stage0_21[42], stage0_21[43], stage0_21[44], stage0_21[45], stage0_21[46], stage0_21[47]},
      {stage1_23[7],stage1_22[22],stage1_21[42],stage1_20[46],stage1_19[57]}
   );
   gpc606_5 gpc265 (
      {stage0_19[148], stage0_19[149], stage0_19[150], stage0_19[151], stage0_19[152], stage0_19[153]},
      {stage0_21[48], stage0_21[49], stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53]},
      {stage1_23[8],stage1_22[23],stage1_21[43],stage1_20[47],stage1_19[58]}
   );
   gpc606_5 gpc266 (
      {stage0_20[94], stage0_20[95], stage0_20[96], stage0_20[97], stage0_20[98], stage0_20[99]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[9],stage1_22[24],stage1_21[44],stage1_20[48]}
   );
   gpc606_5 gpc267 (
      {stage0_20[100], stage0_20[101], stage0_20[102], stage0_20[103], stage0_20[104], stage0_20[105]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[10],stage1_22[25],stage1_21[45],stage1_20[49]}
   );
   gpc606_5 gpc268 (
      {stage0_20[106], stage0_20[107], stage0_20[108], stage0_20[109], stage0_20[110], stage0_20[111]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[11],stage1_22[26],stage1_21[46],stage1_20[50]}
   );
   gpc615_5 gpc269 (
      {stage0_20[112], stage0_20[113], stage0_20[114], stage0_20[115], stage0_20[116]},
      {stage0_21[54]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[12],stage1_22[27],stage1_21[47],stage1_20[51]}
   );
   gpc615_5 gpc270 (
      {stage0_20[117], stage0_20[118], stage0_20[119], stage0_20[120], stage0_20[121]},
      {stage0_21[55]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[13],stage1_22[28],stage1_21[48],stage1_20[52]}
   );
   gpc615_5 gpc271 (
      {stage0_20[122], stage0_20[123], stage0_20[124], stage0_20[125], stage0_20[126]},
      {stage0_21[56]},
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage1_24[5],stage1_23[14],stage1_22[29],stage1_21[49],stage1_20[53]}
   );
   gpc615_5 gpc272 (
      {stage0_20[127], stage0_20[128], stage0_20[129], stage0_20[130], stage0_20[131]},
      {stage0_21[57]},
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage1_24[6],stage1_23[15],stage1_22[30],stage1_21[50],stage1_20[54]}
   );
   gpc615_5 gpc273 (
      {stage0_20[132], stage0_20[133], stage0_20[134], stage0_20[135], stage0_20[136]},
      {stage0_21[58]},
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47]},
      {stage1_24[7],stage1_23[16],stage1_22[31],stage1_21[51],stage1_20[55]}
   );
   gpc615_5 gpc274 (
      {stage0_20[137], stage0_20[138], stage0_20[139], stage0_20[140], stage0_20[141]},
      {stage0_21[59]},
      {stage0_22[48], stage0_22[49], stage0_22[50], stage0_22[51], stage0_22[52], stage0_22[53]},
      {stage1_24[8],stage1_23[17],stage1_22[32],stage1_21[52],stage1_20[56]}
   );
   gpc615_5 gpc275 (
      {stage0_20[142], stage0_20[143], stage0_20[144], stage0_20[145], stage0_20[146]},
      {stage0_21[60]},
      {stage0_22[54], stage0_22[55], stage0_22[56], stage0_22[57], stage0_22[58], stage0_22[59]},
      {stage1_24[9],stage1_23[18],stage1_22[33],stage1_21[53],stage1_20[57]}
   );
   gpc615_5 gpc276 (
      {stage0_20[147], stage0_20[148], stage0_20[149], stage0_20[150], stage0_20[151]},
      {stage0_21[61]},
      {stage0_22[60], stage0_22[61], stage0_22[62], stage0_22[63], stage0_22[64], stage0_22[65]},
      {stage1_24[10],stage1_23[19],stage1_22[34],stage1_21[54],stage1_20[58]}
   );
   gpc615_5 gpc277 (
      {stage0_20[152], stage0_20[153], stage0_20[154], stage0_20[155], stage0_20[156]},
      {stage0_21[62]},
      {stage0_22[66], stage0_22[67], stage0_22[68], stage0_22[69], stage0_22[70], stage0_22[71]},
      {stage1_24[11],stage1_23[20],stage1_22[35],stage1_21[55],stage1_20[59]}
   );
   gpc615_5 gpc278 (
      {stage0_20[157], stage0_20[158], stage0_20[159], stage0_20[160], stage0_20[161]},
      {stage0_21[63]},
      {stage0_22[72], stage0_22[73], stage0_22[74], stage0_22[75], stage0_22[76], stage0_22[77]},
      {stage1_24[12],stage1_23[21],stage1_22[36],stage1_21[56],stage1_20[60]}
   );
   gpc1163_5 gpc279 (
      {stage0_21[64], stage0_21[65], stage0_21[66]},
      {stage0_22[78], stage0_22[79], stage0_22[80], stage0_22[81], stage0_22[82], stage0_22[83]},
      {stage0_23[0]},
      {stage0_24[0]},
      {stage1_25[0],stage1_24[13],stage1_23[22],stage1_22[37],stage1_21[57]}
   );
   gpc1163_5 gpc280 (
      {stage0_21[67], stage0_21[68], stage0_21[69]},
      {stage0_22[84], stage0_22[85], stage0_22[86], stage0_22[87], stage0_22[88], stage0_22[89]},
      {stage0_23[1]},
      {stage0_24[1]},
      {stage1_25[1],stage1_24[14],stage1_23[23],stage1_22[38],stage1_21[58]}
   );
   gpc1163_5 gpc281 (
      {stage0_21[70], stage0_21[71], stage0_21[72]},
      {stage0_22[90], stage0_22[91], stage0_22[92], stage0_22[93], stage0_22[94], stage0_22[95]},
      {stage0_23[2]},
      {stage0_24[2]},
      {stage1_25[2],stage1_24[15],stage1_23[24],stage1_22[39],stage1_21[59]}
   );
   gpc1163_5 gpc282 (
      {stage0_21[73], stage0_21[74], stage0_21[75]},
      {stage0_22[96], stage0_22[97], stage0_22[98], stage0_22[99], stage0_22[100], stage0_22[101]},
      {stage0_23[3]},
      {stage0_24[3]},
      {stage1_25[3],stage1_24[16],stage1_23[25],stage1_22[40],stage1_21[60]}
   );
   gpc1163_5 gpc283 (
      {stage0_21[76], stage0_21[77], stage0_21[78]},
      {stage0_22[102], stage0_22[103], stage0_22[104], stage0_22[105], stage0_22[106], stage0_22[107]},
      {stage0_23[4]},
      {stage0_24[4]},
      {stage1_25[4],stage1_24[17],stage1_23[26],stage1_22[41],stage1_21[61]}
   );
   gpc1163_5 gpc284 (
      {stage0_21[79], stage0_21[80], stage0_21[81]},
      {stage0_22[108], stage0_22[109], stage0_22[110], stage0_22[111], stage0_22[112], stage0_22[113]},
      {stage0_23[5]},
      {stage0_24[5]},
      {stage1_25[5],stage1_24[18],stage1_23[27],stage1_22[42],stage1_21[62]}
   );
   gpc1163_5 gpc285 (
      {stage0_21[82], stage0_21[83], stage0_21[84]},
      {stage0_22[114], stage0_22[115], stage0_22[116], stage0_22[117], stage0_22[118], stage0_22[119]},
      {stage0_23[6]},
      {stage0_24[6]},
      {stage1_25[6],stage1_24[19],stage1_23[28],stage1_22[43],stage1_21[63]}
   );
   gpc1163_5 gpc286 (
      {stage0_21[85], stage0_21[86], stage0_21[87]},
      {stage0_22[120], stage0_22[121], stage0_22[122], stage0_22[123], stage0_22[124], stage0_22[125]},
      {stage0_23[7]},
      {stage0_24[7]},
      {stage1_25[7],stage1_24[20],stage1_23[29],stage1_22[44],stage1_21[64]}
   );
   gpc1163_5 gpc287 (
      {stage0_21[88], stage0_21[89], stage0_21[90]},
      {stage0_22[126], stage0_22[127], stage0_22[128], stage0_22[129], stage0_22[130], stage0_22[131]},
      {stage0_23[8]},
      {stage0_24[8]},
      {stage1_25[8],stage1_24[21],stage1_23[30],stage1_22[45],stage1_21[65]}
   );
   gpc1163_5 gpc288 (
      {stage0_21[91], stage0_21[92], stage0_21[93]},
      {stage0_22[132], stage0_22[133], stage0_22[134], stage0_22[135], stage0_22[136], stage0_22[137]},
      {stage0_23[9]},
      {stage0_24[9]},
      {stage1_25[9],stage1_24[22],stage1_23[31],stage1_22[46],stage1_21[66]}
   );
   gpc606_5 gpc289 (
      {stage0_21[94], stage0_21[95], stage0_21[96], stage0_21[97], stage0_21[98], stage0_21[99]},
      {stage0_23[10], stage0_23[11], stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15]},
      {stage1_25[10],stage1_24[23],stage1_23[32],stage1_22[47],stage1_21[67]}
   );
   gpc606_5 gpc290 (
      {stage0_21[100], stage0_21[101], stage0_21[102], stage0_21[103], stage0_21[104], stage0_21[105]},
      {stage0_23[16], stage0_23[17], stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21]},
      {stage1_25[11],stage1_24[24],stage1_23[33],stage1_22[48],stage1_21[68]}
   );
   gpc606_5 gpc291 (
      {stage0_21[106], stage0_21[107], stage0_21[108], stage0_21[109], stage0_21[110], stage0_21[111]},
      {stage0_23[22], stage0_23[23], stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27]},
      {stage1_25[12],stage1_24[25],stage1_23[34],stage1_22[49],stage1_21[69]}
   );
   gpc606_5 gpc292 (
      {stage0_21[112], stage0_21[113], stage0_21[114], stage0_21[115], stage0_21[116], stage0_21[117]},
      {stage0_23[28], stage0_23[29], stage0_23[30], stage0_23[31], stage0_23[32], stage0_23[33]},
      {stage1_25[13],stage1_24[26],stage1_23[35],stage1_22[50],stage1_21[70]}
   );
   gpc606_5 gpc293 (
      {stage0_21[118], stage0_21[119], stage0_21[120], stage0_21[121], stage0_21[122], stage0_21[123]},
      {stage0_23[34], stage0_23[35], stage0_23[36], stage0_23[37], stage0_23[38], stage0_23[39]},
      {stage1_25[14],stage1_24[27],stage1_23[36],stage1_22[51],stage1_21[71]}
   );
   gpc606_5 gpc294 (
      {stage0_21[124], stage0_21[125], stage0_21[126], stage0_21[127], stage0_21[128], stage0_21[129]},
      {stage0_23[40], stage0_23[41], stage0_23[42], stage0_23[43], stage0_23[44], stage0_23[45]},
      {stage1_25[15],stage1_24[28],stage1_23[37],stage1_22[52],stage1_21[72]}
   );
   gpc606_5 gpc295 (
      {stage0_21[130], stage0_21[131], stage0_21[132], stage0_21[133], stage0_21[134], stage0_21[135]},
      {stage0_23[46], stage0_23[47], stage0_23[48], stage0_23[49], stage0_23[50], stage0_23[51]},
      {stage1_25[16],stage1_24[29],stage1_23[38],stage1_22[53],stage1_21[73]}
   );
   gpc606_5 gpc296 (
      {stage0_21[136], stage0_21[137], stage0_21[138], stage0_21[139], stage0_21[140], stage0_21[141]},
      {stage0_23[52], stage0_23[53], stage0_23[54], stage0_23[55], stage0_23[56], stage0_23[57]},
      {stage1_25[17],stage1_24[30],stage1_23[39],stage1_22[54],stage1_21[74]}
   );
   gpc606_5 gpc297 (
      {stage0_21[142], stage0_21[143], stage0_21[144], stage0_21[145], stage0_21[146], stage0_21[147]},
      {stage0_23[58], stage0_23[59], stage0_23[60], stage0_23[61], stage0_23[62], stage0_23[63]},
      {stage1_25[18],stage1_24[31],stage1_23[40],stage1_22[55],stage1_21[75]}
   );
   gpc606_5 gpc298 (
      {stage0_21[148], stage0_21[149], stage0_21[150], stage0_21[151], stage0_21[152], stage0_21[153]},
      {stage0_23[64], stage0_23[65], stage0_23[66], stage0_23[67], stage0_23[68], stage0_23[69]},
      {stage1_25[19],stage1_24[32],stage1_23[41],stage1_22[56],stage1_21[76]}
   );
   gpc606_5 gpc299 (
      {stage0_21[154], stage0_21[155], stage0_21[156], stage0_21[157], stage0_21[158], stage0_21[159]},
      {stage0_23[70], stage0_23[71], stage0_23[72], stage0_23[73], stage0_23[74], stage0_23[75]},
      {stage1_25[20],stage1_24[33],stage1_23[42],stage1_22[57],stage1_21[77]}
   );
   gpc606_5 gpc300 (
      {stage0_23[76], stage0_23[77], stage0_23[78], stage0_23[79], stage0_23[80], stage0_23[81]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[0],stage1_25[21],stage1_24[34],stage1_23[43]}
   );
   gpc606_5 gpc301 (
      {stage0_23[82], stage0_23[83], stage0_23[84], stage0_23[85], stage0_23[86], stage0_23[87]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[1],stage1_25[22],stage1_24[35],stage1_23[44]}
   );
   gpc606_5 gpc302 (
      {stage0_23[88], stage0_23[89], stage0_23[90], stage0_23[91], stage0_23[92], stage0_23[93]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[2],stage1_25[23],stage1_24[36],stage1_23[45]}
   );
   gpc606_5 gpc303 (
      {stage0_23[94], stage0_23[95], stage0_23[96], stage0_23[97], stage0_23[98], stage0_23[99]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[3],stage1_25[24],stage1_24[37],stage1_23[46]}
   );
   gpc606_5 gpc304 (
      {stage0_23[100], stage0_23[101], stage0_23[102], stage0_23[103], stage0_23[104], stage0_23[105]},
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage1_27[4],stage1_26[4],stage1_25[25],stage1_24[38],stage1_23[47]}
   );
   gpc606_5 gpc305 (
      {stage0_23[106], stage0_23[107], stage0_23[108], stage0_23[109], stage0_23[110], stage0_23[111]},
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage1_27[5],stage1_26[5],stage1_25[26],stage1_24[39],stage1_23[48]}
   );
   gpc615_5 gpc306 (
      {stage0_23[112], stage0_23[113], stage0_23[114], stage0_23[115], stage0_23[116]},
      {stage0_24[10]},
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage1_27[6],stage1_26[6],stage1_25[27],stage1_24[40],stage1_23[49]}
   );
   gpc615_5 gpc307 (
      {stage0_23[117], stage0_23[118], stage0_23[119], stage0_23[120], stage0_23[121]},
      {stage0_24[11]},
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46], stage0_25[47]},
      {stage1_27[7],stage1_26[7],stage1_25[28],stage1_24[41],stage1_23[50]}
   );
   gpc606_5 gpc308 (
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[8],stage1_26[8],stage1_25[29],stage1_24[42]}
   );
   gpc606_5 gpc309 (
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[9],stage1_26[9],stage1_25[30],stage1_24[43]}
   );
   gpc606_5 gpc310 (
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[10],stage1_26[10],stage1_25[31],stage1_24[44]}
   );
   gpc606_5 gpc311 (
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[11],stage1_26[11],stage1_25[32],stage1_24[45]}
   );
   gpc606_5 gpc312 (
      {stage0_24[36], stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[12],stage1_26[12],stage1_25[33],stage1_24[46]}
   );
   gpc606_5 gpc313 (
      {stage0_24[42], stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[13],stage1_26[13],stage1_25[34],stage1_24[47]}
   );
   gpc606_5 gpc314 (
      {stage0_24[48], stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[14],stage1_26[14],stage1_25[35],stage1_24[48]}
   );
   gpc606_5 gpc315 (
      {stage0_24[54], stage0_24[55], stage0_24[56], stage0_24[57], stage0_24[58], stage0_24[59]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[15],stage1_26[15],stage1_25[36],stage1_24[49]}
   );
   gpc606_5 gpc316 (
      {stage0_24[60], stage0_24[61], stage0_24[62], stage0_24[63], stage0_24[64], stage0_24[65]},
      {stage0_26[48], stage0_26[49], stage0_26[50], stage0_26[51], stage0_26[52], stage0_26[53]},
      {stage1_28[8],stage1_27[16],stage1_26[16],stage1_25[37],stage1_24[50]}
   );
   gpc606_5 gpc317 (
      {stage0_24[66], stage0_24[67], stage0_24[68], stage0_24[69], stage0_24[70], stage0_24[71]},
      {stage0_26[54], stage0_26[55], stage0_26[56], stage0_26[57], stage0_26[58], stage0_26[59]},
      {stage1_28[9],stage1_27[17],stage1_26[17],stage1_25[38],stage1_24[51]}
   );
   gpc606_5 gpc318 (
      {stage0_24[72], stage0_24[73], stage0_24[74], stage0_24[75], stage0_24[76], stage0_24[77]},
      {stage0_26[60], stage0_26[61], stage0_26[62], stage0_26[63], stage0_26[64], stage0_26[65]},
      {stage1_28[10],stage1_27[18],stage1_26[18],stage1_25[39],stage1_24[52]}
   );
   gpc606_5 gpc319 (
      {stage0_24[78], stage0_24[79], stage0_24[80], stage0_24[81], stage0_24[82], stage0_24[83]},
      {stage0_26[66], stage0_26[67], stage0_26[68], stage0_26[69], stage0_26[70], stage0_26[71]},
      {stage1_28[11],stage1_27[19],stage1_26[19],stage1_25[40],stage1_24[53]}
   );
   gpc606_5 gpc320 (
      {stage0_24[84], stage0_24[85], stage0_24[86], stage0_24[87], stage0_24[88], stage0_24[89]},
      {stage0_26[72], stage0_26[73], stage0_26[74], stage0_26[75], stage0_26[76], stage0_26[77]},
      {stage1_28[12],stage1_27[20],stage1_26[20],stage1_25[41],stage1_24[54]}
   );
   gpc606_5 gpc321 (
      {stage0_24[90], stage0_24[91], stage0_24[92], stage0_24[93], stage0_24[94], stage0_24[95]},
      {stage0_26[78], stage0_26[79], stage0_26[80], stage0_26[81], stage0_26[82], stage0_26[83]},
      {stage1_28[13],stage1_27[21],stage1_26[21],stage1_25[42],stage1_24[55]}
   );
   gpc606_5 gpc322 (
      {stage0_24[96], stage0_24[97], stage0_24[98], stage0_24[99], stage0_24[100], stage0_24[101]},
      {stage0_26[84], stage0_26[85], stage0_26[86], stage0_26[87], stage0_26[88], stage0_26[89]},
      {stage1_28[14],stage1_27[22],stage1_26[22],stage1_25[43],stage1_24[56]}
   );
   gpc606_5 gpc323 (
      {stage0_24[102], stage0_24[103], stage0_24[104], stage0_24[105], stage0_24[106], stage0_24[107]},
      {stage0_26[90], stage0_26[91], stage0_26[92], stage0_26[93], stage0_26[94], stage0_26[95]},
      {stage1_28[15],stage1_27[23],stage1_26[23],stage1_25[44],stage1_24[57]}
   );
   gpc606_5 gpc324 (
      {stage0_24[108], stage0_24[109], stage0_24[110], stage0_24[111], stage0_24[112], stage0_24[113]},
      {stage0_26[96], stage0_26[97], stage0_26[98], stage0_26[99], stage0_26[100], stage0_26[101]},
      {stage1_28[16],stage1_27[24],stage1_26[24],stage1_25[45],stage1_24[58]}
   );
   gpc606_5 gpc325 (
      {stage0_24[114], stage0_24[115], stage0_24[116], stage0_24[117], stage0_24[118], stage0_24[119]},
      {stage0_26[102], stage0_26[103], stage0_26[104], stage0_26[105], stage0_26[106], stage0_26[107]},
      {stage1_28[17],stage1_27[25],stage1_26[25],stage1_25[46],stage1_24[59]}
   );
   gpc606_5 gpc326 (
      {stage0_24[120], stage0_24[121], stage0_24[122], stage0_24[123], stage0_24[124], stage0_24[125]},
      {stage0_26[108], stage0_26[109], stage0_26[110], stage0_26[111], stage0_26[112], stage0_26[113]},
      {stage1_28[18],stage1_27[26],stage1_26[26],stage1_25[47],stage1_24[60]}
   );
   gpc606_5 gpc327 (
      {stage0_24[126], stage0_24[127], stage0_24[128], stage0_24[129], stage0_24[130], stage0_24[131]},
      {stage0_26[114], stage0_26[115], stage0_26[116], stage0_26[117], stage0_26[118], stage0_26[119]},
      {stage1_28[19],stage1_27[27],stage1_26[27],stage1_25[48],stage1_24[61]}
   );
   gpc606_5 gpc328 (
      {stage0_24[132], stage0_24[133], stage0_24[134], stage0_24[135], stage0_24[136], stage0_24[137]},
      {stage0_26[120], stage0_26[121], stage0_26[122], stage0_26[123], stage0_26[124], stage0_26[125]},
      {stage1_28[20],stage1_27[28],stage1_26[28],stage1_25[49],stage1_24[62]}
   );
   gpc606_5 gpc329 (
      {stage0_24[138], stage0_24[139], stage0_24[140], stage0_24[141], stage0_24[142], stage0_24[143]},
      {stage0_26[126], stage0_26[127], stage0_26[128], stage0_26[129], stage0_26[130], stage0_26[131]},
      {stage1_28[21],stage1_27[29],stage1_26[29],stage1_25[50],stage1_24[63]}
   );
   gpc606_5 gpc330 (
      {stage0_24[144], stage0_24[145], stage0_24[146], stage0_24[147], stage0_24[148], stage0_24[149]},
      {stage0_26[132], stage0_26[133], stage0_26[134], stage0_26[135], stage0_26[136], stage0_26[137]},
      {stage1_28[22],stage1_27[30],stage1_26[30],stage1_25[51],stage1_24[64]}
   );
   gpc606_5 gpc331 (
      {stage0_24[150], stage0_24[151], stage0_24[152], stage0_24[153], stage0_24[154], stage0_24[155]},
      {stage0_26[138], stage0_26[139], stage0_26[140], stage0_26[141], stage0_26[142], stage0_26[143]},
      {stage1_28[23],stage1_27[31],stage1_26[31],stage1_25[52],stage1_24[65]}
   );
   gpc606_5 gpc332 (
      {stage0_24[156], stage0_24[157], stage0_24[158], stage0_24[159], stage0_24[160], stage0_24[161]},
      {stage0_26[144], stage0_26[145], stage0_26[146], stage0_26[147], stage0_26[148], stage0_26[149]},
      {stage1_28[24],stage1_27[32],stage1_26[32],stage1_25[53],stage1_24[66]}
   );
   gpc606_5 gpc333 (
      {stage0_25[48], stage0_25[49], stage0_25[50], stage0_25[51], stage0_25[52], stage0_25[53]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[25],stage1_27[33],stage1_26[33],stage1_25[54]}
   );
   gpc606_5 gpc334 (
      {stage0_25[54], stage0_25[55], stage0_25[56], stage0_25[57], stage0_25[58], stage0_25[59]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[26],stage1_27[34],stage1_26[34],stage1_25[55]}
   );
   gpc606_5 gpc335 (
      {stage0_25[60], stage0_25[61], stage0_25[62], stage0_25[63], stage0_25[64], stage0_25[65]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[27],stage1_27[35],stage1_26[35],stage1_25[56]}
   );
   gpc606_5 gpc336 (
      {stage0_25[66], stage0_25[67], stage0_25[68], stage0_25[69], stage0_25[70], stage0_25[71]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[28],stage1_27[36],stage1_26[36],stage1_25[57]}
   );
   gpc606_5 gpc337 (
      {stage0_25[72], stage0_25[73], stage0_25[74], stage0_25[75], stage0_25[76], stage0_25[77]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[29],stage1_27[37],stage1_26[37],stage1_25[58]}
   );
   gpc606_5 gpc338 (
      {stage0_25[78], stage0_25[79], stage0_25[80], stage0_25[81], stage0_25[82], stage0_25[83]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[30],stage1_27[38],stage1_26[38],stage1_25[59]}
   );
   gpc606_5 gpc339 (
      {stage0_25[84], stage0_25[85], stage0_25[86], stage0_25[87], stage0_25[88], stage0_25[89]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[31],stage1_27[39],stage1_26[39],stage1_25[60]}
   );
   gpc606_5 gpc340 (
      {stage0_25[90], stage0_25[91], stage0_25[92], stage0_25[93], stage0_25[94], stage0_25[95]},
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage1_29[7],stage1_28[32],stage1_27[40],stage1_26[40],stage1_25[61]}
   );
   gpc606_5 gpc341 (
      {stage0_25[96], stage0_25[97], stage0_25[98], stage0_25[99], stage0_25[100], stage0_25[101]},
      {stage0_27[48], stage0_27[49], stage0_27[50], stage0_27[51], stage0_27[52], stage0_27[53]},
      {stage1_29[8],stage1_28[33],stage1_27[41],stage1_26[41],stage1_25[62]}
   );
   gpc606_5 gpc342 (
      {stage0_25[102], stage0_25[103], stage0_25[104], stage0_25[105], stage0_25[106], stage0_25[107]},
      {stage0_27[54], stage0_27[55], stage0_27[56], stage0_27[57], stage0_27[58], stage0_27[59]},
      {stage1_29[9],stage1_28[34],stage1_27[42],stage1_26[42],stage1_25[63]}
   );
   gpc615_5 gpc343 (
      {stage0_25[108], stage0_25[109], stage0_25[110], stage0_25[111], stage0_25[112]},
      {stage0_26[150]},
      {stage0_27[60], stage0_27[61], stage0_27[62], stage0_27[63], stage0_27[64], stage0_27[65]},
      {stage1_29[10],stage1_28[35],stage1_27[43],stage1_26[43],stage1_25[64]}
   );
   gpc615_5 gpc344 (
      {stage0_25[113], stage0_25[114], stage0_25[115], stage0_25[116], stage0_25[117]},
      {stage0_26[151]},
      {stage0_27[66], stage0_27[67], stage0_27[68], stage0_27[69], stage0_27[70], stage0_27[71]},
      {stage1_29[11],stage1_28[36],stage1_27[44],stage1_26[44],stage1_25[65]}
   );
   gpc615_5 gpc345 (
      {stage0_25[118], stage0_25[119], stage0_25[120], stage0_25[121], stage0_25[122]},
      {stage0_26[152]},
      {stage0_27[72], stage0_27[73], stage0_27[74], stage0_27[75], stage0_27[76], stage0_27[77]},
      {stage1_29[12],stage1_28[37],stage1_27[45],stage1_26[45],stage1_25[66]}
   );
   gpc615_5 gpc346 (
      {stage0_25[123], stage0_25[124], stage0_25[125], stage0_25[126], stage0_25[127]},
      {stage0_26[153]},
      {stage0_27[78], stage0_27[79], stage0_27[80], stage0_27[81], stage0_27[82], stage0_27[83]},
      {stage1_29[13],stage1_28[38],stage1_27[46],stage1_26[46],stage1_25[67]}
   );
   gpc615_5 gpc347 (
      {stage0_25[128], stage0_25[129], stage0_25[130], stage0_25[131], stage0_25[132]},
      {stage0_26[154]},
      {stage0_27[84], stage0_27[85], stage0_27[86], stage0_27[87], stage0_27[88], stage0_27[89]},
      {stage1_29[14],stage1_28[39],stage1_27[47],stage1_26[47],stage1_25[68]}
   );
   gpc615_5 gpc348 (
      {stage0_25[133], stage0_25[134], stage0_25[135], stage0_25[136], stage0_25[137]},
      {stage0_26[155]},
      {stage0_27[90], stage0_27[91], stage0_27[92], stage0_27[93], stage0_27[94], stage0_27[95]},
      {stage1_29[15],stage1_28[40],stage1_27[48],stage1_26[48],stage1_25[69]}
   );
   gpc615_5 gpc349 (
      {stage0_25[138], stage0_25[139], stage0_25[140], stage0_25[141], stage0_25[142]},
      {stage0_26[156]},
      {stage0_27[96], stage0_27[97], stage0_27[98], stage0_27[99], stage0_27[100], stage0_27[101]},
      {stage1_29[16],stage1_28[41],stage1_27[49],stage1_26[49],stage1_25[70]}
   );
   gpc615_5 gpc350 (
      {stage0_25[143], stage0_25[144], stage0_25[145], stage0_25[146], stage0_25[147]},
      {stage0_26[157]},
      {stage0_27[102], stage0_27[103], stage0_27[104], stage0_27[105], stage0_27[106], stage0_27[107]},
      {stage1_29[17],stage1_28[42],stage1_27[50],stage1_26[50],stage1_25[71]}
   );
   gpc615_5 gpc351 (
      {stage0_25[148], stage0_25[149], stage0_25[150], stage0_25[151], stage0_25[152]},
      {stage0_26[158]},
      {stage0_27[108], stage0_27[109], stage0_27[110], stage0_27[111], stage0_27[112], stage0_27[113]},
      {stage1_29[18],stage1_28[43],stage1_27[51],stage1_26[51],stage1_25[72]}
   );
   gpc615_5 gpc352 (
      {stage0_25[153], stage0_25[154], stage0_25[155], stage0_25[156], stage0_25[157]},
      {stage0_26[159]},
      {stage0_27[114], stage0_27[115], stage0_27[116], stage0_27[117], stage0_27[118], stage0_27[119]},
      {stage1_29[19],stage1_28[44],stage1_27[52],stage1_26[52],stage1_25[73]}
   );
   gpc615_5 gpc353 (
      {stage0_27[120], stage0_27[121], stage0_27[122], stage0_27[123], stage0_27[124]},
      {stage0_28[0]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[0],stage1_29[20],stage1_28[45],stage1_27[53]}
   );
   gpc615_5 gpc354 (
      {stage0_27[125], stage0_27[126], stage0_27[127], stage0_27[128], stage0_27[129]},
      {stage0_28[1]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[1],stage1_29[21],stage1_28[46],stage1_27[54]}
   );
   gpc615_5 gpc355 (
      {stage0_27[130], stage0_27[131], stage0_27[132], stage0_27[133], stage0_27[134]},
      {stage0_28[2]},
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage1_31[2],stage1_30[2],stage1_29[22],stage1_28[47],stage1_27[55]}
   );
   gpc615_5 gpc356 (
      {stage0_27[135], stage0_27[136], stage0_27[137], stage0_27[138], stage0_27[139]},
      {stage0_28[3]},
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage1_31[3],stage1_30[3],stage1_29[23],stage1_28[48],stage1_27[56]}
   );
   gpc615_5 gpc357 (
      {stage0_27[140], stage0_27[141], stage0_27[142], stage0_27[143], stage0_27[144]},
      {stage0_28[4]},
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage1_31[4],stage1_30[4],stage1_29[24],stage1_28[49],stage1_27[57]}
   );
   gpc615_5 gpc358 (
      {stage0_27[145], stage0_27[146], stage0_27[147], stage0_27[148], stage0_27[149]},
      {stage0_28[5]},
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage1_31[5],stage1_30[5],stage1_29[25],stage1_28[50],stage1_27[58]}
   );
   gpc615_5 gpc359 (
      {stage0_27[150], stage0_27[151], stage0_27[152], stage0_27[153], stage0_27[154]},
      {stage0_28[6]},
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage1_31[6],stage1_30[6],stage1_29[26],stage1_28[51],stage1_27[59]}
   );
   gpc2135_5 gpc360 (
      {stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage0_29[42], stage0_29[43], stage0_29[44]},
      {stage0_30[0]},
      {stage0_31[0], stage0_31[1]},
      {stage1_32[0],stage1_31[7],stage1_30[7],stage1_29[27],stage1_28[52]}
   );
   gpc606_5 gpc361 (
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5], stage0_30[6]},
      {stage1_32[1],stage1_31[8],stage1_30[8],stage1_29[28],stage1_28[53]}
   );
   gpc606_5 gpc362 (
      {stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23]},
      {stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11], stage0_30[12]},
      {stage1_32[2],stage1_31[9],stage1_30[9],stage1_29[29],stage1_28[54]}
   );
   gpc606_5 gpc363 (
      {stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29]},
      {stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17], stage0_30[18]},
      {stage1_32[3],stage1_31[10],stage1_30[10],stage1_29[30],stage1_28[55]}
   );
   gpc606_5 gpc364 (
      {stage0_28[30], stage0_28[31], stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35]},
      {stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23], stage0_30[24]},
      {stage1_32[4],stage1_31[11],stage1_30[11],stage1_29[31],stage1_28[56]}
   );
   gpc606_5 gpc365 (
      {stage0_28[36], stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41]},
      {stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29], stage0_30[30]},
      {stage1_32[5],stage1_31[12],stage1_30[12],stage1_29[32],stage1_28[57]}
   );
   gpc606_5 gpc366 (
      {stage0_28[42], stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47]},
      {stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35], stage0_30[36]},
      {stage1_32[6],stage1_31[13],stage1_30[13],stage1_29[33],stage1_28[58]}
   );
   gpc606_5 gpc367 (
      {stage0_28[48], stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53]},
      {stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41], stage0_30[42]},
      {stage1_32[7],stage1_31[14],stage1_30[14],stage1_29[34],stage1_28[59]}
   );
   gpc606_5 gpc368 (
      {stage0_28[54], stage0_28[55], stage0_28[56], stage0_28[57], stage0_28[58], stage0_28[59]},
      {stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47], stage0_30[48]},
      {stage1_32[8],stage1_31[15],stage1_30[15],stage1_29[35],stage1_28[60]}
   );
   gpc606_5 gpc369 (
      {stage0_28[60], stage0_28[61], stage0_28[62], stage0_28[63], stage0_28[64], stage0_28[65]},
      {stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53], stage0_30[54]},
      {stage1_32[9],stage1_31[16],stage1_30[16],stage1_29[36],stage1_28[61]}
   );
   gpc606_5 gpc370 (
      {stage0_28[66], stage0_28[67], stage0_28[68], stage0_28[69], stage0_28[70], stage0_28[71]},
      {stage0_30[55], stage0_30[56], stage0_30[57], stage0_30[58], stage0_30[59], stage0_30[60]},
      {stage1_32[10],stage1_31[17],stage1_30[17],stage1_29[37],stage1_28[62]}
   );
   gpc606_5 gpc371 (
      {stage0_28[72], stage0_28[73], stage0_28[74], stage0_28[75], stage0_28[76], stage0_28[77]},
      {stage0_30[61], stage0_30[62], stage0_30[63], stage0_30[64], stage0_30[65], stage0_30[66]},
      {stage1_32[11],stage1_31[18],stage1_30[18],stage1_29[38],stage1_28[63]}
   );
   gpc606_5 gpc372 (
      {stage0_28[78], stage0_28[79], stage0_28[80], stage0_28[81], stage0_28[82], stage0_28[83]},
      {stage0_30[67], stage0_30[68], stage0_30[69], stage0_30[70], stage0_30[71], stage0_30[72]},
      {stage1_32[12],stage1_31[19],stage1_30[19],stage1_29[39],stage1_28[64]}
   );
   gpc606_5 gpc373 (
      {stage0_28[84], stage0_28[85], stage0_28[86], stage0_28[87], stage0_28[88], stage0_28[89]},
      {stage0_30[73], stage0_30[74], stage0_30[75], stage0_30[76], stage0_30[77], stage0_30[78]},
      {stage1_32[13],stage1_31[20],stage1_30[20],stage1_29[40],stage1_28[65]}
   );
   gpc606_5 gpc374 (
      {stage0_28[90], stage0_28[91], stage0_28[92], stage0_28[93], stage0_28[94], stage0_28[95]},
      {stage0_30[79], stage0_30[80], stage0_30[81], stage0_30[82], stage0_30[83], stage0_30[84]},
      {stage1_32[14],stage1_31[21],stage1_30[21],stage1_29[41],stage1_28[66]}
   );
   gpc606_5 gpc375 (
      {stage0_28[96], stage0_28[97], stage0_28[98], stage0_28[99], stage0_28[100], stage0_28[101]},
      {stage0_30[85], stage0_30[86], stage0_30[87], stage0_30[88], stage0_30[89], stage0_30[90]},
      {stage1_32[15],stage1_31[22],stage1_30[22],stage1_29[42],stage1_28[67]}
   );
   gpc606_5 gpc376 (
      {stage0_28[102], stage0_28[103], stage0_28[104], stage0_28[105], stage0_28[106], stage0_28[107]},
      {stage0_30[91], stage0_30[92], stage0_30[93], stage0_30[94], stage0_30[95], stage0_30[96]},
      {stage1_32[16],stage1_31[23],stage1_30[23],stage1_29[43],stage1_28[68]}
   );
   gpc606_5 gpc377 (
      {stage0_28[108], stage0_28[109], stage0_28[110], stage0_28[111], stage0_28[112], stage0_28[113]},
      {stage0_30[97], stage0_30[98], stage0_30[99], stage0_30[100], stage0_30[101], stage0_30[102]},
      {stage1_32[17],stage1_31[24],stage1_30[24],stage1_29[44],stage1_28[69]}
   );
   gpc606_5 gpc378 (
      {stage0_28[114], stage0_28[115], stage0_28[116], stage0_28[117], stage0_28[118], stage0_28[119]},
      {stage0_30[103], stage0_30[104], stage0_30[105], stage0_30[106], stage0_30[107], stage0_30[108]},
      {stage1_32[18],stage1_31[25],stage1_30[25],stage1_29[45],stage1_28[70]}
   );
   gpc606_5 gpc379 (
      {stage0_28[120], stage0_28[121], stage0_28[122], stage0_28[123], stage0_28[124], stage0_28[125]},
      {stage0_30[109], stage0_30[110], stage0_30[111], stage0_30[112], stage0_30[113], stage0_30[114]},
      {stage1_32[19],stage1_31[26],stage1_30[26],stage1_29[46],stage1_28[71]}
   );
   gpc606_5 gpc380 (
      {stage0_28[126], stage0_28[127], stage0_28[128], stage0_28[129], stage0_28[130], stage0_28[131]},
      {stage0_30[115], stage0_30[116], stage0_30[117], stage0_30[118], stage0_30[119], stage0_30[120]},
      {stage1_32[20],stage1_31[27],stage1_30[27],stage1_29[47],stage1_28[72]}
   );
   gpc606_5 gpc381 (
      {stage0_28[132], stage0_28[133], stage0_28[134], stage0_28[135], stage0_28[136], stage0_28[137]},
      {stage0_30[121], stage0_30[122], stage0_30[123], stage0_30[124], stage0_30[125], stage0_30[126]},
      {stage1_32[21],stage1_31[28],stage1_30[28],stage1_29[48],stage1_28[73]}
   );
   gpc606_5 gpc382 (
      {stage0_28[138], stage0_28[139], stage0_28[140], stage0_28[141], stage0_28[142], stage0_28[143]},
      {stage0_30[127], stage0_30[128], stage0_30[129], stage0_30[130], stage0_30[131], stage0_30[132]},
      {stage1_32[22],stage1_31[29],stage1_30[29],stage1_29[49],stage1_28[74]}
   );
   gpc606_5 gpc383 (
      {stage0_28[144], stage0_28[145], stage0_28[146], stage0_28[147], stage0_28[148], stage0_28[149]},
      {stage0_30[133], stage0_30[134], stage0_30[135], stage0_30[136], stage0_30[137], stage0_30[138]},
      {stage1_32[23],stage1_31[30],stage1_30[30],stage1_29[50],stage1_28[75]}
   );
   gpc606_5 gpc384 (
      {stage0_28[150], stage0_28[151], stage0_28[152], stage0_28[153], stage0_28[154], stage0_28[155]},
      {stage0_30[139], stage0_30[140], stage0_30[141], stage0_30[142], stage0_30[143], stage0_30[144]},
      {stage1_32[24],stage1_31[31],stage1_30[31],stage1_29[51],stage1_28[76]}
   );
   gpc606_5 gpc385 (
      {stage0_28[156], stage0_28[157], stage0_28[158], stage0_28[159], stage0_28[160], stage0_28[161]},
      {stage0_30[145], stage0_30[146], stage0_30[147], stage0_30[148], stage0_30[149], stage0_30[150]},
      {stage1_32[25],stage1_31[32],stage1_30[32],stage1_29[52],stage1_28[77]}
   );
   gpc606_5 gpc386 (
      {stage0_29[45], stage0_29[46], stage0_29[47], stage0_29[48], stage0_29[49], stage0_29[50]},
      {stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5], stage0_31[6], stage0_31[7]},
      {stage1_33[0],stage1_32[26],stage1_31[33],stage1_30[33],stage1_29[53]}
   );
   gpc606_5 gpc387 (
      {stage0_29[51], stage0_29[52], stage0_29[53], stage0_29[54], stage0_29[55], stage0_29[56]},
      {stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11], stage0_31[12], stage0_31[13]},
      {stage1_33[1],stage1_32[27],stage1_31[34],stage1_30[34],stage1_29[54]}
   );
   gpc606_5 gpc388 (
      {stage0_29[57], stage0_29[58], stage0_29[59], stage0_29[60], stage0_29[61], stage0_29[62]},
      {stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17], stage0_31[18], stage0_31[19]},
      {stage1_33[2],stage1_32[28],stage1_31[35],stage1_30[35],stage1_29[55]}
   );
   gpc606_5 gpc389 (
      {stage0_29[63], stage0_29[64], stage0_29[65], stage0_29[66], stage0_29[67], stage0_29[68]},
      {stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23], stage0_31[24], stage0_31[25]},
      {stage1_33[3],stage1_32[29],stage1_31[36],stage1_30[36],stage1_29[56]}
   );
   gpc606_5 gpc390 (
      {stage0_29[69], stage0_29[70], stage0_29[71], stage0_29[72], stage0_29[73], stage0_29[74]},
      {stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29], stage0_31[30], stage0_31[31]},
      {stage1_33[4],stage1_32[30],stage1_31[37],stage1_30[37],stage1_29[57]}
   );
   gpc606_5 gpc391 (
      {stage0_29[75], stage0_29[76], stage0_29[77], stage0_29[78], stage0_29[79], stage0_29[80]},
      {stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35], stage0_31[36], stage0_31[37]},
      {stage1_33[5],stage1_32[31],stage1_31[38],stage1_30[38],stage1_29[58]}
   );
   gpc606_5 gpc392 (
      {stage0_29[81], stage0_29[82], stage0_29[83], stage0_29[84], stage0_29[85], stage0_29[86]},
      {stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41], stage0_31[42], stage0_31[43]},
      {stage1_33[6],stage1_32[32],stage1_31[39],stage1_30[39],stage1_29[59]}
   );
   gpc606_5 gpc393 (
      {stage0_29[87], stage0_29[88], stage0_29[89], stage0_29[90], stage0_29[91], stage0_29[92]},
      {stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47], stage0_31[48], stage0_31[49]},
      {stage1_33[7],stage1_32[33],stage1_31[40],stage1_30[40],stage1_29[60]}
   );
   gpc606_5 gpc394 (
      {stage0_29[93], stage0_29[94], stage0_29[95], stage0_29[96], stage0_29[97], stage0_29[98]},
      {stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53], stage0_31[54], stage0_31[55]},
      {stage1_33[8],stage1_32[34],stage1_31[41],stage1_30[41],stage1_29[61]}
   );
   gpc606_5 gpc395 (
      {stage0_29[99], stage0_29[100], stage0_29[101], stage0_29[102], stage0_29[103], stage0_29[104]},
      {stage0_31[56], stage0_31[57], stage0_31[58], stage0_31[59], stage0_31[60], stage0_31[61]},
      {stage1_33[9],stage1_32[35],stage1_31[42],stage1_30[42],stage1_29[62]}
   );
   gpc606_5 gpc396 (
      {stage0_29[105], stage0_29[106], stage0_29[107], stage0_29[108], stage0_29[109], stage0_29[110]},
      {stage0_31[62], stage0_31[63], stage0_31[64], stage0_31[65], stage0_31[66], stage0_31[67]},
      {stage1_33[10],stage1_32[36],stage1_31[43],stage1_30[43],stage1_29[63]}
   );
   gpc606_5 gpc397 (
      {stage0_29[111], stage0_29[112], stage0_29[113], stage0_29[114], stage0_29[115], stage0_29[116]},
      {stage0_31[68], stage0_31[69], stage0_31[70], stage0_31[71], stage0_31[72], stage0_31[73]},
      {stage1_33[11],stage1_32[37],stage1_31[44],stage1_30[44],stage1_29[64]}
   );
   gpc606_5 gpc398 (
      {stage0_29[117], stage0_29[118], stage0_29[119], stage0_29[120], stage0_29[121], stage0_29[122]},
      {stage0_31[74], stage0_31[75], stage0_31[76], stage0_31[77], stage0_31[78], stage0_31[79]},
      {stage1_33[12],stage1_32[38],stage1_31[45],stage1_30[45],stage1_29[65]}
   );
   gpc606_5 gpc399 (
      {stage0_29[123], stage0_29[124], stage0_29[125], stage0_29[126], stage0_29[127], stage0_29[128]},
      {stage0_31[80], stage0_31[81], stage0_31[82], stage0_31[83], stage0_31[84], stage0_31[85]},
      {stage1_33[13],stage1_32[39],stage1_31[46],stage1_30[46],stage1_29[66]}
   );
   gpc606_5 gpc400 (
      {stage0_29[129], stage0_29[130], stage0_29[131], stage0_29[132], stage0_29[133], stage0_29[134]},
      {stage0_31[86], stage0_31[87], stage0_31[88], stage0_31[89], stage0_31[90], stage0_31[91]},
      {stage1_33[14],stage1_32[40],stage1_31[47],stage1_30[47],stage1_29[67]}
   );
   gpc606_5 gpc401 (
      {stage0_29[135], stage0_29[136], stage0_29[137], stage0_29[138], stage0_29[139], stage0_29[140]},
      {stage0_31[92], stage0_31[93], stage0_31[94], stage0_31[95], stage0_31[96], stage0_31[97]},
      {stage1_33[15],stage1_32[41],stage1_31[48],stage1_30[48],stage1_29[68]}
   );
   gpc606_5 gpc402 (
      {stage0_29[141], stage0_29[142], stage0_29[143], stage0_29[144], stage0_29[145], stage0_29[146]},
      {stage0_31[98], stage0_31[99], stage0_31[100], stage0_31[101], stage0_31[102], stage0_31[103]},
      {stage1_33[16],stage1_32[42],stage1_31[49],stage1_30[49],stage1_29[69]}
   );
   gpc606_5 gpc403 (
      {stage0_29[147], stage0_29[148], stage0_29[149], stage0_29[150], stage0_29[151], stage0_29[152]},
      {stage0_31[104], stage0_31[105], stage0_31[106], stage0_31[107], stage0_31[108], stage0_31[109]},
      {stage1_33[17],stage1_32[43],stage1_31[50],stage1_30[50],stage1_29[70]}
   );
   gpc606_5 gpc404 (
      {stage0_29[153], stage0_29[154], stage0_29[155], stage0_29[156], stage0_29[157], stage0_29[158]},
      {stage0_31[110], stage0_31[111], stage0_31[112], stage0_31[113], stage0_31[114], stage0_31[115]},
      {stage1_33[18],stage1_32[44],stage1_31[51],stage1_30[51],stage1_29[71]}
   );
   gpc1_1 gpc405 (
      {stage0_0[144]},
      {stage1_0[32]}
   );
   gpc1_1 gpc406 (
      {stage0_0[145]},
      {stage1_0[33]}
   );
   gpc1_1 gpc407 (
      {stage0_0[146]},
      {stage1_0[34]}
   );
   gpc1_1 gpc408 (
      {stage0_0[147]},
      {stage1_0[35]}
   );
   gpc1_1 gpc409 (
      {stage0_0[148]},
      {stage1_0[36]}
   );
   gpc1_1 gpc410 (
      {stage0_0[149]},
      {stage1_0[37]}
   );
   gpc1_1 gpc411 (
      {stage0_0[150]},
      {stage1_0[38]}
   );
   gpc1_1 gpc412 (
      {stage0_0[151]},
      {stage1_0[39]}
   );
   gpc1_1 gpc413 (
      {stage0_0[152]},
      {stage1_0[40]}
   );
   gpc1_1 gpc414 (
      {stage0_0[153]},
      {stage1_0[41]}
   );
   gpc1_1 gpc415 (
      {stage0_0[154]},
      {stage1_0[42]}
   );
   gpc1_1 gpc416 (
      {stage0_0[155]},
      {stage1_0[43]}
   );
   gpc1_1 gpc417 (
      {stage0_0[156]},
      {stage1_0[44]}
   );
   gpc1_1 gpc418 (
      {stage0_0[157]},
      {stage1_0[45]}
   );
   gpc1_1 gpc419 (
      {stage0_0[158]},
      {stage1_0[46]}
   );
   gpc1_1 gpc420 (
      {stage0_0[159]},
      {stage1_0[47]}
   );
   gpc1_1 gpc421 (
      {stage0_0[160]},
      {stage1_0[48]}
   );
   gpc1_1 gpc422 (
      {stage0_0[161]},
      {stage1_0[49]}
   );
   gpc1_1 gpc423 (
      {stage0_1[144]},
      {stage1_1[38]}
   );
   gpc1_1 gpc424 (
      {stage0_1[145]},
      {stage1_1[39]}
   );
   gpc1_1 gpc425 (
      {stage0_1[146]},
      {stage1_1[40]}
   );
   gpc1_1 gpc426 (
      {stage0_1[147]},
      {stage1_1[41]}
   );
   gpc1_1 gpc427 (
      {stage0_1[148]},
      {stage1_1[42]}
   );
   gpc1_1 gpc428 (
      {stage0_1[149]},
      {stage1_1[43]}
   );
   gpc1_1 gpc429 (
      {stage0_1[150]},
      {stage1_1[44]}
   );
   gpc1_1 gpc430 (
      {stage0_1[151]},
      {stage1_1[45]}
   );
   gpc1_1 gpc431 (
      {stage0_1[152]},
      {stage1_1[46]}
   );
   gpc1_1 gpc432 (
      {stage0_1[153]},
      {stage1_1[47]}
   );
   gpc1_1 gpc433 (
      {stage0_1[154]},
      {stage1_1[48]}
   );
   gpc1_1 gpc434 (
      {stage0_1[155]},
      {stage1_1[49]}
   );
   gpc1_1 gpc435 (
      {stage0_1[156]},
      {stage1_1[50]}
   );
   gpc1_1 gpc436 (
      {stage0_1[157]},
      {stage1_1[51]}
   );
   gpc1_1 gpc437 (
      {stage0_1[158]},
      {stage1_1[52]}
   );
   gpc1_1 gpc438 (
      {stage0_1[159]},
      {stage1_1[53]}
   );
   gpc1_1 gpc439 (
      {stage0_1[160]},
      {stage1_1[54]}
   );
   gpc1_1 gpc440 (
      {stage0_1[161]},
      {stage1_1[55]}
   );
   gpc1_1 gpc441 (
      {stage0_3[155]},
      {stage1_3[69]}
   );
   gpc1_1 gpc442 (
      {stage0_3[156]},
      {stage1_3[70]}
   );
   gpc1_1 gpc443 (
      {stage0_3[157]},
      {stage1_3[71]}
   );
   gpc1_1 gpc444 (
      {stage0_3[158]},
      {stage1_3[72]}
   );
   gpc1_1 gpc445 (
      {stage0_3[159]},
      {stage1_3[73]}
   );
   gpc1_1 gpc446 (
      {stage0_3[160]},
      {stage1_3[74]}
   );
   gpc1_1 gpc447 (
      {stage0_3[161]},
      {stage1_3[75]}
   );
   gpc1_1 gpc448 (
      {stage0_4[139]},
      {stage1_4[72]}
   );
   gpc1_1 gpc449 (
      {stage0_4[140]},
      {stage1_4[73]}
   );
   gpc1_1 gpc450 (
      {stage0_4[141]},
      {stage1_4[74]}
   );
   gpc1_1 gpc451 (
      {stage0_4[142]},
      {stage1_4[75]}
   );
   gpc1_1 gpc452 (
      {stage0_4[143]},
      {stage1_4[76]}
   );
   gpc1_1 gpc453 (
      {stage0_4[144]},
      {stage1_4[77]}
   );
   gpc1_1 gpc454 (
      {stage0_4[145]},
      {stage1_4[78]}
   );
   gpc1_1 gpc455 (
      {stage0_4[146]},
      {stage1_4[79]}
   );
   gpc1_1 gpc456 (
      {stage0_4[147]},
      {stage1_4[80]}
   );
   gpc1_1 gpc457 (
      {stage0_4[148]},
      {stage1_4[81]}
   );
   gpc1_1 gpc458 (
      {stage0_4[149]},
      {stage1_4[82]}
   );
   gpc1_1 gpc459 (
      {stage0_4[150]},
      {stage1_4[83]}
   );
   gpc1_1 gpc460 (
      {stage0_4[151]},
      {stage1_4[84]}
   );
   gpc1_1 gpc461 (
      {stage0_4[152]},
      {stage1_4[85]}
   );
   gpc1_1 gpc462 (
      {stage0_4[153]},
      {stage1_4[86]}
   );
   gpc1_1 gpc463 (
      {stage0_4[154]},
      {stage1_4[87]}
   );
   gpc1_1 gpc464 (
      {stage0_4[155]},
      {stage1_4[88]}
   );
   gpc1_1 gpc465 (
      {stage0_4[156]},
      {stage1_4[89]}
   );
   gpc1_1 gpc466 (
      {stage0_4[157]},
      {stage1_4[90]}
   );
   gpc1_1 gpc467 (
      {stage0_4[158]},
      {stage1_4[91]}
   );
   gpc1_1 gpc468 (
      {stage0_4[159]},
      {stage1_4[92]}
   );
   gpc1_1 gpc469 (
      {stage0_4[160]},
      {stage1_4[93]}
   );
   gpc1_1 gpc470 (
      {stage0_4[161]},
      {stage1_4[94]}
   );
   gpc1_1 gpc471 (
      {stage0_6[124]},
      {stage1_6[68]}
   );
   gpc1_1 gpc472 (
      {stage0_6[125]},
      {stage1_6[69]}
   );
   gpc1_1 gpc473 (
      {stage0_6[126]},
      {stage1_6[70]}
   );
   gpc1_1 gpc474 (
      {stage0_6[127]},
      {stage1_6[71]}
   );
   gpc1_1 gpc475 (
      {stage0_6[128]},
      {stage1_6[72]}
   );
   gpc1_1 gpc476 (
      {stage0_6[129]},
      {stage1_6[73]}
   );
   gpc1_1 gpc477 (
      {stage0_6[130]},
      {stage1_6[74]}
   );
   gpc1_1 gpc478 (
      {stage0_6[131]},
      {stage1_6[75]}
   );
   gpc1_1 gpc479 (
      {stage0_6[132]},
      {stage1_6[76]}
   );
   gpc1_1 gpc480 (
      {stage0_6[133]},
      {stage1_6[77]}
   );
   gpc1_1 gpc481 (
      {stage0_6[134]},
      {stage1_6[78]}
   );
   gpc1_1 gpc482 (
      {stage0_6[135]},
      {stage1_6[79]}
   );
   gpc1_1 gpc483 (
      {stage0_6[136]},
      {stage1_6[80]}
   );
   gpc1_1 gpc484 (
      {stage0_6[137]},
      {stage1_6[81]}
   );
   gpc1_1 gpc485 (
      {stage0_6[138]},
      {stage1_6[82]}
   );
   gpc1_1 gpc486 (
      {stage0_6[139]},
      {stage1_6[83]}
   );
   gpc1_1 gpc487 (
      {stage0_6[140]},
      {stage1_6[84]}
   );
   gpc1_1 gpc488 (
      {stage0_6[141]},
      {stage1_6[85]}
   );
   gpc1_1 gpc489 (
      {stage0_6[142]},
      {stage1_6[86]}
   );
   gpc1_1 gpc490 (
      {stage0_6[143]},
      {stage1_6[87]}
   );
   gpc1_1 gpc491 (
      {stage0_6[144]},
      {stage1_6[88]}
   );
   gpc1_1 gpc492 (
      {stage0_6[145]},
      {stage1_6[89]}
   );
   gpc1_1 gpc493 (
      {stage0_6[146]},
      {stage1_6[90]}
   );
   gpc1_1 gpc494 (
      {stage0_6[147]},
      {stage1_6[91]}
   );
   gpc1_1 gpc495 (
      {stage0_6[148]},
      {stage1_6[92]}
   );
   gpc1_1 gpc496 (
      {stage0_6[149]},
      {stage1_6[93]}
   );
   gpc1_1 gpc497 (
      {stage0_6[150]},
      {stage1_6[94]}
   );
   gpc1_1 gpc498 (
      {stage0_6[151]},
      {stage1_6[95]}
   );
   gpc1_1 gpc499 (
      {stage0_6[152]},
      {stage1_6[96]}
   );
   gpc1_1 gpc500 (
      {stage0_6[153]},
      {stage1_6[97]}
   );
   gpc1_1 gpc501 (
      {stage0_6[154]},
      {stage1_6[98]}
   );
   gpc1_1 gpc502 (
      {stage0_6[155]},
      {stage1_6[99]}
   );
   gpc1_1 gpc503 (
      {stage0_6[156]},
      {stage1_6[100]}
   );
   gpc1_1 gpc504 (
      {stage0_6[157]},
      {stage1_6[101]}
   );
   gpc1_1 gpc505 (
      {stage0_6[158]},
      {stage1_6[102]}
   );
   gpc1_1 gpc506 (
      {stage0_6[159]},
      {stage1_6[103]}
   );
   gpc1_1 gpc507 (
      {stage0_6[160]},
      {stage1_6[104]}
   );
   gpc1_1 gpc508 (
      {stage0_6[161]},
      {stage1_6[105]}
   );
   gpc1_1 gpc509 (
      {stage0_7[158]},
      {stage1_7[62]}
   );
   gpc1_1 gpc510 (
      {stage0_7[159]},
      {stage1_7[63]}
   );
   gpc1_1 gpc511 (
      {stage0_7[160]},
      {stage1_7[64]}
   );
   gpc1_1 gpc512 (
      {stage0_7[161]},
      {stage1_7[65]}
   );
   gpc1_1 gpc513 (
      {stage0_9[152]},
      {stage1_9[67]}
   );
   gpc1_1 gpc514 (
      {stage0_9[153]},
      {stage1_9[68]}
   );
   gpc1_1 gpc515 (
      {stage0_9[154]},
      {stage1_9[69]}
   );
   gpc1_1 gpc516 (
      {stage0_9[155]},
      {stage1_9[70]}
   );
   gpc1_1 gpc517 (
      {stage0_9[156]},
      {stage1_9[71]}
   );
   gpc1_1 gpc518 (
      {stage0_9[157]},
      {stage1_9[72]}
   );
   gpc1_1 gpc519 (
      {stage0_9[158]},
      {stage1_9[73]}
   );
   gpc1_1 gpc520 (
      {stage0_9[159]},
      {stage1_9[74]}
   );
   gpc1_1 gpc521 (
      {stage0_9[160]},
      {stage1_9[75]}
   );
   gpc1_1 gpc522 (
      {stage0_9[161]},
      {stage1_9[76]}
   );
   gpc1_1 gpc523 (
      {stage0_10[141]},
      {stage1_10[72]}
   );
   gpc1_1 gpc524 (
      {stage0_10[142]},
      {stage1_10[73]}
   );
   gpc1_1 gpc525 (
      {stage0_10[143]},
      {stage1_10[74]}
   );
   gpc1_1 gpc526 (
      {stage0_10[144]},
      {stage1_10[75]}
   );
   gpc1_1 gpc527 (
      {stage0_10[145]},
      {stage1_10[76]}
   );
   gpc1_1 gpc528 (
      {stage0_10[146]},
      {stage1_10[77]}
   );
   gpc1_1 gpc529 (
      {stage0_10[147]},
      {stage1_10[78]}
   );
   gpc1_1 gpc530 (
      {stage0_10[148]},
      {stage1_10[79]}
   );
   gpc1_1 gpc531 (
      {stage0_10[149]},
      {stage1_10[80]}
   );
   gpc1_1 gpc532 (
      {stage0_10[150]},
      {stage1_10[81]}
   );
   gpc1_1 gpc533 (
      {stage0_10[151]},
      {stage1_10[82]}
   );
   gpc1_1 gpc534 (
      {stage0_10[152]},
      {stage1_10[83]}
   );
   gpc1_1 gpc535 (
      {stage0_10[153]},
      {stage1_10[84]}
   );
   gpc1_1 gpc536 (
      {stage0_10[154]},
      {stage1_10[85]}
   );
   gpc1_1 gpc537 (
      {stage0_10[155]},
      {stage1_10[86]}
   );
   gpc1_1 gpc538 (
      {stage0_10[156]},
      {stage1_10[87]}
   );
   gpc1_1 gpc539 (
      {stage0_10[157]},
      {stage1_10[88]}
   );
   gpc1_1 gpc540 (
      {stage0_10[158]},
      {stage1_10[89]}
   );
   gpc1_1 gpc541 (
      {stage0_10[159]},
      {stage1_10[90]}
   );
   gpc1_1 gpc542 (
      {stage0_10[160]},
      {stage1_10[91]}
   );
   gpc1_1 gpc543 (
      {stage0_10[161]},
      {stage1_10[92]}
   );
   gpc1_1 gpc544 (
      {stage0_11[155]},
      {stage1_11[60]}
   );
   gpc1_1 gpc545 (
      {stage0_11[156]},
      {stage1_11[61]}
   );
   gpc1_1 gpc546 (
      {stage0_11[157]},
      {stage1_11[62]}
   );
   gpc1_1 gpc547 (
      {stage0_11[158]},
      {stage1_11[63]}
   );
   gpc1_1 gpc548 (
      {stage0_11[159]},
      {stage1_11[64]}
   );
   gpc1_1 gpc549 (
      {stage0_11[160]},
      {stage1_11[65]}
   );
   gpc1_1 gpc550 (
      {stage0_11[161]},
      {stage1_11[66]}
   );
   gpc1_1 gpc551 (
      {stage0_13[144]},
      {stage1_13[68]}
   );
   gpc1_1 gpc552 (
      {stage0_13[145]},
      {stage1_13[69]}
   );
   gpc1_1 gpc553 (
      {stage0_13[146]},
      {stage1_13[70]}
   );
   gpc1_1 gpc554 (
      {stage0_13[147]},
      {stage1_13[71]}
   );
   gpc1_1 gpc555 (
      {stage0_13[148]},
      {stage1_13[72]}
   );
   gpc1_1 gpc556 (
      {stage0_13[149]},
      {stage1_13[73]}
   );
   gpc1_1 gpc557 (
      {stage0_13[150]},
      {stage1_13[74]}
   );
   gpc1_1 gpc558 (
      {stage0_13[151]},
      {stage1_13[75]}
   );
   gpc1_1 gpc559 (
      {stage0_13[152]},
      {stage1_13[76]}
   );
   gpc1_1 gpc560 (
      {stage0_13[153]},
      {stage1_13[77]}
   );
   gpc1_1 gpc561 (
      {stage0_13[154]},
      {stage1_13[78]}
   );
   gpc1_1 gpc562 (
      {stage0_13[155]},
      {stage1_13[79]}
   );
   gpc1_1 gpc563 (
      {stage0_13[156]},
      {stage1_13[80]}
   );
   gpc1_1 gpc564 (
      {stage0_13[157]},
      {stage1_13[81]}
   );
   gpc1_1 gpc565 (
      {stage0_13[158]},
      {stage1_13[82]}
   );
   gpc1_1 gpc566 (
      {stage0_13[159]},
      {stage1_13[83]}
   );
   gpc1_1 gpc567 (
      {stage0_13[160]},
      {stage1_13[84]}
   );
   gpc1_1 gpc568 (
      {stage0_13[161]},
      {stage1_13[85]}
   );
   gpc1_1 gpc569 (
      {stage0_14[161]},
      {stage1_14[68]}
   );
   gpc1_1 gpc570 (
      {stage0_16[111]},
      {stage1_16[56]}
   );
   gpc1_1 gpc571 (
      {stage0_16[112]},
      {stage1_16[57]}
   );
   gpc1_1 gpc572 (
      {stage0_16[113]},
      {stage1_16[58]}
   );
   gpc1_1 gpc573 (
      {stage0_16[114]},
      {stage1_16[59]}
   );
   gpc1_1 gpc574 (
      {stage0_16[115]},
      {stage1_16[60]}
   );
   gpc1_1 gpc575 (
      {stage0_16[116]},
      {stage1_16[61]}
   );
   gpc1_1 gpc576 (
      {stage0_16[117]},
      {stage1_16[62]}
   );
   gpc1_1 gpc577 (
      {stage0_16[118]},
      {stage1_16[63]}
   );
   gpc1_1 gpc578 (
      {stage0_16[119]},
      {stage1_16[64]}
   );
   gpc1_1 gpc579 (
      {stage0_16[120]},
      {stage1_16[65]}
   );
   gpc1_1 gpc580 (
      {stage0_16[121]},
      {stage1_16[66]}
   );
   gpc1_1 gpc581 (
      {stage0_16[122]},
      {stage1_16[67]}
   );
   gpc1_1 gpc582 (
      {stage0_16[123]},
      {stage1_16[68]}
   );
   gpc1_1 gpc583 (
      {stage0_16[124]},
      {stage1_16[69]}
   );
   gpc1_1 gpc584 (
      {stage0_16[125]},
      {stage1_16[70]}
   );
   gpc1_1 gpc585 (
      {stage0_16[126]},
      {stage1_16[71]}
   );
   gpc1_1 gpc586 (
      {stage0_16[127]},
      {stage1_16[72]}
   );
   gpc1_1 gpc587 (
      {stage0_16[128]},
      {stage1_16[73]}
   );
   gpc1_1 gpc588 (
      {stage0_16[129]},
      {stage1_16[74]}
   );
   gpc1_1 gpc589 (
      {stage0_16[130]},
      {stage1_16[75]}
   );
   gpc1_1 gpc590 (
      {stage0_16[131]},
      {stage1_16[76]}
   );
   gpc1_1 gpc591 (
      {stage0_16[132]},
      {stage1_16[77]}
   );
   gpc1_1 gpc592 (
      {stage0_16[133]},
      {stage1_16[78]}
   );
   gpc1_1 gpc593 (
      {stage0_16[134]},
      {stage1_16[79]}
   );
   gpc1_1 gpc594 (
      {stage0_16[135]},
      {stage1_16[80]}
   );
   gpc1_1 gpc595 (
      {stage0_16[136]},
      {stage1_16[81]}
   );
   gpc1_1 gpc596 (
      {stage0_16[137]},
      {stage1_16[82]}
   );
   gpc1_1 gpc597 (
      {stage0_16[138]},
      {stage1_16[83]}
   );
   gpc1_1 gpc598 (
      {stage0_16[139]},
      {stage1_16[84]}
   );
   gpc1_1 gpc599 (
      {stage0_16[140]},
      {stage1_16[85]}
   );
   gpc1_1 gpc600 (
      {stage0_16[141]},
      {stage1_16[86]}
   );
   gpc1_1 gpc601 (
      {stage0_16[142]},
      {stage1_16[87]}
   );
   gpc1_1 gpc602 (
      {stage0_16[143]},
      {stage1_16[88]}
   );
   gpc1_1 gpc603 (
      {stage0_16[144]},
      {stage1_16[89]}
   );
   gpc1_1 gpc604 (
      {stage0_16[145]},
      {stage1_16[90]}
   );
   gpc1_1 gpc605 (
      {stage0_16[146]},
      {stage1_16[91]}
   );
   gpc1_1 gpc606 (
      {stage0_16[147]},
      {stage1_16[92]}
   );
   gpc1_1 gpc607 (
      {stage0_16[148]},
      {stage1_16[93]}
   );
   gpc1_1 gpc608 (
      {stage0_16[149]},
      {stage1_16[94]}
   );
   gpc1_1 gpc609 (
      {stage0_16[150]},
      {stage1_16[95]}
   );
   gpc1_1 gpc610 (
      {stage0_16[151]},
      {stage1_16[96]}
   );
   gpc1_1 gpc611 (
      {stage0_16[152]},
      {stage1_16[97]}
   );
   gpc1_1 gpc612 (
      {stage0_16[153]},
      {stage1_16[98]}
   );
   gpc1_1 gpc613 (
      {stage0_16[154]},
      {stage1_16[99]}
   );
   gpc1_1 gpc614 (
      {stage0_16[155]},
      {stage1_16[100]}
   );
   gpc1_1 gpc615 (
      {stage0_16[156]},
      {stage1_16[101]}
   );
   gpc1_1 gpc616 (
      {stage0_16[157]},
      {stage1_16[102]}
   );
   gpc1_1 gpc617 (
      {stage0_16[158]},
      {stage1_16[103]}
   );
   gpc1_1 gpc618 (
      {stage0_16[159]},
      {stage1_16[104]}
   );
   gpc1_1 gpc619 (
      {stage0_16[160]},
      {stage1_16[105]}
   );
   gpc1_1 gpc620 (
      {stage0_16[161]},
      {stage1_16[106]}
   );
   gpc1_1 gpc621 (
      {stage0_18[142]},
      {stage1_18[62]}
   );
   gpc1_1 gpc622 (
      {stage0_18[143]},
      {stage1_18[63]}
   );
   gpc1_1 gpc623 (
      {stage0_18[144]},
      {stage1_18[64]}
   );
   gpc1_1 gpc624 (
      {stage0_18[145]},
      {stage1_18[65]}
   );
   gpc1_1 gpc625 (
      {stage0_18[146]},
      {stage1_18[66]}
   );
   gpc1_1 gpc626 (
      {stage0_18[147]},
      {stage1_18[67]}
   );
   gpc1_1 gpc627 (
      {stage0_18[148]},
      {stage1_18[68]}
   );
   gpc1_1 gpc628 (
      {stage0_18[149]},
      {stage1_18[69]}
   );
   gpc1_1 gpc629 (
      {stage0_18[150]},
      {stage1_18[70]}
   );
   gpc1_1 gpc630 (
      {stage0_18[151]},
      {stage1_18[71]}
   );
   gpc1_1 gpc631 (
      {stage0_18[152]},
      {stage1_18[72]}
   );
   gpc1_1 gpc632 (
      {stage0_18[153]},
      {stage1_18[73]}
   );
   gpc1_1 gpc633 (
      {stage0_18[154]},
      {stage1_18[74]}
   );
   gpc1_1 gpc634 (
      {stage0_18[155]},
      {stage1_18[75]}
   );
   gpc1_1 gpc635 (
      {stage0_18[156]},
      {stage1_18[76]}
   );
   gpc1_1 gpc636 (
      {stage0_18[157]},
      {stage1_18[77]}
   );
   gpc1_1 gpc637 (
      {stage0_18[158]},
      {stage1_18[78]}
   );
   gpc1_1 gpc638 (
      {stage0_18[159]},
      {stage1_18[79]}
   );
   gpc1_1 gpc639 (
      {stage0_18[160]},
      {stage1_18[80]}
   );
   gpc1_1 gpc640 (
      {stage0_18[161]},
      {stage1_18[81]}
   );
   gpc1_1 gpc641 (
      {stage0_19[154]},
      {stage1_19[59]}
   );
   gpc1_1 gpc642 (
      {stage0_19[155]},
      {stage1_19[60]}
   );
   gpc1_1 gpc643 (
      {stage0_19[156]},
      {stage1_19[61]}
   );
   gpc1_1 gpc644 (
      {stage0_19[157]},
      {stage1_19[62]}
   );
   gpc1_1 gpc645 (
      {stage0_19[158]},
      {stage1_19[63]}
   );
   gpc1_1 gpc646 (
      {stage0_19[159]},
      {stage1_19[64]}
   );
   gpc1_1 gpc647 (
      {stage0_19[160]},
      {stage1_19[65]}
   );
   gpc1_1 gpc648 (
      {stage0_19[161]},
      {stage1_19[66]}
   );
   gpc1_1 gpc649 (
      {stage0_21[160]},
      {stage1_21[78]}
   );
   gpc1_1 gpc650 (
      {stage0_21[161]},
      {stage1_21[79]}
   );
   gpc1_1 gpc651 (
      {stage0_22[138]},
      {stage1_22[58]}
   );
   gpc1_1 gpc652 (
      {stage0_22[139]},
      {stage1_22[59]}
   );
   gpc1_1 gpc653 (
      {stage0_22[140]},
      {stage1_22[60]}
   );
   gpc1_1 gpc654 (
      {stage0_22[141]},
      {stage1_22[61]}
   );
   gpc1_1 gpc655 (
      {stage0_22[142]},
      {stage1_22[62]}
   );
   gpc1_1 gpc656 (
      {stage0_22[143]},
      {stage1_22[63]}
   );
   gpc1_1 gpc657 (
      {stage0_22[144]},
      {stage1_22[64]}
   );
   gpc1_1 gpc658 (
      {stage0_22[145]},
      {stage1_22[65]}
   );
   gpc1_1 gpc659 (
      {stage0_22[146]},
      {stage1_22[66]}
   );
   gpc1_1 gpc660 (
      {stage0_22[147]},
      {stage1_22[67]}
   );
   gpc1_1 gpc661 (
      {stage0_22[148]},
      {stage1_22[68]}
   );
   gpc1_1 gpc662 (
      {stage0_22[149]},
      {stage1_22[69]}
   );
   gpc1_1 gpc663 (
      {stage0_22[150]},
      {stage1_22[70]}
   );
   gpc1_1 gpc664 (
      {stage0_22[151]},
      {stage1_22[71]}
   );
   gpc1_1 gpc665 (
      {stage0_22[152]},
      {stage1_22[72]}
   );
   gpc1_1 gpc666 (
      {stage0_22[153]},
      {stage1_22[73]}
   );
   gpc1_1 gpc667 (
      {stage0_22[154]},
      {stage1_22[74]}
   );
   gpc1_1 gpc668 (
      {stage0_22[155]},
      {stage1_22[75]}
   );
   gpc1_1 gpc669 (
      {stage0_22[156]},
      {stage1_22[76]}
   );
   gpc1_1 gpc670 (
      {stage0_22[157]},
      {stage1_22[77]}
   );
   gpc1_1 gpc671 (
      {stage0_22[158]},
      {stage1_22[78]}
   );
   gpc1_1 gpc672 (
      {stage0_22[159]},
      {stage1_22[79]}
   );
   gpc1_1 gpc673 (
      {stage0_22[160]},
      {stage1_22[80]}
   );
   gpc1_1 gpc674 (
      {stage0_22[161]},
      {stage1_22[81]}
   );
   gpc1_1 gpc675 (
      {stage0_23[122]},
      {stage1_23[51]}
   );
   gpc1_1 gpc676 (
      {stage0_23[123]},
      {stage1_23[52]}
   );
   gpc1_1 gpc677 (
      {stage0_23[124]},
      {stage1_23[53]}
   );
   gpc1_1 gpc678 (
      {stage0_23[125]},
      {stage1_23[54]}
   );
   gpc1_1 gpc679 (
      {stage0_23[126]},
      {stage1_23[55]}
   );
   gpc1_1 gpc680 (
      {stage0_23[127]},
      {stage1_23[56]}
   );
   gpc1_1 gpc681 (
      {stage0_23[128]},
      {stage1_23[57]}
   );
   gpc1_1 gpc682 (
      {stage0_23[129]},
      {stage1_23[58]}
   );
   gpc1_1 gpc683 (
      {stage0_23[130]},
      {stage1_23[59]}
   );
   gpc1_1 gpc684 (
      {stage0_23[131]},
      {stage1_23[60]}
   );
   gpc1_1 gpc685 (
      {stage0_23[132]},
      {stage1_23[61]}
   );
   gpc1_1 gpc686 (
      {stage0_23[133]},
      {stage1_23[62]}
   );
   gpc1_1 gpc687 (
      {stage0_23[134]},
      {stage1_23[63]}
   );
   gpc1_1 gpc688 (
      {stage0_23[135]},
      {stage1_23[64]}
   );
   gpc1_1 gpc689 (
      {stage0_23[136]},
      {stage1_23[65]}
   );
   gpc1_1 gpc690 (
      {stage0_23[137]},
      {stage1_23[66]}
   );
   gpc1_1 gpc691 (
      {stage0_23[138]},
      {stage1_23[67]}
   );
   gpc1_1 gpc692 (
      {stage0_23[139]},
      {stage1_23[68]}
   );
   gpc1_1 gpc693 (
      {stage0_23[140]},
      {stage1_23[69]}
   );
   gpc1_1 gpc694 (
      {stage0_23[141]},
      {stage1_23[70]}
   );
   gpc1_1 gpc695 (
      {stage0_23[142]},
      {stage1_23[71]}
   );
   gpc1_1 gpc696 (
      {stage0_23[143]},
      {stage1_23[72]}
   );
   gpc1_1 gpc697 (
      {stage0_23[144]},
      {stage1_23[73]}
   );
   gpc1_1 gpc698 (
      {stage0_23[145]},
      {stage1_23[74]}
   );
   gpc1_1 gpc699 (
      {stage0_23[146]},
      {stage1_23[75]}
   );
   gpc1_1 gpc700 (
      {stage0_23[147]},
      {stage1_23[76]}
   );
   gpc1_1 gpc701 (
      {stage0_23[148]},
      {stage1_23[77]}
   );
   gpc1_1 gpc702 (
      {stage0_23[149]},
      {stage1_23[78]}
   );
   gpc1_1 gpc703 (
      {stage0_23[150]},
      {stage1_23[79]}
   );
   gpc1_1 gpc704 (
      {stage0_23[151]},
      {stage1_23[80]}
   );
   gpc1_1 gpc705 (
      {stage0_23[152]},
      {stage1_23[81]}
   );
   gpc1_1 gpc706 (
      {stage0_23[153]},
      {stage1_23[82]}
   );
   gpc1_1 gpc707 (
      {stage0_23[154]},
      {stage1_23[83]}
   );
   gpc1_1 gpc708 (
      {stage0_23[155]},
      {stage1_23[84]}
   );
   gpc1_1 gpc709 (
      {stage0_23[156]},
      {stage1_23[85]}
   );
   gpc1_1 gpc710 (
      {stage0_23[157]},
      {stage1_23[86]}
   );
   gpc1_1 gpc711 (
      {stage0_23[158]},
      {stage1_23[87]}
   );
   gpc1_1 gpc712 (
      {stage0_23[159]},
      {stage1_23[88]}
   );
   gpc1_1 gpc713 (
      {stage0_23[160]},
      {stage1_23[89]}
   );
   gpc1_1 gpc714 (
      {stage0_23[161]},
      {stage1_23[90]}
   );
   gpc1_1 gpc715 (
      {stage0_25[158]},
      {stage1_25[74]}
   );
   gpc1_1 gpc716 (
      {stage0_25[159]},
      {stage1_25[75]}
   );
   gpc1_1 gpc717 (
      {stage0_25[160]},
      {stage1_25[76]}
   );
   gpc1_1 gpc718 (
      {stage0_25[161]},
      {stage1_25[77]}
   );
   gpc1_1 gpc719 (
      {stage0_26[160]},
      {stage1_26[53]}
   );
   gpc1_1 gpc720 (
      {stage0_26[161]},
      {stage1_26[54]}
   );
   gpc1_1 gpc721 (
      {stage0_27[155]},
      {stage1_27[60]}
   );
   gpc1_1 gpc722 (
      {stage0_27[156]},
      {stage1_27[61]}
   );
   gpc1_1 gpc723 (
      {stage0_27[157]},
      {stage1_27[62]}
   );
   gpc1_1 gpc724 (
      {stage0_27[158]},
      {stage1_27[63]}
   );
   gpc1_1 gpc725 (
      {stage0_27[159]},
      {stage1_27[64]}
   );
   gpc1_1 gpc726 (
      {stage0_27[160]},
      {stage1_27[65]}
   );
   gpc1_1 gpc727 (
      {stage0_27[161]},
      {stage1_27[66]}
   );
   gpc1_1 gpc728 (
      {stage0_29[159]},
      {stage1_29[72]}
   );
   gpc1_1 gpc729 (
      {stage0_29[160]},
      {stage1_29[73]}
   );
   gpc1_1 gpc730 (
      {stage0_29[161]},
      {stage1_29[74]}
   );
   gpc1_1 gpc731 (
      {stage0_30[151]},
      {stage1_30[52]}
   );
   gpc1_1 gpc732 (
      {stage0_30[152]},
      {stage1_30[53]}
   );
   gpc1_1 gpc733 (
      {stage0_30[153]},
      {stage1_30[54]}
   );
   gpc1_1 gpc734 (
      {stage0_30[154]},
      {stage1_30[55]}
   );
   gpc1_1 gpc735 (
      {stage0_30[155]},
      {stage1_30[56]}
   );
   gpc1_1 gpc736 (
      {stage0_30[156]},
      {stage1_30[57]}
   );
   gpc1_1 gpc737 (
      {stage0_30[157]},
      {stage1_30[58]}
   );
   gpc1_1 gpc738 (
      {stage0_30[158]},
      {stage1_30[59]}
   );
   gpc1_1 gpc739 (
      {stage0_30[159]},
      {stage1_30[60]}
   );
   gpc1_1 gpc740 (
      {stage0_30[160]},
      {stage1_30[61]}
   );
   gpc1_1 gpc741 (
      {stage0_30[161]},
      {stage1_30[62]}
   );
   gpc1_1 gpc742 (
      {stage0_31[116]},
      {stage1_31[52]}
   );
   gpc1_1 gpc743 (
      {stage0_31[117]},
      {stage1_31[53]}
   );
   gpc1_1 gpc744 (
      {stage0_31[118]},
      {stage1_31[54]}
   );
   gpc1_1 gpc745 (
      {stage0_31[119]},
      {stage1_31[55]}
   );
   gpc1_1 gpc746 (
      {stage0_31[120]},
      {stage1_31[56]}
   );
   gpc1_1 gpc747 (
      {stage0_31[121]},
      {stage1_31[57]}
   );
   gpc1_1 gpc748 (
      {stage0_31[122]},
      {stage1_31[58]}
   );
   gpc1_1 gpc749 (
      {stage0_31[123]},
      {stage1_31[59]}
   );
   gpc1_1 gpc750 (
      {stage0_31[124]},
      {stage1_31[60]}
   );
   gpc1_1 gpc751 (
      {stage0_31[125]},
      {stage1_31[61]}
   );
   gpc1_1 gpc752 (
      {stage0_31[126]},
      {stage1_31[62]}
   );
   gpc1_1 gpc753 (
      {stage0_31[127]},
      {stage1_31[63]}
   );
   gpc1_1 gpc754 (
      {stage0_31[128]},
      {stage1_31[64]}
   );
   gpc1_1 gpc755 (
      {stage0_31[129]},
      {stage1_31[65]}
   );
   gpc1_1 gpc756 (
      {stage0_31[130]},
      {stage1_31[66]}
   );
   gpc1_1 gpc757 (
      {stage0_31[131]},
      {stage1_31[67]}
   );
   gpc1_1 gpc758 (
      {stage0_31[132]},
      {stage1_31[68]}
   );
   gpc1_1 gpc759 (
      {stage0_31[133]},
      {stage1_31[69]}
   );
   gpc1_1 gpc760 (
      {stage0_31[134]},
      {stage1_31[70]}
   );
   gpc1_1 gpc761 (
      {stage0_31[135]},
      {stage1_31[71]}
   );
   gpc1_1 gpc762 (
      {stage0_31[136]},
      {stage1_31[72]}
   );
   gpc1_1 gpc763 (
      {stage0_31[137]},
      {stage1_31[73]}
   );
   gpc1_1 gpc764 (
      {stage0_31[138]},
      {stage1_31[74]}
   );
   gpc1_1 gpc765 (
      {stage0_31[139]},
      {stage1_31[75]}
   );
   gpc1_1 gpc766 (
      {stage0_31[140]},
      {stage1_31[76]}
   );
   gpc1_1 gpc767 (
      {stage0_31[141]},
      {stage1_31[77]}
   );
   gpc1_1 gpc768 (
      {stage0_31[142]},
      {stage1_31[78]}
   );
   gpc1_1 gpc769 (
      {stage0_31[143]},
      {stage1_31[79]}
   );
   gpc1_1 gpc770 (
      {stage0_31[144]},
      {stage1_31[80]}
   );
   gpc1_1 gpc771 (
      {stage0_31[145]},
      {stage1_31[81]}
   );
   gpc1_1 gpc772 (
      {stage0_31[146]},
      {stage1_31[82]}
   );
   gpc1_1 gpc773 (
      {stage0_31[147]},
      {stage1_31[83]}
   );
   gpc1_1 gpc774 (
      {stage0_31[148]},
      {stage1_31[84]}
   );
   gpc1_1 gpc775 (
      {stage0_31[149]},
      {stage1_31[85]}
   );
   gpc1_1 gpc776 (
      {stage0_31[150]},
      {stage1_31[86]}
   );
   gpc1_1 gpc777 (
      {stage0_31[151]},
      {stage1_31[87]}
   );
   gpc1_1 gpc778 (
      {stage0_31[152]},
      {stage1_31[88]}
   );
   gpc1_1 gpc779 (
      {stage0_31[153]},
      {stage1_31[89]}
   );
   gpc1_1 gpc780 (
      {stage0_31[154]},
      {stage1_31[90]}
   );
   gpc1_1 gpc781 (
      {stage0_31[155]},
      {stage1_31[91]}
   );
   gpc1_1 gpc782 (
      {stage0_31[156]},
      {stage1_31[92]}
   );
   gpc1_1 gpc783 (
      {stage0_31[157]},
      {stage1_31[93]}
   );
   gpc1_1 gpc784 (
      {stage0_31[158]},
      {stage1_31[94]}
   );
   gpc1_1 gpc785 (
      {stage0_31[159]},
      {stage1_31[95]}
   );
   gpc1_1 gpc786 (
      {stage0_31[160]},
      {stage1_31[96]}
   );
   gpc1_1 gpc787 (
      {stage0_31[161]},
      {stage1_31[97]}
   );
   gpc1163_5 gpc788 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc789 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc790 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc606_5 gpc791 (
      {stage1_0[9], stage1_0[10], stage1_0[11], stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6], stage1_2[7], stage1_2[8]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc615_5 gpc792 (
      {stage1_0[15], stage1_0[16], stage1_0[17], stage1_0[18], stage1_0[19]},
      {stage1_1[18]},
      {stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12], stage1_2[13], stage1_2[14]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc615_5 gpc793 (
      {stage1_0[20], stage1_0[21], stage1_0[22], stage1_0[23], stage1_0[24]},
      {stage1_1[19]},
      {stage1_2[15], stage1_2[16], stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc615_5 gpc794 (
      {stage1_0[25], stage1_0[26], stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_1[20]},
      {stage1_2[21], stage1_2[22], stage1_2[23], stage1_2[24], stage1_2[25], stage1_2[26]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc615_5 gpc795 (
      {stage1_0[30], stage1_0[31], stage1_0[32], stage1_0[33], stage1_0[34]},
      {stage1_1[21]},
      {stage1_2[27], stage1_2[28], stage1_2[29], stage1_2[30], stage1_2[31], stage1_2[32]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc615_5 gpc796 (
      {stage1_0[35], stage1_0[36], stage1_0[37], stage1_0[38], stage1_0[39]},
      {stage1_1[22]},
      {stage1_2[33], stage1_2[34], stage1_2[35], stage1_2[36], stage1_2[37], stage1_2[38]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc615_5 gpc797 (
      {stage1_0[40], stage1_0[41], stage1_0[42], stage1_0[43], stage1_0[44]},
      {stage1_1[23]},
      {stage1_2[39], stage1_2[40], stage1_2[41], stage1_2[42], stage1_2[43], stage1_2[44]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc615_5 gpc798 (
      {stage1_0[45], stage1_0[46], stage1_0[47], stage1_0[48], stage1_0[49]},
      {stage1_1[24]},
      {stage1_2[45], stage1_2[46], stage1_2[47], stage1_2[48], stage1_2[49], stage1_2[50]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc606_5 gpc799 (
      {stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29], stage1_1[30]},
      {stage1_3[3], stage1_3[4], stage1_3[5], stage1_3[6], stage1_3[7], stage1_3[8]},
      {stage2_5[0],stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11]}
   );
   gpc606_5 gpc800 (
      {stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35], stage1_1[36]},
      {stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12], stage1_3[13], stage1_3[14]},
      {stage2_5[1],stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12]}
   );
   gpc606_5 gpc801 (
      {stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41], stage1_1[42]},
      {stage1_3[15], stage1_3[16], stage1_3[17], stage1_3[18], stage1_3[19], stage1_3[20]},
      {stage2_5[2],stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13]}
   );
   gpc606_5 gpc802 (
      {stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47], stage1_1[48]},
      {stage1_3[21], stage1_3[22], stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26]},
      {stage2_5[3],stage2_4[14],stage2_3[14],stage2_2[14],stage2_1[14]}
   );
   gpc606_5 gpc803 (
      {stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53], stage1_1[54]},
      {stage1_3[27], stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31], stage1_3[32]},
      {stage2_5[4],stage2_4[15],stage2_3[15],stage2_2[15],stage2_1[15]}
   );
   gpc615_5 gpc804 (
      {stage1_2[51], stage1_2[52], stage1_2[53], stage1_2[54], stage1_2[55]},
      {stage1_3[33]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[5],stage2_4[16],stage2_3[16],stage2_2[16]}
   );
   gpc615_5 gpc805 (
      {stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37], stage1_3[38]},
      {stage1_4[6]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[1],stage2_5[6],stage2_4[17],stage2_3[17]}
   );
   gpc615_5 gpc806 (
      {stage1_3[39], stage1_3[40], stage1_3[41], stage1_3[42], stage1_3[43]},
      {stage1_4[7]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[2],stage2_5[7],stage2_4[18],stage2_3[18]}
   );
   gpc615_5 gpc807 (
      {stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47], stage1_3[48]},
      {stage1_4[8]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[3],stage2_5[8],stage2_4[19],stage2_3[19]}
   );
   gpc615_5 gpc808 (
      {stage1_3[49], stage1_3[50], stage1_3[51], stage1_3[52], stage1_3[53]},
      {stage1_4[9]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[4],stage2_5[9],stage2_4[20],stage2_3[20]}
   );
   gpc615_5 gpc809 (
      {stage1_3[54], stage1_3[55], stage1_3[56], stage1_3[57], stage1_3[58]},
      {stage1_4[10]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[5],stage2_5[10],stage2_4[21],stage2_3[21]}
   );
   gpc615_5 gpc810 (
      {stage1_3[59], stage1_3[60], stage1_3[61], stage1_3[62], stage1_3[63]},
      {stage1_4[11]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[6],stage2_5[11],stage2_4[22],stage2_3[22]}
   );
   gpc606_5 gpc811 (
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[6],stage2_6[7],stage2_5[12],stage2_4[23]}
   );
   gpc606_5 gpc812 (
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[7],stage2_6[8],stage2_5[13],stage2_4[24]}
   );
   gpc606_5 gpc813 (
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[8],stage2_6[9],stage2_5[14],stage2_4[25]}
   );
   gpc606_5 gpc814 (
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[9],stage2_6[10],stage2_5[15],stage2_4[26]}
   );
   gpc606_5 gpc815 (
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage2_8[4],stage2_7[10],stage2_6[11],stage2_5[16],stage2_4[27]}
   );
   gpc606_5 gpc816 (
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage2_8[5],stage2_7[11],stage2_6[12],stage2_5[17],stage2_4[28]}
   );
   gpc606_5 gpc817 (
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage2_8[6],stage2_7[12],stage2_6[13],stage2_5[18],stage2_4[29]}
   );
   gpc606_5 gpc818 (
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47]},
      {stage2_8[7],stage2_7[13],stage2_6[14],stage2_5[19],stage2_4[30]}
   );
   gpc606_5 gpc819 (
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage1_6[48], stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53]},
      {stage2_8[8],stage2_7[14],stage2_6[15],stage2_5[20],stage2_4[31]}
   );
   gpc606_5 gpc820 (
      {stage1_4[66], stage1_4[67], stage1_4[68], stage1_4[69], stage1_4[70], stage1_4[71]},
      {stage1_6[54], stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59]},
      {stage2_8[9],stage2_7[15],stage2_6[16],stage2_5[21],stage2_4[32]}
   );
   gpc606_5 gpc821 (
      {stage1_4[72], stage1_4[73], stage1_4[74], stage1_4[75], stage1_4[76], stage1_4[77]},
      {stage1_6[60], stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65]},
      {stage2_8[10],stage2_7[16],stage2_6[17],stage2_5[22],stage2_4[33]}
   );
   gpc606_5 gpc822 (
      {stage1_4[78], stage1_4[79], stage1_4[80], stage1_4[81], stage1_4[82], stage1_4[83]},
      {stage1_6[66], stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71]},
      {stage2_8[11],stage2_7[17],stage2_6[18],stage2_5[23],stage2_4[34]}
   );
   gpc606_5 gpc823 (
      {stage1_4[84], stage1_4[85], stage1_4[86], stage1_4[87], stage1_4[88], stage1_4[89]},
      {stage1_6[72], stage1_6[73], stage1_6[74], stage1_6[75], stage1_6[76], stage1_6[77]},
      {stage2_8[12],stage2_7[18],stage2_6[19],stage2_5[24],stage2_4[35]}
   );
   gpc606_5 gpc824 (
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[13],stage2_7[19],stage2_6[20],stage2_5[25]}
   );
   gpc606_5 gpc825 (
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[14],stage2_7[20],stage2_6[21],stage2_5[26]}
   );
   gpc606_5 gpc826 (
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[15],stage2_7[21],stage2_6[22],stage2_5[27]}
   );
   gpc606_5 gpc827 (
      {stage1_6[78], stage1_6[79], stage1_6[80], stage1_6[81], stage1_6[82], stage1_6[83]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[3],stage2_8[16],stage2_7[22],stage2_6[23]}
   );
   gpc606_5 gpc828 (
      {stage1_6[84], stage1_6[85], stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[4],stage2_8[17],stage2_7[23],stage2_6[24]}
   );
   gpc606_5 gpc829 (
      {stage1_6[90], stage1_6[91], stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[5],stage2_8[18],stage2_7[24],stage2_6[25]}
   );
   gpc606_5 gpc830 (
      {stage1_6[96], stage1_6[97], stage1_6[98], stage1_6[99], stage1_6[100], stage1_6[101]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[6],stage2_8[19],stage2_7[25],stage2_6[26]}
   );
   gpc606_5 gpc831 (
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[4],stage2_9[7],stage2_8[20],stage2_7[26]}
   );
   gpc606_5 gpc832 (
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[5],stage2_9[8],stage2_8[21],stage2_7[27]}
   );
   gpc606_5 gpc833 (
      {stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[6],stage2_9[9],stage2_8[22],stage2_7[28]}
   );
   gpc606_5 gpc834 (
      {stage1_7[36], stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[7],stage2_9[10],stage2_8[23],stage2_7[29]}
   );
   gpc606_5 gpc835 (
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[8],stage2_9[11],stage2_8[24],stage2_7[30]}
   );
   gpc606_5 gpc836 (
      {stage1_7[48], stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[9],stage2_9[12],stage2_8[25],stage2_7[31]}
   );
   gpc606_5 gpc837 (
      {stage1_7[54], stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58], stage1_7[59]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[10],stage2_9[13],stage2_8[26],stage2_7[32]}
   );
   gpc606_5 gpc838 (
      {stage1_7[60], stage1_7[61], stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[11],stage2_9[14],stage2_8[27],stage2_7[33]}
   );
   gpc606_5 gpc839 (
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[8],stage2_10[12],stage2_9[15],stage2_8[28]}
   );
   gpc606_5 gpc840 (
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[9],stage2_10[13],stage2_9[16],stage2_8[29]}
   );
   gpc606_5 gpc841 (
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[10],stage2_10[14],stage2_9[17],stage2_8[30]}
   );
   gpc606_5 gpc842 (
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[11],stage2_10[15],stage2_9[18],stage2_8[31]}
   );
   gpc606_5 gpc843 (
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[12],stage2_10[16],stage2_9[19],stage2_8[32]}
   );
   gpc606_5 gpc844 (
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[5],stage2_11[13],stage2_10[17],stage2_9[20]}
   );
   gpc615_5 gpc845 (
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58]},
      {stage1_10[30]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[6],stage2_11[14],stage2_10[18],stage2_9[21]}
   );
   gpc615_5 gpc846 (
      {stage1_9[59], stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63]},
      {stage1_10[31]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[7],stage2_11[15],stage2_10[19],stage2_9[22]}
   );
   gpc615_5 gpc847 (
      {stage1_9[64], stage1_9[65], stage1_9[66], stage1_9[67], stage1_9[68]},
      {stage1_10[32]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[8],stage2_11[16],stage2_10[20],stage2_9[23]}
   );
   gpc606_5 gpc848 (
      {stage1_10[33], stage1_10[34], stage1_10[35], stage1_10[36], stage1_10[37], stage1_10[38]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[4],stage2_12[9],stage2_11[17],stage2_10[21]}
   );
   gpc606_5 gpc849 (
      {stage1_10[39], stage1_10[40], stage1_10[41], stage1_10[42], stage1_10[43], stage1_10[44]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[5],stage2_12[10],stage2_11[18],stage2_10[22]}
   );
   gpc606_5 gpc850 (
      {stage1_10[45], stage1_10[46], stage1_10[47], stage1_10[48], stage1_10[49], stage1_10[50]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[6],stage2_12[11],stage2_11[19],stage2_10[23]}
   );
   gpc606_5 gpc851 (
      {stage1_10[51], stage1_10[52], stage1_10[53], stage1_10[54], stage1_10[55], stage1_10[56]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[7],stage2_12[12],stage2_11[20],stage2_10[24]}
   );
   gpc606_5 gpc852 (
      {stage1_10[57], stage1_10[58], stage1_10[59], stage1_10[60], stage1_10[61], stage1_10[62]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[8],stage2_12[13],stage2_11[21],stage2_10[25]}
   );
   gpc606_5 gpc853 (
      {stage1_10[63], stage1_10[64], stage1_10[65], stage1_10[66], stage1_10[67], stage1_10[68]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[9],stage2_12[14],stage2_11[22],stage2_10[26]}
   );
   gpc606_5 gpc854 (
      {stage1_10[69], stage1_10[70], stage1_10[71], stage1_10[72], stage1_10[73], stage1_10[74]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[10],stage2_12[15],stage2_11[23],stage2_10[27]}
   );
   gpc606_5 gpc855 (
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[7],stage2_13[11],stage2_12[16],stage2_11[24]}
   );
   gpc606_5 gpc856 (
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[8],stage2_13[12],stage2_12[17],stage2_11[25]}
   );
   gpc606_5 gpc857 (
      {stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[9],stage2_13[13],stage2_12[18],stage2_11[26]}
   );
   gpc606_5 gpc858 (
      {stage1_11[42], stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[10],stage2_13[14],stage2_12[19],stage2_11[27]}
   );
   gpc615_5 gpc859 (
      {stage1_11[48], stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52]},
      {stage1_12[42]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[11],stage2_13[15],stage2_12[20],stage2_11[28]}
   );
   gpc615_5 gpc860 (
      {stage1_11[53], stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57]},
      {stage1_12[43]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[12],stage2_13[16],stage2_12[21],stage2_11[29]}
   );
   gpc606_5 gpc861 (
      {stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47], stage1_12[48], stage1_12[49]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[6],stage2_14[13],stage2_13[17],stage2_12[22]}
   );
   gpc606_5 gpc862 (
      {stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53], stage1_12[54], stage1_12[55]},
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage2_16[1],stage2_15[7],stage2_14[14],stage2_13[18],stage2_12[23]}
   );
   gpc1415_5 gpc863 (
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40]},
      {stage1_14[12]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3]},
      {stage1_16[0]},
      {stage2_17[0],stage2_16[2],stage2_15[8],stage2_14[15],stage2_13[19]}
   );
   gpc615_5 gpc864 (
      {stage1_13[41], stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45]},
      {stage1_14[13]},
      {stage1_15[4], stage1_15[5], stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9]},
      {stage2_17[1],stage2_16[3],stage2_15[9],stage2_14[16],stage2_13[20]}
   );
   gpc615_5 gpc865 (
      {stage1_13[46], stage1_13[47], stage1_13[48], stage1_13[49], stage1_13[50]},
      {stage1_14[14]},
      {stage1_15[10], stage1_15[11], stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15]},
      {stage2_17[2],stage2_16[4],stage2_15[10],stage2_14[17],stage2_13[21]}
   );
   gpc615_5 gpc866 (
      {stage1_13[51], stage1_13[52], stage1_13[53], stage1_13[54], stage1_13[55]},
      {stage1_14[15]},
      {stage1_15[16], stage1_15[17], stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21]},
      {stage2_17[3],stage2_16[5],stage2_15[11],stage2_14[18],stage2_13[22]}
   );
   gpc615_5 gpc867 (
      {stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59], stage1_13[60]},
      {stage1_14[16]},
      {stage1_15[22], stage1_15[23], stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27]},
      {stage2_17[4],stage2_16[6],stage2_15[12],stage2_14[19],stage2_13[23]}
   );
   gpc615_5 gpc868 (
      {stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage1_14[17]},
      {stage1_15[28], stage1_15[29], stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33]},
      {stage2_17[5],stage2_16[7],stage2_15[13],stage2_14[20],stage2_13[24]}
   );
   gpc606_5 gpc869 (
      {stage1_14[18], stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23]},
      {stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5], stage1_16[6]},
      {stage2_18[0],stage2_17[6],stage2_16[8],stage2_15[14],stage2_14[21]}
   );
   gpc606_5 gpc870 (
      {stage1_14[24], stage1_14[25], stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29]},
      {stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11], stage1_16[12]},
      {stage2_18[1],stage2_17[7],stage2_16[9],stage2_15[15],stage2_14[22]}
   );
   gpc606_5 gpc871 (
      {stage1_14[30], stage1_14[31], stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35]},
      {stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17], stage1_16[18]},
      {stage2_18[2],stage2_17[8],stage2_16[10],stage2_15[16],stage2_14[23]}
   );
   gpc606_5 gpc872 (
      {stage1_14[36], stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41]},
      {stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23], stage1_16[24]},
      {stage2_18[3],stage2_17[9],stage2_16[11],stage2_15[17],stage2_14[24]}
   );
   gpc606_5 gpc873 (
      {stage1_14[42], stage1_14[43], stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47]},
      {stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29], stage1_16[30]},
      {stage2_18[4],stage2_17[10],stage2_16[12],stage2_15[18],stage2_14[25]}
   );
   gpc606_5 gpc874 (
      {stage1_14[48], stage1_14[49], stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53]},
      {stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35], stage1_16[36]},
      {stage2_18[5],stage2_17[11],stage2_16[13],stage2_15[19],stage2_14[26]}
   );
   gpc606_5 gpc875 (
      {stage1_14[54], stage1_14[55], stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59]},
      {stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41], stage1_16[42]},
      {stage2_18[6],stage2_17[12],stage2_16[14],stage2_15[20],stage2_14[27]}
   );
   gpc1406_5 gpc876 (
      {stage1_15[34], stage1_15[35], stage1_15[36], stage1_15[37], stage1_15[38], stage1_15[39]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3]},
      {stage1_18[0]},
      {stage2_19[0],stage2_18[7],stage2_17[13],stage2_16[15],stage2_15[21]}
   );
   gpc615_5 gpc877 (
      {stage1_15[40], stage1_15[41], stage1_15[42], stage1_15[43], stage1_15[44]},
      {stage1_16[43]},
      {stage1_17[4], stage1_17[5], stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9]},
      {stage2_19[1],stage2_18[8],stage2_17[14],stage2_16[16],stage2_15[22]}
   );
   gpc615_5 gpc878 (
      {stage1_15[45], stage1_15[46], stage1_15[47], stage1_15[48], stage1_15[49]},
      {stage1_16[44]},
      {stage1_17[10], stage1_17[11], stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15]},
      {stage2_19[2],stage2_18[9],stage2_17[15],stage2_16[17],stage2_15[23]}
   );
   gpc615_5 gpc879 (
      {stage1_16[45], stage1_16[46], stage1_16[47], stage1_16[48], stage1_16[49]},
      {stage1_17[16]},
      {stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5], stage1_18[6]},
      {stage2_20[0],stage2_19[3],stage2_18[10],stage2_17[16],stage2_16[18]}
   );
   gpc615_5 gpc880 (
      {stage1_16[50], stage1_16[51], stage1_16[52], stage1_16[53], stage1_16[54]},
      {stage1_17[17]},
      {stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11], stage1_18[12]},
      {stage2_20[1],stage2_19[4],stage2_18[11],stage2_17[17],stage2_16[19]}
   );
   gpc615_5 gpc881 (
      {stage1_16[55], stage1_16[56], stage1_16[57], stage1_16[58], stage1_16[59]},
      {stage1_17[18]},
      {stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17], stage1_18[18]},
      {stage2_20[2],stage2_19[5],stage2_18[12],stage2_17[18],stage2_16[20]}
   );
   gpc615_5 gpc882 (
      {stage1_16[60], stage1_16[61], stage1_16[62], stage1_16[63], stage1_16[64]},
      {stage1_17[19]},
      {stage1_18[19], stage1_18[20], stage1_18[21], stage1_18[22], stage1_18[23], stage1_18[24]},
      {stage2_20[3],stage2_19[6],stage2_18[13],stage2_17[19],stage2_16[21]}
   );
   gpc615_5 gpc883 (
      {stage1_16[65], stage1_16[66], stage1_16[67], stage1_16[68], stage1_16[69]},
      {stage1_17[20]},
      {stage1_18[25], stage1_18[26], stage1_18[27], stage1_18[28], stage1_18[29], stage1_18[30]},
      {stage2_20[4],stage2_19[7],stage2_18[14],stage2_17[20],stage2_16[22]}
   );
   gpc615_5 gpc884 (
      {stage1_16[70], stage1_16[71], stage1_16[72], stage1_16[73], stage1_16[74]},
      {stage1_17[21]},
      {stage1_18[31], stage1_18[32], stage1_18[33], stage1_18[34], stage1_18[35], stage1_18[36]},
      {stage2_20[5],stage2_19[8],stage2_18[15],stage2_17[21],stage2_16[23]}
   );
   gpc615_5 gpc885 (
      {stage1_16[75], stage1_16[76], stage1_16[77], stage1_16[78], stage1_16[79]},
      {stage1_17[22]},
      {stage1_18[37], stage1_18[38], stage1_18[39], stage1_18[40], stage1_18[41], stage1_18[42]},
      {stage2_20[6],stage2_19[9],stage2_18[16],stage2_17[22],stage2_16[24]}
   );
   gpc615_5 gpc886 (
      {stage1_16[80], stage1_16[81], stage1_16[82], stage1_16[83], stage1_16[84]},
      {stage1_17[23]},
      {stage1_18[43], stage1_18[44], stage1_18[45], stage1_18[46], stage1_18[47], stage1_18[48]},
      {stage2_20[7],stage2_19[10],stage2_18[17],stage2_17[23],stage2_16[25]}
   );
   gpc615_5 gpc887 (
      {stage1_16[85], stage1_16[86], stage1_16[87], stage1_16[88], stage1_16[89]},
      {stage1_17[24]},
      {stage1_18[49], stage1_18[50], stage1_18[51], stage1_18[52], stage1_18[53], stage1_18[54]},
      {stage2_20[8],stage2_19[11],stage2_18[18],stage2_17[24],stage2_16[26]}
   );
   gpc606_5 gpc888 (
      {stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29], stage1_17[30]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[9],stage2_19[12],stage2_18[19],stage2_17[25]}
   );
   gpc606_5 gpc889 (
      {stage1_17[31], stage1_17[32], stage1_17[33], stage1_17[34], stage1_17[35], stage1_17[36]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[10],stage2_19[13],stage2_18[20],stage2_17[26]}
   );
   gpc606_5 gpc890 (
      {stage1_17[37], stage1_17[38], stage1_17[39], stage1_17[40], stage1_17[41], stage1_17[42]},
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17]},
      {stage2_21[2],stage2_20[11],stage2_19[14],stage2_18[21],stage2_17[27]}
   );
   gpc615_5 gpc891 (
      {stage1_17[43], stage1_17[44], stage1_17[45], stage1_17[46], stage1_17[47]},
      {stage1_18[55]},
      {stage1_19[18], stage1_19[19], stage1_19[20], stage1_19[21], stage1_19[22], stage1_19[23]},
      {stage2_21[3],stage2_20[12],stage2_19[15],stage2_18[22],stage2_17[28]}
   );
   gpc615_5 gpc892 (
      {stage1_17[48], stage1_17[49], stage1_17[50], stage1_17[51], stage1_17[52]},
      {stage1_18[56]},
      {stage1_19[24], stage1_19[25], stage1_19[26], stage1_19[27], stage1_19[28], stage1_19[29]},
      {stage2_21[4],stage2_20[13],stage2_19[16],stage2_18[23],stage2_17[29]}
   );
   gpc615_5 gpc893 (
      {stage1_17[53], stage1_17[54], stage1_17[55], stage1_17[56], stage1_17[57]},
      {stage1_18[57]},
      {stage1_19[30], stage1_19[31], stage1_19[32], stage1_19[33], stage1_19[34], stage1_19[35]},
      {stage2_21[5],stage2_20[14],stage2_19[17],stage2_18[24],stage2_17[30]}
   );
   gpc606_5 gpc894 (
      {stage1_18[58], stage1_18[59], stage1_18[60], stage1_18[61], stage1_18[62], stage1_18[63]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[6],stage2_20[15],stage2_19[18],stage2_18[25]}
   );
   gpc606_5 gpc895 (
      {stage1_18[64], stage1_18[65], stage1_18[66], stage1_18[67], stage1_18[68], stage1_18[69]},
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage2_22[1],stage2_21[7],stage2_20[16],stage2_19[19],stage2_18[26]}
   );
   gpc606_5 gpc896 (
      {stage1_18[70], stage1_18[71], stage1_18[72], stage1_18[73], stage1_18[74], stage1_18[75]},
      {stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15], stage1_20[16], stage1_20[17]},
      {stage2_22[2],stage2_21[8],stage2_20[17],stage2_19[20],stage2_18[27]}
   );
   gpc606_5 gpc897 (
      {stage1_18[76], stage1_18[77], stage1_18[78], stage1_18[79], stage1_18[80], stage1_18[81]},
      {stage1_20[18], stage1_20[19], stage1_20[20], stage1_20[21], stage1_20[22], stage1_20[23]},
      {stage2_22[3],stage2_21[9],stage2_20[18],stage2_19[21],stage2_18[28]}
   );
   gpc606_5 gpc898 (
      {stage1_19[36], stage1_19[37], stage1_19[38], stage1_19[39], stage1_19[40], stage1_19[41]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[4],stage2_21[10],stage2_20[19],stage2_19[22]}
   );
   gpc606_5 gpc899 (
      {stage1_19[42], stage1_19[43], stage1_19[44], stage1_19[45], stage1_19[46], stage1_19[47]},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[5],stage2_21[11],stage2_20[20],stage2_19[23]}
   );
   gpc606_5 gpc900 (
      {stage1_19[48], stage1_19[49], stage1_19[50], stage1_19[51], stage1_19[52], stage1_19[53]},
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage2_23[2],stage2_22[6],stage2_21[12],stage2_20[21],stage2_19[24]}
   );
   gpc606_5 gpc901 (
      {stage1_19[54], stage1_19[55], stage1_19[56], stage1_19[57], stage1_19[58], stage1_19[59]},
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage2_23[3],stage2_22[7],stage2_21[13],stage2_20[22],stage2_19[25]}
   );
   gpc606_5 gpc902 (
      {stage1_19[60], stage1_19[61], stage1_19[62], stage1_19[63], stage1_19[64], stage1_19[65]},
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage2_23[4],stage2_22[8],stage2_21[14],stage2_20[23],stage2_19[26]}
   );
   gpc606_5 gpc903 (
      {stage1_20[24], stage1_20[25], stage1_20[26], stage1_20[27], stage1_20[28], stage1_20[29]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[5],stage2_22[9],stage2_21[15],stage2_20[24]}
   );
   gpc606_5 gpc904 (
      {stage1_20[30], stage1_20[31], stage1_20[32], stage1_20[33], stage1_20[34], stage1_20[35]},
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage2_24[1],stage2_23[6],stage2_22[10],stage2_21[16],stage2_20[25]}
   );
   gpc606_5 gpc905 (
      {stage1_20[36], stage1_20[37], stage1_20[38], stage1_20[39], stage1_20[40], stage1_20[41]},
      {stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage2_24[2],stage2_23[7],stage2_22[11],stage2_21[17],stage2_20[26]}
   );
   gpc615_5 gpc906 (
      {stage1_20[42], stage1_20[43], stage1_20[44], stage1_20[45], stage1_20[46]},
      {stage1_21[30]},
      {stage1_22[18], stage1_22[19], stage1_22[20], stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage2_24[3],stage2_23[8],stage2_22[12],stage2_21[18],stage2_20[27]}
   );
   gpc615_5 gpc907 (
      {stage1_20[47], stage1_20[48], stage1_20[49], stage1_20[50], stage1_20[51]},
      {stage1_21[31]},
      {stage1_22[24], stage1_22[25], stage1_22[26], stage1_22[27], stage1_22[28], stage1_22[29]},
      {stage2_24[4],stage2_23[9],stage2_22[13],stage2_21[19],stage2_20[28]}
   );
   gpc606_5 gpc908 (
      {stage1_21[32], stage1_21[33], stage1_21[34], stage1_21[35], stage1_21[36], stage1_21[37]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[5],stage2_23[10],stage2_22[14],stage2_21[20]}
   );
   gpc606_5 gpc909 (
      {stage1_21[38], stage1_21[39], stage1_21[40], stage1_21[41], stage1_21[42], stage1_21[43]},
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage2_25[1],stage2_24[6],stage2_23[11],stage2_22[15],stage2_21[21]}
   );
   gpc606_5 gpc910 (
      {stage1_21[44], stage1_21[45], stage1_21[46], stage1_21[47], stage1_21[48], stage1_21[49]},
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage2_25[2],stage2_24[7],stage2_23[12],stage2_22[16],stage2_21[22]}
   );
   gpc606_5 gpc911 (
      {stage1_21[50], stage1_21[51], stage1_21[52], stage1_21[53], stage1_21[54], stage1_21[55]},
      {stage1_23[18], stage1_23[19], stage1_23[20], stage1_23[21], stage1_23[22], stage1_23[23]},
      {stage2_25[3],stage2_24[8],stage2_23[13],stage2_22[17],stage2_21[23]}
   );
   gpc606_5 gpc912 (
      {stage1_21[56], stage1_21[57], stage1_21[58], stage1_21[59], stage1_21[60], stage1_21[61]},
      {stage1_23[24], stage1_23[25], stage1_23[26], stage1_23[27], stage1_23[28], stage1_23[29]},
      {stage2_25[4],stage2_24[9],stage2_23[14],stage2_22[18],stage2_21[24]}
   );
   gpc606_5 gpc913 (
      {stage1_21[62], stage1_21[63], stage1_21[64], stage1_21[65], stage1_21[66], stage1_21[67]},
      {stage1_23[30], stage1_23[31], stage1_23[32], stage1_23[33], stage1_23[34], stage1_23[35]},
      {stage2_25[5],stage2_24[10],stage2_23[15],stage2_22[19],stage2_21[25]}
   );
   gpc606_5 gpc914 (
      {stage1_21[68], stage1_21[69], stage1_21[70], stage1_21[71], stage1_21[72], stage1_21[73]},
      {stage1_23[36], stage1_23[37], stage1_23[38], stage1_23[39], stage1_23[40], stage1_23[41]},
      {stage2_25[6],stage2_24[11],stage2_23[16],stage2_22[20],stage2_21[26]}
   );
   gpc606_5 gpc915 (
      {stage1_21[74], stage1_21[75], stage1_21[76], stage1_21[77], stage1_21[78], stage1_21[79]},
      {stage1_23[42], stage1_23[43], stage1_23[44], stage1_23[45], stage1_23[46], stage1_23[47]},
      {stage2_25[7],stage2_24[12],stage2_23[17],stage2_22[21],stage2_21[27]}
   );
   gpc606_5 gpc916 (
      {stage1_22[30], stage1_22[31], stage1_22[32], stage1_22[33], stage1_22[34], stage1_22[35]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5]},
      {stage2_26[0],stage2_25[8],stage2_24[13],stage2_23[18],stage2_22[22]}
   );
   gpc606_5 gpc917 (
      {stage1_22[36], stage1_22[37], stage1_22[38], stage1_22[39], stage1_22[40], stage1_22[41]},
      {stage1_24[6], stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11]},
      {stage2_26[1],stage2_25[9],stage2_24[14],stage2_23[19],stage2_22[23]}
   );
   gpc606_5 gpc918 (
      {stage1_22[42], stage1_22[43], stage1_22[44], stage1_22[45], stage1_22[46], stage1_22[47]},
      {stage1_24[12], stage1_24[13], stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17]},
      {stage2_26[2],stage2_25[10],stage2_24[15],stage2_23[20],stage2_22[24]}
   );
   gpc606_5 gpc919 (
      {stage1_22[48], stage1_22[49], stage1_22[50], stage1_22[51], stage1_22[52], stage1_22[53]},
      {stage1_24[18], stage1_24[19], stage1_24[20], stage1_24[21], stage1_24[22], stage1_24[23]},
      {stage2_26[3],stage2_25[11],stage2_24[16],stage2_23[21],stage2_22[25]}
   );
   gpc606_5 gpc920 (
      {stage1_22[54], stage1_22[55], stage1_22[56], stage1_22[57], stage1_22[58], stage1_22[59]},
      {stage1_24[24], stage1_24[25], stage1_24[26], stage1_24[27], stage1_24[28], stage1_24[29]},
      {stage2_26[4],stage2_25[12],stage2_24[17],stage2_23[22],stage2_22[26]}
   );
   gpc606_5 gpc921 (
      {stage1_22[60], stage1_22[61], stage1_22[62], stage1_22[63], stage1_22[64], stage1_22[65]},
      {stage1_24[30], stage1_24[31], stage1_24[32], stage1_24[33], stage1_24[34], stage1_24[35]},
      {stage2_26[5],stage2_25[13],stage2_24[18],stage2_23[23],stage2_22[27]}
   );
   gpc606_5 gpc922 (
      {stage1_22[66], stage1_22[67], stage1_22[68], stage1_22[69], stage1_22[70], stage1_22[71]},
      {stage1_24[36], stage1_24[37], stage1_24[38], stage1_24[39], stage1_24[40], stage1_24[41]},
      {stage2_26[6],stage2_25[14],stage2_24[19],stage2_23[24],stage2_22[28]}
   );
   gpc606_5 gpc923 (
      {stage1_22[72], stage1_22[73], stage1_22[74], stage1_22[75], stage1_22[76], stage1_22[77]},
      {stage1_24[42], stage1_24[43], stage1_24[44], stage1_24[45], stage1_24[46], stage1_24[47]},
      {stage2_26[7],stage2_25[15],stage2_24[20],stage2_23[25],stage2_22[29]}
   );
   gpc606_5 gpc924 (
      {stage1_23[48], stage1_23[49], stage1_23[50], stage1_23[51], stage1_23[52], stage1_23[53]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[8],stage2_25[16],stage2_24[21],stage2_23[26]}
   );
   gpc606_5 gpc925 (
      {stage1_23[54], stage1_23[55], stage1_23[56], stage1_23[57], stage1_23[58], stage1_23[59]},
      {stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11]},
      {stage2_27[1],stage2_26[9],stage2_25[17],stage2_24[22],stage2_23[27]}
   );
   gpc606_5 gpc926 (
      {stage1_23[60], stage1_23[61], stage1_23[62], stage1_23[63], stage1_23[64], stage1_23[65]},
      {stage1_25[12], stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {stage2_27[2],stage2_26[10],stage2_25[18],stage2_24[23],stage2_23[28]}
   );
   gpc606_5 gpc927 (
      {stage1_23[66], stage1_23[67], stage1_23[68], stage1_23[69], stage1_23[70], stage1_23[71]},
      {stage1_25[18], stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23]},
      {stage2_27[3],stage2_26[11],stage2_25[19],stage2_24[24],stage2_23[29]}
   );
   gpc606_5 gpc928 (
      {stage1_23[72], stage1_23[73], stage1_23[74], stage1_23[75], stage1_23[76], stage1_23[77]},
      {stage1_25[24], stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29]},
      {stage2_27[4],stage2_26[12],stage2_25[20],stage2_24[25],stage2_23[30]}
   );
   gpc606_5 gpc929 (
      {stage1_24[48], stage1_24[49], stage1_24[50], stage1_24[51], stage1_24[52], stage1_24[53]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[5],stage2_26[13],stage2_25[21],stage2_24[26]}
   );
   gpc606_5 gpc930 (
      {stage1_24[54], stage1_24[55], stage1_24[56], stage1_24[57], stage1_24[58], stage1_24[59]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[6],stage2_26[14],stage2_25[22],stage2_24[27]}
   );
   gpc606_5 gpc931 (
      {stage1_25[30], stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[2],stage2_27[7],stage2_26[15],stage2_25[23]}
   );
   gpc606_5 gpc932 (
      {stage1_25[36], stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41]},
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage2_29[1],stage2_28[3],stage2_27[8],stage2_26[16],stage2_25[24]}
   );
   gpc606_5 gpc933 (
      {stage1_25[42], stage1_25[43], stage1_25[44], stage1_25[45], stage1_25[46], stage1_25[47]},
      {stage1_27[12], stage1_27[13], stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17]},
      {stage2_29[2],stage2_28[4],stage2_27[9],stage2_26[17],stage2_25[25]}
   );
   gpc606_5 gpc934 (
      {stage1_25[48], stage1_25[49], stage1_25[50], stage1_25[51], stage1_25[52], stage1_25[53]},
      {stage1_27[18], stage1_27[19], stage1_27[20], stage1_27[21], stage1_27[22], stage1_27[23]},
      {stage2_29[3],stage2_28[5],stage2_27[10],stage2_26[18],stage2_25[26]}
   );
   gpc606_5 gpc935 (
      {stage1_25[54], stage1_25[55], stage1_25[56], stage1_25[57], stage1_25[58], stage1_25[59]},
      {stage1_27[24], stage1_27[25], stage1_27[26], stage1_27[27], stage1_27[28], stage1_27[29]},
      {stage2_29[4],stage2_28[6],stage2_27[11],stage2_26[19],stage2_25[27]}
   );
   gpc606_5 gpc936 (
      {stage1_25[60], stage1_25[61], stage1_25[62], stage1_25[63], stage1_25[64], stage1_25[65]},
      {stage1_27[30], stage1_27[31], stage1_27[32], stage1_27[33], stage1_27[34], stage1_27[35]},
      {stage2_29[5],stage2_28[7],stage2_27[12],stage2_26[20],stage2_25[28]}
   );
   gpc606_5 gpc937 (
      {stage1_25[66], stage1_25[67], stage1_25[68], stage1_25[69], stage1_25[70], stage1_25[71]},
      {stage1_27[36], stage1_27[37], stage1_27[38], stage1_27[39], stage1_27[40], stage1_27[41]},
      {stage2_29[6],stage2_28[8],stage2_27[13],stage2_26[21],stage2_25[29]}
   );
   gpc606_5 gpc938 (
      {stage1_25[72], stage1_25[73], stage1_25[74], stage1_25[75], stage1_25[76], stage1_25[77]},
      {stage1_27[42], stage1_27[43], stage1_27[44], stage1_27[45], stage1_27[46], stage1_27[47]},
      {stage2_29[7],stage2_28[9],stage2_27[14],stage2_26[22],stage2_25[30]}
   );
   gpc606_5 gpc939 (
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[8],stage2_28[10],stage2_27[15],stage2_26[23]}
   );
   gpc606_5 gpc940 (
      {stage1_26[18], stage1_26[19], stage1_26[20], stage1_26[21], stage1_26[22], stage1_26[23]},
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11]},
      {stage2_30[1],stage2_29[9],stage2_28[11],stage2_27[16],stage2_26[24]}
   );
   gpc606_5 gpc941 (
      {stage1_26[24], stage1_26[25], stage1_26[26], stage1_26[27], stage1_26[28], stage1_26[29]},
      {stage1_28[12], stage1_28[13], stage1_28[14], stage1_28[15], stage1_28[16], stage1_28[17]},
      {stage2_30[2],stage2_29[10],stage2_28[12],stage2_27[17],stage2_26[25]}
   );
   gpc606_5 gpc942 (
      {stage1_26[30], stage1_26[31], stage1_26[32], stage1_26[33], stage1_26[34], stage1_26[35]},
      {stage1_28[18], stage1_28[19], stage1_28[20], stage1_28[21], stage1_28[22], stage1_28[23]},
      {stage2_30[3],stage2_29[11],stage2_28[13],stage2_27[18],stage2_26[26]}
   );
   gpc606_5 gpc943 (
      {stage1_26[36], stage1_26[37], stage1_26[38], stage1_26[39], stage1_26[40], stage1_26[41]},
      {stage1_28[24], stage1_28[25], stage1_28[26], stage1_28[27], stage1_28[28], stage1_28[29]},
      {stage2_30[4],stage2_29[12],stage2_28[14],stage2_27[19],stage2_26[27]}
   );
   gpc606_5 gpc944 (
      {stage1_26[42], stage1_26[43], stage1_26[44], stage1_26[45], stage1_26[46], stage1_26[47]},
      {stage1_28[30], stage1_28[31], stage1_28[32], stage1_28[33], stage1_28[34], stage1_28[35]},
      {stage2_30[5],stage2_29[13],stage2_28[15],stage2_27[20],stage2_26[28]}
   );
   gpc606_5 gpc945 (
      {stage1_26[48], stage1_26[49], stage1_26[50], stage1_26[51], stage1_26[52], stage1_26[53]},
      {stage1_28[36], stage1_28[37], stage1_28[38], stage1_28[39], stage1_28[40], stage1_28[41]},
      {stage2_30[6],stage2_29[14],stage2_28[16],stage2_27[21],stage2_26[29]}
   );
   gpc615_5 gpc946 (
      {stage1_27[48], stage1_27[49], stage1_27[50], stage1_27[51], stage1_27[52]},
      {stage1_28[42]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[7],stage2_29[15],stage2_28[17],stage2_27[22]}
   );
   gpc615_5 gpc947 (
      {stage1_27[53], stage1_27[54], stage1_27[55], stage1_27[56], stage1_27[57]},
      {stage1_28[43]},
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage2_31[1],stage2_30[8],stage2_29[16],stage2_28[18],stage2_27[23]}
   );
   gpc606_5 gpc948 (
      {stage1_28[44], stage1_28[45], stage1_28[46], stage1_28[47], stage1_28[48], stage1_28[49]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[2],stage2_30[9],stage2_29[17],stage2_28[19]}
   );
   gpc606_5 gpc949 (
      {stage1_28[50], stage1_28[51], stage1_28[52], stage1_28[53], stage1_28[54], stage1_28[55]},
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage2_32[1],stage2_31[3],stage2_30[10],stage2_29[18],stage2_28[20]}
   );
   gpc606_5 gpc950 (
      {stage1_28[56], stage1_28[57], stage1_28[58], stage1_28[59], stage1_28[60], stage1_28[61]},
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage2_32[2],stage2_31[4],stage2_30[11],stage2_29[19],stage2_28[21]}
   );
   gpc615_5 gpc951 (
      {stage1_28[62], stage1_28[63], stage1_28[64], stage1_28[65], stage1_28[66]},
      {stage1_29[12]},
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22], stage1_30[23]},
      {stage2_32[3],stage2_31[5],stage2_30[12],stage2_29[20],stage2_28[22]}
   );
   gpc615_5 gpc952 (
      {stage1_28[67], stage1_28[68], stage1_28[69], stage1_28[70], stage1_28[71]},
      {stage1_29[13]},
      {stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27], stage1_30[28], stage1_30[29]},
      {stage2_32[4],stage2_31[6],stage2_30[13],stage2_29[21],stage2_28[23]}
   );
   gpc606_5 gpc953 (
      {stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17], stage1_29[18], stage1_29[19]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[5],stage2_31[7],stage2_30[14],stage2_29[22]}
   );
   gpc606_5 gpc954 (
      {stage1_29[20], stage1_29[21], stage1_29[22], stage1_29[23], stage1_29[24], stage1_29[25]},
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10], stage1_31[11]},
      {stage2_33[1],stage2_32[6],stage2_31[8],stage2_30[15],stage2_29[23]}
   );
   gpc606_5 gpc955 (
      {stage1_29[26], stage1_29[27], stage1_29[28], stage1_29[29], stage1_29[30], stage1_29[31]},
      {stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15], stage1_31[16], stage1_31[17]},
      {stage2_33[2],stage2_32[7],stage2_31[9],stage2_30[16],stage2_29[24]}
   );
   gpc606_5 gpc956 (
      {stage1_29[32], stage1_29[33], stage1_29[34], stage1_29[35], stage1_29[36], stage1_29[37]},
      {stage1_31[18], stage1_31[19], stage1_31[20], stage1_31[21], stage1_31[22], stage1_31[23]},
      {stage2_33[3],stage2_32[8],stage2_31[10],stage2_30[17],stage2_29[25]}
   );
   gpc606_5 gpc957 (
      {stage1_29[38], stage1_29[39], stage1_29[40], stage1_29[41], stage1_29[42], stage1_29[43]},
      {stage1_31[24], stage1_31[25], stage1_31[26], stage1_31[27], stage1_31[28], stage1_31[29]},
      {stage2_33[4],stage2_32[9],stage2_31[11],stage2_30[18],stage2_29[26]}
   );
   gpc606_5 gpc958 (
      {stage1_29[44], stage1_29[45], stage1_29[46], stage1_29[47], stage1_29[48], stage1_29[49]},
      {stage1_31[30], stage1_31[31], stage1_31[32], stage1_31[33], stage1_31[34], stage1_31[35]},
      {stage2_33[5],stage2_32[10],stage2_31[12],stage2_30[19],stage2_29[27]}
   );
   gpc615_5 gpc959 (
      {stage1_29[50], stage1_29[51], stage1_29[52], stage1_29[53], stage1_29[54]},
      {stage1_30[30]},
      {stage1_31[36], stage1_31[37], stage1_31[38], stage1_31[39], stage1_31[40], stage1_31[41]},
      {stage2_33[6],stage2_32[11],stage2_31[13],stage2_30[20],stage2_29[28]}
   );
   gpc615_5 gpc960 (
      {stage1_29[55], stage1_29[56], stage1_29[57], stage1_29[58], stage1_29[59]},
      {stage1_30[31]},
      {stage1_31[42], stage1_31[43], stage1_31[44], stage1_31[45], stage1_31[46], stage1_31[47]},
      {stage2_33[7],stage2_32[12],stage2_31[14],stage2_30[21],stage2_29[29]}
   );
   gpc615_5 gpc961 (
      {stage1_29[60], stage1_29[61], stage1_29[62], stage1_29[63], stage1_29[64]},
      {stage1_30[32]},
      {stage1_31[48], stage1_31[49], stage1_31[50], stage1_31[51], stage1_31[52], stage1_31[53]},
      {stage2_33[8],stage2_32[13],stage2_31[15],stage2_30[22],stage2_29[30]}
   );
   gpc615_5 gpc962 (
      {stage1_29[65], stage1_29[66], stage1_29[67], stage1_29[68], stage1_29[69]},
      {stage1_30[33]},
      {stage1_31[54], stage1_31[55], stage1_31[56], stage1_31[57], stage1_31[58], stage1_31[59]},
      {stage2_33[9],stage2_32[14],stage2_31[16],stage2_30[23],stage2_29[31]}
   );
   gpc615_5 gpc963 (
      {stage1_29[70], stage1_29[71], stage1_29[72], stage1_29[73], stage1_29[74]},
      {stage1_30[34]},
      {stage1_31[60], stage1_31[61], stage1_31[62], stage1_31[63], stage1_31[64], stage1_31[65]},
      {stage2_33[10],stage2_32[15],stage2_31[17],stage2_30[24],stage2_29[32]}
   );
   gpc615_5 gpc964 (
      {stage1_30[35], stage1_30[36], stage1_30[37], stage1_30[38], stage1_30[39]},
      {stage1_31[66]},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[11],stage2_32[16],stage2_31[18],stage2_30[25]}
   );
   gpc615_5 gpc965 (
      {stage1_30[40], stage1_30[41], stage1_30[42], stage1_30[43], stage1_30[44]},
      {stage1_31[67]},
      {stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11]},
      {stage2_34[1],stage2_33[12],stage2_32[17],stage2_31[19],stage2_30[26]}
   );
   gpc615_5 gpc966 (
      {stage1_30[45], stage1_30[46], stage1_30[47], stage1_30[48], stage1_30[49]},
      {stage1_31[68]},
      {stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16], stage1_32[17]},
      {stage2_34[2],stage2_33[13],stage2_32[18],stage2_31[20],stage2_30[27]}
   );
   gpc615_5 gpc967 (
      {stage1_30[50], stage1_30[51], stage1_30[52], stage1_30[53], stage1_30[54]},
      {stage1_31[69]},
      {stage1_32[18], stage1_32[19], stage1_32[20], stage1_32[21], stage1_32[22], stage1_32[23]},
      {stage2_34[3],stage2_33[14],stage2_32[19],stage2_31[21],stage2_30[28]}
   );
   gpc135_4 gpc968 (
      {stage1_31[70], stage1_31[71], stage1_31[72], stage1_31[73], stage1_31[74]},
      {stage1_32[24], stage1_32[25], stage1_32[26]},
      {stage1_33[0]},
      {stage2_34[4],stage2_33[15],stage2_32[20],stage2_31[22]}
   );
   gpc606_5 gpc969 (
      {stage1_31[75], stage1_31[76], stage1_31[77], stage1_31[78], stage1_31[79], stage1_31[80]},
      {stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5], stage1_33[6]},
      {stage2_35[0],stage2_34[5],stage2_33[16],stage2_32[21],stage2_31[23]}
   );
   gpc606_5 gpc970 (
      {stage1_31[81], stage1_31[82], stage1_31[83], stage1_31[84], stage1_31[85], stage1_31[86]},
      {stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11], stage1_33[12]},
      {stage2_35[1],stage2_34[6],stage2_33[17],stage2_32[22],stage2_31[24]}
   );
   gpc1_1 gpc971 (
      {stage1_1[55]},
      {stage2_1[16]}
   );
   gpc1_1 gpc972 (
      {stage1_3[64]},
      {stage2_3[23]}
   );
   gpc1_1 gpc973 (
      {stage1_3[65]},
      {stage2_3[24]}
   );
   gpc1_1 gpc974 (
      {stage1_3[66]},
      {stage2_3[25]}
   );
   gpc1_1 gpc975 (
      {stage1_3[67]},
      {stage2_3[26]}
   );
   gpc1_1 gpc976 (
      {stage1_3[68]},
      {stage2_3[27]}
   );
   gpc1_1 gpc977 (
      {stage1_3[69]},
      {stage2_3[28]}
   );
   gpc1_1 gpc978 (
      {stage1_3[70]},
      {stage2_3[29]}
   );
   gpc1_1 gpc979 (
      {stage1_3[71]},
      {stage2_3[30]}
   );
   gpc1_1 gpc980 (
      {stage1_3[72]},
      {stage2_3[31]}
   );
   gpc1_1 gpc981 (
      {stage1_3[73]},
      {stage2_3[32]}
   );
   gpc1_1 gpc982 (
      {stage1_3[74]},
      {stage2_3[33]}
   );
   gpc1_1 gpc983 (
      {stage1_3[75]},
      {stage2_3[34]}
   );
   gpc1_1 gpc984 (
      {stage1_4[90]},
      {stage2_4[36]}
   );
   gpc1_1 gpc985 (
      {stage1_4[91]},
      {stage2_4[37]}
   );
   gpc1_1 gpc986 (
      {stage1_4[92]},
      {stage2_4[38]}
   );
   gpc1_1 gpc987 (
      {stage1_4[93]},
      {stage2_4[39]}
   );
   gpc1_1 gpc988 (
      {stage1_4[94]},
      {stage2_4[40]}
   );
   gpc1_1 gpc989 (
      {stage1_6[102]},
      {stage2_6[27]}
   );
   gpc1_1 gpc990 (
      {stage1_6[103]},
      {stage2_6[28]}
   );
   gpc1_1 gpc991 (
      {stage1_6[104]},
      {stage2_6[29]}
   );
   gpc1_1 gpc992 (
      {stage1_6[105]},
      {stage2_6[30]}
   );
   gpc1_1 gpc993 (
      {stage1_9[69]},
      {stage2_9[24]}
   );
   gpc1_1 gpc994 (
      {stage1_9[70]},
      {stage2_9[25]}
   );
   gpc1_1 gpc995 (
      {stage1_9[71]},
      {stage2_9[26]}
   );
   gpc1_1 gpc996 (
      {stage1_9[72]},
      {stage2_9[27]}
   );
   gpc1_1 gpc997 (
      {stage1_9[73]},
      {stage2_9[28]}
   );
   gpc1_1 gpc998 (
      {stage1_9[74]},
      {stage2_9[29]}
   );
   gpc1_1 gpc999 (
      {stage1_9[75]},
      {stage2_9[30]}
   );
   gpc1_1 gpc1000 (
      {stage1_9[76]},
      {stage2_9[31]}
   );
   gpc1_1 gpc1001 (
      {stage1_10[75]},
      {stage2_10[28]}
   );
   gpc1_1 gpc1002 (
      {stage1_10[76]},
      {stage2_10[29]}
   );
   gpc1_1 gpc1003 (
      {stage1_10[77]},
      {stage2_10[30]}
   );
   gpc1_1 gpc1004 (
      {stage1_10[78]},
      {stage2_10[31]}
   );
   gpc1_1 gpc1005 (
      {stage1_10[79]},
      {stage2_10[32]}
   );
   gpc1_1 gpc1006 (
      {stage1_10[80]},
      {stage2_10[33]}
   );
   gpc1_1 gpc1007 (
      {stage1_10[81]},
      {stage2_10[34]}
   );
   gpc1_1 gpc1008 (
      {stage1_10[82]},
      {stage2_10[35]}
   );
   gpc1_1 gpc1009 (
      {stage1_10[83]},
      {stage2_10[36]}
   );
   gpc1_1 gpc1010 (
      {stage1_10[84]},
      {stage2_10[37]}
   );
   gpc1_1 gpc1011 (
      {stage1_10[85]},
      {stage2_10[38]}
   );
   gpc1_1 gpc1012 (
      {stage1_10[86]},
      {stage2_10[39]}
   );
   gpc1_1 gpc1013 (
      {stage1_10[87]},
      {stage2_10[40]}
   );
   gpc1_1 gpc1014 (
      {stage1_10[88]},
      {stage2_10[41]}
   );
   gpc1_1 gpc1015 (
      {stage1_10[89]},
      {stage2_10[42]}
   );
   gpc1_1 gpc1016 (
      {stage1_10[90]},
      {stage2_10[43]}
   );
   gpc1_1 gpc1017 (
      {stage1_10[91]},
      {stage2_10[44]}
   );
   gpc1_1 gpc1018 (
      {stage1_10[92]},
      {stage2_10[45]}
   );
   gpc1_1 gpc1019 (
      {stage1_11[58]},
      {stage2_11[30]}
   );
   gpc1_1 gpc1020 (
      {stage1_11[59]},
      {stage2_11[31]}
   );
   gpc1_1 gpc1021 (
      {stage1_11[60]},
      {stage2_11[32]}
   );
   gpc1_1 gpc1022 (
      {stage1_11[61]},
      {stage2_11[33]}
   );
   gpc1_1 gpc1023 (
      {stage1_11[62]},
      {stage2_11[34]}
   );
   gpc1_1 gpc1024 (
      {stage1_11[63]},
      {stage2_11[35]}
   );
   gpc1_1 gpc1025 (
      {stage1_11[64]},
      {stage2_11[36]}
   );
   gpc1_1 gpc1026 (
      {stage1_11[65]},
      {stage2_11[37]}
   );
   gpc1_1 gpc1027 (
      {stage1_11[66]},
      {stage2_11[38]}
   );
   gpc1_1 gpc1028 (
      {stage1_13[66]},
      {stage2_13[25]}
   );
   gpc1_1 gpc1029 (
      {stage1_13[67]},
      {stage2_13[26]}
   );
   gpc1_1 gpc1030 (
      {stage1_13[68]},
      {stage2_13[27]}
   );
   gpc1_1 gpc1031 (
      {stage1_13[69]},
      {stage2_13[28]}
   );
   gpc1_1 gpc1032 (
      {stage1_13[70]},
      {stage2_13[29]}
   );
   gpc1_1 gpc1033 (
      {stage1_13[71]},
      {stage2_13[30]}
   );
   gpc1_1 gpc1034 (
      {stage1_13[72]},
      {stage2_13[31]}
   );
   gpc1_1 gpc1035 (
      {stage1_13[73]},
      {stage2_13[32]}
   );
   gpc1_1 gpc1036 (
      {stage1_13[74]},
      {stage2_13[33]}
   );
   gpc1_1 gpc1037 (
      {stage1_13[75]},
      {stage2_13[34]}
   );
   gpc1_1 gpc1038 (
      {stage1_13[76]},
      {stage2_13[35]}
   );
   gpc1_1 gpc1039 (
      {stage1_13[77]},
      {stage2_13[36]}
   );
   gpc1_1 gpc1040 (
      {stage1_13[78]},
      {stage2_13[37]}
   );
   gpc1_1 gpc1041 (
      {stage1_13[79]},
      {stage2_13[38]}
   );
   gpc1_1 gpc1042 (
      {stage1_13[80]},
      {stage2_13[39]}
   );
   gpc1_1 gpc1043 (
      {stage1_13[81]},
      {stage2_13[40]}
   );
   gpc1_1 gpc1044 (
      {stage1_13[82]},
      {stage2_13[41]}
   );
   gpc1_1 gpc1045 (
      {stage1_13[83]},
      {stage2_13[42]}
   );
   gpc1_1 gpc1046 (
      {stage1_13[84]},
      {stage2_13[43]}
   );
   gpc1_1 gpc1047 (
      {stage1_13[85]},
      {stage2_13[44]}
   );
   gpc1_1 gpc1048 (
      {stage1_14[60]},
      {stage2_14[28]}
   );
   gpc1_1 gpc1049 (
      {stage1_14[61]},
      {stage2_14[29]}
   );
   gpc1_1 gpc1050 (
      {stage1_14[62]},
      {stage2_14[30]}
   );
   gpc1_1 gpc1051 (
      {stage1_14[63]},
      {stage2_14[31]}
   );
   gpc1_1 gpc1052 (
      {stage1_14[64]},
      {stage2_14[32]}
   );
   gpc1_1 gpc1053 (
      {stage1_14[65]},
      {stage2_14[33]}
   );
   gpc1_1 gpc1054 (
      {stage1_14[66]},
      {stage2_14[34]}
   );
   gpc1_1 gpc1055 (
      {stage1_14[67]},
      {stage2_14[35]}
   );
   gpc1_1 gpc1056 (
      {stage1_14[68]},
      {stage2_14[36]}
   );
   gpc1_1 gpc1057 (
      {stage1_15[50]},
      {stage2_15[24]}
   );
   gpc1_1 gpc1058 (
      {stage1_15[51]},
      {stage2_15[25]}
   );
   gpc1_1 gpc1059 (
      {stage1_15[52]},
      {stage2_15[26]}
   );
   gpc1_1 gpc1060 (
      {stage1_15[53]},
      {stage2_15[27]}
   );
   gpc1_1 gpc1061 (
      {stage1_15[54]},
      {stage2_15[28]}
   );
   gpc1_1 gpc1062 (
      {stage1_15[55]},
      {stage2_15[29]}
   );
   gpc1_1 gpc1063 (
      {stage1_15[56]},
      {stage2_15[30]}
   );
   gpc1_1 gpc1064 (
      {stage1_15[57]},
      {stage2_15[31]}
   );
   gpc1_1 gpc1065 (
      {stage1_15[58]},
      {stage2_15[32]}
   );
   gpc1_1 gpc1066 (
      {stage1_15[59]},
      {stage2_15[33]}
   );
   gpc1_1 gpc1067 (
      {stage1_16[90]},
      {stage2_16[27]}
   );
   gpc1_1 gpc1068 (
      {stage1_16[91]},
      {stage2_16[28]}
   );
   gpc1_1 gpc1069 (
      {stage1_16[92]},
      {stage2_16[29]}
   );
   gpc1_1 gpc1070 (
      {stage1_16[93]},
      {stage2_16[30]}
   );
   gpc1_1 gpc1071 (
      {stage1_16[94]},
      {stage2_16[31]}
   );
   gpc1_1 gpc1072 (
      {stage1_16[95]},
      {stage2_16[32]}
   );
   gpc1_1 gpc1073 (
      {stage1_16[96]},
      {stage2_16[33]}
   );
   gpc1_1 gpc1074 (
      {stage1_16[97]},
      {stage2_16[34]}
   );
   gpc1_1 gpc1075 (
      {stage1_16[98]},
      {stage2_16[35]}
   );
   gpc1_1 gpc1076 (
      {stage1_16[99]},
      {stage2_16[36]}
   );
   gpc1_1 gpc1077 (
      {stage1_16[100]},
      {stage2_16[37]}
   );
   gpc1_1 gpc1078 (
      {stage1_16[101]},
      {stage2_16[38]}
   );
   gpc1_1 gpc1079 (
      {stage1_16[102]},
      {stage2_16[39]}
   );
   gpc1_1 gpc1080 (
      {stage1_16[103]},
      {stage2_16[40]}
   );
   gpc1_1 gpc1081 (
      {stage1_16[104]},
      {stage2_16[41]}
   );
   gpc1_1 gpc1082 (
      {stage1_16[105]},
      {stage2_16[42]}
   );
   gpc1_1 gpc1083 (
      {stage1_16[106]},
      {stage2_16[43]}
   );
   gpc1_1 gpc1084 (
      {stage1_17[58]},
      {stage2_17[31]}
   );
   gpc1_1 gpc1085 (
      {stage1_17[59]},
      {stage2_17[32]}
   );
   gpc1_1 gpc1086 (
      {stage1_17[60]},
      {stage2_17[33]}
   );
   gpc1_1 gpc1087 (
      {stage1_17[61]},
      {stage2_17[34]}
   );
   gpc1_1 gpc1088 (
      {stage1_17[62]},
      {stage2_17[35]}
   );
   gpc1_1 gpc1089 (
      {stage1_17[63]},
      {stage2_17[36]}
   );
   gpc1_1 gpc1090 (
      {stage1_19[66]},
      {stage2_19[27]}
   );
   gpc1_1 gpc1091 (
      {stage1_20[52]},
      {stage2_20[29]}
   );
   gpc1_1 gpc1092 (
      {stage1_20[53]},
      {stage2_20[30]}
   );
   gpc1_1 gpc1093 (
      {stage1_20[54]},
      {stage2_20[31]}
   );
   gpc1_1 gpc1094 (
      {stage1_20[55]},
      {stage2_20[32]}
   );
   gpc1_1 gpc1095 (
      {stage1_20[56]},
      {stage2_20[33]}
   );
   gpc1_1 gpc1096 (
      {stage1_20[57]},
      {stage2_20[34]}
   );
   gpc1_1 gpc1097 (
      {stage1_20[58]},
      {stage2_20[35]}
   );
   gpc1_1 gpc1098 (
      {stage1_20[59]},
      {stage2_20[36]}
   );
   gpc1_1 gpc1099 (
      {stage1_20[60]},
      {stage2_20[37]}
   );
   gpc1_1 gpc1100 (
      {stage1_22[78]},
      {stage2_22[30]}
   );
   gpc1_1 gpc1101 (
      {stage1_22[79]},
      {stage2_22[31]}
   );
   gpc1_1 gpc1102 (
      {stage1_22[80]},
      {stage2_22[32]}
   );
   gpc1_1 gpc1103 (
      {stage1_22[81]},
      {stage2_22[33]}
   );
   gpc1_1 gpc1104 (
      {stage1_23[78]},
      {stage2_23[31]}
   );
   gpc1_1 gpc1105 (
      {stage1_23[79]},
      {stage2_23[32]}
   );
   gpc1_1 gpc1106 (
      {stage1_23[80]},
      {stage2_23[33]}
   );
   gpc1_1 gpc1107 (
      {stage1_23[81]},
      {stage2_23[34]}
   );
   gpc1_1 gpc1108 (
      {stage1_23[82]},
      {stage2_23[35]}
   );
   gpc1_1 gpc1109 (
      {stage1_23[83]},
      {stage2_23[36]}
   );
   gpc1_1 gpc1110 (
      {stage1_23[84]},
      {stage2_23[37]}
   );
   gpc1_1 gpc1111 (
      {stage1_23[85]},
      {stage2_23[38]}
   );
   gpc1_1 gpc1112 (
      {stage1_23[86]},
      {stage2_23[39]}
   );
   gpc1_1 gpc1113 (
      {stage1_23[87]},
      {stage2_23[40]}
   );
   gpc1_1 gpc1114 (
      {stage1_23[88]},
      {stage2_23[41]}
   );
   gpc1_1 gpc1115 (
      {stage1_23[89]},
      {stage2_23[42]}
   );
   gpc1_1 gpc1116 (
      {stage1_23[90]},
      {stage2_23[43]}
   );
   gpc1_1 gpc1117 (
      {stage1_24[60]},
      {stage2_24[28]}
   );
   gpc1_1 gpc1118 (
      {stage1_24[61]},
      {stage2_24[29]}
   );
   gpc1_1 gpc1119 (
      {stage1_24[62]},
      {stage2_24[30]}
   );
   gpc1_1 gpc1120 (
      {stage1_24[63]},
      {stage2_24[31]}
   );
   gpc1_1 gpc1121 (
      {stage1_24[64]},
      {stage2_24[32]}
   );
   gpc1_1 gpc1122 (
      {stage1_24[65]},
      {stage2_24[33]}
   );
   gpc1_1 gpc1123 (
      {stage1_24[66]},
      {stage2_24[34]}
   );
   gpc1_1 gpc1124 (
      {stage1_26[54]},
      {stage2_26[30]}
   );
   gpc1_1 gpc1125 (
      {stage1_27[58]},
      {stage2_27[24]}
   );
   gpc1_1 gpc1126 (
      {stage1_27[59]},
      {stage2_27[25]}
   );
   gpc1_1 gpc1127 (
      {stage1_27[60]},
      {stage2_27[26]}
   );
   gpc1_1 gpc1128 (
      {stage1_27[61]},
      {stage2_27[27]}
   );
   gpc1_1 gpc1129 (
      {stage1_27[62]},
      {stage2_27[28]}
   );
   gpc1_1 gpc1130 (
      {stage1_27[63]},
      {stage2_27[29]}
   );
   gpc1_1 gpc1131 (
      {stage1_27[64]},
      {stage2_27[30]}
   );
   gpc1_1 gpc1132 (
      {stage1_27[65]},
      {stage2_27[31]}
   );
   gpc1_1 gpc1133 (
      {stage1_27[66]},
      {stage2_27[32]}
   );
   gpc1_1 gpc1134 (
      {stage1_28[72]},
      {stage2_28[24]}
   );
   gpc1_1 gpc1135 (
      {stage1_28[73]},
      {stage2_28[25]}
   );
   gpc1_1 gpc1136 (
      {stage1_28[74]},
      {stage2_28[26]}
   );
   gpc1_1 gpc1137 (
      {stage1_28[75]},
      {stage2_28[27]}
   );
   gpc1_1 gpc1138 (
      {stage1_28[76]},
      {stage2_28[28]}
   );
   gpc1_1 gpc1139 (
      {stage1_28[77]},
      {stage2_28[29]}
   );
   gpc1_1 gpc1140 (
      {stage1_30[55]},
      {stage2_30[29]}
   );
   gpc1_1 gpc1141 (
      {stage1_30[56]},
      {stage2_30[30]}
   );
   gpc1_1 gpc1142 (
      {stage1_30[57]},
      {stage2_30[31]}
   );
   gpc1_1 gpc1143 (
      {stage1_30[58]},
      {stage2_30[32]}
   );
   gpc1_1 gpc1144 (
      {stage1_30[59]},
      {stage2_30[33]}
   );
   gpc1_1 gpc1145 (
      {stage1_30[60]},
      {stage2_30[34]}
   );
   gpc1_1 gpc1146 (
      {stage1_30[61]},
      {stage2_30[35]}
   );
   gpc1_1 gpc1147 (
      {stage1_30[62]},
      {stage2_30[36]}
   );
   gpc1_1 gpc1148 (
      {stage1_31[87]},
      {stage2_31[25]}
   );
   gpc1_1 gpc1149 (
      {stage1_31[88]},
      {stage2_31[26]}
   );
   gpc1_1 gpc1150 (
      {stage1_31[89]},
      {stage2_31[27]}
   );
   gpc1_1 gpc1151 (
      {stage1_31[90]},
      {stage2_31[28]}
   );
   gpc1_1 gpc1152 (
      {stage1_31[91]},
      {stage2_31[29]}
   );
   gpc1_1 gpc1153 (
      {stage1_31[92]},
      {stage2_31[30]}
   );
   gpc1_1 gpc1154 (
      {stage1_31[93]},
      {stage2_31[31]}
   );
   gpc1_1 gpc1155 (
      {stage1_31[94]},
      {stage2_31[32]}
   );
   gpc1_1 gpc1156 (
      {stage1_31[95]},
      {stage2_31[33]}
   );
   gpc1_1 gpc1157 (
      {stage1_31[96]},
      {stage2_31[34]}
   );
   gpc1_1 gpc1158 (
      {stage1_31[97]},
      {stage2_31[35]}
   );
   gpc1_1 gpc1159 (
      {stage1_32[27]},
      {stage2_32[23]}
   );
   gpc1_1 gpc1160 (
      {stage1_32[28]},
      {stage2_32[24]}
   );
   gpc1_1 gpc1161 (
      {stage1_32[29]},
      {stage2_32[25]}
   );
   gpc1_1 gpc1162 (
      {stage1_32[30]},
      {stage2_32[26]}
   );
   gpc1_1 gpc1163 (
      {stage1_32[31]},
      {stage2_32[27]}
   );
   gpc1_1 gpc1164 (
      {stage1_32[32]},
      {stage2_32[28]}
   );
   gpc1_1 gpc1165 (
      {stage1_32[33]},
      {stage2_32[29]}
   );
   gpc1_1 gpc1166 (
      {stage1_32[34]},
      {stage2_32[30]}
   );
   gpc1_1 gpc1167 (
      {stage1_32[35]},
      {stage2_32[31]}
   );
   gpc1_1 gpc1168 (
      {stage1_32[36]},
      {stage2_32[32]}
   );
   gpc1_1 gpc1169 (
      {stage1_32[37]},
      {stage2_32[33]}
   );
   gpc1_1 gpc1170 (
      {stage1_32[38]},
      {stage2_32[34]}
   );
   gpc1_1 gpc1171 (
      {stage1_32[39]},
      {stage2_32[35]}
   );
   gpc1_1 gpc1172 (
      {stage1_32[40]},
      {stage2_32[36]}
   );
   gpc1_1 gpc1173 (
      {stage1_32[41]},
      {stage2_32[37]}
   );
   gpc1_1 gpc1174 (
      {stage1_32[42]},
      {stage2_32[38]}
   );
   gpc1_1 gpc1175 (
      {stage1_32[43]},
      {stage2_32[39]}
   );
   gpc1_1 gpc1176 (
      {stage1_32[44]},
      {stage2_32[40]}
   );
   gpc1_1 gpc1177 (
      {stage1_33[13]},
      {stage2_33[18]}
   );
   gpc1_1 gpc1178 (
      {stage1_33[14]},
      {stage2_33[19]}
   );
   gpc1_1 gpc1179 (
      {stage1_33[15]},
      {stage2_33[20]}
   );
   gpc1_1 gpc1180 (
      {stage1_33[16]},
      {stage2_33[21]}
   );
   gpc1_1 gpc1181 (
      {stage1_33[17]},
      {stage2_33[22]}
   );
   gpc1_1 gpc1182 (
      {stage1_33[18]},
      {stage2_33[23]}
   );
   gpc135_4 gpc1183 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4]},
      {stage2_1[0], stage2_1[1], stage2_1[2]},
      {stage2_2[0]},
      {stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc1184 (
      {stage2_1[3], stage2_1[4], stage2_1[5], stage2_1[6], stage2_1[7], stage2_1[8]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[0],stage3_3[1],stage3_2[1],stage3_1[1]}
   );
   gpc615_5 gpc1185 (
      {stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage2_3[6]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[1],stage3_4[1],stage3_3[2],stage3_2[2]}
   );
   gpc615_5 gpc1186 (
      {stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10]},
      {stage2_3[7]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[2],stage3_4[2],stage3_3[3],stage3_2[3]}
   );
   gpc1163_5 gpc1187 (
      {stage2_3[8], stage2_3[9], stage2_3[10]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage2_5[0]},
      {stage2_6[0]},
      {stage3_7[0],stage3_6[2],stage3_5[3],stage3_4[3],stage3_3[4]}
   );
   gpc1163_5 gpc1188 (
      {stage2_3[11], stage2_3[12], stage2_3[13]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage2_5[1]},
      {stage2_6[1]},
      {stage3_7[1],stage3_6[3],stage3_5[4],stage3_4[4],stage3_3[5]}
   );
   gpc1163_5 gpc1189 (
      {stage2_3[14], stage2_3[15], stage2_3[16]},
      {stage2_4[24], stage2_4[25], stage2_4[26], stage2_4[27], stage2_4[28], stage2_4[29]},
      {stage2_5[2]},
      {stage2_6[2]},
      {stage3_7[2],stage3_6[4],stage3_5[5],stage3_4[5],stage3_3[6]}
   );
   gpc623_5 gpc1190 (
      {stage2_3[17], stage2_3[18], stage2_3[19]},
      {stage2_4[30], stage2_4[31]},
      {stage2_5[3], stage2_5[4], stage2_5[5], stage2_5[6], stage2_5[7], stage2_5[8]},
      {stage3_7[3],stage3_6[5],stage3_5[6],stage3_4[6],stage3_3[7]}
   );
   gpc615_5 gpc1191 (
      {stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35], stage2_4[36]},
      {stage2_5[9]},
      {stage2_6[3], stage2_6[4], stage2_6[5], stage2_6[6], stage2_6[7], stage2_6[8]},
      {stage3_8[0],stage3_7[4],stage3_6[6],stage3_5[7],stage3_4[7]}
   );
   gpc615_5 gpc1192 (
      {stage2_4[37], stage2_4[38], stage2_4[39], stage2_4[40], 1'b0},
      {stage2_5[10]},
      {stage2_6[9], stage2_6[10], stage2_6[11], stage2_6[12], stage2_6[13], stage2_6[14]},
      {stage3_8[1],stage3_7[5],stage3_6[7],stage3_5[8],stage3_4[8]}
   );
   gpc606_5 gpc1193 (
      {stage2_5[11], stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[2],stage3_7[6],stage3_6[8],stage3_5[9]}
   );
   gpc606_5 gpc1194 (
      {stage2_5[17], stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[3],stage3_7[7],stage3_6[9],stage3_5[10]}
   );
   gpc606_5 gpc1195 (
      {stage2_5[23], stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], 1'b0},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[4],stage3_7[8],stage3_6[10],stage3_5[11]}
   );
   gpc606_5 gpc1196 (
      {stage2_6[15], stage2_6[16], stage2_6[17], stage2_6[18], stage2_6[19], stage2_6[20]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[3],stage3_8[5],stage3_7[9],stage3_6[11]}
   );
   gpc606_5 gpc1197 (
      {stage2_6[21], stage2_6[22], stage2_6[23], stage2_6[24], stage2_6[25], stage2_6[26]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[4],stage3_8[6],stage3_7[10],stage3_6[12]}
   );
   gpc615_5 gpc1198 (
      {stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22]},
      {stage2_8[12]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[2],stage3_9[5],stage3_8[7],stage3_7[11]}
   );
   gpc615_5 gpc1199 (
      {stage2_7[23], stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27]},
      {stage2_8[13]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[3],stage3_9[6],stage3_8[8],stage3_7[12]}
   );
   gpc606_5 gpc1200 (
      {stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17], stage2_8[18], stage2_8[19]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[2],stage3_10[4],stage3_9[7],stage3_8[9]}
   );
   gpc606_5 gpc1201 (
      {stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23], stage2_8[24], stage2_8[25]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[3],stage3_10[5],stage3_9[8],stage3_8[10]}
   );
   gpc1343_5 gpc1202 (
      {stage2_9[12], stage2_9[13], stage2_9[14]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15]},
      {stage2_11[0], stage2_11[1], stage2_11[2]},
      {stage2_12[0]},
      {stage3_13[0],stage3_12[2],stage3_11[4],stage3_10[6],stage3_9[9]}
   );
   gpc1343_5 gpc1203 (
      {stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage2_10[16], stage2_10[17], stage2_10[18], stage2_10[19]},
      {stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage2_12[1]},
      {stage3_13[1],stage3_12[3],stage3_11[5],stage3_10[7],stage3_9[10]}
   );
   gpc1343_5 gpc1204 (
      {stage2_9[18], stage2_9[19], stage2_9[20]},
      {stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage2_11[6], stage2_11[7], stage2_11[8]},
      {stage2_12[2]},
      {stage3_13[2],stage3_12[4],stage3_11[6],stage3_10[8],stage3_9[11]}
   );
   gpc1343_5 gpc1205 (
      {stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27]},
      {stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage2_12[3]},
      {stage3_13[3],stage3_12[5],stage3_11[7],stage3_10[9],stage3_9[12]}
   );
   gpc1343_5 gpc1206 (
      {stage2_9[24], stage2_9[25], stage2_9[26]},
      {stage2_10[28], stage2_10[29], stage2_10[30], stage2_10[31]},
      {stage2_11[12], stage2_11[13], stage2_11[14]},
      {stage2_12[4]},
      {stage3_13[4],stage3_12[6],stage3_11[8],stage3_10[10],stage3_9[13]}
   );
   gpc606_5 gpc1207 (
      {stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35], stage2_10[36], stage2_10[37]},
      {stage2_12[5], stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10]},
      {stage3_14[0],stage3_13[5],stage3_12[7],stage3_11[9],stage3_10[11]}
   );
   gpc606_5 gpc1208 (
      {stage2_10[38], stage2_10[39], stage2_10[40], stage2_10[41], stage2_10[42], stage2_10[43]},
      {stage2_12[11], stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16]},
      {stage3_14[1],stage3_13[6],stage3_12[8],stage3_11[10],stage3_10[12]}
   );
   gpc606_5 gpc1209 (
      {stage2_11[15], stage2_11[16], stage2_11[17], stage2_11[18], stage2_11[19], stage2_11[20]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[2],stage3_13[7],stage3_12[9],stage3_11[11]}
   );
   gpc606_5 gpc1210 (
      {stage2_11[21], stage2_11[22], stage2_11[23], stage2_11[24], stage2_11[25], stage2_11[26]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[3],stage3_13[8],stage3_12[10],stage3_11[12]}
   );
   gpc606_5 gpc1211 (
      {stage2_11[27], stage2_11[28], stage2_11[29], stage2_11[30], stage2_11[31], stage2_11[32]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[4],stage3_13[9],stage3_12[11],stage3_11[13]}
   );
   gpc606_5 gpc1212 (
      {stage2_11[33], stage2_11[34], stage2_11[35], stage2_11[36], stage2_11[37], stage2_11[38]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[5],stage3_13[10],stage3_12[12],stage3_11[14]}
   );
   gpc606_5 gpc1213 (
      {stage2_12[17], stage2_12[18], stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[4],stage3_14[6],stage3_13[11],stage3_12[13]}
   );
   gpc606_5 gpc1214 (
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[1],stage3_15[5],stage3_14[7],stage3_13[12]}
   );
   gpc606_5 gpc1215 (
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage3_17[1],stage3_16[2],stage3_15[6],stage3_14[8],stage3_13[13]}
   );
   gpc606_5 gpc1216 (
      {stage2_13[36], stage2_13[37], stage2_13[38], stage2_13[39], stage2_13[40], stage2_13[41]},
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17]},
      {stage3_17[2],stage3_16[3],stage3_15[7],stage3_14[9],stage3_13[14]}
   );
   gpc615_5 gpc1217 (
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10]},
      {stage2_15[18]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[3],stage3_16[4],stage3_15[8],stage3_14[10]}
   );
   gpc615_5 gpc1218 (
      {stage2_14[11], stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15]},
      {stage2_15[19]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[4],stage3_16[5],stage3_15[9],stage3_14[11]}
   );
   gpc615_5 gpc1219 (
      {stage2_14[16], stage2_14[17], stage2_14[18], stage2_14[19], stage2_14[20]},
      {stage2_15[20]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[5],stage3_16[6],stage3_15[10],stage3_14[12]}
   );
   gpc615_5 gpc1220 (
      {stage2_14[21], stage2_14[22], stage2_14[23], stage2_14[24], stage2_14[25]},
      {stage2_15[21]},
      {stage2_16[18], stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23]},
      {stage3_18[3],stage3_17[6],stage3_16[7],stage3_15[11],stage3_14[13]}
   );
   gpc615_5 gpc1221 (
      {stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29], stage2_14[30]},
      {stage2_15[22]},
      {stage2_16[24], stage2_16[25], stage2_16[26], stage2_16[27], stage2_16[28], stage2_16[29]},
      {stage3_18[4],stage3_17[7],stage3_16[8],stage3_15[12],stage3_14[14]}
   );
   gpc615_5 gpc1222 (
      {stage2_14[31], stage2_14[32], stage2_14[33], stage2_14[34], stage2_14[35]},
      {stage2_15[23]},
      {stage2_16[30], stage2_16[31], stage2_16[32], stage2_16[33], stage2_16[34], stage2_16[35]},
      {stage3_18[5],stage3_17[8],stage3_16[9],stage3_15[13],stage3_14[15]}
   );
   gpc615_5 gpc1223 (
      {stage2_15[24], stage2_15[25], stage2_15[26], stage2_15[27], stage2_15[28]},
      {stage2_16[36]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[6],stage3_17[9],stage3_16[10],stage3_15[14]}
   );
   gpc615_5 gpc1224 (
      {stage2_15[29], stage2_15[30], stage2_15[31], stage2_15[32], stage2_15[33]},
      {stage2_16[37]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[7],stage3_17[10],stage3_16[11],stage3_15[15]}
   );
   gpc606_5 gpc1225 (
      {stage2_16[38], stage2_16[39], stage2_16[40], stage2_16[41], stage2_16[42], stage2_16[43]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[2],stage3_18[8],stage3_17[11],stage3_16[12]}
   );
   gpc606_5 gpc1226 (
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[1],stage3_19[3],stage3_18[9],stage3_17[12]}
   );
   gpc606_5 gpc1227 (
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23]},
      {stage2_19[6], stage2_19[7], stage2_19[8], stage2_19[9], stage2_19[10], stage2_19[11]},
      {stage3_21[1],stage3_20[2],stage3_19[4],stage3_18[10],stage3_17[13]}
   );
   gpc606_5 gpc1228 (
      {stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29]},
      {stage2_19[12], stage2_19[13], stage2_19[14], stage2_19[15], stage2_19[16], stage2_19[17]},
      {stage3_21[2],stage3_20[3],stage3_19[5],stage3_18[11],stage3_17[14]}
   );
   gpc606_5 gpc1229 (
      {stage2_17[30], stage2_17[31], stage2_17[32], stage2_17[33], stage2_17[34], stage2_17[35]},
      {stage2_19[18], stage2_19[19], stage2_19[20], stage2_19[21], stage2_19[22], stage2_19[23]},
      {stage3_21[3],stage3_20[4],stage3_19[6],stage3_18[12],stage3_17[15]}
   );
   gpc606_5 gpc1230 (
      {stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10], stage2_18[11]},
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage3_22[0],stage3_21[4],stage3_20[5],stage3_19[7],stage3_18[13]}
   );
   gpc606_5 gpc1231 (
      {stage2_18[12], stage2_18[13], stage2_18[14], stage2_18[15], stage2_18[16], stage2_18[17]},
      {stage2_20[6], stage2_20[7], stage2_20[8], stage2_20[9], stage2_20[10], stage2_20[11]},
      {stage3_22[1],stage3_21[5],stage3_20[6],stage3_19[8],stage3_18[14]}
   );
   gpc606_5 gpc1232 (
      {stage2_18[18], stage2_18[19], stage2_18[20], stage2_18[21], stage2_18[22], stage2_18[23]},
      {stage2_20[12], stage2_20[13], stage2_20[14], stage2_20[15], stage2_20[16], stage2_20[17]},
      {stage3_22[2],stage3_21[6],stage3_20[7],stage3_19[9],stage3_18[15]}
   );
   gpc615_5 gpc1233 (
      {stage2_18[24], stage2_18[25], stage2_18[26], stage2_18[27], stage2_18[28]},
      {stage2_19[24]},
      {stage2_20[18], stage2_20[19], stage2_20[20], stage2_20[21], stage2_20[22], stage2_20[23]},
      {stage3_22[3],stage3_21[7],stage3_20[8],stage3_19[10],stage3_18[16]}
   );
   gpc615_5 gpc1234 (
      {stage2_19[25], stage2_19[26], stage2_19[27], 1'b0, 1'b0},
      {stage2_20[24]},
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3], stage2_21[4], stage2_21[5]},
      {stage3_23[0],stage3_22[4],stage3_21[8],stage3_20[9],stage3_19[11]}
   );
   gpc606_5 gpc1235 (
      {stage2_20[25], stage2_20[26], stage2_20[27], stage2_20[28], stage2_20[29], stage2_20[30]},
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage3_24[0],stage3_23[1],stage3_22[5],stage3_21[9],stage3_20[10]}
   );
   gpc615_5 gpc1236 (
      {stage2_21[6], stage2_21[7], stage2_21[8], stage2_21[9], stage2_21[10]},
      {stage2_22[6]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[1],stage3_23[2],stage3_22[6],stage3_21[10]}
   );
   gpc615_5 gpc1237 (
      {stage2_21[11], stage2_21[12], stage2_21[13], stage2_21[14], stage2_21[15]},
      {stage2_22[7]},
      {stage2_23[6], stage2_23[7], stage2_23[8], stage2_23[9], stage2_23[10], stage2_23[11]},
      {stage3_25[1],stage3_24[2],stage3_23[3],stage3_22[7],stage3_21[11]}
   );
   gpc615_5 gpc1238 (
      {stage2_21[16], stage2_21[17], stage2_21[18], stage2_21[19], stage2_21[20]},
      {stage2_22[8]},
      {stage2_23[12], stage2_23[13], stage2_23[14], stage2_23[15], stage2_23[16], stage2_23[17]},
      {stage3_25[2],stage3_24[3],stage3_23[4],stage3_22[8],stage3_21[12]}
   );
   gpc615_5 gpc1239 (
      {stage2_21[21], stage2_21[22], stage2_21[23], stage2_21[24], stage2_21[25]},
      {stage2_22[9]},
      {stage2_23[18], stage2_23[19], stage2_23[20], stage2_23[21], stage2_23[22], stage2_23[23]},
      {stage3_25[3],stage3_24[4],stage3_23[5],stage3_22[9],stage3_21[13]}
   );
   gpc615_5 gpc1240 (
      {stage2_21[26], stage2_21[27], 1'b0, 1'b0, 1'b0},
      {stage2_22[10]},
      {stage2_23[24], stage2_23[25], stage2_23[26], stage2_23[27], stage2_23[28], stage2_23[29]},
      {stage3_25[4],stage3_24[5],stage3_23[6],stage3_22[10],stage3_21[14]}
   );
   gpc207_4 gpc1241 (
      {stage2_22[11], stage2_22[12], stage2_22[13], stage2_22[14], stage2_22[15], stage2_22[16], stage2_22[17]},
      {stage2_24[0], stage2_24[1]},
      {stage3_25[5],stage3_24[6],stage3_23[7],stage3_22[11]}
   );
   gpc606_5 gpc1242 (
      {stage2_22[18], stage2_22[19], stage2_22[20], stage2_22[21], stage2_22[22], stage2_22[23]},
      {stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5], stage2_24[6], stage2_24[7]},
      {stage3_26[0],stage3_25[6],stage3_24[7],stage3_23[8],stage3_22[12]}
   );
   gpc606_5 gpc1243 (
      {stage2_23[30], stage2_23[31], stage2_23[32], stage2_23[33], stage2_23[34], stage2_23[35]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage3_27[0],stage3_26[1],stage3_25[7],stage3_24[8],stage3_23[9]}
   );
   gpc606_5 gpc1244 (
      {stage2_23[36], stage2_23[37], stage2_23[38], stage2_23[39], stage2_23[40], stage2_23[41]},
      {stage2_25[6], stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11]},
      {stage3_27[1],stage3_26[2],stage3_25[8],stage3_24[9],stage3_23[10]}
   );
   gpc606_5 gpc1245 (
      {stage2_24[8], stage2_24[9], stage2_24[10], stage2_24[11], stage2_24[12], stage2_24[13]},
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage3_28[0],stage3_27[2],stage3_26[3],stage3_25[9],stage3_24[10]}
   );
   gpc606_5 gpc1246 (
      {stage2_24[14], stage2_24[15], stage2_24[16], stage2_24[17], stage2_24[18], stage2_24[19]},
      {stage2_26[6], stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11]},
      {stage3_28[1],stage3_27[3],stage3_26[4],stage3_25[10],stage3_24[11]}
   );
   gpc606_5 gpc1247 (
      {stage2_24[20], stage2_24[21], stage2_24[22], stage2_24[23], stage2_24[24], stage2_24[25]},
      {stage2_26[12], stage2_26[13], stage2_26[14], stage2_26[15], stage2_26[16], stage2_26[17]},
      {stage3_28[2],stage3_27[4],stage3_26[5],stage3_25[11],stage3_24[12]}
   );
   gpc606_5 gpc1248 (
      {stage2_24[26], stage2_24[27], stage2_24[28], stage2_24[29], stage2_24[30], stage2_24[31]},
      {stage2_26[18], stage2_26[19], stage2_26[20], stage2_26[21], stage2_26[22], stage2_26[23]},
      {stage3_28[3],stage3_27[5],stage3_26[6],stage3_25[12],stage3_24[13]}
   );
   gpc606_5 gpc1249 (
      {stage2_25[12], stage2_25[13], stage2_25[14], stage2_25[15], stage2_25[16], stage2_25[17]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage3_29[0],stage3_28[4],stage3_27[6],stage3_26[7],stage3_25[13]}
   );
   gpc606_5 gpc1250 (
      {stage2_25[18], stage2_25[19], stage2_25[20], stage2_25[21], stage2_25[22], stage2_25[23]},
      {stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11]},
      {stage3_29[1],stage3_28[5],stage3_27[7],stage3_26[8],stage3_25[14]}
   );
   gpc606_5 gpc1251 (
      {stage2_25[24], stage2_25[25], stage2_25[26], stage2_25[27], stage2_25[28], stage2_25[29]},
      {stage2_27[12], stage2_27[13], stage2_27[14], stage2_27[15], stage2_27[16], stage2_27[17]},
      {stage3_29[2],stage3_28[6],stage3_27[8],stage3_26[9],stage3_25[15]}
   );
   gpc606_5 gpc1252 (
      {stage2_26[24], stage2_26[25], stage2_26[26], stage2_26[27], stage2_26[28], stage2_26[29]},
      {stage2_28[0], stage2_28[1], stage2_28[2], stage2_28[3], stage2_28[4], stage2_28[5]},
      {stage3_30[0],stage3_29[3],stage3_28[7],stage3_27[9],stage3_26[10]}
   );
   gpc615_5 gpc1253 (
      {stage2_27[18], stage2_27[19], stage2_27[20], stage2_27[21], stage2_27[22]},
      {stage2_28[6]},
      {stage2_29[0], stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5]},
      {stage3_31[0],stage3_30[1],stage3_29[4],stage3_28[8],stage3_27[10]}
   );
   gpc615_5 gpc1254 (
      {stage2_27[23], stage2_27[24], stage2_27[25], stage2_27[26], stage2_27[27]},
      {stage2_28[7]},
      {stage2_29[6], stage2_29[7], stage2_29[8], stage2_29[9], stage2_29[10], stage2_29[11]},
      {stage3_31[1],stage3_30[2],stage3_29[5],stage3_28[9],stage3_27[11]}
   );
   gpc615_5 gpc1255 (
      {stage2_27[28], stage2_27[29], stage2_27[30], stage2_27[31], stage2_27[32]},
      {stage2_28[8]},
      {stage2_29[12], stage2_29[13], stage2_29[14], stage2_29[15], stage2_29[16], stage2_29[17]},
      {stage3_31[2],stage3_30[3],stage3_29[6],stage3_28[10],stage3_27[12]}
   );
   gpc135_4 gpc1256 (
      {stage2_28[9], stage2_28[10], stage2_28[11], stage2_28[12], stage2_28[13]},
      {stage2_29[18], stage2_29[19], stage2_29[20]},
      {stage2_30[0]},
      {stage3_31[3],stage3_30[4],stage3_29[7],stage3_28[11]}
   );
   gpc606_5 gpc1257 (
      {stage2_28[14], stage2_28[15], stage2_28[16], stage2_28[17], stage2_28[18], stage2_28[19]},
      {stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5], stage2_30[6]},
      {stage3_32[0],stage3_31[4],stage3_30[5],stage3_29[8],stage3_28[12]}
   );
   gpc606_5 gpc1258 (
      {stage2_29[21], stage2_29[22], stage2_29[23], stage2_29[24], stage2_29[25], stage2_29[26]},
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage3_33[0],stage3_32[1],stage3_31[5],stage3_30[6],stage3_29[9]}
   );
   gpc606_5 gpc1259 (
      {stage2_29[27], stage2_29[28], stage2_29[29], stage2_29[30], stage2_29[31], stage2_29[32]},
      {stage2_31[6], stage2_31[7], stage2_31[8], stage2_31[9], stage2_31[10], stage2_31[11]},
      {stage3_33[1],stage3_32[2],stage3_31[6],stage3_30[7],stage3_29[10]}
   );
   gpc615_5 gpc1260 (
      {stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage2_31[12]},
      {stage2_32[0], stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5]},
      {stage3_34[0],stage3_33[2],stage3_32[3],stage3_31[7],stage3_30[8]}
   );
   gpc615_5 gpc1261 (
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16]},
      {stage2_31[13]},
      {stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10], stage2_32[11]},
      {stage3_34[1],stage3_33[3],stage3_32[4],stage3_31[8],stage3_30[9]}
   );
   gpc615_5 gpc1262 (
      {stage2_30[17], stage2_30[18], stage2_30[19], stage2_30[20], stage2_30[21]},
      {stage2_31[14]},
      {stage2_32[12], stage2_32[13], stage2_32[14], stage2_32[15], stage2_32[16], stage2_32[17]},
      {stage3_34[2],stage3_33[4],stage3_32[5],stage3_31[9],stage3_30[10]}
   );
   gpc615_5 gpc1263 (
      {stage2_30[22], stage2_30[23], stage2_30[24], stage2_30[25], stage2_30[26]},
      {stage2_31[15]},
      {stage2_32[18], stage2_32[19], stage2_32[20], stage2_32[21], stage2_32[22], stage2_32[23]},
      {stage3_34[3],stage3_33[5],stage3_32[6],stage3_31[10],stage3_30[11]}
   );
   gpc615_5 gpc1264 (
      {stage2_30[27], stage2_30[28], stage2_30[29], stage2_30[30], stage2_30[31]},
      {stage2_31[16]},
      {stage2_32[24], stage2_32[25], stage2_32[26], stage2_32[27], stage2_32[28], stage2_32[29]},
      {stage3_34[4],stage3_33[6],stage3_32[7],stage3_31[11],stage3_30[12]}
   );
   gpc615_5 gpc1265 (
      {stage2_30[32], stage2_30[33], stage2_30[34], stage2_30[35], stage2_30[36]},
      {stage2_31[17]},
      {stage2_32[30], stage2_32[31], stage2_32[32], stage2_32[33], stage2_32[34], stage2_32[35]},
      {stage3_34[5],stage3_33[7],stage3_32[8],stage3_31[12],stage3_30[13]}
   );
   gpc606_5 gpc1266 (
      {stage2_31[18], stage2_31[19], stage2_31[20], stage2_31[21], stage2_31[22], stage2_31[23]},
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5]},
      {stage3_35[0],stage3_34[6],stage3_33[8],stage3_32[9],stage3_31[13]}
   );
   gpc606_5 gpc1267 (
      {stage2_31[24], stage2_31[25], stage2_31[26], stage2_31[27], stage2_31[28], stage2_31[29]},
      {stage2_33[6], stage2_33[7], stage2_33[8], stage2_33[9], stage2_33[10], stage2_33[11]},
      {stage3_35[1],stage3_34[7],stage3_33[9],stage3_32[10],stage3_31[14]}
   );
   gpc615_5 gpc1268 (
      {stage2_31[30], stage2_31[31], stage2_31[32], stage2_31[33], stage2_31[34]},
      {stage2_32[36]},
      {stage2_33[12], stage2_33[13], stage2_33[14], stage2_33[15], stage2_33[16], stage2_33[17]},
      {stage3_35[2],stage3_34[8],stage3_33[10],stage3_32[11],stage3_31[15]}
   );
   gpc1_1 gpc1269 (
      {stage2_0[5]},
      {stage3_0[1]}
   );
   gpc1_1 gpc1270 (
      {stage2_0[6]},
      {stage3_0[2]}
   );
   gpc1_1 gpc1271 (
      {stage2_0[7]},
      {stage3_0[3]}
   );
   gpc1_1 gpc1272 (
      {stage2_0[8]},
      {stage3_0[4]}
   );
   gpc1_1 gpc1273 (
      {stage2_0[9]},
      {stage3_0[5]}
   );
   gpc1_1 gpc1274 (
      {stage2_0[10]},
      {stage3_0[6]}
   );
   gpc1_1 gpc1275 (
      {stage2_1[9]},
      {stage3_1[2]}
   );
   gpc1_1 gpc1276 (
      {stage2_1[10]},
      {stage3_1[3]}
   );
   gpc1_1 gpc1277 (
      {stage2_1[11]},
      {stage3_1[4]}
   );
   gpc1_1 gpc1278 (
      {stage2_1[12]},
      {stage3_1[5]}
   );
   gpc1_1 gpc1279 (
      {stage2_1[13]},
      {stage3_1[6]}
   );
   gpc1_1 gpc1280 (
      {stage2_1[14]},
      {stage3_1[7]}
   );
   gpc1_1 gpc1281 (
      {stage2_1[15]},
      {stage3_1[8]}
   );
   gpc1_1 gpc1282 (
      {stage2_1[16]},
      {stage3_1[9]}
   );
   gpc1_1 gpc1283 (
      {stage2_2[11]},
      {stage3_2[4]}
   );
   gpc1_1 gpc1284 (
      {stage2_2[12]},
      {stage3_2[5]}
   );
   gpc1_1 gpc1285 (
      {stage2_2[13]},
      {stage3_2[6]}
   );
   gpc1_1 gpc1286 (
      {stage2_2[14]},
      {stage3_2[7]}
   );
   gpc1_1 gpc1287 (
      {stage2_2[15]},
      {stage3_2[8]}
   );
   gpc1_1 gpc1288 (
      {stage2_2[16]},
      {stage3_2[9]}
   );
   gpc1_1 gpc1289 (
      {stage2_3[20]},
      {stage3_3[8]}
   );
   gpc1_1 gpc1290 (
      {stage2_3[21]},
      {stage3_3[9]}
   );
   gpc1_1 gpc1291 (
      {stage2_3[22]},
      {stage3_3[10]}
   );
   gpc1_1 gpc1292 (
      {stage2_3[23]},
      {stage3_3[11]}
   );
   gpc1_1 gpc1293 (
      {stage2_3[24]},
      {stage3_3[12]}
   );
   gpc1_1 gpc1294 (
      {stage2_3[25]},
      {stage3_3[13]}
   );
   gpc1_1 gpc1295 (
      {stage2_3[26]},
      {stage3_3[14]}
   );
   gpc1_1 gpc1296 (
      {stage2_3[27]},
      {stage3_3[15]}
   );
   gpc1_1 gpc1297 (
      {stage2_3[28]},
      {stage3_3[16]}
   );
   gpc1_1 gpc1298 (
      {stage2_3[29]},
      {stage3_3[17]}
   );
   gpc1_1 gpc1299 (
      {stage2_3[30]},
      {stage3_3[18]}
   );
   gpc1_1 gpc1300 (
      {stage2_3[31]},
      {stage3_3[19]}
   );
   gpc1_1 gpc1301 (
      {stage2_3[32]},
      {stage3_3[20]}
   );
   gpc1_1 gpc1302 (
      {stage2_3[33]},
      {stage3_3[21]}
   );
   gpc1_1 gpc1303 (
      {stage2_3[34]},
      {stage3_3[22]}
   );
   gpc1_1 gpc1304 (
      {stage2_6[27]},
      {stage3_6[13]}
   );
   gpc1_1 gpc1305 (
      {stage2_6[28]},
      {stage3_6[14]}
   );
   gpc1_1 gpc1306 (
      {stage2_6[29]},
      {stage3_6[15]}
   );
   gpc1_1 gpc1307 (
      {stage2_6[30]},
      {stage3_6[16]}
   );
   gpc1_1 gpc1308 (
      {stage2_7[28]},
      {stage3_7[13]}
   );
   gpc1_1 gpc1309 (
      {stage2_7[29]},
      {stage3_7[14]}
   );
   gpc1_1 gpc1310 (
      {stage2_7[30]},
      {stage3_7[15]}
   );
   gpc1_1 gpc1311 (
      {stage2_7[31]},
      {stage3_7[16]}
   );
   gpc1_1 gpc1312 (
      {stage2_7[32]},
      {stage3_7[17]}
   );
   gpc1_1 gpc1313 (
      {stage2_7[33]},
      {stage3_7[18]}
   );
   gpc1_1 gpc1314 (
      {stage2_8[26]},
      {stage3_8[11]}
   );
   gpc1_1 gpc1315 (
      {stage2_8[27]},
      {stage3_8[12]}
   );
   gpc1_1 gpc1316 (
      {stage2_8[28]},
      {stage3_8[13]}
   );
   gpc1_1 gpc1317 (
      {stage2_8[29]},
      {stage3_8[14]}
   );
   gpc1_1 gpc1318 (
      {stage2_8[30]},
      {stage3_8[15]}
   );
   gpc1_1 gpc1319 (
      {stage2_8[31]},
      {stage3_8[16]}
   );
   gpc1_1 gpc1320 (
      {stage2_8[32]},
      {stage3_8[17]}
   );
   gpc1_1 gpc1321 (
      {stage2_9[27]},
      {stage3_9[14]}
   );
   gpc1_1 gpc1322 (
      {stage2_9[28]},
      {stage3_9[15]}
   );
   gpc1_1 gpc1323 (
      {stage2_9[29]},
      {stage3_9[16]}
   );
   gpc1_1 gpc1324 (
      {stage2_9[30]},
      {stage3_9[17]}
   );
   gpc1_1 gpc1325 (
      {stage2_9[31]},
      {stage3_9[18]}
   );
   gpc1_1 gpc1326 (
      {stage2_10[44]},
      {stage3_10[13]}
   );
   gpc1_1 gpc1327 (
      {stage2_10[45]},
      {stage3_10[14]}
   );
   gpc1_1 gpc1328 (
      {stage2_12[23]},
      {stage3_12[14]}
   );
   gpc1_1 gpc1329 (
      {stage2_13[42]},
      {stage3_13[15]}
   );
   gpc1_1 gpc1330 (
      {stage2_13[43]},
      {stage3_13[16]}
   );
   gpc1_1 gpc1331 (
      {stage2_13[44]},
      {stage3_13[17]}
   );
   gpc1_1 gpc1332 (
      {stage2_14[36]},
      {stage3_14[16]}
   );
   gpc1_1 gpc1333 (
      {stage2_17[36]},
      {stage3_17[16]}
   );
   gpc1_1 gpc1334 (
      {stage2_20[31]},
      {stage3_20[11]}
   );
   gpc1_1 gpc1335 (
      {stage2_20[32]},
      {stage3_20[12]}
   );
   gpc1_1 gpc1336 (
      {stage2_20[33]},
      {stage3_20[13]}
   );
   gpc1_1 gpc1337 (
      {stage2_20[34]},
      {stage3_20[14]}
   );
   gpc1_1 gpc1338 (
      {stage2_20[35]},
      {stage3_20[15]}
   );
   gpc1_1 gpc1339 (
      {stage2_20[36]},
      {stage3_20[16]}
   );
   gpc1_1 gpc1340 (
      {stage2_20[37]},
      {stage3_20[17]}
   );
   gpc1_1 gpc1341 (
      {stage2_22[24]},
      {stage3_22[13]}
   );
   gpc1_1 gpc1342 (
      {stage2_22[25]},
      {stage3_22[14]}
   );
   gpc1_1 gpc1343 (
      {stage2_22[26]},
      {stage3_22[15]}
   );
   gpc1_1 gpc1344 (
      {stage2_22[27]},
      {stage3_22[16]}
   );
   gpc1_1 gpc1345 (
      {stage2_22[28]},
      {stage3_22[17]}
   );
   gpc1_1 gpc1346 (
      {stage2_22[29]},
      {stage3_22[18]}
   );
   gpc1_1 gpc1347 (
      {stage2_22[30]},
      {stage3_22[19]}
   );
   gpc1_1 gpc1348 (
      {stage2_22[31]},
      {stage3_22[20]}
   );
   gpc1_1 gpc1349 (
      {stage2_22[32]},
      {stage3_22[21]}
   );
   gpc1_1 gpc1350 (
      {stage2_22[33]},
      {stage3_22[22]}
   );
   gpc1_1 gpc1351 (
      {stage2_23[42]},
      {stage3_23[11]}
   );
   gpc1_1 gpc1352 (
      {stage2_23[43]},
      {stage3_23[12]}
   );
   gpc1_1 gpc1353 (
      {stage2_24[32]},
      {stage3_24[14]}
   );
   gpc1_1 gpc1354 (
      {stage2_24[33]},
      {stage3_24[15]}
   );
   gpc1_1 gpc1355 (
      {stage2_24[34]},
      {stage3_24[16]}
   );
   gpc1_1 gpc1356 (
      {stage2_25[30]},
      {stage3_25[16]}
   );
   gpc1_1 gpc1357 (
      {stage2_26[30]},
      {stage3_26[11]}
   );
   gpc1_1 gpc1358 (
      {stage2_28[20]},
      {stage3_28[13]}
   );
   gpc1_1 gpc1359 (
      {stage2_28[21]},
      {stage3_28[14]}
   );
   gpc1_1 gpc1360 (
      {stage2_28[22]},
      {stage3_28[15]}
   );
   gpc1_1 gpc1361 (
      {stage2_28[23]},
      {stage3_28[16]}
   );
   gpc1_1 gpc1362 (
      {stage2_28[24]},
      {stage3_28[17]}
   );
   gpc1_1 gpc1363 (
      {stage2_28[25]},
      {stage3_28[18]}
   );
   gpc1_1 gpc1364 (
      {stage2_28[26]},
      {stage3_28[19]}
   );
   gpc1_1 gpc1365 (
      {stage2_28[27]},
      {stage3_28[20]}
   );
   gpc1_1 gpc1366 (
      {stage2_28[28]},
      {stage3_28[21]}
   );
   gpc1_1 gpc1367 (
      {stage2_28[29]},
      {stage3_28[22]}
   );
   gpc1_1 gpc1368 (
      {stage2_31[35]},
      {stage3_31[16]}
   );
   gpc1_1 gpc1369 (
      {stage2_32[37]},
      {stage3_32[12]}
   );
   gpc1_1 gpc1370 (
      {stage2_32[38]},
      {stage3_32[13]}
   );
   gpc1_1 gpc1371 (
      {stage2_32[39]},
      {stage3_32[14]}
   );
   gpc1_1 gpc1372 (
      {stage2_32[40]},
      {stage3_32[15]}
   );
   gpc1_1 gpc1373 (
      {stage2_33[18]},
      {stage3_33[11]}
   );
   gpc1_1 gpc1374 (
      {stage2_33[19]},
      {stage3_33[12]}
   );
   gpc1_1 gpc1375 (
      {stage2_33[20]},
      {stage3_33[13]}
   );
   gpc1_1 gpc1376 (
      {stage2_33[21]},
      {stage3_33[14]}
   );
   gpc1_1 gpc1377 (
      {stage2_33[22]},
      {stage3_33[15]}
   );
   gpc1_1 gpc1378 (
      {stage2_33[23]},
      {stage3_33[16]}
   );
   gpc1_1 gpc1379 (
      {stage2_34[0]},
      {stage3_34[9]}
   );
   gpc1_1 gpc1380 (
      {stage2_34[1]},
      {stage3_34[10]}
   );
   gpc1_1 gpc1381 (
      {stage2_34[2]},
      {stage3_34[11]}
   );
   gpc1_1 gpc1382 (
      {stage2_34[3]},
      {stage3_34[12]}
   );
   gpc1_1 gpc1383 (
      {stage2_34[4]},
      {stage3_34[13]}
   );
   gpc1_1 gpc1384 (
      {stage2_34[5]},
      {stage3_34[14]}
   );
   gpc1_1 gpc1385 (
      {stage2_34[6]},
      {stage3_34[15]}
   );
   gpc1_1 gpc1386 (
      {stage2_35[0]},
      {stage3_35[3]}
   );
   gpc1_1 gpc1387 (
      {stage2_35[1]},
      {stage3_35[4]}
   );
   gpc606_5 gpc1388 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc606_5 gpc1389 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc615_5 gpc1390 (
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10]},
      {stage3_4[0]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[0],stage4_5[1],stage4_4[2],stage4_3[2]}
   );
   gpc615_5 gpc1391 (
      {stage3_3[11], stage3_3[12], stage3_3[13], stage3_3[14], stage3_3[15]},
      {stage3_4[1]},
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage4_7[1],stage4_6[1],stage4_5[2],stage4_4[3],stage4_3[3]}
   );
   gpc606_5 gpc1392 (
      {stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5], stage3_4[6], stage3_4[7]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[2],stage4_6[2],stage4_5[3],stage4_4[4]}
   );
   gpc615_5 gpc1393 (
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10]},
      {stage3_7[0]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[1],stage4_7[3],stage4_6[3]}
   );
   gpc615_5 gpc1394 (
      {stage3_6[11], stage3_6[12], stage3_6[13], stage3_6[14], stage3_6[15]},
      {stage3_7[1]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[1],stage4_8[2],stage4_7[4],stage4_6[4]}
   );
   gpc1406_5 gpc1395 (
      {stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5], stage3_7[6], stage3_7[7]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3]},
      {stage3_10[0]},
      {stage4_11[0],stage4_10[2],stage4_9[2],stage4_8[3],stage4_7[5]}
   );
   gpc606_5 gpc1396 (
      {stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11], stage3_7[12], stage3_7[13]},
      {stage3_9[4], stage3_9[5], stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9]},
      {stage4_11[1],stage4_10[3],stage4_9[3],stage4_8[4],stage4_7[6]}
   );
   gpc615_5 gpc1397 (
      {stage3_7[14], stage3_7[15], stage3_7[16], stage3_7[17], stage3_7[18]},
      {stage3_8[12]},
      {stage3_9[10], stage3_9[11], stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15]},
      {stage4_11[2],stage4_10[4],stage4_9[4],stage4_8[5],stage4_7[7]}
   );
   gpc615_5 gpc1398 (
      {stage3_8[13], stage3_8[14], stage3_8[15], stage3_8[16], stage3_8[17]},
      {stage3_9[16]},
      {stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5], stage3_10[6]},
      {stage4_12[0],stage4_11[3],stage4_10[5],stage4_9[5],stage4_8[6]}
   );
   gpc7_3 gpc1399 (
      {stage3_10[7], stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11], stage3_10[12], stage3_10[13]},
      {stage4_12[1],stage4_11[4],stage4_10[6]}
   );
   gpc606_5 gpc1400 (
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage4_15[0],stage4_14[0],stage4_13[0],stage4_12[2],stage4_11[5]}
   );
   gpc606_5 gpc1401 (
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11]},
      {stage4_15[1],stage4_14[1],stage4_13[1],stage4_12[3],stage4_11[6]}
   );
   gpc606_5 gpc1402 (
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[2],stage4_14[2],stage4_13[2],stage4_12[4]}
   );
   gpc606_5 gpc1403 (
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10], stage3_14[11]},
      {stage4_16[1],stage4_15[3],stage4_14[3],stage4_13[3],stage4_12[5]}
   );
   gpc606_5 gpc1404 (
      {stage3_13[12], stage3_13[13], stage3_13[14], stage3_13[15], stage3_13[16], stage3_13[17]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[2],stage4_15[4],stage4_14[4],stage4_13[4]}
   );
   gpc615_5 gpc1405 (
      {stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15], stage3_14[16]},
      {stage3_15[6]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[1],stage4_16[3],stage4_15[5],stage4_14[5]}
   );
   gpc606_5 gpc1406 (
      {stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11], stage3_15[12]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage4_19[0],stage4_18[1],stage4_17[2],stage4_16[4],stage4_15[6]}
   );
   gpc606_5 gpc1407 (
      {stage3_16[6], stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[1],stage4_18[2],stage4_17[3],stage4_16[5]}
   );
   gpc1163_5 gpc1408 (
      {stage3_17[6], stage3_17[7], stage3_17[8]},
      {stage3_18[6], stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11]},
      {stage3_19[0]},
      {stage3_20[0]},
      {stage4_21[0],stage4_20[1],stage4_19[2],stage4_18[3],stage4_17[4]}
   );
   gpc1343_5 gpc1409 (
      {stage3_19[1], stage3_19[2], stage3_19[3]},
      {stage3_20[1], stage3_20[2], stage3_20[3], stage3_20[4]},
      {stage3_21[0], stage3_21[1], stage3_21[2]},
      {stage3_22[0]},
      {stage4_23[0],stage4_22[0],stage4_21[1],stage4_20[2],stage4_19[3]}
   );
   gpc606_5 gpc1410 (
      {stage3_20[5], stage3_20[6], stage3_20[7], stage3_20[8], stage3_20[9], stage3_20[10]},
      {stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5], stage3_22[6]},
      {stage4_24[0],stage4_23[1],stage4_22[1],stage4_21[2],stage4_20[3]}
   );
   gpc606_5 gpc1411 (
      {stage3_20[11], stage3_20[12], stage3_20[13], stage3_20[14], stage3_20[15], stage3_20[16]},
      {stage3_22[7], stage3_22[8], stage3_22[9], stage3_22[10], stage3_22[11], stage3_22[12]},
      {stage4_24[1],stage4_23[2],stage4_22[2],stage4_21[3],stage4_20[4]}
   );
   gpc606_5 gpc1412 (
      {stage3_21[3], stage3_21[4], stage3_21[5], stage3_21[6], stage3_21[7], stage3_21[8]},
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5]},
      {stage4_25[0],stage4_24[2],stage4_23[3],stage4_22[3],stage4_21[4]}
   );
   gpc606_5 gpc1413 (
      {stage3_21[9], stage3_21[10], stage3_21[11], stage3_21[12], stage3_21[13], stage3_21[14]},
      {stage3_23[6], stage3_23[7], stage3_23[8], stage3_23[9], stage3_23[10], stage3_23[11]},
      {stage4_25[1],stage4_24[3],stage4_23[4],stage4_22[4],stage4_21[5]}
   );
   gpc207_4 gpc1414 (
      {stage3_22[13], stage3_22[14], stage3_22[15], stage3_22[16], stage3_22[17], stage3_22[18], stage3_22[19]},
      {stage3_24[0], stage3_24[1]},
      {stage4_25[2],stage4_24[4],stage4_23[5],stage4_22[5]}
   );
   gpc2135_5 gpc1415 (
      {stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5], stage3_24[6]},
      {stage3_25[0], stage3_25[1], stage3_25[2]},
      {stage3_26[0]},
      {stage3_27[0], stage3_27[1]},
      {stage4_28[0],stage4_27[0],stage4_26[0],stage4_25[3],stage4_24[5]}
   );
   gpc2135_5 gpc1416 (
      {stage3_24[7], stage3_24[8], stage3_24[9], stage3_24[10], stage3_24[11]},
      {stage3_25[3], stage3_25[4], stage3_25[5]},
      {stage3_26[1]},
      {stage3_27[2], stage3_27[3]},
      {stage4_28[1],stage4_27[1],stage4_26[1],stage4_25[4],stage4_24[6]}
   );
   gpc2135_5 gpc1417 (
      {stage3_24[12], stage3_24[13], stage3_24[14], stage3_24[15], stage3_24[16]},
      {stage3_25[6], stage3_25[7], stage3_25[8]},
      {stage3_26[2]},
      {stage3_27[4], stage3_27[5]},
      {stage4_28[2],stage4_27[2],stage4_26[2],stage4_25[5],stage4_24[7]}
   );
   gpc606_5 gpc1418 (
      {stage3_25[9], stage3_25[10], stage3_25[11], stage3_25[12], stage3_25[13], stage3_25[14]},
      {stage3_27[6], stage3_27[7], stage3_27[8], stage3_27[9], stage3_27[10], stage3_27[11]},
      {stage4_29[0],stage4_28[3],stage4_27[3],stage4_26[3],stage4_25[6]}
   );
   gpc615_5 gpc1419 (
      {stage3_26[3], stage3_26[4], stage3_26[5], stage3_26[6], stage3_26[7]},
      {stage3_27[12]},
      {stage3_28[0], stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4], stage3_28[5]},
      {stage4_30[0],stage4_29[1],stage4_28[4],stage4_27[4],stage4_26[4]}
   );
   gpc2135_5 gpc1420 (
      {stage3_28[6], stage3_28[7], stage3_28[8], stage3_28[9], stage3_28[10]},
      {stage3_29[0], stage3_29[1], stage3_29[2]},
      {stage3_30[0]},
      {stage3_31[0], stage3_31[1]},
      {stage4_32[0],stage4_31[0],stage4_30[1],stage4_29[2],stage4_28[5]}
   );
   gpc2135_5 gpc1421 (
      {stage3_28[11], stage3_28[12], stage3_28[13], stage3_28[14], stage3_28[15]},
      {stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage3_30[1]},
      {stage3_31[2], stage3_31[3]},
      {stage4_32[1],stage4_31[1],stage4_30[2],stage4_29[3],stage4_28[6]}
   );
   gpc606_5 gpc1422 (
      {stage3_28[16], stage3_28[17], stage3_28[18], stage3_28[19], stage3_28[20], stage3_28[21]},
      {stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5], stage3_30[6], stage3_30[7]},
      {stage4_32[2],stage4_31[2],stage4_30[3],stage4_29[4],stage4_28[7]}
   );
   gpc615_5 gpc1423 (
      {stage3_29[6], stage3_29[7], stage3_29[8], stage3_29[9], stage3_29[10]},
      {stage3_30[8]},
      {stage3_31[4], stage3_31[5], stage3_31[6], stage3_31[7], stage3_31[8], stage3_31[9]},
      {stage4_33[0],stage4_32[3],stage4_31[3],stage4_30[4],stage4_29[5]}
   );
   gpc615_5 gpc1424 (
      {stage3_30[9], stage3_30[10], stage3_30[11], stage3_30[12], stage3_30[13]},
      {stage3_31[10]},
      {stage3_32[0], stage3_32[1], stage3_32[2], stage3_32[3], stage3_32[4], stage3_32[5]},
      {stage4_34[0],stage4_33[1],stage4_32[4],stage4_31[4],stage4_30[5]}
   );
   gpc606_5 gpc1425 (
      {stage3_31[11], stage3_31[12], stage3_31[13], stage3_31[14], stage3_31[15], stage3_31[16]},
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4], stage3_33[5]},
      {stage4_35[0],stage4_34[1],stage4_33[2],stage4_32[5],stage4_31[5]}
   );
   gpc606_5 gpc1426 (
      {stage3_32[6], stage3_32[7], stage3_32[8], stage3_32[9], stage3_32[10], stage3_32[11]},
      {stage3_34[0], stage3_34[1], stage3_34[2], stage3_34[3], stage3_34[4], stage3_34[5]},
      {stage4_36[0],stage4_35[1],stage4_34[2],stage4_33[3],stage4_32[6]}
   );
   gpc1163_5 gpc1427 (
      {stage3_33[6], stage3_33[7], stage3_33[8]},
      {stage3_34[6], stage3_34[7], stage3_34[8], stage3_34[9], stage3_34[10], stage3_34[11]},
      {stage3_35[0]},
      {1'b0},
      {stage4_37[0],stage4_36[1],stage4_35[2],stage4_34[3],stage4_33[4]}
   );
   gpc606_5 gpc1428 (
      {stage3_33[9], stage3_33[10], stage3_33[11], stage3_33[12], stage3_33[13], stage3_33[14]},
      {stage3_35[1], stage3_35[2], stage3_35[3], stage3_35[4], 1'b0, 1'b0},
      {stage4_37[1],stage4_36[2],stage4_35[3],stage4_34[4],stage4_33[5]}
   );
   gpc1_1 gpc1429 (
      {stage3_0[6]},
      {stage4_0[1]}
   );
   gpc1_1 gpc1430 (
      {stage3_1[6]},
      {stage4_1[2]}
   );
   gpc1_1 gpc1431 (
      {stage3_1[7]},
      {stage4_1[3]}
   );
   gpc1_1 gpc1432 (
      {stage3_1[8]},
      {stage4_1[4]}
   );
   gpc1_1 gpc1433 (
      {stage3_1[9]},
      {stage4_1[5]}
   );
   gpc1_1 gpc1434 (
      {stage3_2[6]},
      {stage4_2[2]}
   );
   gpc1_1 gpc1435 (
      {stage3_2[7]},
      {stage4_2[3]}
   );
   gpc1_1 gpc1436 (
      {stage3_2[8]},
      {stage4_2[4]}
   );
   gpc1_1 gpc1437 (
      {stage3_2[9]},
      {stage4_2[5]}
   );
   gpc1_1 gpc1438 (
      {stage3_3[16]},
      {stage4_3[4]}
   );
   gpc1_1 gpc1439 (
      {stage3_3[17]},
      {stage4_3[5]}
   );
   gpc1_1 gpc1440 (
      {stage3_3[18]},
      {stage4_3[6]}
   );
   gpc1_1 gpc1441 (
      {stage3_3[19]},
      {stage4_3[7]}
   );
   gpc1_1 gpc1442 (
      {stage3_3[20]},
      {stage4_3[8]}
   );
   gpc1_1 gpc1443 (
      {stage3_3[21]},
      {stage4_3[9]}
   );
   gpc1_1 gpc1444 (
      {stage3_3[22]},
      {stage4_3[10]}
   );
   gpc1_1 gpc1445 (
      {stage3_4[8]},
      {stage4_4[5]}
   );
   gpc1_1 gpc1446 (
      {stage3_6[16]},
      {stage4_6[5]}
   );
   gpc1_1 gpc1447 (
      {stage3_9[17]},
      {stage4_9[6]}
   );
   gpc1_1 gpc1448 (
      {stage3_9[18]},
      {stage4_9[7]}
   );
   gpc1_1 gpc1449 (
      {stage3_10[14]},
      {stage4_10[7]}
   );
   gpc1_1 gpc1450 (
      {stage3_11[12]},
      {stage4_11[7]}
   );
   gpc1_1 gpc1451 (
      {stage3_11[13]},
      {stage4_11[8]}
   );
   gpc1_1 gpc1452 (
      {stage3_11[14]},
      {stage4_11[9]}
   );
   gpc1_1 gpc1453 (
      {stage3_12[12]},
      {stage4_12[6]}
   );
   gpc1_1 gpc1454 (
      {stage3_12[13]},
      {stage4_12[7]}
   );
   gpc1_1 gpc1455 (
      {stage3_12[14]},
      {stage4_12[8]}
   );
   gpc1_1 gpc1456 (
      {stage3_15[13]},
      {stage4_15[7]}
   );
   gpc1_1 gpc1457 (
      {stage3_15[14]},
      {stage4_15[8]}
   );
   gpc1_1 gpc1458 (
      {stage3_15[15]},
      {stage4_15[9]}
   );
   gpc1_1 gpc1459 (
      {stage3_16[12]},
      {stage4_16[6]}
   );
   gpc1_1 gpc1460 (
      {stage3_17[9]},
      {stage4_17[5]}
   );
   gpc1_1 gpc1461 (
      {stage3_17[10]},
      {stage4_17[6]}
   );
   gpc1_1 gpc1462 (
      {stage3_17[11]},
      {stage4_17[7]}
   );
   gpc1_1 gpc1463 (
      {stage3_17[12]},
      {stage4_17[8]}
   );
   gpc1_1 gpc1464 (
      {stage3_17[13]},
      {stage4_17[9]}
   );
   gpc1_1 gpc1465 (
      {stage3_17[14]},
      {stage4_17[10]}
   );
   gpc1_1 gpc1466 (
      {stage3_17[15]},
      {stage4_17[11]}
   );
   gpc1_1 gpc1467 (
      {stage3_17[16]},
      {stage4_17[12]}
   );
   gpc1_1 gpc1468 (
      {stage3_18[12]},
      {stage4_18[4]}
   );
   gpc1_1 gpc1469 (
      {stage3_18[13]},
      {stage4_18[5]}
   );
   gpc1_1 gpc1470 (
      {stage3_18[14]},
      {stage4_18[6]}
   );
   gpc1_1 gpc1471 (
      {stage3_18[15]},
      {stage4_18[7]}
   );
   gpc1_1 gpc1472 (
      {stage3_18[16]},
      {stage4_18[8]}
   );
   gpc1_1 gpc1473 (
      {stage3_19[4]},
      {stage4_19[4]}
   );
   gpc1_1 gpc1474 (
      {stage3_19[5]},
      {stage4_19[5]}
   );
   gpc1_1 gpc1475 (
      {stage3_19[6]},
      {stage4_19[6]}
   );
   gpc1_1 gpc1476 (
      {stage3_19[7]},
      {stage4_19[7]}
   );
   gpc1_1 gpc1477 (
      {stage3_19[8]},
      {stage4_19[8]}
   );
   gpc1_1 gpc1478 (
      {stage3_19[9]},
      {stage4_19[9]}
   );
   gpc1_1 gpc1479 (
      {stage3_19[10]},
      {stage4_19[10]}
   );
   gpc1_1 gpc1480 (
      {stage3_19[11]},
      {stage4_19[11]}
   );
   gpc1_1 gpc1481 (
      {stage3_20[17]},
      {stage4_20[5]}
   );
   gpc1_1 gpc1482 (
      {stage3_22[20]},
      {stage4_22[6]}
   );
   gpc1_1 gpc1483 (
      {stage3_22[21]},
      {stage4_22[7]}
   );
   gpc1_1 gpc1484 (
      {stage3_22[22]},
      {stage4_22[8]}
   );
   gpc1_1 gpc1485 (
      {stage3_23[12]},
      {stage4_23[6]}
   );
   gpc1_1 gpc1486 (
      {stage3_25[15]},
      {stage4_25[7]}
   );
   gpc1_1 gpc1487 (
      {stage3_25[16]},
      {stage4_25[8]}
   );
   gpc1_1 gpc1488 (
      {stage3_26[8]},
      {stage4_26[5]}
   );
   gpc1_1 gpc1489 (
      {stage3_26[9]},
      {stage4_26[6]}
   );
   gpc1_1 gpc1490 (
      {stage3_26[10]},
      {stage4_26[7]}
   );
   gpc1_1 gpc1491 (
      {stage3_26[11]},
      {stage4_26[8]}
   );
   gpc1_1 gpc1492 (
      {stage3_28[22]},
      {stage4_28[8]}
   );
   gpc1_1 gpc1493 (
      {stage3_32[12]},
      {stage4_32[7]}
   );
   gpc1_1 gpc1494 (
      {stage3_32[13]},
      {stage4_32[8]}
   );
   gpc1_1 gpc1495 (
      {stage3_32[14]},
      {stage4_32[9]}
   );
   gpc1_1 gpc1496 (
      {stage3_32[15]},
      {stage4_32[10]}
   );
   gpc1_1 gpc1497 (
      {stage3_33[15]},
      {stage4_33[6]}
   );
   gpc1_1 gpc1498 (
      {stage3_33[16]},
      {stage4_33[7]}
   );
   gpc1_1 gpc1499 (
      {stage3_34[12]},
      {stage4_34[5]}
   );
   gpc1_1 gpc1500 (
      {stage3_34[13]},
      {stage4_34[6]}
   );
   gpc1_1 gpc1501 (
      {stage3_34[14]},
      {stage4_34[7]}
   );
   gpc1_1 gpc1502 (
      {stage3_34[15]},
      {stage4_34[8]}
   );
   gpc623_5 gpc1503 (
      {stage4_1[0], stage4_1[1], stage4_1[2]},
      {stage4_2[0], stage4_2[1]},
      {stage4_3[0], stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5]},
      {stage5_5[0],stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0]}
   );
   gpc1163_5 gpc1504 (
      {stage4_3[6], stage4_3[7], stage4_3[8]},
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5]},
      {stage4_5[0]},
      {stage4_6[0]},
      {stage5_7[0],stage5_6[0],stage5_5[1],stage5_4[1],stage5_3[1]}
   );
   gpc1415_5 gpc1505 (
      {stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage4_7[0]},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3]},
      {stage4_9[0]},
      {stage5_10[0],stage5_9[0],stage5_8[0],stage5_7[1],stage5_6[1]}
   );
   gpc223_4 gpc1506 (
      {stage4_7[1], stage4_7[2], stage4_7[3]},
      {stage4_8[4], stage4_8[5]},
      {stage4_9[1], stage4_9[2]},
      {stage5_10[1],stage5_9[1],stage5_8[1],stage5_7[2]}
   );
   gpc2135_5 gpc1507 (
      {stage4_9[3], stage4_9[4], stage4_9[5], stage4_9[6], stage4_9[7]},
      {stage4_10[0], stage4_10[1], stage4_10[2]},
      {stage4_11[0]},
      {stage4_12[0], stage4_12[1]},
      {stage5_13[0],stage5_12[0],stage5_11[0],stage5_10[2],stage5_9[2]}
   );
   gpc615_5 gpc1508 (
      {stage4_10[3], stage4_10[4], stage4_10[5], stage4_10[6], stage4_10[7]},
      {stage4_11[1]},
      {stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5], stage4_12[6], stage4_12[7]},
      {stage5_14[0],stage5_13[1],stage5_12[1],stage5_11[1],stage5_10[3]}
   );
   gpc615_5 gpc1509 (
      {stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5], stage4_11[6]},
      {stage4_12[8]},
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3], stage4_13[4], 1'b0},
      {stage5_15[0],stage5_14[1],stage5_13[2],stage5_12[2],stage5_11[2]}
   );
   gpc1163_5 gpc1510 (
      {stage4_14[0], stage4_14[1], stage4_14[2]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5]},
      {stage4_16[0]},
      {stage4_17[0]},
      {stage5_18[0],stage5_17[0],stage5_16[0],stage5_15[1],stage5_14[2]}
   );
   gpc606_5 gpc1511 (
      {stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5], stage4_16[6]},
      {stage4_18[0], stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5]},
      {stage5_20[0],stage5_19[0],stage5_18[1],stage5_17[1],stage5_16[1]}
   );
   gpc615_5 gpc1512 (
      {stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage4_18[6]},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage5_21[0],stage5_20[1],stage5_19[1],stage5_18[2],stage5_17[2]}
   );
   gpc615_5 gpc1513 (
      {stage4_17[6], stage4_17[7], stage4_17[8], stage4_17[9], stage4_17[10]},
      {stage4_18[7]},
      {stage4_19[6], stage4_19[7], stage4_19[8], stage4_19[9], stage4_19[10], stage4_19[11]},
      {stage5_21[1],stage5_20[2],stage5_19[2],stage5_18[3],stage5_17[3]}
   );
   gpc606_5 gpc1514 (
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], stage4_20[4], stage4_20[5]},
      {stage4_22[0], stage4_22[1], stage4_22[2], stage4_22[3], stage4_22[4], stage4_22[5]},
      {stage5_24[0],stage5_23[0],stage5_22[0],stage5_21[2],stage5_20[3]}
   );
   gpc135_4 gpc1515 (
      {stage4_21[0], stage4_21[1], stage4_21[2], stage4_21[3], stage4_21[4]},
      {stage4_22[6], stage4_22[7], stage4_22[8]},
      {stage4_23[0]},
      {stage5_24[1],stage5_23[1],stage5_22[1],stage5_21[3]}
   );
   gpc615_5 gpc1516 (
      {stage4_23[1], stage4_23[2], stage4_23[3], stage4_23[4], stage4_23[5]},
      {stage4_24[0]},
      {stage4_25[0], stage4_25[1], stage4_25[2], stage4_25[3], stage4_25[4], stage4_25[5]},
      {stage5_27[0],stage5_26[0],stage5_25[0],stage5_24[2],stage5_23[2]}
   );
   gpc2135_5 gpc1517 (
      {stage4_24[1], stage4_24[2], stage4_24[3], stage4_24[4], stage4_24[5]},
      {stage4_25[6], stage4_25[7], stage4_25[8]},
      {stage4_26[0]},
      {stage4_27[0], stage4_27[1]},
      {stage5_28[0],stage5_27[1],stage5_26[1],stage5_25[1],stage5_24[3]}
   );
   gpc2223_5 gpc1518 (
      {stage4_26[1], stage4_26[2], stage4_26[3]},
      {stage4_27[2], stage4_27[3]},
      {stage4_28[0], stage4_28[1]},
      {stage4_29[0], stage4_29[1]},
      {stage5_30[0],stage5_29[0],stage5_28[1],stage5_27[2],stage5_26[2]}
   );
   gpc615_5 gpc1519 (
      {stage4_26[4], stage4_26[5], stage4_26[6], stage4_26[7], stage4_26[8]},
      {stage4_27[4]},
      {stage4_28[2], stage4_28[3], stage4_28[4], stage4_28[5], stage4_28[6], stage4_28[7]},
      {stage5_30[1],stage5_29[1],stage5_28[2],stage5_27[3],stage5_26[3]}
   );
   gpc606_5 gpc1520 (
      {stage4_30[0], stage4_30[1], stage4_30[2], stage4_30[3], stage4_30[4], stage4_30[5]},
      {stage4_32[0], stage4_32[1], stage4_32[2], stage4_32[3], stage4_32[4], stage4_32[5]},
      {stage5_34[0],stage5_33[0],stage5_32[0],stage5_31[0],stage5_30[2]}
   );
   gpc606_5 gpc1521 (
      {stage4_31[0], stage4_31[1], stage4_31[2], stage4_31[3], stage4_31[4], stage4_31[5]},
      {stage4_33[0], stage4_33[1], stage4_33[2], stage4_33[3], stage4_33[4], stage4_33[5]},
      {stage5_35[0],stage5_34[1],stage5_33[1],stage5_32[1],stage5_31[1]}
   );
   gpc606_5 gpc1522 (
      {stage4_32[6], stage4_32[7], stage4_32[8], stage4_32[9], stage4_32[10], 1'b0},
      {stage4_34[0], stage4_34[1], stage4_34[2], stage4_34[3], stage4_34[4], stage4_34[5]},
      {stage5_36[0],stage5_35[1],stage5_34[2],stage5_33[2],stage5_32[2]}
   );
   gpc2116_5 gpc1523 (
      {stage4_34[6], stage4_34[7], stage4_34[8], 1'b0, 1'b0, 1'b0},
      {stage4_35[0]},
      {stage4_36[0]},
      {stage4_37[0], stage4_37[1]},
      {stage5_38[0],stage5_37[0],stage5_36[1],stage5_35[2],stage5_34[3]}
   );
   gpc1_1 gpc1524 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc1525 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc1526 (
      {stage4_1[3]},
      {stage5_1[1]}
   );
   gpc1_1 gpc1527 (
      {stage4_1[4]},
      {stage5_1[2]}
   );
   gpc1_1 gpc1528 (
      {stage4_1[5]},
      {stage5_1[3]}
   );
   gpc1_1 gpc1529 (
      {stage4_2[2]},
      {stage5_2[1]}
   );
   gpc1_1 gpc1530 (
      {stage4_2[3]},
      {stage5_2[2]}
   );
   gpc1_1 gpc1531 (
      {stage4_2[4]},
      {stage5_2[3]}
   );
   gpc1_1 gpc1532 (
      {stage4_2[5]},
      {stage5_2[4]}
   );
   gpc1_1 gpc1533 (
      {stage4_3[9]},
      {stage5_3[2]}
   );
   gpc1_1 gpc1534 (
      {stage4_3[10]},
      {stage5_3[3]}
   );
   gpc1_1 gpc1535 (
      {stage4_5[1]},
      {stage5_5[2]}
   );
   gpc1_1 gpc1536 (
      {stage4_5[2]},
      {stage5_5[3]}
   );
   gpc1_1 gpc1537 (
      {stage4_5[3]},
      {stage5_5[4]}
   );
   gpc1_1 gpc1538 (
      {stage4_7[4]},
      {stage5_7[3]}
   );
   gpc1_1 gpc1539 (
      {stage4_7[5]},
      {stage5_7[4]}
   );
   gpc1_1 gpc1540 (
      {stage4_7[6]},
      {stage5_7[5]}
   );
   gpc1_1 gpc1541 (
      {stage4_7[7]},
      {stage5_7[6]}
   );
   gpc1_1 gpc1542 (
      {stage4_8[6]},
      {stage5_8[2]}
   );
   gpc1_1 gpc1543 (
      {stage4_11[7]},
      {stage5_11[3]}
   );
   gpc1_1 gpc1544 (
      {stage4_11[8]},
      {stage5_11[4]}
   );
   gpc1_1 gpc1545 (
      {stage4_11[9]},
      {stage5_11[5]}
   );
   gpc1_1 gpc1546 (
      {stage4_14[3]},
      {stage5_14[3]}
   );
   gpc1_1 gpc1547 (
      {stage4_14[4]},
      {stage5_14[4]}
   );
   gpc1_1 gpc1548 (
      {stage4_14[5]},
      {stage5_14[5]}
   );
   gpc1_1 gpc1549 (
      {stage4_15[6]},
      {stage5_15[2]}
   );
   gpc1_1 gpc1550 (
      {stage4_15[7]},
      {stage5_15[3]}
   );
   gpc1_1 gpc1551 (
      {stage4_15[8]},
      {stage5_15[4]}
   );
   gpc1_1 gpc1552 (
      {stage4_15[9]},
      {stage5_15[5]}
   );
   gpc1_1 gpc1553 (
      {stage4_17[11]},
      {stage5_17[4]}
   );
   gpc1_1 gpc1554 (
      {stage4_17[12]},
      {stage5_17[5]}
   );
   gpc1_1 gpc1555 (
      {stage4_18[8]},
      {stage5_18[4]}
   );
   gpc1_1 gpc1556 (
      {stage4_21[5]},
      {stage5_21[4]}
   );
   gpc1_1 gpc1557 (
      {stage4_23[6]},
      {stage5_23[3]}
   );
   gpc1_1 gpc1558 (
      {stage4_24[6]},
      {stage5_24[4]}
   );
   gpc1_1 gpc1559 (
      {stage4_24[7]},
      {stage5_24[5]}
   );
   gpc1_1 gpc1560 (
      {stage4_28[8]},
      {stage5_28[3]}
   );
   gpc1_1 gpc1561 (
      {stage4_29[2]},
      {stage5_29[2]}
   );
   gpc1_1 gpc1562 (
      {stage4_29[3]},
      {stage5_29[3]}
   );
   gpc1_1 gpc1563 (
      {stage4_29[4]},
      {stage5_29[4]}
   );
   gpc1_1 gpc1564 (
      {stage4_29[5]},
      {stage5_29[5]}
   );
   gpc1_1 gpc1565 (
      {stage4_33[6]},
      {stage5_33[3]}
   );
   gpc1_1 gpc1566 (
      {stage4_33[7]},
      {stage5_33[4]}
   );
   gpc1_1 gpc1567 (
      {stage4_35[1]},
      {stage5_35[3]}
   );
   gpc1_1 gpc1568 (
      {stage4_35[2]},
      {stage5_35[4]}
   );
   gpc1_1 gpc1569 (
      {stage4_35[3]},
      {stage5_35[5]}
   );
   gpc1_1 gpc1570 (
      {stage4_36[1]},
      {stage5_36[2]}
   );
   gpc1_1 gpc1571 (
      {stage4_36[2]},
      {stage5_36[3]}
   );
   gpc1343_5 gpc1572 (
      {stage5_1[0], stage5_1[1], stage5_1[2]},
      {stage5_2[0], stage5_2[1], stage5_2[2], stage5_2[3]},
      {stage5_3[0], stage5_3[1], stage5_3[2]},
      {stage5_4[0]},
      {stage6_5[0],stage6_4[0],stage6_3[0],stage6_2[0],stage6_1[0]}
   );
   gpc615_5 gpc1573 (
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4]},
      {stage5_6[0]},
      {stage5_7[0], stage5_7[1], stage5_7[2], stage5_7[3], stage5_7[4], stage5_7[5]},
      {stage6_9[0],stage6_8[0],stage6_7[0],stage6_6[0],stage6_5[1]}
   );
   gpc1343_5 gpc1574 (
      {stage5_8[0], stage5_8[1], stage5_8[2]},
      {stage5_9[0], stage5_9[1], stage5_9[2], 1'b0},
      {stage5_10[0], stage5_10[1], stage5_10[2]},
      {stage5_11[0]},
      {stage6_12[0],stage6_11[0],stage6_10[0],stage6_9[1],stage6_8[1]}
   );
   gpc135_4 gpc1575 (
      {stage5_11[1], stage5_11[2], stage5_11[3], stage5_11[4], stage5_11[5]},
      {stage5_12[0], stage5_12[1], stage5_12[2]},
      {stage5_13[0]},
      {stage6_14[0],stage6_13[0],stage6_12[1],stage6_11[1]}
   );
   gpc1163_5 gpc1576 (
      {stage5_13[1], stage5_13[2], 1'b0},
      {stage5_14[0], stage5_14[1], stage5_14[2], stage5_14[3], stage5_14[4], stage5_14[5]},
      {stage5_15[0]},
      {stage5_16[0]},
      {stage6_17[0],stage6_16[0],stage6_15[0],stage6_14[1],stage6_13[1]}
   );
   gpc615_5 gpc1577 (
      {stage5_15[1], stage5_15[2], stage5_15[3], stage5_15[4], stage5_15[5]},
      {stage5_16[1]},
      {stage5_17[0], stage5_17[1], stage5_17[2], stage5_17[3], stage5_17[4], stage5_17[5]},
      {stage6_19[0],stage6_18[0],stage6_17[1],stage6_16[1],stage6_15[1]}
   );
   gpc135_4 gpc1578 (
      {stage5_18[0], stage5_18[1], stage5_18[2], stage5_18[3], stage5_18[4]},
      {stage5_19[0], stage5_19[1], stage5_19[2]},
      {stage5_20[0]},
      {stage6_21[0],stage6_20[0],stage6_19[1],stage6_18[1]}
   );
   gpc1163_5 gpc1579 (
      {stage5_20[1], stage5_20[2], stage5_20[3]},
      {stage5_21[0], stage5_21[1], stage5_21[2], stage5_21[3], stage5_21[4], 1'b0},
      {stage5_22[0]},
      {stage5_23[0]},
      {stage6_24[0],stage6_23[0],stage6_22[0],stage6_21[1],stage6_20[1]}
   );
   gpc1163_5 gpc1580 (
      {stage5_23[1], stage5_23[2], stage5_23[3]},
      {stage5_24[0], stage5_24[1], stage5_24[2], stage5_24[3], stage5_24[4], stage5_24[5]},
      {stage5_25[0]},
      {stage5_26[0]},
      {stage6_27[0],stage6_26[0],stage6_25[0],stage6_24[1],stage6_23[1]}
   );
   gpc1343_5 gpc1581 (
      {stage5_26[1], stage5_26[2], stage5_26[3]},
      {stage5_27[0], stage5_27[1], stage5_27[2], stage5_27[3]},
      {stage5_28[0], stage5_28[1], stage5_28[2]},
      {stage5_29[0]},
      {stage6_30[0],stage6_29[0],stage6_28[0],stage6_27[1],stage6_26[1]}
   );
   gpc2135_5 gpc1582 (
      {stage5_29[1], stage5_29[2], stage5_29[3], stage5_29[4], stage5_29[5]},
      {stage5_30[0], stage5_30[1], stage5_30[2]},
      {stage5_31[0]},
      {stage5_32[0], stage5_32[1]},
      {stage6_33[0],stage6_32[0],stage6_31[0],stage6_30[1],stage6_29[1]}
   );
   gpc606_5 gpc1583 (
      {stage5_33[0], stage5_33[1], stage5_33[2], stage5_33[3], stage5_33[4], 1'b0},
      {stage5_35[0], stage5_35[1], stage5_35[2], stage5_35[3], stage5_35[4], stage5_35[5]},
      {stage6_37[0],stage6_36[0],stage6_35[0],stage6_34[0],stage6_33[1]}
   );
   gpc1415_5 gpc1584 (
      {stage5_34[0], stage5_34[1], stage5_34[2], stage5_34[3], 1'b0},
      {1'b0},
      {stage5_36[0], stage5_36[1], stage5_36[2], stage5_36[3]},
      {stage5_37[0]},
      {stage6_38[0],stage6_37[1],stage6_36[1],stage6_35[1],stage6_34[1]}
   );
   gpc1_1 gpc1585 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc1586 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc1587 (
      {stage5_1[3]},
      {stage6_1[1]}
   );
   gpc1_1 gpc1588 (
      {stage5_2[4]},
      {stage6_2[1]}
   );
   gpc1_1 gpc1589 (
      {stage5_3[3]},
      {stage6_3[1]}
   );
   gpc1_1 gpc1590 (
      {stage5_4[1]},
      {stage6_4[1]}
   );
   gpc1_1 gpc1591 (
      {stage5_6[1]},
      {stage6_6[1]}
   );
   gpc1_1 gpc1592 (
      {stage5_7[6]},
      {stage6_7[1]}
   );
   gpc1_1 gpc1593 (
      {stage5_10[3]},
      {stage6_10[1]}
   );
   gpc1_1 gpc1594 (
      {stage5_22[1]},
      {stage6_22[1]}
   );
   gpc1_1 gpc1595 (
      {stage5_25[1]},
      {stage6_25[1]}
   );
   gpc1_1 gpc1596 (
      {stage5_28[3]},
      {stage6_28[1]}
   );
   gpc1_1 gpc1597 (
      {stage5_31[1]},
      {stage6_31[1]}
   );
   gpc1_1 gpc1598 (
      {stage5_32[2]},
      {stage6_32[1]}
   );
   gpc1_1 gpc1599 (
      {stage5_38[0]},
      {stage6_38[1]}
   );
endmodule

module testbench();
    reg [161:0] src0;
    reg [161:0] src1;
    reg [161:0] src2;
    reg [161:0] src3;
    reg [161:0] src4;
    reg [161:0] src5;
    reg [161:0] src6;
    reg [161:0] src7;
    reg [161:0] src8;
    reg [161:0] src9;
    reg [161:0] src10;
    reg [161:0] src11;
    reg [161:0] src12;
    reg [161:0] src13;
    reg [161:0] src14;
    reg [161:0] src15;
    reg [161:0] src16;
    reg [161:0] src17;
    reg [161:0] src18;
    reg [161:0] src19;
    reg [161:0] src20;
    reg [161:0] src21;
    reg [161:0] src22;
    reg [161:0] src23;
    reg [161:0] src24;
    reg [161:0] src25;
    reg [161:0] src26;
    reg [161:0] src27;
    reg [161:0] src28;
    reg [161:0] src29;
    reg [161:0] src30;
    reg [161:0] src31;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [39:0] srcsum;
    wire [39:0] dstsum;
    wire test;
    compressor_CLA162_32 compressor_CLA162_32(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63] + src16[64] + src16[65] + src16[66] + src16[67] + src16[68] + src16[69] + src16[70] + src16[71] + src16[72] + src16[73] + src16[74] + src16[75] + src16[76] + src16[77] + src16[78] + src16[79] + src16[80] + src16[81] + src16[82] + src16[83] + src16[84] + src16[85] + src16[86] + src16[87] + src16[88] + src16[89] + src16[90] + src16[91] + src16[92] + src16[93] + src16[94] + src16[95] + src16[96] + src16[97] + src16[98] + src16[99] + src16[100] + src16[101] + src16[102] + src16[103] + src16[104] + src16[105] + src16[106] + src16[107] + src16[108] + src16[109] + src16[110] + src16[111] + src16[112] + src16[113] + src16[114] + src16[115] + src16[116] + src16[117] + src16[118] + src16[119] + src16[120] + src16[121] + src16[122] + src16[123] + src16[124] + src16[125] + src16[126] + src16[127] + src16[128] + src16[129] + src16[130] + src16[131] + src16[132] + src16[133] + src16[134] + src16[135] + src16[136] + src16[137] + src16[138] + src16[139] + src16[140] + src16[141] + src16[142] + src16[143] + src16[144] + src16[145] + src16[146] + src16[147] + src16[148] + src16[149] + src16[150] + src16[151] + src16[152] + src16[153] + src16[154] + src16[155] + src16[156] + src16[157] + src16[158] + src16[159] + src16[160] + src16[161])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63] + src17[64] + src17[65] + src17[66] + src17[67] + src17[68] + src17[69] + src17[70] + src17[71] + src17[72] + src17[73] + src17[74] + src17[75] + src17[76] + src17[77] + src17[78] + src17[79] + src17[80] + src17[81] + src17[82] + src17[83] + src17[84] + src17[85] + src17[86] + src17[87] + src17[88] + src17[89] + src17[90] + src17[91] + src17[92] + src17[93] + src17[94] + src17[95] + src17[96] + src17[97] + src17[98] + src17[99] + src17[100] + src17[101] + src17[102] + src17[103] + src17[104] + src17[105] + src17[106] + src17[107] + src17[108] + src17[109] + src17[110] + src17[111] + src17[112] + src17[113] + src17[114] + src17[115] + src17[116] + src17[117] + src17[118] + src17[119] + src17[120] + src17[121] + src17[122] + src17[123] + src17[124] + src17[125] + src17[126] + src17[127] + src17[128] + src17[129] + src17[130] + src17[131] + src17[132] + src17[133] + src17[134] + src17[135] + src17[136] + src17[137] + src17[138] + src17[139] + src17[140] + src17[141] + src17[142] + src17[143] + src17[144] + src17[145] + src17[146] + src17[147] + src17[148] + src17[149] + src17[150] + src17[151] + src17[152] + src17[153] + src17[154] + src17[155] + src17[156] + src17[157] + src17[158] + src17[159] + src17[160] + src17[161])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63] + src18[64] + src18[65] + src18[66] + src18[67] + src18[68] + src18[69] + src18[70] + src18[71] + src18[72] + src18[73] + src18[74] + src18[75] + src18[76] + src18[77] + src18[78] + src18[79] + src18[80] + src18[81] + src18[82] + src18[83] + src18[84] + src18[85] + src18[86] + src18[87] + src18[88] + src18[89] + src18[90] + src18[91] + src18[92] + src18[93] + src18[94] + src18[95] + src18[96] + src18[97] + src18[98] + src18[99] + src18[100] + src18[101] + src18[102] + src18[103] + src18[104] + src18[105] + src18[106] + src18[107] + src18[108] + src18[109] + src18[110] + src18[111] + src18[112] + src18[113] + src18[114] + src18[115] + src18[116] + src18[117] + src18[118] + src18[119] + src18[120] + src18[121] + src18[122] + src18[123] + src18[124] + src18[125] + src18[126] + src18[127] + src18[128] + src18[129] + src18[130] + src18[131] + src18[132] + src18[133] + src18[134] + src18[135] + src18[136] + src18[137] + src18[138] + src18[139] + src18[140] + src18[141] + src18[142] + src18[143] + src18[144] + src18[145] + src18[146] + src18[147] + src18[148] + src18[149] + src18[150] + src18[151] + src18[152] + src18[153] + src18[154] + src18[155] + src18[156] + src18[157] + src18[158] + src18[159] + src18[160] + src18[161])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63] + src19[64] + src19[65] + src19[66] + src19[67] + src19[68] + src19[69] + src19[70] + src19[71] + src19[72] + src19[73] + src19[74] + src19[75] + src19[76] + src19[77] + src19[78] + src19[79] + src19[80] + src19[81] + src19[82] + src19[83] + src19[84] + src19[85] + src19[86] + src19[87] + src19[88] + src19[89] + src19[90] + src19[91] + src19[92] + src19[93] + src19[94] + src19[95] + src19[96] + src19[97] + src19[98] + src19[99] + src19[100] + src19[101] + src19[102] + src19[103] + src19[104] + src19[105] + src19[106] + src19[107] + src19[108] + src19[109] + src19[110] + src19[111] + src19[112] + src19[113] + src19[114] + src19[115] + src19[116] + src19[117] + src19[118] + src19[119] + src19[120] + src19[121] + src19[122] + src19[123] + src19[124] + src19[125] + src19[126] + src19[127] + src19[128] + src19[129] + src19[130] + src19[131] + src19[132] + src19[133] + src19[134] + src19[135] + src19[136] + src19[137] + src19[138] + src19[139] + src19[140] + src19[141] + src19[142] + src19[143] + src19[144] + src19[145] + src19[146] + src19[147] + src19[148] + src19[149] + src19[150] + src19[151] + src19[152] + src19[153] + src19[154] + src19[155] + src19[156] + src19[157] + src19[158] + src19[159] + src19[160] + src19[161])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63] + src20[64] + src20[65] + src20[66] + src20[67] + src20[68] + src20[69] + src20[70] + src20[71] + src20[72] + src20[73] + src20[74] + src20[75] + src20[76] + src20[77] + src20[78] + src20[79] + src20[80] + src20[81] + src20[82] + src20[83] + src20[84] + src20[85] + src20[86] + src20[87] + src20[88] + src20[89] + src20[90] + src20[91] + src20[92] + src20[93] + src20[94] + src20[95] + src20[96] + src20[97] + src20[98] + src20[99] + src20[100] + src20[101] + src20[102] + src20[103] + src20[104] + src20[105] + src20[106] + src20[107] + src20[108] + src20[109] + src20[110] + src20[111] + src20[112] + src20[113] + src20[114] + src20[115] + src20[116] + src20[117] + src20[118] + src20[119] + src20[120] + src20[121] + src20[122] + src20[123] + src20[124] + src20[125] + src20[126] + src20[127] + src20[128] + src20[129] + src20[130] + src20[131] + src20[132] + src20[133] + src20[134] + src20[135] + src20[136] + src20[137] + src20[138] + src20[139] + src20[140] + src20[141] + src20[142] + src20[143] + src20[144] + src20[145] + src20[146] + src20[147] + src20[148] + src20[149] + src20[150] + src20[151] + src20[152] + src20[153] + src20[154] + src20[155] + src20[156] + src20[157] + src20[158] + src20[159] + src20[160] + src20[161])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63] + src21[64] + src21[65] + src21[66] + src21[67] + src21[68] + src21[69] + src21[70] + src21[71] + src21[72] + src21[73] + src21[74] + src21[75] + src21[76] + src21[77] + src21[78] + src21[79] + src21[80] + src21[81] + src21[82] + src21[83] + src21[84] + src21[85] + src21[86] + src21[87] + src21[88] + src21[89] + src21[90] + src21[91] + src21[92] + src21[93] + src21[94] + src21[95] + src21[96] + src21[97] + src21[98] + src21[99] + src21[100] + src21[101] + src21[102] + src21[103] + src21[104] + src21[105] + src21[106] + src21[107] + src21[108] + src21[109] + src21[110] + src21[111] + src21[112] + src21[113] + src21[114] + src21[115] + src21[116] + src21[117] + src21[118] + src21[119] + src21[120] + src21[121] + src21[122] + src21[123] + src21[124] + src21[125] + src21[126] + src21[127] + src21[128] + src21[129] + src21[130] + src21[131] + src21[132] + src21[133] + src21[134] + src21[135] + src21[136] + src21[137] + src21[138] + src21[139] + src21[140] + src21[141] + src21[142] + src21[143] + src21[144] + src21[145] + src21[146] + src21[147] + src21[148] + src21[149] + src21[150] + src21[151] + src21[152] + src21[153] + src21[154] + src21[155] + src21[156] + src21[157] + src21[158] + src21[159] + src21[160] + src21[161])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63] + src22[64] + src22[65] + src22[66] + src22[67] + src22[68] + src22[69] + src22[70] + src22[71] + src22[72] + src22[73] + src22[74] + src22[75] + src22[76] + src22[77] + src22[78] + src22[79] + src22[80] + src22[81] + src22[82] + src22[83] + src22[84] + src22[85] + src22[86] + src22[87] + src22[88] + src22[89] + src22[90] + src22[91] + src22[92] + src22[93] + src22[94] + src22[95] + src22[96] + src22[97] + src22[98] + src22[99] + src22[100] + src22[101] + src22[102] + src22[103] + src22[104] + src22[105] + src22[106] + src22[107] + src22[108] + src22[109] + src22[110] + src22[111] + src22[112] + src22[113] + src22[114] + src22[115] + src22[116] + src22[117] + src22[118] + src22[119] + src22[120] + src22[121] + src22[122] + src22[123] + src22[124] + src22[125] + src22[126] + src22[127] + src22[128] + src22[129] + src22[130] + src22[131] + src22[132] + src22[133] + src22[134] + src22[135] + src22[136] + src22[137] + src22[138] + src22[139] + src22[140] + src22[141] + src22[142] + src22[143] + src22[144] + src22[145] + src22[146] + src22[147] + src22[148] + src22[149] + src22[150] + src22[151] + src22[152] + src22[153] + src22[154] + src22[155] + src22[156] + src22[157] + src22[158] + src22[159] + src22[160] + src22[161])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63] + src23[64] + src23[65] + src23[66] + src23[67] + src23[68] + src23[69] + src23[70] + src23[71] + src23[72] + src23[73] + src23[74] + src23[75] + src23[76] + src23[77] + src23[78] + src23[79] + src23[80] + src23[81] + src23[82] + src23[83] + src23[84] + src23[85] + src23[86] + src23[87] + src23[88] + src23[89] + src23[90] + src23[91] + src23[92] + src23[93] + src23[94] + src23[95] + src23[96] + src23[97] + src23[98] + src23[99] + src23[100] + src23[101] + src23[102] + src23[103] + src23[104] + src23[105] + src23[106] + src23[107] + src23[108] + src23[109] + src23[110] + src23[111] + src23[112] + src23[113] + src23[114] + src23[115] + src23[116] + src23[117] + src23[118] + src23[119] + src23[120] + src23[121] + src23[122] + src23[123] + src23[124] + src23[125] + src23[126] + src23[127] + src23[128] + src23[129] + src23[130] + src23[131] + src23[132] + src23[133] + src23[134] + src23[135] + src23[136] + src23[137] + src23[138] + src23[139] + src23[140] + src23[141] + src23[142] + src23[143] + src23[144] + src23[145] + src23[146] + src23[147] + src23[148] + src23[149] + src23[150] + src23[151] + src23[152] + src23[153] + src23[154] + src23[155] + src23[156] + src23[157] + src23[158] + src23[159] + src23[160] + src23[161])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63] + src24[64] + src24[65] + src24[66] + src24[67] + src24[68] + src24[69] + src24[70] + src24[71] + src24[72] + src24[73] + src24[74] + src24[75] + src24[76] + src24[77] + src24[78] + src24[79] + src24[80] + src24[81] + src24[82] + src24[83] + src24[84] + src24[85] + src24[86] + src24[87] + src24[88] + src24[89] + src24[90] + src24[91] + src24[92] + src24[93] + src24[94] + src24[95] + src24[96] + src24[97] + src24[98] + src24[99] + src24[100] + src24[101] + src24[102] + src24[103] + src24[104] + src24[105] + src24[106] + src24[107] + src24[108] + src24[109] + src24[110] + src24[111] + src24[112] + src24[113] + src24[114] + src24[115] + src24[116] + src24[117] + src24[118] + src24[119] + src24[120] + src24[121] + src24[122] + src24[123] + src24[124] + src24[125] + src24[126] + src24[127] + src24[128] + src24[129] + src24[130] + src24[131] + src24[132] + src24[133] + src24[134] + src24[135] + src24[136] + src24[137] + src24[138] + src24[139] + src24[140] + src24[141] + src24[142] + src24[143] + src24[144] + src24[145] + src24[146] + src24[147] + src24[148] + src24[149] + src24[150] + src24[151] + src24[152] + src24[153] + src24[154] + src24[155] + src24[156] + src24[157] + src24[158] + src24[159] + src24[160] + src24[161])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63] + src25[64] + src25[65] + src25[66] + src25[67] + src25[68] + src25[69] + src25[70] + src25[71] + src25[72] + src25[73] + src25[74] + src25[75] + src25[76] + src25[77] + src25[78] + src25[79] + src25[80] + src25[81] + src25[82] + src25[83] + src25[84] + src25[85] + src25[86] + src25[87] + src25[88] + src25[89] + src25[90] + src25[91] + src25[92] + src25[93] + src25[94] + src25[95] + src25[96] + src25[97] + src25[98] + src25[99] + src25[100] + src25[101] + src25[102] + src25[103] + src25[104] + src25[105] + src25[106] + src25[107] + src25[108] + src25[109] + src25[110] + src25[111] + src25[112] + src25[113] + src25[114] + src25[115] + src25[116] + src25[117] + src25[118] + src25[119] + src25[120] + src25[121] + src25[122] + src25[123] + src25[124] + src25[125] + src25[126] + src25[127] + src25[128] + src25[129] + src25[130] + src25[131] + src25[132] + src25[133] + src25[134] + src25[135] + src25[136] + src25[137] + src25[138] + src25[139] + src25[140] + src25[141] + src25[142] + src25[143] + src25[144] + src25[145] + src25[146] + src25[147] + src25[148] + src25[149] + src25[150] + src25[151] + src25[152] + src25[153] + src25[154] + src25[155] + src25[156] + src25[157] + src25[158] + src25[159] + src25[160] + src25[161])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63] + src26[64] + src26[65] + src26[66] + src26[67] + src26[68] + src26[69] + src26[70] + src26[71] + src26[72] + src26[73] + src26[74] + src26[75] + src26[76] + src26[77] + src26[78] + src26[79] + src26[80] + src26[81] + src26[82] + src26[83] + src26[84] + src26[85] + src26[86] + src26[87] + src26[88] + src26[89] + src26[90] + src26[91] + src26[92] + src26[93] + src26[94] + src26[95] + src26[96] + src26[97] + src26[98] + src26[99] + src26[100] + src26[101] + src26[102] + src26[103] + src26[104] + src26[105] + src26[106] + src26[107] + src26[108] + src26[109] + src26[110] + src26[111] + src26[112] + src26[113] + src26[114] + src26[115] + src26[116] + src26[117] + src26[118] + src26[119] + src26[120] + src26[121] + src26[122] + src26[123] + src26[124] + src26[125] + src26[126] + src26[127] + src26[128] + src26[129] + src26[130] + src26[131] + src26[132] + src26[133] + src26[134] + src26[135] + src26[136] + src26[137] + src26[138] + src26[139] + src26[140] + src26[141] + src26[142] + src26[143] + src26[144] + src26[145] + src26[146] + src26[147] + src26[148] + src26[149] + src26[150] + src26[151] + src26[152] + src26[153] + src26[154] + src26[155] + src26[156] + src26[157] + src26[158] + src26[159] + src26[160] + src26[161])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63] + src27[64] + src27[65] + src27[66] + src27[67] + src27[68] + src27[69] + src27[70] + src27[71] + src27[72] + src27[73] + src27[74] + src27[75] + src27[76] + src27[77] + src27[78] + src27[79] + src27[80] + src27[81] + src27[82] + src27[83] + src27[84] + src27[85] + src27[86] + src27[87] + src27[88] + src27[89] + src27[90] + src27[91] + src27[92] + src27[93] + src27[94] + src27[95] + src27[96] + src27[97] + src27[98] + src27[99] + src27[100] + src27[101] + src27[102] + src27[103] + src27[104] + src27[105] + src27[106] + src27[107] + src27[108] + src27[109] + src27[110] + src27[111] + src27[112] + src27[113] + src27[114] + src27[115] + src27[116] + src27[117] + src27[118] + src27[119] + src27[120] + src27[121] + src27[122] + src27[123] + src27[124] + src27[125] + src27[126] + src27[127] + src27[128] + src27[129] + src27[130] + src27[131] + src27[132] + src27[133] + src27[134] + src27[135] + src27[136] + src27[137] + src27[138] + src27[139] + src27[140] + src27[141] + src27[142] + src27[143] + src27[144] + src27[145] + src27[146] + src27[147] + src27[148] + src27[149] + src27[150] + src27[151] + src27[152] + src27[153] + src27[154] + src27[155] + src27[156] + src27[157] + src27[158] + src27[159] + src27[160] + src27[161])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63] + src28[64] + src28[65] + src28[66] + src28[67] + src28[68] + src28[69] + src28[70] + src28[71] + src28[72] + src28[73] + src28[74] + src28[75] + src28[76] + src28[77] + src28[78] + src28[79] + src28[80] + src28[81] + src28[82] + src28[83] + src28[84] + src28[85] + src28[86] + src28[87] + src28[88] + src28[89] + src28[90] + src28[91] + src28[92] + src28[93] + src28[94] + src28[95] + src28[96] + src28[97] + src28[98] + src28[99] + src28[100] + src28[101] + src28[102] + src28[103] + src28[104] + src28[105] + src28[106] + src28[107] + src28[108] + src28[109] + src28[110] + src28[111] + src28[112] + src28[113] + src28[114] + src28[115] + src28[116] + src28[117] + src28[118] + src28[119] + src28[120] + src28[121] + src28[122] + src28[123] + src28[124] + src28[125] + src28[126] + src28[127] + src28[128] + src28[129] + src28[130] + src28[131] + src28[132] + src28[133] + src28[134] + src28[135] + src28[136] + src28[137] + src28[138] + src28[139] + src28[140] + src28[141] + src28[142] + src28[143] + src28[144] + src28[145] + src28[146] + src28[147] + src28[148] + src28[149] + src28[150] + src28[151] + src28[152] + src28[153] + src28[154] + src28[155] + src28[156] + src28[157] + src28[158] + src28[159] + src28[160] + src28[161])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63] + src29[64] + src29[65] + src29[66] + src29[67] + src29[68] + src29[69] + src29[70] + src29[71] + src29[72] + src29[73] + src29[74] + src29[75] + src29[76] + src29[77] + src29[78] + src29[79] + src29[80] + src29[81] + src29[82] + src29[83] + src29[84] + src29[85] + src29[86] + src29[87] + src29[88] + src29[89] + src29[90] + src29[91] + src29[92] + src29[93] + src29[94] + src29[95] + src29[96] + src29[97] + src29[98] + src29[99] + src29[100] + src29[101] + src29[102] + src29[103] + src29[104] + src29[105] + src29[106] + src29[107] + src29[108] + src29[109] + src29[110] + src29[111] + src29[112] + src29[113] + src29[114] + src29[115] + src29[116] + src29[117] + src29[118] + src29[119] + src29[120] + src29[121] + src29[122] + src29[123] + src29[124] + src29[125] + src29[126] + src29[127] + src29[128] + src29[129] + src29[130] + src29[131] + src29[132] + src29[133] + src29[134] + src29[135] + src29[136] + src29[137] + src29[138] + src29[139] + src29[140] + src29[141] + src29[142] + src29[143] + src29[144] + src29[145] + src29[146] + src29[147] + src29[148] + src29[149] + src29[150] + src29[151] + src29[152] + src29[153] + src29[154] + src29[155] + src29[156] + src29[157] + src29[158] + src29[159] + src29[160] + src29[161])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63] + src30[64] + src30[65] + src30[66] + src30[67] + src30[68] + src30[69] + src30[70] + src30[71] + src30[72] + src30[73] + src30[74] + src30[75] + src30[76] + src30[77] + src30[78] + src30[79] + src30[80] + src30[81] + src30[82] + src30[83] + src30[84] + src30[85] + src30[86] + src30[87] + src30[88] + src30[89] + src30[90] + src30[91] + src30[92] + src30[93] + src30[94] + src30[95] + src30[96] + src30[97] + src30[98] + src30[99] + src30[100] + src30[101] + src30[102] + src30[103] + src30[104] + src30[105] + src30[106] + src30[107] + src30[108] + src30[109] + src30[110] + src30[111] + src30[112] + src30[113] + src30[114] + src30[115] + src30[116] + src30[117] + src30[118] + src30[119] + src30[120] + src30[121] + src30[122] + src30[123] + src30[124] + src30[125] + src30[126] + src30[127] + src30[128] + src30[129] + src30[130] + src30[131] + src30[132] + src30[133] + src30[134] + src30[135] + src30[136] + src30[137] + src30[138] + src30[139] + src30[140] + src30[141] + src30[142] + src30[143] + src30[144] + src30[145] + src30[146] + src30[147] + src30[148] + src30[149] + src30[150] + src30[151] + src30[152] + src30[153] + src30[154] + src30[155] + src30[156] + src30[157] + src30[158] + src30[159] + src30[160] + src30[161])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63] + src31[64] + src31[65] + src31[66] + src31[67] + src31[68] + src31[69] + src31[70] + src31[71] + src31[72] + src31[73] + src31[74] + src31[75] + src31[76] + src31[77] + src31[78] + src31[79] + src31[80] + src31[81] + src31[82] + src31[83] + src31[84] + src31[85] + src31[86] + src31[87] + src31[88] + src31[89] + src31[90] + src31[91] + src31[92] + src31[93] + src31[94] + src31[95] + src31[96] + src31[97] + src31[98] + src31[99] + src31[100] + src31[101] + src31[102] + src31[103] + src31[104] + src31[105] + src31[106] + src31[107] + src31[108] + src31[109] + src31[110] + src31[111] + src31[112] + src31[113] + src31[114] + src31[115] + src31[116] + src31[117] + src31[118] + src31[119] + src31[120] + src31[121] + src31[122] + src31[123] + src31[124] + src31[125] + src31[126] + src31[127] + src31[128] + src31[129] + src31[130] + src31[131] + src31[132] + src31[133] + src31[134] + src31[135] + src31[136] + src31[137] + src31[138] + src31[139] + src31[140] + src31[141] + src31[142] + src31[143] + src31[144] + src31[145] + src31[146] + src31[147] + src31[148] + src31[149] + src31[150] + src31[151] + src31[152] + src31[153] + src31[154] + src31[155] + src31[156] + src31[157] + src31[158] + src31[159] + src31[160] + src31[161])<<31);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h9fada86f7cf08268cd685be5c34ed4d5c822daa365239cdb148b53253c50c506e60e8ee99f2e33b5c5d3e8428ae3613f34575ea49e8aa7d22e4e6bbaefd82a51916ddca8e1af7b32e9c810d475b5573b825e99d7fd30186cf7cf43e9054133d0396dea222fc69c0b95239c6285453f8948a284fe4a639365548284b228102c9b556734d3f64a18c1e8b812795a336a7c48af1abba0ec404dd69a57bdb51b7c982e159b15262a50729bb90d90287d30e3fe8e1e2f9679291e56c71c827302a14ef05e181074dfc70ecb4e105c96a752069e9e7b6a565d425bf1e6d8347bd666ac8a38f1ced053bed6daad59150e7f92a1873909f63899ed6353f2b175d21a734f191422898568e82a4a344403c458e3c753580fc97e0b2062c71245855665c29987a72bf4ebed1b2ae27cf12ba791c52f037e00d1d13ff78cabbbcefd9669012acd4c94e23ecc642c751970d2d11d2b2011a61aeaabf43ae54f8d54bfa69291f014e837120e06d9e268d1d87c9c4f26a42962c24403b8b4be6fe03ecc6bdb561f20c434165931a292fde79222163033016fc28d7bcb6dc8014c2b7d04328044d01c6dddd7792b340acc1afdf5510a0109b184638b05e05e3676cd6c17c6b2ab161b050baf48e2b098916aaf23a1b85aa8efcc562147348c26d13daa5847b727d37d43d3d97837a646dd63d837a5fd65368268b884acfcd10fadd473eb6d54606df1274a006401404ba06c376e11144c7b62c7bb7cac135fd91a14badcfd0d6f17a566f8365f037a7afb4b69b66480bf6760078229b25278bce3adbc570efd1cd2d06c89da20f7a1bffe751bdf6c92982634d60a4eaf448653cd92824e255e35d7ef56e390f6519f7e057378bbf33cb26cdd48f6b4029b36ca13bfa70b38fabfe40fab0b56dcc00450;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'ha26e647ed2f151b245b821f245c5a7ba3109a33f43270711c15a34108f77dcdc9840e8690607f25944bbcd8d25d1a0213af94244cc3a4ee0a48f43e607d5a865d6a01b5c99efa59b25bbf3d894a71042e256c19ef95487b28d283a7266937d2f2a8bf8906afd925253ab27e454c3a6daa32eb4af4e4bed97964b27c8e77fcdd917c2f2ef6a071496d630e88886cb8a4ed319dea04bba9b8b0787e4b0a472926a5f14033a71d7c29490f67933be104f466b512361f59d49e27b36f298caf559493d7423e6c1a8c57194cf34ce5d03922d1b75adf384105f9ee143161af004d1efb8e4d27a3e601d51e0a97bf43bc97210a9fb0e9c9be15510579b1e511eb7a6629e61948644924a698feab8bc3a57d17c0a9c6a90833a098b722cc1f6b95a4ce92789beb402e6c6ae806e98e8779ebd15d982a64e3086053a9a360330630dffe3fcfab7cdbe9460722eec538bd7d58e8efdb0c452ebd5aa3b37a28862f2aa9ce6c874a4a5233ea72bd17a889d917c099922e67c7a5c1728025ebff7fb1feb888b9064f170632cded639952f69b9cbfe1b1f5552ca0f057c3b1697354d4d9e28dd1b049b72aae7bb501325bf71dcddf1090b881bcfed56af424db78d510870f380cb4c372824fde883794f2ffc7cdd14ceaca20761de9c8e5e133fe8246e462d9d5e87dcb3ad0929a66cfed0790517e71d5e2cfd74709a6ba813fc9de771c456544482ee4a9ff662bdeede41771ff6ed98bd77c586d2c5e48c1a0b4b38e73cb10e67c1e27dadadb77d0be796ca63da61edb5679d1e9f44fb1acdb9578984d6ccc58dd4013bf41ccb48757c6b5b0bc676a00efaeedf2808cfe5b4f0b207170b2ffcde1be4e9767f647120d1edac4f81053cb7c6503788d1afad9b84fb5477c073f0e67c7b823fe926db;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h914907606994782607d979a82840ed77af4796fc71cda0cdd407419171b3485182d102fa0059b4ca1e486b45163ac0dae3329948ef50f72a6d85f2f9c5b0c81a4328e198d4d2100494e05e7bbd6021367eeb7d60a041b5dd441c59e690703944bd75f6a7d5a56e3b9b642b9b848845c4bd759ee4eebb412e3d3e4e89565de4a3d7d05c47c982243c38efc8906be4b0c02c93a7b2c7143437385a19176cb9fd85d141adbddcf8c6203a6b60936775ea883a9349d557b996eb273eccdd61fa9dbb57ee3868ee216b978559d02f4843cb7f3dbd44ece0075049dcd04ae2fbdf547c6deb166a1d71dc533d7e665bd2aeee486b1a7b73bb390862adab281ed8d2c44ca188915fbc70366d1f227ff2a431704a952389baea9f9e80269e3ff677be7b08579f6d1efe879e2a59f85d096e1f8122d5592e956ad42a1f2148d39709aa9451c0c23fa380e8b1e5ff690b69256198f645f71b6b715ee533ade87422559e0aea61754e71dc8457a69f277cdd29251feb22b7c4a250b005edf8ec7f4093df93ff7073d527d8e323648a368797e8dcb97d521d19e4847244bbdcbcb09fc486eaa7450b6f54181c5b8faee0acff43e2677157f57019a1ebd1d29ca06a4826c21d168dda7ff684ac0bcf5147aa461b43264601317d2b2156f238c4075bb14bb882e9218fb55951d644a837d75ff4f2be55e2c95d6b435f5813dfc6029e0396dcc1ae6781ae0e872cb354c361da39efe2013f723fc91abf114d1013d235dab8d8dfccac711b403ef89d3a5fa9704c22cef1c2797b2723d20195c141188af64e898777f0efd5314cb2787ad17807fb411e9c1e87b8bd130b2304e5c73111e4bc9e91d10e17521f7da2de799ad4a586694aa60419f7578b54c549d0085f4802bb4fa4a9bb6b69d68a3e0dbc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hf89c8688c663f360083a47db48f2fe77c0deb176650e4f7f9160b2062e00e5db648813157bdeff3be44580940fcf5bccf4acf8b1ab70dc2b87df3ef53c9d30d246ca95f590ef4a37b9564ef902a1b94b4929acb4a550e7ba288eff0e54663d7b34bab90dd9843d171f5af4c24a0dcead2a3b8711621b28daa473b3e8f91598e93f6bf28ffb570313eb9b44cf1b1e357ec08fde1413923aeb67635dd9d0263fe6c3bdf405471ab4ce1435674d83f8d666831924bfeecf1f840b0fc7ae12b1cd7b529586a88bac2926c51603398dd5781854f0ec088896b3f27c6173d28c144f7acb100fba6f9695c97ec3e8713a7106a1e525f957d18355b9f9638bd6ff91930fa0cc45e77093a293f04909941b071aaaed219b633776452537bc1e6458f71b2f8832eefa4d752d9b222bce240d9aa2d3212ccf7dade6b6ae16f477dfa5930200193026ff595a2470ba4e37de0549b0ff0206554db9b19d949cd0e49b68a3e405ff42978aac8613c0d7ab611fd0dc9e32b1c43cefdf63081ddca24058b67517f299ce92d5b55c53425cb0f4adcea0fbd7081f1f5a049348553ddffb6fb68e953770723db2e70b604e8c7d88ccb07a707732b52dbe2b015e954241d7a7af01f8761fad485b57b031c387f8e8f2eb7dbe91f935040fec4ab8909d9448c34d82d290c455baee84620de4f108ea9a1536338910945c78fe5791b45dc10222ace590dba1a3cd59f8887bd9f13d532dcd29c47445da04192fb1b9a0ecc7728d2ee8501829c1c210f4c7b327742c40914b6af128aa4abe46466a245decf7f1606de866a7ee03dc0049f02bb770fc423622da597f463e37d39ee604c678d78c32696598fb0c6353059d9a197802ff3b631404ec6e06e6a1c653de9185700eb93ec65e39a55b7c86551a9c3b66;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h8f2230b04a054b0cca70c9b99da3c4f4287584beb3ebcb90c0f7a4868ac534698a7f2e5861dfa3ffbef8696618ca02be140dca47783a70b311c2d933d7695dc1785de479ce2ec65ee78788a9eafbbb8e685871c45ba1840b10c6506cb3c385ed4957ac7d79282b11605ba18c4b09cd7ab1c92a77571c225243bfb337f3ceaf33ef8f853661d304fe979ee0f05790969a19d4493faa2536163ae615cf2cdd900843da06f2d4948822dd0d1226a9bee6ca1985d300bce15744aa33666a78ac55b55b5647d27929bf88f9d368de7fde72c0090b62ac7729db7c31874fa7787289cd78e74b780e4b6ebbcbf77965dad7845ba810128a2cc9dd0ab085275d1edd8289b3f065d83116ba751154c007e194a49bbedec14deb121d3ed359952c03c8195d3f5e4b5def95bf42c35618c4ad09eeb9caa96095817b479034359fd64a68ebbb1856a1ab8bcb2b716bfa359a8742ee3b602b8bd3dd9dd6902e93c0ad1d41f0709571d5b946aa522e38c55af2285c3fc213a414e3af259f65abbf2a636d8ef68548a8aaca45d3c64c78400b20d4b152f281d21bda8a398182c6521e9266e53d5be39f7a94f8b4f4134571bfc5bcbdefee4bf58bc5d7a869b8a67c41ab60c1b85e0edcf5c7a03a0cd645a0794c1684163f67003c4565e6c5ac667fb995679d4b94d6fb44944b688186286e7c8f45fd32acd8e790b616719e71275425c21a987c5bad4f19e42b31319741c13d373f147a84ea0fa2d7449b1d8e3a12b16ee6b1b00aabd811d243c65b4d97b30b6602fdb715e626d679de010e745efe17afdefbbaf03f49b605eb95a1dfb61a294ebd82be9b2873497e16c60b9a70578a24417ec81a0b82344720b34ea0ab852ddaa3dcb6aab46695fa03e8eff39957eac4c89fafa742811c7cac5d2f9a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hc4bb7ee84b48af8ecc0c340aaf2f1b9e8183522a7e995381cd228593ec6df8034db0b52a4171dcac16188c8b8e1d9f0ef923c86f672b99ba5e0a4bb88ee17445ecd486e8367dd3cce256dc0ab3f98b05cbdb47e41b26d5b947995ee5a94accce1a8288408b028dc394716bd41238813ea523eb51161785d0cca4fba991e706c1f091934fb50ff7ae3603e4e12b8ebb2decbf1c202d5c917e9276b806990949ac6c38bb3829841a1b83d2218c6934c7b22cac04974352f185cccc954343f1c914ad462ca06ba9c4df8ad9e63a38dc76d9d751ebd82f3c1aa5be2230c8705ee000ef9cad593f60f0e4a080c2e94e766615a020c23d1079c5895a822d0d72558627e56ee90d57dd79b841d1163c0c5e2cd8e33d9c846ad470b37a41736aebe1f61adb60df3692a514966bee1b6810793cf5863bb7a967989f382fb414b3dd5de0cae871772962e2021be0bd653bf39e101b55dff64e31007ba29e439dab8d0f0425e9a37bbbf42d8b3939d53d3077c6793232d5f7b5064e3f8f160ee7c341c75bd82018d44537988eb02ecf45b3467d6cad11483b3c3edddd0f543293531a722e7491e9610e704c3b645663ad38e6e1d4ac5f774d970cc7dcdd7eb46cc260ac7aa1867ed42fd84ad4ff98dd65a3f91bc4c60877a5535c99ade785073de9edcd9d2c5b7035b15e47c6edc6d12562e2f5f165b1aa5611f09e1fe40bae0cb865b7e1d5acc8f18c1bd5b5a7dc65695b4fa8cf432b8d88828b1281dc4dc2a4c2df57beeede7f921d4963c4bf1d49d347f53d473916cc4b2df7d850f0615999f5415576430acb46cd694a1bb67e52212feca5c9756d9f675fa8a36bade035e00a0f35ab2e2327c5e34e454ce67a4624bf972aed523b2d218cf92e6de0ba0fa4c1b2cd39c4cdbcd16244432ee7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h1c35cbcc0d54ff025e0bedfae0d2d5703e45e19739ad691461f90aee52a246205c23fbc1966e7e0a0ef844a456eb617481d06c5ef1d21747082e1b7b66f3a25ec3e3950e5100e732e709e9988d03c07a0d80ddfe8861588d09cdd5b7e593d572818e8b2785cc9fd890337f8cf03dc3255f08ccdeb473803f59e599f7a404b5d40719b78d25f1ff8b609537b128151978d1d6d53d47ba85a7fa37914d1fbfd46a267bdd0af6d1d3d5c7239e7213895a56f0ca25335126f33cab2b9600830ca2457a4b36ef45e3a84dcfc25ffd53141581876049c5d20a8d5d00f52d7d7ccd4650f24865cea8c1a47d6675b7af6b2cac4fec47b0edcb7b77bce7870d30985f62d37da2f4c112916e1d636e542d08470f1fdb74b3be66d4804447f7e89e0939b202236bf6a04ef17074b8dfac65cb07839a054fd8f6703228d2b46cfe053f31e5ecbdc094ed4c5a0e79dd7540062ad83ba01bc140fe3e6c4554ce6740407eae03dae108b0e744e80f5c14415788ca2d9b1943012600ef0a3f1847a0ace15f7360f29a54f3957f5c8684fd1480f8a05f2712ba04c675903a935ca8136f6b8e341ea7dab00761a3b7797f143600117681a09d32ad7a9f8a988bde1b1299f3afb8b07e87c1e3fc7c9c427702468e2133d4f330ad4850673ff9062687d28c28e463712e1836ba95bf731069631993c8b2534674175f1be7457d2639dba9918bd9bcb9c9b89130d76a1539d76ad7cf0f1071831f5a8b11e2cfe4e0a05841bb649b4b6fa09daf2455a11ae596f07ef1def54317cfcf28ab0383e13c3139177507502c45629fff492c84fd5a528e8b96bab9554a1c71b19753aeae667b76759e2786a48143c6585d48a2cc7c0ddba1162b1229727bccc6968e490ce4e897b55007cacb7611e4e4c0c6bbcb2307;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hc5874d5770779880a92a7376a1bf0ad6fb657fad4cbbba39f0fa544810fe9b6e6d241a63c475f43a9264c97c6eee0669a67fc6a9b062e1f02cb396d404c2b5e52cf0a9932af559b2abf3f993da62064fc614a5d2d8edadd1034ffe552ba5b5ff9c9a3707a2106ece16b444cd04870eac094d40e0bfc71a4536024777281a747dff7e3152aeccc44bc27f52d5b72d38dc18a3c6110e06c8d0129b27d4699060dccd0541ba206bf3315e6c20ffa091b1b2d3c1a47fb9b15f4f06645760f663ebb48d57be2b30ea4a8faa22dc716b9c450a834e4c51f6184ea0eed8f6108cd78c191666f43ed1f3f4f235f37bc8a993b3992b83edbdc898105e30823d1f27de286c6b8ddf76c68475ea50c2b0b6f9e1ea6d2959dce7aa3065f1b8996d6d3bcf966eefa7d8a6959adf44367c896cb3879d7f3fef0edc64489af1837966972062a1f7b9a547c4b7788ff89442c62b065a5d1eb159f133d246b3c051f5993976845d0de13b36f8a51412ac429ff4fc8875b234f443e8420889cee88e697f37eb324961640d1d74b188fa0c1c4eefb3d6cd550f2ad3b3f4d344cc6c445137c3bbe725fec475e85fef7f78d9a1f6b8921e7d36fba6efb3b3aa0653c430ecbcf481a622f108a9162cc7b7b531eb682c03e4081930490787ea8337c4ecb2605a297405ac7701f5e00b8657fed49487ef28f877e15613c8b52aa37d172f4bf79f022bbb422347d9aff38f680d4aca313edf59f3f63411fb5878b0094b263fafa1403d683d1e12f460d428eb2566d1aa080f3b5ae358ab47d84e3fee1230ecbf96beb396ddbf94867b52648af66a2d60f2f4a90307f115fefcfa35f0442df312f46748fa64692f0fa27c5ad83c381ffeca2a852a9e945f256cf387a0ce08deea6853036bb90c1d66dd92e6b0011e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h81f27d0a051c0f836339784f36508dd05097cb5b1f31b9d8f552e4334e0c7cfb81c3c9e81d4b6bda2446224c28a4e644ffff0cf0516ac78ad33aa29c4584f3c2c244df30c323847b5be11c67b7853feff71f561549e22c41803b7ed8f122204e62ff2be5c80d02c596d897bfd79c36b9b2bb572b2d5d761b5084a1fbabac2aac6c0b4a91431b2b16506be0c7117f8195203bd5a7a43068d0f212e9278b791ab6c033263128ddaddedcf6da7b3891053258e58b50311f460e0555f052fc87dd9e8714266adcabe791788141efcf27ea3729df6c377ed13ddfcc8531df95dde45eae7b7fda6471a415e42626b9a2605e4e81b7e03bf53c89b04ed0bc495581415cfd2ee3c5f697daad3eee2424773c6a3137864c588352181c365ab003a4cacc7221ba44ffcd9f9265702607808b09dff3123673c4a332eb1475b6bd0d733f7156184344f5bb36f22cc6750534a12f7a45c3640704cdaae97c75f42d7a86f29760174f5de58b819d095570c8a8ff475be343629bb5125068a7e2020d99e772056b7d2cec1319d2ae74dc61fc5d4239a810e5a965b193a1fec89b652a1695552d80d308046942897958b6f11f2f3acc21826754ec68c0b92c8b79d853a562f27fce9e0364b583b0be9abe3c0592fbbe3a6479719b4e10d9fcc6306736df68ea1c0952166afe654c64e960bcce5bcd5c1fc133c76f30be25d8a15ce6a1977ba9c062afd5a2fdad8463c116270719ea5bbefd1ec5eed97e8f4807e1713e64f497e1309381cf688ad1d45e76b71ca6f9cc715c82326b54e19a9f26dd331df66c68e14140b5970e50f70f10792b608dbe3e2f7551f452f550f932a2e73b0b924accc8c9357136a190fe07d1126ed8c4a200cfb72f4bac53b878c061e9f4e141eb328e215c9b997d6b45fb0b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hdc086f89959e876fc218f891b71ebae6b6da7844a0ad04d8a24b328acc4fde81dc13ecf4d3b17361cac7fe15f4974afb62c4ab6f2f93cfe58ccafff2c0dc975269bde855bb07afd7eb65f78b0b1ab4a1afc0d947e8077700778ab8f2bfaee82540895a44cac36b9e192212f014a8e521b6c6fde350db1ed7e2231fd67def971bb7574391f3eabc09d3c34efe79938f416dffa905c373a2e9da36b1116e743cfaf01ea38c3b41dd316ed5e29b5203894d1b2f6915e317a9be0aeb872edee2c0bdc940a98793501000438f5ac2584d19127a5bd4c66693144d383f076cdca049ab1b696b6e8809276850e23596a135e929770c7dff8631d0a28219489de6d993d2a981996a8ae6730c6f8a089a81d269262423f13c5a79e487e5317f68d6377e6376965f665aeffc9fa8b02e3f5a5dbbcd42256c0e58d6224aed64eab0bee5b2de64df3deb752dc5ee787610c9868efb43ac3cf3115c8cd5e5de03c41bce987f86e1a847600c0d734a312edd286b0b5de3aed70d702cab42df2869168a4b8ad5cc64465800156ad6d1369883b7fb1a938c910ceb09ee3ebb653c139f14955dff70c8c31bb66c63e5a06df621e45a80b362a103f9689901080d810a012b37ec02d9dbe06bd78a5ce525e91f0862853c3a45834affd7e4befd0dc7d5598e5ed7ccd844fab0c2859736bada33f7b66d930793ad5bf0724ab34b0483d77caeda1c293749a9eb5f16491ad7f7858731b3aac446af2fe35c0fd57af13b99450cb07cb8bebe51c858e4506d97dde46b395f98aefe815b3bc73abddb2c36da0a3dd578002b56f0b3b4991861f40feff004fda16bb9ebb197a2b977282113e6ace3f1d780842fcd01d5d191fe9d5f97786c2f61e0bb651b0e0668539ef5a4a1b7aa59b077d4c9ed86ad20007f87;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'ha950fafc2d15fac8b5dedaec3fd69c964479eba5dc7d9dc2f558f557768d3909d93d724f71538005d58f63c797894b9240b760b025cfdbb46f13adc5090e688853d0e4e27e8a911f3d2bd0aa2a153f92b64dd65f855fb80a409d4856c329bb5194e9a2c7eaf11431f899be09ee38f7892e37756da983ff2eead1575b828e955eab847271be88853f8a2c67d333475a197c5e3632cb740440d9ee3fb1153735b514e90788067da85fccc710c54105bc384c49657be427aa2667f261bbe261e56ea868f6ec8d5b4e2adcf9f1ea91bca80f72bf99aedc833d720227f2fd3aaba37e46d1bebb0bba8530b7660d62c597b0a71519c7b390c9ed6a1ef32a2ac661df4f621f636f47833e35df2082307ce99a6d0ae5f14baff5165ab1126ecd885678fd52b74bc9dc1cd6b80e9510b0d1555cb420bed8d0c4e0b2f90cb269d4411f84e259a57c98c06ab7b5f7b5ba2ea2f3419966f85fe5b97200f4c279130acf6f24179d937d08993a5b41f9c49c475f05f3b5f70b492e380f4ca89388a4cbedee10b2fb77f49badba251b55b0a33cf1cd94e8d41cafa879e43502a68642db199b338f3166daa3cb26b519b2175a1ed6bd1afe230869070c180d97bc6b44a14ae39242690292c803676c25d2458c5f3b70346e5986e30ca5032aace0d244686a1f66e6293f1f4d15df2441e087efd357231bdd2d3baa374fe5cc4e1d2b97492deca44a9c0f2facc8387f4d4cdd46572c0de1a927fb4cc7ea86847679e045e68d487e13f2b0cbaf436dbc78f54e4d0845ce280ed0ca9677a85b996dfba98ef5928097c79985eabf2dab16ccc3002f5fd77cf173f98662f8e5ac7b12c2a3a3774a838f600f080019424639313f217316c30ff02810144f94934d2ba2601f19e5ea3663d103497d65f6bbcae7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h9c0abfb1d24db7dd8b3d74d254080804ddf15fea781ee0bb8915fdd749a1f5a218c0eac947fbdcb3e30b2dcc726dff08c6599eac876f2b1aabb695523ddf4f740bfaafbc7322414cae243cd69af164af9f18621c5703c58d81b6f228926f4b589d048056409ffaace2f64235d4cbca982429d9748bdaf2f3fc4c51c0ee1da13c156cfdee19722934b12ceb7237e8af5e1d04b35c0f4bfd58fbcff8ddecf12de1e3174baae11ce2c8f76835d1e8edca15a704152bb0a35d633129ad959556668af32749fa2cbe22dd6824f19670248e899a33a9c5b79793dfd5df79b275164548e03bd999783c9c0fd76daedc816c5d718eda50c6dee413a5ca5f289bfe8f491a4513d78aa35fd7eaec40ab850e2147f9609018d61f3c0171480c6eec24e034ef1e0b2f5bc8205841f9298f5d2a5890ef35134552d3776bfaad7e1a0e37fae47c42e8ec38c730c97509c3360599bfd36f8d565c16d770487afed4f4a2c2f246b840dd42e61c5ec9703f8a7ef63e31b6f375680cf0b07acc9fed29c787d7330df6599bf4f103b7afb6f8f1d2cfa883dbfe1c07a54671537ec6f641da4d2b811e6a987070f88882d8150e91461c5636be3ec210495d26fe80895b1ce51bdf6a7547347435950c8a6e96886c57ae4f6e7ef9c4b8a10fa62385810971f4d2804e7fdbf241e9b953f6ffd83598db6490250080a7af9bbd7112e0975812140eb78058246e241483a11a5d2f9fa435c9f061a4573bbcef0a7d1e181af10e64750a8f7da532f1e685be7bb8a9d4611e7b0414024c81e24bbcc5eaa4a9d8894fa933488d9539b38f9552d32341a21354409d2c7dcca4c9614752d7cf1c81d3150293315e507d475d9ac454962e3311eb6c6a506223c0ddbc6b9d95415e3bf31c467e6bf5894a9cfcafc8eb2080;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h73ef7787337cbcdfbab181a8d23d32d7edf48bac45ffcea3f2459c81ae6888a6c647fd828c4b3497a58c91ec34bb5f50d09cebcc4ee7dab72eb5ddd3d76ec4f005e5c9549863631a0f3c0100043344faffb07df78dd6a3d5982cbf5b1fb4450eef2b26d51ae7f46cc447449b40353194007eab80f2c9269d8c270af51544a88fe0838e6ed1d6f0db217b45ca1def3df3167d9c6548f7f16428a2e1c94f64fc54218feef450109b3c7203698a56f4b5acdaa2963a6b35c2e25464424951a8586da9edc165407fcf0bdd24e17c2aa199f5a965df9e94b653299a7e116fc72f3357209183185dac13efa2010ac72b8465873437dfed6d469ed82eb849041e4364d426f58a6f2f1d03006764f8a16439514a604338b7cc8dc16cfdbf47879afe5b047966c2c1944a3630d2cf7993a87f46689f90756f77e296a2b2ed40ffd45d8ab4135d5582a482c6d7f8864d23891849edbe8dd88fd001c593352677e8866480ac8bc219b3ffa601dc90f621fdd8fd62193d005a96fd41fdd8bb962d764a9c4abf76ec2f0d8eb202282f43c1bc5290649ef26a573fd96d757f67e888d7bde95b8314b15b8d77de2883e005ce6b6f662c5485fc566a7bc3d189814d4f6ce53b32a7d72f3b420742177081dd86af85823fb32ba5a9b239bb04f6b4a956c517a5199f49c52f58cd01eb5515bdcf8cafb4fab4e42a30906f279fa23212101955c53a681f8af4f930aca411e7c0a7753b7de3a0457fb95325187707e07e37485bb636b18cd1838a3b478c4951d9ac6f588a47dd6152fa1faa49421c426c80adad497d8c4438c0f131074ff38ff4be27e04945087194f7fe0a081356f9998c060c543f3f25deb625e3c214e1b6e0b93ea64d4287b87ef6a66400a39153f6660772ad7ceb3481a85d0c5cfeec;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'ha2a3c55683de9be0a41b3b78f7b94ae02f770a00a383d3af95ffaf1eb0b29cbdb666cee650c1b1370ec0924cc6888329b7ab291f675e0ae34700e63d40dd81090942d711871a690942c6fd0b029672578e2822373f636d753505b52bdacf7d7496e909de06e2669da2509686530fef411cc550f972f13ab4f9f98edacd0594af7aac39e6c65fb879cced809d25140535dc7639bff5ef5de562315ec97f1529a70f049c59a252a1d35de0d354bef553fadae41e3b34f9bc40e011f1577106f38c3a7c01f8c415ff5e2f8f1027e2d7b3e84c56af3cf69b1d3626a46367eeaaf357165ba8e5276f068d6e659754ac4174a43f4590c0cc45542cf06ef5785918a2c6d1118bc51034036923083296ca835c1c7d527b3c344b6ad4ee9947f84821f3c8826a0397dcbb6374ec362e264d124dc4d9bd6f75768a6e7cd0b31de46c8f22b7db5c08a91d25bc8b2b9fa84103db7c56ac5daf6f9bfb10077b97d7dfe53e4e119e39216ccab7b5aab6ed7f1d950a39137035127755eff429dc524486783685886ea514f6423669c9f2fbe383198dcc75150afbacb59d141a485d746331f5e8962de21413e86fbd80028f9510aaba98b34bcd9e5303e9f37bc582765d5c51f1bcf68f786a44af8a65fe99de9af856ed09d8fc2a55c9a55eb16f3f07f3453ae4e84be9d6f05aa22e16dcd32b4994c71c8e7797418e20de9ab2754777a5d8729141a6bc7fcfc4dd785e8b169931e0d82913c071ba68e44899617d201aca9a597b62c2bc0044b6ba744e3d43fdbda35e9efff1cacf3bad8e834a33713e89ba7544e2d3d59b1de8956d390d9931a3423f4a2dac1467c25a81fefc8b074d127516b4b9a6e6fd5dbdd6d89020fc0bdbc57d5dc2db2857c5fa24ba88d5b41637a0a3e75de4ff1c10b5bee1a6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h85d07f0dbf2bc9ca7439965ab3bb31c24fa8b2ce1306f00b10068f6eb3988e9e8c6fa8a1b84ca81320e4cf040659499f42864f5931fdd22bc1db4df4dcc41c20fa1f276008c2ec44ced410b5805dbbf5bf12eec0109f6f9e8fc7c9a6fb13b59474368f9b0e56ad07cf90b707f69a1efd4f48083a759b76772d2ae2cee2f52c402066f12bae749785c3b46c6dbbab3bcde16817de5273af06248dfad4470bb8d0ca9db3da517fe6dca74b164defbb891139d766ae4c4dfb8117685cbe17f71f6b1524a3c24c7738ceb596a799bb852274b7ceeb8b74635060d9029c388d0bbde12924fc681d8f9ec1cda55307f187d41f3c34d25914bb2068153af40f7836353f7659c675fc38ffada6387b11ee4ea29b003c67fc19d9e4627883f2d173e08ce508fd86cc7c4e66389c0d14c7f8025d55a7bbe16a034dff54533b353f2a44be9102f5156b91593303bddafe38a2e86c92d0f8c7a6fa4d62e4d11b8fe4bfa4e06f8dbc9592a392bfd5ab48dddc255d05116758ee63804952724d9e8d641bcc33b00baf308f61a03ba1168adb0d5bd67f7f335fc5dd33b18197f5cbde24e68ad6efcbec97065947b5b5f1a59dd52d0b4f1fd4a5073f6863560ecb897f1b703061f8b5379625a67f6cf444893c1565f42c65b9155b50ce62660a37d24d5cebeb49a7aed33fc3fd770d15b56fa7d8b8c6475c4e2d89ebd053bedd52784b97c1df9b89c4e523ac397fc269fe3da5ba3a610803f708c759b918efb995e1bbfb3c04e2161662eac94bc20a7f14cd7de4de7aa710d2fab5041b4290b13dec506c1a16c96b95415aceed20823fbd6d61da7ccc212afb1fb66e08e03a6151785649f045a8c0a7f2c0c9e04f3290ed56dc14a56a5a6e48043bd2a0d36cfd45eec31bcbaee3f8cc0b0a09897a3e3b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h462e7d60b2a4eab91506576b9eb9ea56b19b7eea68497e5ba5c6cc64ec95d76c415838cfdaac12362c6a4263bc5da2cc35564df360b86278b3d5efeeefa4bb8e5b1f3571de4d0938f328bef6f3058f126db79007c5c4de08795121f83d1177cbc52ac29a4a6c1f5021e60420ce8f9c88b0cef6d7e42d1c27d9c822cdfca58b15a64cee124fef34141787ce7510de27aaae13c6cf4dd4225a998cf876e1d88bf9fb4502d05a90466cd2326725c218ecedca0b4806207253b136e33dc94e391cd1991e4c76e2a3ed3ceeeba3e493af990ff7829ee9850f65afc3766ea67c376c2c4fb002ef8e01ba4cd125bb2e0931db36b2076e7578ce98712b1c8bbbfe885b23d6c5ded2eebc5b5674a701a925dd39827280d9bf9c0c9f7c68a9cee042b7faf1a6c1f3b810a22e47936f9075d5eec266913ebe382e6884b04605c60fa5657a0de7f308fbca497f3a92fcb0768f77af9c7f77b025da8546dede5413f1788f04591ad69e2a5e839270509d46764dc24b540025654029ea0b259db10862c80a01ad4a16b6642603851e6bf3f66d908541e7c4c5878ad62bee914513c98612484e1683256bc5628c705a912ccdfa47185b37d98f1b4aa7e386b5aca085b871f76e21f0efdaff10a2f37d30e6f9152581928c84fef8016ce6ba2a9dddc44448fe466be242e40c4f8789d07c641c259f8f1e259d541de6f6e34e5becd1690e11117447fb9a63f07a4913a8157f02675a2c19c7f5122df3e0b0556d98ec90b4d0ee14d0342eacea386011563ed9cd4016d9d56a41b49011949571f1304faaeba1518e5e2d6e1e2c3785676501f4c9d96ee76bd4428ae010f220f437f09fa414f447aafd9af588e3f53797a44fafda1e9e8b8ac23c3ad31045ee9214c83d52bce0eb75bcc4351d055920933f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h563b4868cc72d7f525654d0faea86e4a17c93f5f38c8217880085afa92a1c96cd5ae5122053fe1fee307a547c85053daaeb7ff3ed08025cb1fb96ba6a0d48ff8f5d4496ebd32edb4d85b5220ca13c38f52dc4b9270db0a6a3314d3bdfd3818e952bd091bc8983f4ecf57d8bb9170a23f29e45c9e59a2db5f37c0f31ddabd054fdf1fb869dd86909df54e2f41f9de4cf554a6f2eefc07c8bcf918f5ddf15d6a2cc3f8cc3c3f3fef7bac9100530a536a0cfcce30eb46352f61555f861d509ca60bb5ade0ff52a65943d687133c43dabc1fcd342b598dfadfc012491229a610d81b343e5ae89b01568720adbd93d31c082fca93d075af1ef28129e1feabced914f1e654b2296230531ea55d05b4b468a9f69cae4a39c54918bb7b2af66a44cabc26a6cf2402d19e17b04503c64b0a6ed487eaf4d42dfed9128d08b2ed08195bc15a71528fda03aec25f0ea8fd74908b7686d9648d85b59783979dff49bc9f3a959754fcd49a18d413275d0775ef3592319f2f15af244001d8c706e89d07106c2840a704e6e8868b59d92d0e32274fb03021cc8d6a464f92b3ddf1847e1a77a7e8c53c4c4650951d95cc851b219a08af0ea470c9937379f1d3fca6d53d5b72c837155a9c2f78926f87009d58a9134af267ea2d266019452dde4fb544f808db6195a33cebc18709d0f21111be21beaf027b366c3df0df0c0b3dd40382947ef03e06b89f79114165df4a21cecc804bf92b579c9f4130985ce2e384505af77d82f7f1f323860bee2babc93877cc577afac6e9efb88257b0bb13a77175d61c3c6c74b9cfa95a4c413e4f1046a84f0edeb753eaa8f22af2ed2cc38b78ac171b77182384b00c357268a41b3e4452bf1d77076f6813fee5a1a4d9a6cc304a0089b8af90fe692dffe18581cca1bc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h18f4024f74308b620eca27e1d613ef4fd98f878a9520d1cf93dd9169b932c97bfc7cddd2a2c10dabea699aea5987543fe6920faf4d23bf05dfa4595d9e835c7acdeb402dd114440794b5195c87056b18aabbfd81a5e7dc72ef82ebe5813caa613f9e72db25d50e6d488033c38fe8f5330b873a4b7278126c83c54f4c7dc076c822c5d5478d7642b41cdaa1fe284015aa566501c050e4c8148015f43707f8fa0c07fd19b11bf8e589d7d2cf02af3f2c489a220d480082cdda230376145635bae3ce7f6a78795f9c4e8036829d35616dacc59e1ed6947c5399c6264250a6e1d072dce549a07ed14f6c96f5d1a4d21c71b32df5a2daf2c6327e099eccf597ce11041ee2073dc4cfc1ee31bcd3934e30de616bbd48e7ed06a74a5faad849fbbd35ae859ee6d7a4be4a50f33b73c79a698476891126566dc1c140f103fc206f20c1649828165e558ba0c2fee8e1cba5e3727159f2cac31fe601a8500a8021aca00027df9e7a743ca1f689be23e57343cda49290a7366459d0591c304cffbabbf1d7fe6f72fda222a6e65fbfd530f1de15f385786c77e9d483d6cd6153cd28a0368f700f45a3d7ac862cca4b99d43459d7b9b80dd5d11a6de9d2c75a02c62822118f72e51eacd82505d2c55b6a3ea58d23498a03421f2d8702617da3765f89013895106e53a0a5a423cf59f8bbd3e97e8b9fc83183fd43508a9bcfaa98352636020f9eb6e22694e6635f91a26c35f628142581606c9284f1bd866ef365d9d47e489db65862835bf615ca8f89d3fe8588441f6d7cc3ab09ec3f13903c7ab924fa00b8a4f98b000a045145e98010d30504963f05b2e35a9d07c52e799252f2e98b1fca5b33eeba65a38e917be41be3ff50aecf7b02623c7bff4323e2f32a1fc54c39b6d973f08a74d3f7a23d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h7bc5c505a6b548fe389bddd4109741762e46bafd0dc07fc70f6e0d53b3892dfe9d5f0c26d9579b81fd080da1567dc4db2dc6ff9ef802fc1731d03ff9695b872b46683aa2f33ebdc1f67fc1543c5a1e502373ad9755445740cb3bfd021917042c5663ad63d77edb29a0ede58a328550bd1effb39e05a2b5fc7e228b2921aad0fd0e287f08c15583ac4cf18e5c675bca1cdb049957f809cde39020e67ae21a124ebc251d22a5c42749160d3eb3e65113148be15c2d010ce0ec3e4648ac1ca0ccc02dd013c246a382502639ff44672f50962d2e7c78f98ca67fad220a39f4ca4f49a4ee2d5f1858617ce6a40ff8e99d68db45f43740ca234bac5711153a9f46a50528b780c60588e10e38df620d36f56873435657046c9aca2eef9213c432e1ef08270cca755abb7de6a951923381a1b96cb7806bb67e3e2e489339c877539a4b6d82cfb929acb78b5db4a990141074fc89cfe741453cda9db6af41404bc9f66492f39fef0d8db7d3c63d0b53532f0dcd2d771e13248cdc673d46401ea360d013a31aa4c052a34d6c15e496a5b551b046268409f08cb437845fe022511f10a7cd53f8920fa0c4603b1bf1f7deacaa7a11d9400fd9512e2f6f4e23c972a155564eabf11e0e857f030d3d2144ff2af76897bab62cab8754f73884e151aafe9b0931c613a937a47d99d7b3901876ceceb12d56977c78a03dd4ae2b90a641858783850f8e1ef89a2171f465c7468b7c325c5fd87d1e69b07f503c09b131a3bb8cb92938ae2a3046b8451b5e6c803ef40abe8d25f9cea7a0076fe8ce4830a137b693c4a3eceeb12132d7bee0d91bb023d42f65c647d3b67d0dbebbf522af451afd9cbea432c61d6c168502835306d126bf9d08d43756301a94282ef09c76d1e8483fea0bd79c6f4e4185e129;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'ha572aac210958827775ac4e2b57308b2eb825835879b1b881e7577752070b77fe17f8b0d2fdd05563139a2e2f4217ea69f9937dff6b5679db7cf9fb926c45357130819e18fadbb8eb92d87ce6ab9391bdb06b491b658aebbbf937b78308313a3ce2e34b43d66d47446a5510c7f351d4df2049c813ec31f0be7b24cc82de051a103a47422ad5d177aee0b23c9c45fdf006d01e2e652cdf11bb9d52071f3addb7a559e760bbd0f748cdef085c527e314d2f3e506c4374f421fa5c06735614915643b592fb63720263dcae5f70bb20db1eb047ba64dcde9f49f113ade8c3d084a69a30e3d9f171bb0ba8c0c3cdbd21b4a7abcaeb095f0720bb1c8dd2de7718e357729ca2a50f4b86dc72412d45249f8e1f8afc56b7216e8af63290c7bdc37b076021aaf9a80f30bcaf27f67fcd2cd410665810637366c12a1621420aedfd24af8251e33cc9ebd6a3b88a945136446a4109de5371923f0847115fee752eb8ecea9c1cf6fb605e8345ea90722370966dcf7cfe6f1705b0f062d813922bea5a657d063ca8675fbce971fa780a46388bf998986c6f7c589d16c1d6d4dbcd20e8fb07b45ba46770cee34731a71d5a87cfaffd6f168f1aa533d48f6039cc710aa49c3ac204fa8a56241f4c1eb126bb00ec18ee2388ccf43945100a597292b32a7f3bc5ddcc404b76f1040dd173a1ddcb3669b59dab4b02e4f361b378725e6377c721fe197a9a8e45ef913406dd2c0c4417950d2225013a7b8ce86082c2123316ec3ee39c4956a4e1119219d1f7021b0f22d8db999942367cef673788c1df2f309842fba308ba4518ab2a0f3d8a40c4cb13bd6cc2f4fa464dbe3c0e6c88e2319ed24f802debfd2eb5dbe0e93b69b9190214139cf0f5590de4349ca888bc84789154294760a7493628b0ca37548;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hf8518df06522d4fa72d3fb830c824ba3f4ba8f9525c5e01648d195f7a6d7169da3e13607082abe28ffb78e9b6ccb447045b1ca92d84c4e2c01d839f3420dfeb95cb78a417562d8c4fe67786368f523c5e53b3d55d8fa97eb7e34746e22a10043a7bc093fbe65cc1679c243f580bf35372c7610c44ff0eacfb21c231741278b5d0b6dca38cf508bc02a820e24ffbb98f26eac687d57a4ebf2c0bf0d56c8e8c5d06b0f023978bbb83060fdfc031da69c4aa20d4f038feec467f14d83fd11acd0e9ebd6c171300e4e0e0f14fc3619a532c78e3a193ac86160155bfaa5ee77e4d0fd12ccf92ca7541728e32be1a5a9600c12944912c8284f9e454527d4fb25eb2caa48a7c5dc329950ac425e56f89f151ff7a4f90d7f00a7a00c0fa632dc30f9ed7a70723252b06711eb82082a0e0155fec332441e41c8aaf4f0db439cd0f1c931476acb27e5eea2389bc0a9d30e8901b24e31f946435226b8826b757c12322d64fe8166c284d9db6f6bca7a6c317b02fa61c4ad186fe1605f361a39fcc39058cc0863b61c3480b5f10d54cbbf2f4bda955279776c848d5a3a3c0dbd0217c5b8de0ef0ddfbc7de8dbf2a48243c01982ae6a0ccd4e92ee67023382eb843f9ecd585354c79841206e2cf92674e6f571e658b004580284b938f24f33beb84fcb986c6b4a7f4bc188bb927124adb3035d518cea3f4892470c44df376250ed5a2906400c35353e0e6a26f69c8b1405dd2d031803a863f21e0c20a2cca759d16283eabc01bd5229467ade18ba3957f5c1e67369811f5c36f5bf2b39bfa793d748b60e9c5c4be37754060d4ebe9b29294879f56218f9e6f191eeedb2762e7ee31d4145d348c9e7f7f31fb329e556538c1de4e65ad7b863783359ce25aaf4a3869508286236093519c9bdd26395a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hc9db8d9ce1f592a4444212e973ab429fc43088d468ae246bda04a0fa6827da9b13150af8c77e59e324649d78039dd97f65b6a9473a27990998e4344360fa39d13706795bff11fcbed44e20fe87ba192af7b15c7b3a4f7a6a23863d2bb6f65cb54f163bbf2a4811e211da59687bb604ba436edf00198c0e3a06ff18b87a073cc4e8619cce0fb787be9d2ade905751f3fcd0cdd59bbab97d5ce3923d0854a1ca0c4323cf2607e8b839380fa79b015dc36e04871d2893e09854d4292d54ac3374fa8dfb253e0bc45e7025b853cc33d8e429c1d271779c5c4a9aea8a86ebb49f4dc29a58b6b513f984a763b23fff8fb6f989b240a0b98d9f3631d21387c5a639ca9867f95bf6f653ce048bf385cd367dc320e3a8bbfa4596ca2685f4fcf0fc7ca9402098ae9f91a973e7b60fd7d6616dbab8688dc2c912de9575f3d414575b75c6ff2284c9378c64ea0f8a8049ef99a4a5d553b66f05e7186a3fd66dc6ec6dd5957bdecae44c3bac50bfec3f10aad892ffc9e879cc067678dce91bb134619b6b91fbc9bc75b801bafef8c13d9a273702dce32937a302abff38e1d62941b6b9077cc1dde0c7999db8e96f6203f10e7e98bf0707bed03f492a6aa627dfe270edde8bdf5dca8140976ee4597856dab4d625797c3512ed8965e4765b2050816f8b5d116364b487d1945114919ff8d2033ece314ec2fa25c5d74a262b235e0f7f606a7ba1c015d7d2e7b9bf904055fe81e2a6eef3edb9817bea6dfab9c57cddafa8929b8bca3229f8eac2f575322b95d72aeb19d35a1648b54c706811cf1e7662dba6267a0634f2332a6fc74bf462ab107aa7db70118e578b7ab821a57e9b79d9d5b6909c1ab6e2451209b3af371df6a6628d5a3c7cebaca979a5904e2198143e7a4a11846af4943e9eacc402;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h5ae9088baa4ca9c2e5f4296e7ffc26e729047950b2803cb73466ce69ee3f214edddb0bc129940d48a400d05bc1b8f924f104753caea73225c9879535db578cb26ae0f19d95d52f882abeb89af9f0f05cc2644681b4deea89e58a80625fe3d7e16b6b2c4654fc6b3bcee8b29f9ad92abf6d48b4379c99bfbb72882bd26e4ee70a3f43a5e8becc5dc7e360823f5a3b8368bc57be0e13927af2212c4ac3b4835131729324925a9c96023ec4a77a11fc2f67f5042952e97af8a01ba64687456239f9ba87cd4bb87af37083b0c34579f971810fa302b0a04e5ae0ab3096c1f1b6ec433116bdd5a85817da20e70bc5594a43adde66ff240e439d688092e836c52aea967824ffb8961b1ee1087c25dae5751f6f6deae7c446adf7850e017daa3126180afc314699a3a3566901958591cc39cfe5e328123e7c90f00bec099f2c8fa16ffd51af305febfdd949fcd7613b039eaa3bfbeab80d62ec4c7e156e758cc633ba78072b710e67bfbc330b2dde3cd06fd636bfcb65b7020be5b2356ec062008fd5a7d4e5069f07946ce6dacfb5edf56f014cb31185b85807c92398a27213481f79aca43928b629a744cb2a3664a0a08e83a061947b4269b0dbac9de9968bdc026e9845b74935c07bb82446f24da7301acfe5b076549d2055cdbfc337aabc5247b518f1ca2e1bc2f7fdf34a78d1eae1d73533cd970742e86c91bcac0dbf3d8658a5495d91d8b003c0a7a1e29ee1cc52d7110591e13f711e12bfca4495bb9ab1ceafcc0f9b91882775a524ead8df3b4cc62adc0488685da274d4ff52e9ecf71b6c1787e7b9fcd5b69a4d244af90a1e7a0193425ac5abee00f91086d29fa2d53412d5f78d47e2906e4a6c698018ac856d88dde7344b0068dfd21ff9b8abec135b4e7d455244454895505631;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hc68a49c82319fc980c050249772fcda9dbc7c600027adf0ef7d9246a151b6212c9a792b5d094b5af5e4c33c26fbc307e28faf6f9c08a25df147149ac8f510d7b5d3aac5a10f5db568bf8870afef64fd7a30b91be9e821a2be2f2a5c397cbda6d1701d3e6686949353fea64130019e93f7260f56c377b323695e9ef6a69a4b75a5e245cdb3c053d1f61d5317dc799bbddb7bd3a5daafd14716f296f6f1eeecc3c04a1f3e1565d374b41495c813bc336b30d24facbbe1fddd0eb0429b2f6f4634228c5c2b1e7ed17131d3a585e912bd66f3f565c7555647194fb9e375c35cb752d0fe20162622413a7e736f072881e051547b92a2a3f5b147007ab77de5b558f24b5c4c39bc6dd6c1298cb4ef99b654d60ec1035eaa43fa71826aa4755ec2b9f92c7c404b32328c93bceb081ebc69800e0beb91e5496422f7485aa31c9e8d6915fb95a7562f08fda919679968ab4245adc620db3f1bf0be7f3ecf34659b5dc6d854ee0f71b14921b0cdff68c3d27b39ff1c24f465e2fd47ee5012ca60ca209057b61527725b400ce1c8dfbbb112b003b77ce07ce3f2ab445a25619c618a0ac935079e912950f62145dca88100294dcf0187bc12c056c98327f21f5e03cc0073d1bacffcb2485f6c3dd41e7dfa224bb6670f25cf0edfc16994fc0a6116a3647725208932d65a41dba424eb2cece7992b0fea3f9e52ac343c7de11cb52b0f66b8a824d6f5ede07e893ed13eba1a5894a3f749b7008a16317175b87c5f35761951c39b0d60a33b3e8a7d3d6bd4cc8dba7badca2ebd84bba52148f698b313b6028b340b0c880bf04be2067d9ca61c22c4605cfd4e11c8ceaf5ab6a276f6aef0bd5f15abe8e5f6e3799c7964d2843918001fa44d906a3d927b8ac39e5f3b23c1ad4c90be7e4d8ac79792e06;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hf456de294668956954efad47cdd192f19cf2cf1de3fff35ed2a13328fd63fd71500c396eae0462977097f5766da2efa6e260787bd6188903e328564fa996255319f98af39fcf64b197ddf30a8c62e6b94fd42b4f8fd689c68810855cfc399ff37b86e2577f4d84f9b0773e38cd1ae5a9ab360ba22aaff9dcec195ee747898b4f246c53a14a473ce9f6da2a73fd9f51d995446ab1e0af115b2d620a4f354b675468addd7e3bce1ebed468dffa6ccf796938c0f3c99abb217eaa16e9305c20540676449f4a8707d4b5ca6ff3511302cc16b48c61e274428b8e15495afb780d03a9dbc3b04cd94e314222b601cfa56c1b644c702930918acabf90b4fd682cf744837b2700ba6973375c4bd9f0332d566d3dc99a2737443a8a7cded8d7a83e6b0b2ac6953c1a84317ef8757bfd9e94752a46532f0ac5179e65aa10d68ac2bbd03844afbc17f11a77fd204cd0dcd5cc3a1daeef08499feaae18ed2b1c209d10dba5b13a1e645f1236f8aa06405293daf29ad645e8832eec835b0e048520214af71868f2f3091eae235ffb6555b5f17567faa6eb6de42b2eba49a9393f36249dd869e35a536ebfeb70411904d6be07641971d2c388011bd8a3e50f8f1326ecf0f36256cc20e850b5121e2c000ddd9958939a2ca52ab5dc990948d433aa1e60d9acc4551701436f5c50d46255f3d23639501e6e4e50f4d6fd3b6c31397d428476e50adbfbe6eda22ba175a9d8572cdd36b8601e2308f1c389b754dc300efa76bed301f8e9d6558d5f4d3a6ccb4e854c9ac85b740f18b6162bef34fe933c4325e9254e15f72d32666e316d166d9a04064762b4a8710da43e1c684bc24909ec4af69c8b2fa7ac192bce7704a64b649d7f2b75e4db582f26713cc68b2edbe0344099048886dc9ac39a6e2dba5c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h4ddbcca3c1230262ea3a74cdc719ad3453e7c8cd0ca11bc31e7c8348b89bd8d900461a3f74cb195b036d7996b9ee6e9917d55d32f6dd9d620a38c81091f20bf5371f951dc59c87232f6cc79fc99376571c9d8a86ebe3c0e4eed19444d202b5a0b9aa4dfccca8ae5d739b21dbb207d6a1247f4d056a760ca2a8973ecd2d512d48720b71ac7d3ae3bc82d774933c7700133e4f990a8db8f2f2b573aaa8bbbe6817fa62a7df6afd3884e0366af9a377c6a3c44f3150786704a508de9f21d686cad873e2a8b062abc187e8afe9ee7d6b5a9b897f7a85e309e81a11cf28fbcae9e956f2e0091ae158009b372fd6c664184e84e6e1a4f6fa3cb4ecd9998bce0616525416bdb0cec176e35136d6f8bf9e919e1920c76b78c1a6020a0c49bc7520fb62d7d826087d5e04c1bea036c36d0dc24701a2038140eafb588761f248a143ed5d33f9a6dbfb4264b2af56d6fa25dcc9ed045d27cea343e8b5a383896445ce5279e2886bb0ac34d35311784cb78002555b5354353d9969c0a2f7333eea044084290d89f39c107a8039e1d4faa9b0634702678ac5394765b534e613d3bedf5c878d631cabeb46d17205ba51306d4fb6c256fb044303d0fd1e840c650fae89d14a661214d270a799d6e1379981e6a4fae77d4fca73550db653d44b072b0307d45daa99fe14da58c803ee5468725b1b908f2d9073301168bce9b4807b99a19e1975aecf2d8c5a0952d18253cbcaed99ff2ea70d0f6f1999fa6a2e07d1a03182fd2d36afbee7d13f5e3dee30bca1210694c686099cf24d2c049320928d18d398540433070ac2c9d6d30aeeb8509ec08d43e0290058d17d11ba4f40f7d9a3736a8ec099e3dd4c84bdae1b44a7edb65f215989d36716da8c7ea2f973ebbbc22e0a49143df4f384c99f83de6e4e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h1e75b5bfb16bce0deb31ba8dc062503dd2a94ee8c2e309f737b3dbdf93b1894875cd85b6e52beaf65181f2a91d2e92fe4ad18ac9b8b7f1182a7a44a1452dfbff13f3858148e73a8928e4fca6a4dfee74cff874224484a36501a66229cb472f473816d836618cab6c9bb75f9372267f81ee2fa4db6f111cd5ee8fc1594c26adf61ffaeac327b46929aee9884834f046d197107505f0517d820da3ac6ec51b02cc5d8717d3e55303166d90993a45341a2c90c44c97acc1e13f3e5a4bbbf825ae412a73b84120b7490a09ffaaa8247074f460d4930f6aed95594767fe1ba3dc149f05b6c9e46eec5d56327e49196fdbbcf34453be535d7353a57fa392f20680d74497e44e869394bac055a61b17f60d64112c3d1484e7f90bfb51dcb4db8cf26ae60e5d249d849ebdae65f5933e4fa97dce165eeab546fd953372effaee2772908738377078e89c8b3c745752c389ae81b08adc95ce47f93be4d0bceb93f416f2b4d58d34f941b136fe0a421ee02386e8ef1b8ec9b965d5fa378c17bfc74f0cc6d79390cef56d68c884d597af65a9bc99a6ef46b96e123b05f8d3e25fb890a9eccc6fa193151e35b4cee201bdbc52460db6d3a41a73636fc3294ef64df01c07be4885aa7a6e2dcf4346cff313207772541cf5a23322de6ada60142b3d6cdd62fa61934a69deead82c7ae8b8e4d118d52758743b1de8fe0c8ec5e9566c77c668276df8fd8e5ebc289e30a5f8ccdd0952ace2f617fe367a535029246d93153d124b54c14ddb844b3ab2385eac384a36937f3b82f2add56e8083c8b965456f48c959c972f34842a4956a97415602ebd0b4eeca60cf0d191d33bc2aedabe5952141a02d4d8308867795cacb312080ff78a3e18ecbdc245b1927768a0a5b0c96b0373db2b2e17202d65f63;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'he175984c482ce2d8e118bc87d87284b6b9d67eeb3b6271e783d8d24a68c4978edb338f298fd03696e4b1be92e19bbd504f974a8b52c805d6791e3a8af568ff2279d0387a042e79b89faa8220f1e1f0e6ca9fb0b2f96278e5194bdfff79168b58109be789b2a3facc064f05fa76691ca364b1c604802762d288b837c237f77af736407d1951e1fc40b1c6b8a4091904eced24e332491aac9be35b2cde02f4e14a042bce6c5f144fdeca06a70ed443cce4b9d1b87a30a0d2f9ea52548ef13f0e3c43c4215771cc6f093c534455f956b39869077dc29bdf16b0b10b3f39a6c9fce8aa4c993f6c0d77a24c4e68c092ee1a37de45a44c61ec6f63a79f6c756bb5f1a2f4b3e4d7ea4c379da50e54e9a4b9784d1d646e5505ac8959668eb000fc05ddb8ad93894b9a57d2aea6922d11a0b38cd84ce64641355c0b8a0a3a121a809d032ce23c44be506510db1799d7f5f460dbec040ed15ae100e23b65f056de684528cb4ffd8435f998405b0ce300fd109cb786c25d5d89106e8b6d38aae3e353831baae7fe0af20e67eaa7750668afd898e3522238e2f4215924c0a4f7bae795e74323a739d6d321f4dda5f8426c528cd9a615ed391a45905f56b71fb1b3a72730d864f617874ac23495e417db00ffd14c2cf61973857e9589e2b8f75c9c43d1a7986fdddff5f0274f3f92045bf5dc287add889db53674f91a606eec386a1d43c83536ef9e675606c1bd3b6247fde5295269ccdcfc9195b6da8fc94eb79d44ed120c4df6d3ecdf52edd328ccea66932c547581a74ef99cf6dc4450c14c4b6ccbd877d305d0f633fa7400d2be13b61fb390b39af18beffcc6f86601d4ee86340df68c9aba11111fa488aee5a66cf2515acd35165ccbc40c072d77637bbd0ce8ea4a3dd0232735954dd18579;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h8708371f1705be4fa70aed948333172d0474aec1b56d6ff030000d0289ceee5c11fc2dbca9d9887a83a5b7730b474c5bf415d091c3765baec61d0021cbb5fc3835ed5160da5e25640bad73d6134165760c3f36b628671d5fbbc57c95502f5de48c386f794362682158138a87f2360d735f9c843e46a893ab8aa067f1230349ae7698d9f440a8cd178aa508ca3f890d42935995e54027914494e1d2c152acd9f8c5b9fa24e35ef6fa071f3416c4e5d92baf92d4eed5ece5ce6f67909cfafa8c3b097376589414304b9726c78061d9cd4e0d2211e8c73c36799457b369e967cb812796e03e5136f64a10001b299ae06cd4c41288a88e3e558d0d23b13351c7a58df543d63107b04725d89ad09b879829ff232a3d10e919676bd73302b6cfe4b958b3b739e2862a53704c79ed5e8169d6b42ae0e829a7ee7f3034603bf1c0ef40f4874d530e51b9bc8803c22e32ff40c60f57243e86794ed895f31660b34d02fce94f7d394259bc11ec11a0b6c7e1f8707c17428d97b9da9d9cabc0b26c7994d4ce6c34f433e3123793baa4b725e472a57423f29a2b9fe698ab27af92afe99e857c24949ced9710980f69e6cea4d6ec6104cf4de67dc8c74619657c0438207199dc7876f888698e4b357b1ec4239e6ac3f2178d459798f073b6f2226e25db3def14d8e197f5bda098cb5df63771becd017b1104fca68666bfe5013c3a36aa8f0a4644bfddcd351defaa5856711fbc545c200a2e0c1e57616849967a278d50ccf40a032a3b92e076540b1681391a9f7b9337e0abe4e4ef3a46ac15c2f3a9873e6e91198e809f26de21e324d9333359ca7248f291a278a5843f2f117b4e913b89fa8779ecf38561335db7218d1f685e728772620b3b48a8b61e8695a6683d830e502c909e4d0198a9d190;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hc7ca3c7fecc0e8acd4e7b6e1467cd08eb09f61ce66a4bda130368c5f06771df0c0690506be357671b0460d96e72745e33749a1db5aca75de728a037e493a5832ad6ec953884bd230d9782bab1549042ced8767ea4b97f105dff60377ea096f14309a64767efd4dedd3770da2058f09d3a64b6d1a2d62d9e806b7eeb42b778b7decf52464d476dd0078da22bbc0b71b7f3ab7757d24b4fcad7f842e56af94a904869a030620756b66f3df1b0b2124280998dfb50f54c242dbb9c61abe07fcca9f887fc449c24fce4df15f1077620c5c7fd629d8bb267e00679d1a3fde4057788598909e2593893920035c17cd7bfe9988c1a2df4fd9c6365a5bef6988499f46ece2d57d8f6eadd5dcb3d999e2fa318e1706376cc0c0ab5969b9e0cb2940018e0ce6943bfe523af03a6724999aaad09aeea0a7d000be4e7cb0727f30588a2f46b26d6b5f71a5c78cef9db648e0afd4cf631b4a32ddea55c9e5ccee240f610899e658ad66ea35bff922695a0d372d4b3f428539b695995e8023b656d9566d03d333dbab44faf9c65a3b7f966db667c3f7268b9ca82be0e90d0fb63d5780b98c19b9e5d25ba9e85a6fb6c661a97af3d31c6d42df259866ed86c47489e2395682f1e4650dad0917712d99a83fd020ee7999df0374224dd310474e9895ca6f7b4dc3d017ec5f171470b67c21baa692f074a736ba23a3b44a49ad79bc32a0a85156161e9b359ec259428e99314a2b32439f2e7f55dd7912faff1746cb60dead9e23f56bc3927207a331a6aa1c7d25eb5ebdbbbe145962d2527c1375aab82518add158e1a2a38119041e62c4af10007521bd4784f526bc8a1ce7c31f480be2c28f59084768b30e150bf945449267b5c4c53a75e4f36fa5af249d33066a8d7c635f54f0786842edab26ea0d71;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h3283daa5ebdd1d1c9801f73489c6f49806d4fb173c7fa0fd5811c9043c2983ed0d6c20daf49df0b0bab71cb69e8271acbf837497ee56be61914e704d5f58646c3670643b7080192e86fefe84ee223495d5c9b95f574c98a57c375e9590890d6acbc665b5422d9b91b15bdab014878f5344c73626b543e54189626c2a3d124d6df27b3d85942d7aa37b8737272fdb2a8bf083c7c0f3af3afacbc980a964870af642db38928d32f5e0ad7edc35ed2f905bce95c4f3c068929f129964f64601e60575e01d6667a7d6e65160c52f0e067d9a112d008d26850b13d695467d8cb3d24b048140029b904620c023a95358c2960736619d795c97d69da993314e13efa23776fe7d0e49b0a91023ff1abb51eb5d8540a4a2b25592cb4425940d8fa5e870c48c4c7f7aa1d291f2d4c9b9db52bb6b955813eb6358df77371eebc5b28e88d8f1cd7499056744e56f75722ea6659e58d4b438e54e7aeaecda50e9c38b444767b0c292d68e9e698a692bbfe5004c4fd3e493b2a9af6bd0212d5d6c9df87b588ce4f275845b4868c8e0e55fe8a2e65d40a313c52cabf8ef389031d1eedae2b7b3558808f9c98fcf7cb22987ec23935254fd86f4f20bff8a1fe61b15b8c725a112ba8f4192b4ca74446d79f38e3eb2c6ab04f0ae7cc02173e929910c8e322dce7b74a7bacf81e33949639ac084110896aef14a22f7e4ce07dd519590f0a358847d47084c6a22d0521c2648e7ddda487293f7507ff750dfc4349e06a5258aaea52d3b3978a37b7b01d8542ace71dfc361b13bf8cfafdee458c0f2632f3a72a393dab228e27c1f7ddc52ec3b9ff83f97382361d71efe7d0f184cfd5ca4eb972e3b9b025ba19cb9fb8f74fb25a8a769ee186ba9c23e4f3378edc1cda5a7bb8aa6011b024e13c5084aa2bba8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'ha1c41c31cb48e409e0d830d1223bf5669e810409cd23fe69cd1f75677036b04c1cb5badba00cdf6e6aeb374061629457ef9398757a8a671b4a497d0a015ffe29620a0313a2ee6a90b4f413c5735fee1e9094b70ddcbee6aba428f7527fce7bac247655d0c32e3cd8a62c2046b430d0f129fd2b0dbb5d55cdafc404d1d914622b71a66f36dace97221b9c04e77ee770141345e202c021d8b0f78578402779f0806c5c77135a7f5c351b6c835db6e18fb159049435b8a616466f7d85f2892172763cba764614de540f71bde3f05e7d7fd2bc12c504f671c4caf8c2c50205f4b6468e09439a90ca0ae2a0ee0f31586cefab552515ae0a4d36a4b522052805d3eac11bf415cfe10123116629cee17634b9b13922bae9381254501f4e9e57a6e34974e01eded4a746b505633e5fd2b2a42f41f662de9f1d0c4488421c63a6cbdba72bb7c22029236e1774a4805aef7886cb56982de96ea6931b1b66db6f0f80adf15d03c6b68ba427c435554f446b4fc776000b7ba6f370c6689d92ba98229d5deecfe7b4d7a19c4eeaf62ae0818c42c145d33b19eaf268d84a1e561c2274312066c5a23421ad064387af17b11a4c173674203441e91f9532e8554956ca4e69e862212f74206f001c4ded6359a620fcc3781b7b6c588d65adca24c9dc858771778c1282d0948f0378e799caa9894233b31806b253602960cff6de52177fa8d6adec68945d68bd9a099bb80c72c79851c276f1ae1d3ad48d0d8776d377601c13b61d23f9a92ca2f15739b48982e31152a696947d130303d264b94300370e1834e50f90a6c5112c3a6b4b212f23aadd3671d82a49ec24453f7ab369dfa5234e0d8f0413f46ccd0c6fcaa7b6eab451428fca59f0460f3c768e82a7571d0932922f55ab73848d61df5cb85358;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h41f49d7ca2c0c2500d18ed9c1658aa50b02134d31f72afc0274b52b4e3ad235202358c05f70488d6f57e3793575b771fe25357425e377e3a814f4353f8c69536add83b86cdecfd5c6dd21bae0e1619af2da379e33f79e2fda7c3cef3dcf95318cf37d39ecf0b3121e42d8a672dcda96ed46a27addd093bee6c55c7444decf2da377c3887cf874dc1a71c10094be2817d4e2a4794e23e7031986daed4146bb2172860c2135d1871f86aed02ec0834e814e340d4ec2177f54c56c710076453a10bec43ff0f979f355703a35a2f792346fd26fc408318b02527e63404a9e52e639eb21fa945f201658ea89411bd75e84096536b40de000ff183924659c9a08c0920bd812557c0fb7c27a3e2ce7e11c0d4639540f0656580a91035c11113adc57843f355938e52e28c2de46265f22080c5159da2d6d6bdacbec54c918b9c7f92bd3b5d3744430a5b1e346678d052a8c122910e1558e4753dd9fed12abd4adc1665e1075fa0b0dd8b46a8c1eb2c8380cf6f94a2a8419732803fc161dbb55f3ab9b31e7a23383a4ddd987ad45db2f5c533a449cbf26875d8449fd742c26b51cf5adac06133dba1aa1391adc05d48f9f52ab7cc79799922afef679e952f11b468cfd42e6c48b9c6ab7bdcaec733afcfea12ee76f452120449e6699a4e13fe49efa18a044cde6c5eb8f4efdcf982fedb2368098e96ffb980919e40e5819637527487785cd058ae1799feafd1ff44fd8e1d0c42d33971463c85b6074d385477c5aa71729ed46edd30a56e8921e25ddcbbc61d0184ed51fd31cff2dc804a80392a47c1e974bec0b2c5682d60334bbb182c41cea731e2d3a259489cf6220588a556e8b2e395811bfb2d622191691eef6db1e18e890906f1510205d8a5b4ededd56d568a04889c91f75d4bc5c6fd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'he0c6d939562328a923f26907b43f327df749e53337a57ec7fd70341249d043ac03704a9d45ffbd8d551ece19b2d6f90c052e9a1d1dd25cb144dbe6cc7196296a01cfd4a2115c3b0f3cf6f581bfb3ffc04a77740f45d9b4b29a0962243a4312d6813efefea5e8471bd2203e60a629b16bc451d4d75f0e975eebcd1062b5e1d30b9e218d0158e2854a0955c4db7abd56ceee34fce33050609e1fb2065533e0e675eb60441be4e87b351667d7735384d47213c8edd73dddd54b805d5850aa62fcd2a3ab64569e7549ddbc17bab12d4792964c35bc50297f336c3d51b7f650c5361a563283b9c046872f39c3e45d5b75ce415fd71f02998c76ebdfa0fa2d745501a4c19cb1216cd2c58293a9f55f8163222dc54df6cd7cb1715905edbb198968134d2c5de62b7a0c065e074d1af035265e28ac96b82fbea0b04d14ed515ed42576d1836fe219088bcfed8df787df2ee459983baa50e0efefed4a298462fef6bf05bc79327add524cb40f36ca64292d1755d32fd7f6a67c5b2c8a862751eab176ff28a63e5fcb1d4e28859eeeb6eb73d97e4bbac450477ea3324fd3fd7333124fc27c8ae159f9faa1e2bd9ec519c1b46f95de0726bdb7c4e27ad84129f4157b1e146c8f04266f7afedcd63d9c1019cb2750e80ce0ab46d76b4e952264988ae3303139f81cfbd603e0d19a493f3fc5e5c394b2dc5ca52421db83b0ab280c6325c77b358630dcbab6f97142cbec8d86f0ddd1b8834ae70e31d5ddd75e188eaa4f19a479a61f716da85aa682e52f9f44d117f68632b6937ae7f375507e2af2ebffc6de25e3061e03e260059b544f20f6a2fb85d9c8b13b5fff08fabb2786a0c25b03d3a58e6463f8f49c2bb544ab8897968e9b42968fc5d75c2be1838407647449caf947716920a6d890cb1b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h130f1824bab85c998eeb7b93bbafb56ac2c5d9702c7808e33d646f49ca2e2922f167a420f8782ec8598debf3a2b91f9a96b10347113845c3a907aa1211ddc1a48f86be3920db302c33983d315e610c403f07e44e7dc8c9f63991e324360b577047bb87f45ac1f639dd395fe074537dcdf96b3feb452efdbe4248ca150c79cdd815a1f5d8e92ecc098bd53d7540c6d99c866d390d42ae9e370f4d93a07b5be70d9434ecc2f7e4746475a186cd53faaabec67e6f5e7cdec8165096f9af18cdfaad18a43fea129cc75ac8ddf1c2f99af22237c2a2611aeb42d3872d93113592847e3a8c3d859ec5efa3fbc7ea768c2bd158e88f9ba7d75227345154f33dab09598682f0231c16986bbae3fa5fdfec2f3c14b28942514de0f5d8dc5af6a6a5f6bd812457a0bb49fdc2d1f8afbdd3cf0dc21fa57b1316f1a3c1392a4e562752d09a2635ac7b86db44ab9b4e088f4c356c9125743723236518683390ca7b308b2361e124c38cc005678e78d8d81850b5024ad8edf16392180260d9dd918bf9bf2182c1c25653779c81880f4e3ea7981ab79b89f89281db492979feb179416d98310408091a53f30a684a45b68bdf0ebcff99e12721371189953ef0d94cdf7c094781ed5e604e9374e5122e86f45ca06c6c799fcf63a64ead0e81136b3c08fce71f24b283270b17c19610edc272361cd98a39f26b5b52110782b179c01781d96d6c7e987aeeb82d250f57be73bde1eee2535dd7ec837a9fe6a8759504102e771527da2f96c0e70765be60b73838619e6e3f263a9d3762cdb36545d85fbcb9f2b780705994d60648af19d903597cc6d6e6ccb4e9069f75fc61fbac19ecc4d7650eea935c041ce8394d383d7d6aae71470e2f086c05e22bb5386c90e40460d4d476646a34aaa384c65850ac04;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hf0b997accb0ed5ae99a846414e0b15655dfecb88e93e165d40653b9e1b54ef0e47438cdb144f023fe45eefaed4544cf33a6f7166dcb0e3d8f2561be0790ae1a46856716a32cfd9530ad96e43d0e7c138686dd7f45ae1578ec5fa085e401b0228ff4d5ee16b5e873cfba26ebab4b55f393ef8a488280c47306d8382a56d25c820d26126feba4b8b59424cba47151c8eb9e8a76395885f1d2bc56c85f5c171f51491fb925f8316da9006c9d0e103d46e13ab0e0396cbed158a42087afc887a4cb51334546a2dbc97354936688d1469186d9fd377b519e3585cc17da37e46af997e786c5e32c74dee47ab0574c4b56c91446102d5d7d206d944013fd01087ee39731adef1773b886de5674a264bd0e5de869bbfb27171979e0590b349c295c661201fd9bac20b9388261f065b63f4f125139b5e74cccf1ff896b5fca10abe98e49fe668bacd66646c5ff4ece98102dbc07a8a5e0e05e4016c98e42470ec963b7c7fdf14b61031d254bee593855dc3d990492ceef2060f4efbcea016b924092fad38358c46ef1a5babcbb4d1b680a89765d4892763495be8cf5f27efe3ed356384f807b4b96fa4ae34d811bad408360ad3a412a30234b7fc7e07e1a11265698947bb48addda1fcfffcd3740670f9eb92bf56f21e2d6a28288d558aaf4b634f87198855b0c4c5fb8b57365aff334fb9676e3cc01da53a37f70b606489888e252bfb200b090a2a632a14ce602cc765284f9d9eb06ebb1d7a3c3a2dc18778bf6d33b152fe96cc1a5574125b41f206b98c98a7496c0c9278d266f1cc7a32ea6a175e1d9125830ae02e6d4000950f73f81bbc70df0053d2cc1a4d4c0d5b63876610581d1113d88d0468417a3fc4b6a65ce1d42a1b4eaa8698ca882930f367e7e109201f16aebe7fcad3821312;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hfd88a3db737f1ca282e0a6f3059ca3346e8ddcf5c0b8b49d45176b22dae97362bd30e036c8f20f2b65f82922e364c8d41967e90fc117e9399ae8f16b589c3eedd235d4f0abc82ec7b302142cef11c0d11eaa67cee16264bae67e745cc3423b9ee22da2b80c46fc0408bea5e8f2d7c50227df95b769020790669d7e56d3bd22e8f9ca738efae567d4d35a5f756a64014f90e339d469cd03ffb951fbf2da8c526556dc5ee07249cc0360e8b4fe21ab51313e26a71b16107d1d1e096623d6eaed74c2c51e2d422844af74f3d3269c60fc30b0f4a27396be14a1e7ce8a02f8a509346731c91c93643a65e1f5588344afc046a71caa4a1a72004c088b53fe35c83ddfaa55be0dee490da11ef91b5c563ace9ff185df611cf60c3e30b244357ac0655b500883348f2cec56de23c153f26ae05f4c5a3481c5147f4e311a5f8000576ac01deb99d92b48e3a787f15257b6d97a1e32616795cd7ecad27f324d24fc852f3995fab08b8b4ddb4772cf56cfd980c6e5f2a62b8301270af8a85666bf64e1a1fcb692c5bbc16191e5c1944928e05140b2285ed77cfc116a056cc2e3fa69b393b320f761c0e5800511de3d2fd973ad12ef34c32be3fae661e706d9ebbf900186006e7c63dc5e85ed8817fedb25acff1f07541fb8726ba73143f3b88b25bd2878ee4c5b7f4daa1bc87e9ab0b024ba31490e88caa62f6d3224759221f9dfbf3b1a4cae1bd78190f6d72bcfcec76d436152f68901ef75c3c5cd414ebeb1f2db991ef44795513727fa183970e657ab04fe364160c39f11809440c5d888fd4150304ca957c1710493591fdc81b38e136670fc821be43c989ba72644c47225a10cb40e24ce4afb4a6b03f49bf689c14b0540c5d4ba34a2bcfa357109a4d56fb3e4746bb49392b89fb9f1eb17;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h5dd6653e542e1cd0dfec1f7d86ac1b54bcc6e4a3c85fcde3b3f58e60477b1175345e0e9952d7b413e1c7036cb07cb4fd009b82cc4a997744467707ad31f1856dd86b9f26c3431d0ce15c365d4edd0e05011c04123ce5d8aec62c20aebba6cbaa1865a32d34c80be39b203839bb38bbf1fd8d63d9ecdc737c17d088cc9b81cf392158b8801019011bc212c03e4b688b3dc0747dabe5834954da8bf383af7b38c999ae990cbdb898aa759064b4524d3b377fe65a4a40bb759ccc7a419abba0c1c313e5501f164a9ef53d139bdcfb92793506f43d31cf96d7c2fd5fadd15fdfdd845b590be8ca95c98cc42719f2ce4e38922f2a8c7dd7790bf6b74e9b2526740696fde3eee96f20945cfb06a811ddbb81b9c27a5586da132b5a4273d34faed5527cbfc22002987f08f82d21430a01772166c97dbbf8403be986ffd3c82975dc2c214a20d417273e214d4146245a492dcff15d5cf872a9a87ad44d6ee76f981915c51aa323d9da4abc42d190f9fd314d362adba1527b5d7d310bc91193853d09063bfbc7918c1d54bccedacbe5176810bd5e136894c95acf1e86b8bce91f61aaac28162a713f865a8735522b77b9fc5c740f80e69195fcb9cba1869c466481302056db61b193fb115a6f45147e1001e10406ba41e7ed742ccf061e7988065542d60c955be6e5d1f64de34fa626eb331563b05cf43c12e9692379d48ef960a8852b95bb6b3132199248d7e2963316df0c2ab53a523b5d2274c7d3485fa84682fc7c1c14fdd4ec7c4df5d82f0390cbaea15597e7286f4131244416b16e75bfffec982922fa3f8d0164c56ce0c4c2fb1961a66f76ac720bff52a57b128dfcd93a527d9504903cc82f232d4a5ce2c3e192651c17fc1457f9dfaf1f2590c3ff5864fe4a6807ef2e5f528b29e2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h38b0fafa677ae398171d7611c5be8894a01c432c6c5dc508d06bfd8f358fbe6a6c7c29dcb822a90a557d84d4eaeb2dd81b5fd58a739352c2ad4ee6f0f710d4ea496b6ac0b10c9cfa23d269f96a1c808acbdd4f4a10ce5ad80c58dc7ffe47068c30fae0dd2b61a45581d3376cb1c242d8c0e8a839da7be517e371974f880e3a8b4b3e82b553da71b2168711b9852418860511c81b355e583fbd8e4e7f68c10f14a770fff056da18cdfdf1cac803ff47a3c489bcbd69260d08f7dec12c279be8a7ded21bfaeaf5e23fcb8e63cf33107b22c21d6c8d44bbeb57225a130bcef5c7972f6f6581882e2999c00623ad4333afd900b9d20c5a18c20696dbc691ea326eb48964e9c1bc8e6024ea24ce4dd2b9f7a00315aaebe62c30d28ae1056e1ba088c6b9f935fd3b35c8227108b7ecc651c225d4f425b2a64eb001593177055cccfbf1113bbf780ec576249bc073fa99ec668890cb29a677d0a0d953e265d428a055a37acd2759267ce9083f9ba1baf5e45c7f64a2c7eb48af68e82dbf65fc64491e63c5f35953a1f5f041b8bb7eb51c18473464dbf65122f9ac6a64c9cf683c704ac24f1fdf852f5c733b1f8b6e04f27628ff5d8f840d78f0a5666f23074dc7193ba038bd036bedda1048882e7b5d0ceaa4c75e900b20458c0aab7772153218d4b39f5945fa13534ca5eb60811efbbdf0700d07f63d60a67f73f261cdd0ed93ec99d5f02734c548bca8c29dd29642297ffad1dffec52146058c3875de5feffbc546961d0b4f07d5c57b53ab9efb5ccd7fef5dbdc6b5b3fb09dc10a79f2e99df84ab25947e473a12c57a1ff02ea7151a256ae5edc213d481681aaaca21842ff6cebb29f026a8d8679175c8e05433917c439afb0ac6479fffd99ed6b38b9187503b7bd55b4bdf02bbd2dd81;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h28ccdd5fffc06e70292defa77f6dfc558b5311a67001367e9463a1fc44174f9c5d8f12a2d10fe3c988943c6c0bb7ad90838a2d1070e00b09550ac4df7c49c088821aef33898072a9c57c1eb41c47b9f98665067012905ebac0d3f6eab7d798e0e2b3463c33da6c5180abd314fcc0728270c31a22a48c5a0500d9ebc1ff53d82f6d5da68eb3c720cdd68c328bf1787d2bbc119dbf5a27d21a86730e15cf935bbde7e454034c564745e0384ed0fc567926c8d6d4da6e62395c92aa0e8824f504de813a1a1a5ededeaa1d962571b2723ffa0834c9a18e0c72985ba5dc66b4f55ee65f3b099ae8ec09dee33affb9c23e656212b74dd5348e3aa5f643c78943be2c55fad0234be67e1d60b18e284f0a05ad967e9e0132e82181c2e1848552a023188722896b7ca155dd271bb8dc45b7e3e9b8de7cb2086f9a6ac7addecd336a06bd40470b044f601b8ca7369b1822655b9df9365429811883ffcf524137e3bfa4f4871f0c239b46c17387d1eaa8ea2239eb9ed231c3ae8b23fa293304936e0abbc754a75b2eadcde463c9d62f4b44e5d0f3d919c37cb269a944b1027065a21bab1ad73a5d1d57a7cf9296f0baa6c6b46a7694e21354163e0ef04bf3a74a4135eca422c169dc7cf1b121e35f608681ce58084ad19ff2119f50973bf1c78b821d69672a30bb7f77bf06720e42e982380fbfb0788fd81edafe5dfbf30e7bc5a3bd8d93653c4e5d5f97127caa9c7d0a286ef8350aaebfae0971ff5deb801a581f4a07476a023d5c3007b9e81e4cfa7cbbc1da42604227f9dee3e8aa937ae12b2bb9642c771f50d716e14afa3c7cc3a818d3724665f2a3607c766f387d1d31512ad6b50252b5fe83b96e13eb86c10ba2acee9218817633e6659d7103ad155e787b1629bc0c44cc8defb114665f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h84b420294fe9770ace0d215b0d0814a69fa48d0cde305b82174e34e1d64ce0619968738f7b9d9ddcf97bf080585498bf9a4ff428a38f152bd7538ef05ec3acbc64f43287c6d99b90a614bbc64b0460545a0da8e21288269002dbaf6097a7e6b7431b219c0a3e0b4f80002470cf130ea5e1dc180216acf813c2cef66ab1c77ef7c8830ab6a4a97dee716d2f041991858a28d45fcbf4a414582b3357ff92180d515d34ce5ec92353fabf2fdb7fb280a7c046d034fc16e52943db41454da852e99d12b300d9d89f1e0183563fc12c5cc8d482db7b4c398c96526a50b2892662ff7c83922f4e76221da3e0c033cf0b5eaa31dfeb37ef39bad849c8b65903b56edd0c6d7be38853fcad7ef6503055ab3c95deca0cbe05ec0514433e2e372b2a3d178fac4e02b06acc3e08ed1c72c594568bc2cc02286b9cbdad142bf214d6513cff7c858890f63ada2747b7c6d1f7107a4c02bc561a9048a3d938d1e2c00ecb057c1902209f0638c79bfbaedc92f73636cb0f30d630512d39d2281dea1b4189f176833c868dcee7c855773885388a7299edb9fbf26bd67824cf53e240eaea15699c2d37b9ee6c514344b4608b7aeecd33ca16f78f7817ea97428dd11e52943978c68af867ee49d3d986b1cd1178553d70d1d3350cd79408456d43d8fac61b3796ea4516df71cb6a016e1cd8135e059323da754c3a79ac270561b5ee54e0455e8ab8848a5abe18779708d99bd744c22c812678279de7c16039c499fe84b164109df90ebe3eff41a55214ff18acbd9e2692adb441452c1a1b9188e685d13bfd33f61f2c746778c6992f17e578d89f9f399b1188f4a2713885564c0d088f287c1d48db4c2cef6653b3f87a91734705867a42892bd31a6333b967b816b434674df9a61988a454c8a76e626616;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h7c6c25ec117a605b3fddca226f94104e3369ac8c506a7c4dc5a99666f96fbb1afd870b2729cdc434c0a691298f041e1ee41ecc0971946bcd7cf36c5e83661e1c40e7828af9c90f69338b57ed1b3ca6026e0ccc938027ec5350e83aa25ddb8b22f660127a3b847058b614e7e5b2da242c59ab34e86bab89209e06380429e31c62dbdc3561fe6687c4969318f1220f7e76f7065d3fd27cef19a62cce5842cc732358a1f39beed566a28aa502dfe7ae9ef7e91cde4b242f8583e2f5154b98c74cb071b8cdb891fbe04913e504a900963bb7b40bb5296e500da3029c4786625d1f590cae5f9ecb574933c2ebb19f02c2ff8ac395c21a91946c4715806addb543c8a0c3ecdab2d2ee9a3b39c457d801b8db9fcfa138a95d683000fc24385d01d106e7b14130bbc275c45b9b2c5b64a674882b3cd2c194334f0f42ba0cdc3081225658ba051e4a75109fe69adf6b6a67463688682c7e13d1d51801672f72e2989880220506f8f001c568d433fdda7dbd15af7a210925ba8a1066ec9643666d0d263c8014060e54bfccc9eae9b312e501d8512a5dd99924051d9f6e71d847f2690c4c78ec3046385a3fa480e0dbcbef641e7199db362b99d0f2deeedb1cd63b332cf096211d024b7cce37223682cf362fcf47de98374f68f2fd07d28446f049bde218a4ce33f667f05f5e3d93eaa1cb471bf907f7fd3eead6a8136dba941f552b00a2b47da0c5ff9f72a3a773f501fb64c7e190e16ead815d7507bbff439685b1edafc37c1b623449ed32f2bdcac5b2a100b58b4aac2f4923303f20016f18513a1c539aed70ec2c435276bd79a8f8bcbd05d0d5281e2d5996ab869ecce7022cae66b1a5441d5e01d4d72f004e280f25576d690a03521424a361cdbe3890a8beb59406d201963f8c5a8780d1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hda3a5fac658a2136108dd1243bf38318c567ffcbc0854173b54351a8b7e439a2b583bc8f4cbd6f08ed7574942e858e099f2134b5d579c0b829540fa7a41f3dbbff9dafc379c3f75de9329925f1fb01d057cf5dc9f1afc24b661f04145eda4b55f99927be4eb630b81893ccff0a5008a5dbc4a701def51a89adc3c12ff5f62c1d0f727c8fd2383326186dbf32ee7d46cf0dfec7df446b411df2becc7a0e22648dd509c84a8f0eadd291ccf17eed736b0de1a4b8434910e45a24306500458db18537f5e59398d8851724efc889959a113a86ce79395affab855ba0b3064c6fc7ea235e14183ba4151e4bfc60d6fe5b6b55345cac84d02bc414c900873dbf05ad9756f132d036bddeb4ff3e6bdecbc4baf64b5ffa867312fe21e00246ed70cb843b82e07e4c38e74df410338a98f9a03c6ae4f536f5558167200e2ffa6f2e4d7b49300780cecf4daaf297e9e733f6885feaceb3b8f3d404d074efdd8963cd9a67004d6b5cc621a721746b36782bea84d3a3380e528b396fe2d0231cf47ffcab7253a3d01d93ccca27f85eecf4c8eb30a088214eadd8b9658ff41fa3fd814e17bb8eaffc3162c36d0d7f3c5f5fb53b230a0725226dd75212317acb41c478f056a795adf5aee50845e38fb2d99559af45663617e0767eb6552725bb582212b8a41c0738dfb27ab875b9343ddeab561d28edd146ba00c927f731e3c0b2c998d7a5d5108f699571c266041b7fc07e75f1420d619ae1318917b879c6c98d46e9c17dd04ef40d9001a6aa539ee67c72b34c035cb5120b83b1a76e3416cf15338424bd8ecfc926bdc44097082c12a28d4006e9ad5381b6d287be78631b995c6f6f646cde5694924040ac57c0cb2506bf3343fb4430b725807876bd4ca8e36ec3aab88b66eae3c9baa57c6de2f2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'ha9a9821e578c984a9cdf3e5f7935ac7045688a8a484e5fb3283c4823ddbd0608c58a35c6276eab6bd9dbd28d012c634fe7760d8392e311a70bcd8dc91f9a3bf6556f24ffd19b23859766e0b04e03ccc05fdad79784453753a1b23ded3686f4ff53d2c0b0c103d32f44bc76bfbca848c96e159239ba53215be65cab687ba4a910739af4c01767062f87f4f33430adf67768a6c08c7870899f27c1a10cb5e513ab59244227bd885b4227b5a2ee1859b92a93bc6e0f715d7d7af24af38a872c64c57dcf891c8ec165d3940fd46f6a83c3f37fbbecdd752b886498930b6a98b6c5ab5ac6d6e44640cb64217cfcba8e974804bb243861c5c70514ccd1c8f087480797de72d8daf631d6b518464ddae8685c67f4dee599c889fe81bf8c7a316685d970f4aebbc2f3bf78e468275f8b9b93fc9da7b8534aedb939d0c51b7dca3248e950923af85523c436b4b2d0b83ef154921c19014d31a55428b1a622fae3b271d4b977d685e903eb5d54fe75eca753070d7aa559dbdd78700adcdfac59ecd085b9873fb6caa2a5a5b5ba0195d532bac372f984c3d61cf800d71e1d099488f463cc282589b7ee89941b234b16ee588c114f88651633bf4fabc76d6b230657a558ed67c2e4fca9286ab4c111d18f3739d26411bf0b40528815ef782e4e87a0c1038fbc076c696bc9b2bef4f2502b198a7a0f984bd60bcf7be2ce9e2b9e1aaadd33b8c834c1a00eff9c7e9a560a5e6f0277bbd298c795198c4276517dfc6188f09eb8010d1613928b08ef66cc84b054b75e05e92c15c56f4c0e4a537ff309f83d09afdfe73c5c42adeab9369e42b203ff664bd2606882abc3f988b36a0a80e19a8b5e13d889b010c5e9ac7236877820b2093614b9bf55370612607ad9f2e276ff2a126e6f2b5c918f540de6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hdec69e6401cad509a0127d2893afc1117673a547680997bf805bd6c85ec471d67d96b75eb7c5ad4fea889c5395b2c9346a6c2bda6da86320f2c2603969da0df963bbf0cee7b95bc339ff06799f003f0c9678661a8ace819065b6b68c7b2dd133f430561aa9e99dee59fdef73a36de4ab468414688eaccf03972265c2697f2af0757bc63e57a3a1e6f3f91fb4dfe0b8bfd00bd336a6ff2fcffeaaf25fe1e62ccd63250b43beadc3ea35ddc580283de3338f5904eb6d3093e8c99f8538fa90cf15eb043bfe51937167bcb5c7cec977b309bec06f0cc9acfda7f5d50dd101928e46413681fe52001e12967004d5143c216974dc43a30482ad28f0c5f3ada582eb7a332ce97fcbc983bf767082562f1619bd7e35b233476061905a61679ea3f33730482c2afb27c149512f1a34c6ceb4f707accc36cd1deeb32be732953fcd1f89283ca76686b68a4133c65dc20a5107d558cfe46f8a8bacbab8613bebc4e5c907fd10534e907426a5d3ad351e2f13f7d52d8978af84d3bafd9ac46cdce604f355669491c3cb50b15a3f31cc49eeaee90c88cc9152438bb40d9b02c26adffb2712fcc51021cd06969d0a0ee86838cb600ef442b95cbaa4540b98c0d1cf8f465c2276f81e59ec1450d8c651813de575932ddcb35b7ad390a2f6991efcc3e8c9db26c3fd6735ae2ee7823734c4af0221601dbb4a4ca391537412a169b670bfb0b086342203d5f06b1a17d637068672f68abae14a6b63383ee34147fdb61f2e405d9b6a79a552e65d0cc36829d07d057b3634ee6c67f55dc8e5f3dc407f30d2509ac045b4ee2b5011f006979df217f4c8c869ff44d348e52618cba3979d4c08bd6afd152fbe0ca3eb3b879fcb60e05e437615a3fe8ad42f6f5a5c0e9186d6cc3812c4b5b4cbff2fb1b60daa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'ha76ae12778ee124a6fec451268ce123ea0bd8916dc8e45769ca4ae27f8b7d7361e67f071f9f990472cc53a505eb0a16e472c65c73b1643bc7e9fb2e14f7fa6224ee5e47114cdaef0a2c5fb5b3aa18bf88c19a2992907b409ebc92803ebe25ed93f7985b20fcf294e54c59c9228c008a2c80f5d60a06da905faf3b635fa68d0c64985461536c3bfbc6a7471ba2d889a1e8ae9e940d6422365cfe33ad99e76046a8a8da821aaf51ea2bcb97453944293a34aa16319c428c4bf8e45252f5eefaff521140b00895d97b8074cfcb98ecf34f6f50af16d0339a3bfe646e0aa8e4a01462551b405b0283659325dac1d9d80aa0566de06202e976052e8fb6d2c36ef46d65ff8f0f24ed4b5734a787d3f2efc5f85b726867f1822827235965e33010ac9a048ef8384b9905c407bdec904cad329bc11ec27b8ffab7dfa46f2d94447bc31fd9116972a2a15e0882b6c9ec9cb5762d0b4a88335b01713e2dbe128a6c6fe28d391e5f93b0ae9339657a8a1c0b93c19c9ba762c5540c5bb49e5bf465cac2f11a6417e5feed954977548784f1711f231f27f6fabb6340a6c0e04ee9f45e12902c6a8152076d7572fce1eeb7eb3416f70d68f87bf1a277380ba98e6ce23edf1133caedbe2046b5196ab0d9f294c098acfedd5effe1e91119949ca4e6345aa8ce93eac2328c7aa2e029cabe5338ae6dbd0ee492258ac7a58f6dd84e63a7210d4f3c5ac84697dd39e16c9a2f636481d557f2b60ee150e55e7ff0aacdccb7b18a1e92435064f9a069298a3125db8b53daf9ee268bd333e6ec6b53e139d726d2e02a867a2a667c411da6421088de0bab6e67ba01c3c593d72057b40ac04091a2597a3a6676cc8d44e851eed0bb668ad9f83e0bfa8c1f74ef8206436b62f21193c3d309fa008f46115b1d96b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h5e6c053f2f5ac0a7894e3f3c6c85d88741cafc3c2f6bb271871694b164febc2694eee0eb31aaf9f67971f25a77d4ca01d4ad2eac67f4274b9d2d171bbe069288453c9a5e3949bcb81632c3381d74fdb0c751d70857f6a06cf4a0c2b908f74cbd91b7893929e987070a607afcd40643a4bd2c33a929a1bd6345ecb59559caf86b4d4e7df56a69571ba262ee0891fd39e7487f924838e1912f1ccde4152087095917927f150ab6c2502a4f8cd537e7e669f5536eee267571298ecb189908e2308c88f781660c14d70a6a6a7e592ffb8cf1c5cc067048d6015327b90506db6177c4160f6d7dac3baac79e2fe8df232f606506f44ce560f958af22a0ef9837a95677d97a49655dc984078219e03bb035684444f562a86524c08d6808c85ea301728d0505d104c36eb4ac86fa444ae43c8b0a997a6c48ced06fcc5eb5fad652bc16feee01ec84ac7c0b58d5f954f0a4f36d4bc739aaf6d4c3079b6eb4bc85dca72b91b402d4d6f9b0c53df8c4f703b477b3e9397cf143b2ea50a77511880acde479ccd331e6d1c2827c39ab36d938e1a83c7a49ca8215f8dba281696bfc615fbc04d673d4f913e6937a7f1e7f76018eafa6fa5faea52659f1676bde36fee1ff2e1b320c8910a41a2f12c98352dca83ade7921806fc46940c17910e4529de42a4769e59deccbb38507e5179b594a66d505078e8d42964a0cf99bd041377604b1314c463c5697576bc45f83d0f36f3f854dd9c24f8a3c547bac1bf62a3060e1edd74682dab9f2e8c8ec07624a7d865dfb29d2cf423e2756795cf90e51d59ce7ada8d3aed8d3fa1c85bf8bcd2573f0beb1f942f25bf79c3b3ee68698edd548a697635c9627f7e762be85eec151dc18f2601543894070e36e79a0802e96bad7a2bfb27808eeeb573572404829;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h48bc189d9cdf55678c92c829062945fe6280f1be77d0357dcd5ed690ef49946df033d1791eadc0dd35e5bed598b9531c35ad1df2cde0edb1bafaee9bc0f4c38f98e3c7f7c272770e2c959d3224870d88fe0ae38a360462ce8532f0af06e818031c9f6ab5b6db65b3ae923710f2e8626527bf0289ca516872d3a29a0c7f599a044b006c76b084937bd73e8d121cb768be36441d19b3e43bba9e304f2dbc6fce5f57eac66f201180d017e03cc379efbf27d0c62133092dddbc6de68a651d3cea0db09fa19a824d18cabff956528978ae7d22937bd58b6aca88fa858f2556202e0f805a93869271847bbf2b26ea1b26dbd67e8377dd748ed7571c2ac358cf8c9784edea2c372fbe732cd00ebc292f5ff8e2375325b36ad151d9e1ef587fe4e0227e5c1718aa6aeb0ba76300a9790c425ee7e4c449805564d4f1e7991699da9996414e09cb81c849fa711177ee169db1e12c589567d6be6fe192e1cb38006983acf20b8958a60c4a6fe37c87ffe017be6b3d1e061fc846a25a77f60330390fb00170f379f78f8ccb4d738463d83583da4e8232a3838631ba908142c1c9faa68c12940e792c737fc72e5420ad214d769e6eb28c6e04edc4cb47e1cc3fe5eafa682b117065b828173085b14bdf77ee604dbb9d7a1d9e466e6837af1dbfde82628d5bfd9497d2e60a0bfee9bd3cedae46f619b06bc7df1d097b182661222641476e119e9c0621f175167d0009e05add1d2ddcdd11da3c044bf60626b6a29bd378898d3bcf77b3f8104e0803d4a6f41b52a936a40147af4a1c52d276363c886cff20af9ed7889fe2f2bff167d3a12a5487f8527516617596d43d20055dd08bd0c7cc6b4d28ca66fcf1893a2aaa5b65c8c1528e88250b98481d52019e6a42104d5257f76b140b89e359781503;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'he24a13c7e87fceecb109a910e789f8aff7ae4ad0e0fc7f146e84125698dce01c45a73386a6c609d8ce79e077737a6f1ee9b1a4bf9e95b0937f46fb396425df464e3d88e918893e736f5cc3d84cb9b6dee1f6759f0258698a98c0ecc916d92c5906307f9a58954af7dd8191c7594a9ea876fa899e2aad61263497cc2d0e5ba3349cedb1706ed51253f914537de3f451333c68b6f846419b974f0e000e934fe8678e9e1ab01f6d2f3423bfc61b3f0cf0fe38d71707826b7781d7c302e04b639c40abc4eaf6e39d7ef4373fa317499c5f289053f6dc3a8b7474c9eb852066ae7fc7332dc91acee7f923b80b82ef24516aeeb5136ead09a8d3886724c14084db663bc9590b2348dc8799da70113b04adb7e7a915ce8bbd1ecfed3f6cc49ec8d8a6c51495c181d90bff0f67249ce8918926700f8398a1aedd5bb89cc03c5de67a5e20f38434a62901bcc9309497e3c816fffae25b785f58d58ac0f04d30134af32fe1f4b6cc349ded539f7484233ee836bb49a27f8452e3b6b833fc9b810110460af16e8ed06f78a034b60d097676d5bb8647780b1a4311d42c81f1e878a0de50a613e93626d3726e60d53ab0ee5b6e0277e0cb401145441f1ce30ecbb09948ad3521d357fb2da2b105334a1b74c6c6e946618a8937ea42bfff873b0ada1b1189cc0c4931fb615a35cd26d4fe1744b6a0f16a7ab6d31cececfb05913c10c27ebb60bd280f060f686be6ada1bf753d669eff9b092473624d31a149d3b09bbb7c4b6187c4365dbfdb2f7aef240bd9494cc93ee7cd9aed3562d64fd0f5ea459e43ae9a5c95e386107f55bfd2d6f94d72be2fbff866da0b23d6b0725b0dbaca8508d3e709a27a31def9127090276ca0e258c3cb60b1ed2176ae313ac16c9989921a6bf129b3eef0f9e263dd6b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h276b0f8a4d030f32a8a663b8bdf32a32a17ef20902a05196ad27fb07cba0b4da5af0db91cd7d0dfb4068c9424f906a6544f3ff80d33e4d239172d1bddd5d603dee3d3e8cdf3e17ad7f4cdb4e830fc2c186409609b9e6690cb40ed4788ba94dbff0637b65133edae455c1366d0d212d8121b346206f89a7d3eb18b88e6a842b14272337e1abdf1d0a08ffeb3638ce6bf5e29e6351a6957641b2c30c1509c68b4058d1033b5c029cab1dd6d8b27ed47345eb43cffd6fefb786b3de08a7626fa6d2598f7b823acdfb091256def13d467fcdce2da3644a73451e48a75d202a9c82395031a58035dfbe715b1192ed64473dc38c4147b9288066ca263427530413b54f6b706e6f6313d970fe27dd27af5464522fc7a1d340df8bb32db45d67079227c8d820af19e3c4779d854f99f6328b5f8e10fbd6505ff96febb84489fc9a6927fbf59cb178f55e965e489441112923ceeffedd7edbbebe5f202dd835644bff82f9e503ecec61cd0a0cb858c400b99f5c5027bd2751448665d8fbbe7ce662ec3b318826edbac9ad3fa7793200ca7abab613e852ce2b6900f40cac50cb63d16210c7abfdf46e3b739afb3d04fe99d7dfae86cd8359884786f4e8f8d965faa6d2dae6e03efca9c281a843e895964286ee6df9aeb65d2347f8bc7fd1eb526b50c4ffddf7ba212d114ad647150b23d19edd4a1921f13bd42b1a666be8adea872c3c80d94c4e366ee051a5d60c8dbdf9f0ddad2b96ac730988b6e91de637d8cba0b6485135ba7f687911e202e7d66ca7456b7f8736a40e1103880aa7eb5e93705416a38d6b2969df96dd2a40894b4369e7368fee6c41eb1edb717620b0b78fa47bca9d6a3c1ec33c49f377144f408994d141b3ad304cfe6f3c29120d08c3ccff9d7ceb7cf680c1b1c70e24ba;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hd42c55786fc988e4e2d1877b3fd6170f468bb2126ca02b1ec760b13dfd4f6a1ba76adbd943137cb9b361e21a056edddaf1c5bf71fe2d3a106baca8d5037df6920f036383d4871cd308d8db99eef7038c327838aa01fe7af9ebd91b80ca6a0ca5e8dd221bc2bb10a5540f43f6c361dd4ec1e14526e2c69318101079a006af176a06d927806425e2272f41fb1559457b367f2412f77217083ff088626341c23abcca441959c592c1eff3946d795dc076a24a702c61e88654ce0dda8387e0a2f3145f90249cbbdb2be17701e7dd18ab4bbfc5f77ee36fe8fc514990c6bb89a105f8f982ec1eeb5d9652be3a869c94dc85f6c6622dcc55b994b21d45586548d4a874a0d530a0f5eee31abe92220c83ef4db1eeec2d0e5a20d04d791d01c6c54a2d7009a670bebcc27784993042e81b70bc2b1c4f8e71b275349a8ec4faf353b652bf1454064bb157d24f842ce185b42863b80e0d535d77e189415b31821080a0b25087da3c6c782ef955cb04aa470e0e95865049eb498d45c19f95640ef57507c20ae80b3b4d20fa08c76474f82a2d93b5f3ef3ceef90810501d49fb4605d972282c57fff8cd60f01adbb5fd79f37c34b51ebc1374c8a5fd469e76ec748ea5ee7419b469ee296d36c590cbb54e5803eba29a0176dbd6ed82c7394608ab76a0e6e3807200bd8f8132fa476d8d1b5c47cefeada955fcd543e78b4a4b48e390d2e5a14a2b91cc45ef1d2df152ab73a68fe022eaef51ac866be7a0067788830ca74be15f8c155657f9527dbb8a86c5779ea00339fa51cdd2d4af8259f7a0681fcdb12edc319403dc82f8c82a483f1c38143c553cc5f9e06e6a8e81ea0a9372e8e77046664245edb017986ed8555a81ebfa7bebf57d261d9adee1a2f25b5ed2c4d93816109f61fc96083282a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hc0aa53c8eac46d5dc11422464ba5ae662b9cc220a2e9df7caeb295bd74b6f61dd35383c2e643b9c90a5d4820a764f3b5740491b8f75349e4a7b3953bb61e3bd9e1d5ad3c56d9d98994f58995ac6ca99ad6f72d2592a9b349c4c91ef0ca94172d54b385e688fc9e1a85b512640b9a8cf6f03043baaef47848ca32345769b2675e37892acc67a769a0c18d76748d30c6cfe3106388193fac9420b43751ab7cafee357f3595daf58e9f47bd9783aa172576f4f725d84d6891ca34b3b4f647fef7abdfa505cec7f3c35ce2fa29122a7fa088074504f50879e792f611c2202af05d5de42309b7fd9027beb40ca0bafe3e8f08c965ed58fad941d6e30f41b30fa1c6d03c831d0a83ebcddd7788d4f31243f5d82dec4ee501499a3ee86f5a9f854508cd4a0c29319aa181de6af63fb2c12bf6c4d9defe2b3c15a2a5b3d5708f639b35a2e848f171117daa67e0c880783d8786e966bb3df50c19ef7a154706af4eff2d9d18504a89aab725601f3223f4e946ddae4bfad86926824212cc072ea85ae91d63f7fcb491166e4d2bae494e3fe2925abfc038705fcbd1603b3b13e6442bfac434ff7e1dda3eee3ea49712ab22cf63148af478ca09b2063918d84146297335e2dd41de9abbde4c264bff5f7ab0fe8b73514db4198f99048bb7969ced9d3d9358dd72d75829f09ff938bc98e515815378fcfd4c107f7bcc794fb6595176f5b633be6df38d772e35d29b520da7c8ac31a900d4c67297efe01c4714136419ac1c688bdcc8e15513094a1cc3c0c321f15fdb6afec12b57fcd01eabc2e6f47e66203a69f590215e15d0f10430db5c6c825c2d8977d61c607bc56fb4aaa19cc1d9abdfb5060ca60e03c5d40eb6af34092a3a8446cdf9b11af6315394b5dadd8f1d8246dbc451d5b5bb1700a2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hba699d938325e0d03184fdf3c327fb6b0944ecafb3431492f99ee6768b9a3f18d368127b54a51c52dbf81a72242215bd32b718ac7ce11400b01b5cb21306b4fb4c9349c34d0c98b7a921d8dfc07186691a387ef7b3238b4377cbaf7b31b8dd0fc4e28b029af4b2e87d5c6127d8c2727a8b0b0e071ca7f93813732a85ae01b670418edda26fe2d15c7e7f31671328eaa30c3e088bbbe3f4807ae0de4c4d41b967f263577d2de734867f3d1732224065b6209cf89e45ec45989313fc95ff6759472f09fabf6ec28150d2640070eefd0e7022b3cf79b9dc6c4332b05e7f49129f6e6a3bf3a6e3d56ab3386ae5e66ba8e2c6f2b1eb51a9c2b62911d750afcebd92a997fd23daadc4035fdac1b471771fc76d357154e902705e681eceeb19b344b5277a69da23f9a4b0ae653925d2d8addbd7a3790a3cec5b5b4a5cfb8179ac21eb85ea1d71dac6791c8aaa79f22f6bd24d8e54103ea70b47c53c2083aacdefb2c84c254063a0b6fc00f422acd431242d3e8e281d4aa59d1d7decf7e5ee572044c6f06c81c0ae554b2d9b3f43fde38640263cd44b0fd3b9f93b99a5dbf11f1a557f376e4a9518c40dbcedc0f368aff29a1e39dce97ba2eaa737a66bd60439490d5e1028a9300596b88be0325a14c88edc9bb3923164b44ced5b24c730e53db432a480b9adf061cc0942331d370408ab33199d00257430cd8cc6ea8e111592d687ed6e51d60252090342b3722811d501fdacf1f5bcbe97d7981d252970672d3ef73ad52d259d7b4a1a2aa1aaa0fbf6b031efe5164fdd9e958312ccc07c144493328c03b41f758dc891788f58704c7297e048e3a19d80c8c9cbb405a35dd85200fc653b66ecc52077cbeb6eb206aa2edf2f21ea6a26230842f0e06224af00bcbcf03999a8a9fc29e391e00b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hcf180494737387ffbf31b8aeb90db03f08b792af988092f9858cc81a810cbdce800181d6e727752385c1b9511fafe05a86752287c01ac21bf8f5cffb45e7016765dd49e19f3110ac8d9879f713bd4945915f6ed8bd71759a02ebb101345f66545c2d6ad26c130b447a7f7496dfa498e9a90e0d21ecb323e6643d8d512c3e702f352ed0ab0f0343a24946857d8a22dc83b5ff58278c35ec7537c1b682545f54191827214ac46cb3e20acf1fd63424d86fe280524404763b1a4589071f5c21e91c76ded619060b65098724676d653da13626ea8b68d959a0b75d45847521c77533d180b807fedc2de923c5f9ec559f77120e4222331287467c01c42590c7c5a8b3fe586ad294ab35a28d41f8fd28a2eafdbb7e50b688a1e1ac4f24a6e48acf29f8bcfe663c161aae777077f37486c531394855f0356369148fe1568a5356aac957f2117940f1c6a76dcfa9a2c582318a53a18ce103a055c2ed3ac4b37e94d37f2d17337fbe50448dd0202c80515f4a231c9148227f93ab37e44b3c43cbb7b536d60f70b3dcaa982fd8f8d035104420596fa28c6559c83a08c5915ce66e63b8053b4c3d045f53a18f07aed28c8713e76c10536f6c7235ec2403d8e60cd8e75bd1f5611b87e54a5b82be25b026b56c7795dd1858d6e3b96ad46d04d7374b47ac79f82d3cdd3e4c608605ea63392cc173749b53f2d99c5fefdaa2547f6ce95f5a46a3b7b9f24c31f65d79b796e3b8a5cc43a63a6cbc1486658c868070264c63099a2bf0f1f256c4d7833dce80711c4baf238e57f755bf08fc1ac9ec8a352982ced7a5c4cd8502939e52b30f08f316bbd48b9ae205139eba5af4d2207fee42112496e444ebfea8cbd13c848d519eeaeceb1f9a53d93c4724b6eb6adbd3ed5b587522f1ca0d152455a6ba81;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h96172f093f66c532e70a62fa75392f1f4eb0edf4591586035b4ada55a94ab3f6afc0a664b37daccc8559de8eebdfacdcbb53f449e578dadef6be8c204d6305301a4a2047cf8caeea0cac2f98a197cae5d28e5831fb54f1b21ca7a78a4a980c84f819f39c4673834d307d13c2f58bd8c56a227b8915fb5466d5180c043d7b545322e3995cfc5156cd85f7a0fb0ae7ece15d43db8bb94a06305734fdf7584d17d9fe624a9cc080d77e6b6af01b78824d584c9919baf73d0c2c50ae107c3ebebc9b5d46a7f229f988604b1aafaa8b79827abeef4af36b1032c61195354aedf24cd758be50735e7894c51405fc53d0a32c09855f5243c820a6df664ff299ff9a486e21179f7f961e143aff77d82f045055ce7febf0a667e25224da9c77dc3f8b483e5dacb5607bc2cfd5bae1c6c26f2c70bc7e0125f7031aec3b715a15e563637e3223d2436d42e58d9f05982d5a855d6a84c78269ab1bdaaec1972ca25effe5294526bd6e0c88a5592514c48988731e5d742c414eadd823868205cc02d326545073fdfb787075c19358c347e5f61d71d903177164e939f3bc773347fd01f8be03e955fac3da937e7ef92c72f076884f37194423124f7e67f7ca2eb57bdee159538ab3a2c1c66c7ab183c9ec489b5b26ad06a29503468fbf7c7731aa376f9e39407240ed5725d57fd873b82162886d6e500b354187bcb68806e6ae153d9c1ba0f642f1fa0765a16411ec6796fc5a832d76f10c0768ba6d9012c4c910099aed433ec0b89edcba41e01de7af18f422a459c78d61fb2560b288612a56f0e3ea78ba16d365d2730c4031bc7e6c70d6bd4c87c4f2dc2dfecd630e8202b65489463456f17ac461a48681764f7f44bb4acecec66c6780ffff2652b4f55e446ddb411fa24d18160edaece07a3f4d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h63bbecd4fc9d3774af7c5574b4e704edc7e97d4469bf3c659622737fa4ef0c297f5763906e2d9b4331147738590ad01f14d7daa8c39a34845787d91fdf3a97ebdec1016a790c97b62d7fddc5795d46afc5c3dec55725c85a58a50339f0ce946ab5791776d7ee8d28a12e90506c7a3005b890c00bf48aa826d83462326fec14e6efe0b89620ca55425ab1b3fe8ec984f909e7cbd4c209b4c52e86c807cd4d1a2990603d303d0d811624ff121928b6b65632b43a4afe17e6b8baf42e7afdeb04a8dd3baa6906a490adc1b0ec0143c0f7c8227abfe9297fbc4dd914cba85d69d48c1630325dd7b4c8c529b4831ac65568f42f48920e6b8d31d9aa49728936ca91423d1eb3fbbabf75c5674cb7ff62906a761db7be3910e232258b997654f48d61597e74800ef936d0e04020a0f925db56b99873e4c58b19e72a01bbd99d4ab8e8a347f1b10b37c64e69448addc0b4d3e85a8bfc37e74b5cd4dbac0e164ae950866c28d435e88d7915d9e0df87576ecccf7000091f51dd75f74fe1f9f821d90d7625b89b798383b8e8882b43fdc7998bdf50211ed9616f44e71bf5cfbaf95da39a90d11292eee18ad8684376d40554b7dec705c5953f2ab6109689cb87e1c45d664a6a54dcc866a20a6e894f9eff3dbd9489d926c48c600d583e807713831339435db7b9c361fbd21e66c428a23c25301a2bc0687b7243e72ebfe7017f5d54f7b71b8204882a30ac1c0809e017720e13af57fb462dd32a5f35f77e17658496672fc44aacf4bed6d8809a2b6cdf0190920f47d95d962a9fcf3ffb1d7a97cff1221df494345be8c36bcf216097a3feacefcb6b36ecf86197ebff21cacbb9f8a64cd29ca58d2a5506863b721d2883eda1c865a4d1420e9a0c3edb84a51e3f8eb4a5e8b2a231f9e8d94f9d55;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h93b65194d4204237250bc25aefd8fe0bb377577e62e80a2acbf10305c8f5ff315e0380791c60df54f943e3080531da3a355614ad871c3c56f4111f61988485ee85984422ef05d2a1719b299e1137d471e6a7c73b2d5b041a61dd9477498a1af0e857cb65ecf707562064bafeddf41f6db11f8c1947cd75a7e590848e6481ed937e8c30270a4974918ca80d9ea3f5b64ca8b70b9065241300390d6d00179ed6ba360548fe68bc122b0bc2d7e8d329e627c46be329dda1fe308f3fa898e6faa1334988d036c70b30cde4114e92a82e697c01b72070f84ffc63555d2ea82020953521a55df548dcb72cd7de9f049469af1500c152d7ba0fa137ef1f9df677dd1e9204c94ab504dbe3b8c08f29980660009ffd10dc238160b1f32d2a5764b440426d8d71b0f560a30d4ae3922d0f8b8feb226fa7af0ec233ad5c627c99c8089bf1659999a1d18013e81262c262a3b2e3e8f68772725a6321f43d1c83b90762a79ec64c46b477912337586575c251fd1dc794b9b09a2b3e59500052bc57f87ada54547d75d0d4820d292bb9b653c15e7dead756400c3b284d8f59328c31e74471145cf3f622087f48239763ce1a4381f79d8f7cff5d65af7fde4f06a1ffd16200d7fdcb9c25ac4b446eaca5aa4a6bd50ef132ab428519cf829dd7aeec5f6cb2d0e0c82daeed2636941d985200b488ea98e8498547795f5ae59b94b30bade945c48859199c69b197c53976c3d9367ac98a641b0cf58f3d41293da5987849886172129a4c1ffd56d66c229d83a4cf1cd69d1453806da395edb86ccd8969a3757456af8ceafa4649e0b9239be7e1efd22a48f44b802e0f6978aa83a3a6ccf5477f9ba62e014746ae9f521362910114b3ab36d87f8d081948bd84b88e0e2c3606ceca59db560d7225b48615bc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'ha0703ca5ef1966f53bd189292bf9dceb7a20140d2d10cf4557dc5a4124d760d93a84e5214022bd057a52a22edd53bf5ab494e78492869e6e6605c83294255d0418561e71931f60411290b41d67eaa177f764284bcd3eb725412d3defc9f539648fe6190add6b75fa41233018821a785c56289a3455d20b64b95a9157436d268c025aae4a7d02bb3dad3e965fb1ac7209e46d938846b8d9e17c473729133e81b8fc9483be24fb29fd1cee946fa307a05c4a99776adf44ee757fd6aa4c0faf152645ca7992986782b3f2b5c37ba72f3d93871b29c7bd2c7b3e6842e3999678b8a80999a47ab91bf0c8412f0752e0ab6a50b955d3b9b98b3f33967115670e3f37e2eb84b6a6c7b5595e32f6162cf496358eeceb2495797d1f67f27a3bf0f1ddb6c7ce007eec8b048d0ef0728525a34b80073d76825d5e74f80acba76502aa42d12c1ebbd79d3120dad8927f2a82f8fbad7c5987f6bb9aa2ac0a45726eaff9ec138815889422cdf36ad90c74c034651541ea0c1c02beb77ae897b7e40d5cca29188f4dab2ac4b50667669a19e62bf22d59a4bd4a891df4c3cacc168bf5c0cf0c2883e2afb177df9edd7e2bf0156c7d2dd5a7fe34787fe98e051c6a0321992eeb908252ffd1d997e4a334261017b819adbe2213f8759b1329680f85311409abbd96745396d5e8281527c0c2442e0df89c7f2d088e810a486b132abff0e299631b978c219de77458672551c689cce21b86a2846086957d60e3aadf5c6dab1131698c7b880cbb4c7475c18c8beb0d7f92cd00aa6d71d6f905e61cb852deee8a704c479903669155165563c820903598fd2b529e73feff3a6f35feddac253d06191faefbdd03a37806abe6e44d5fc9bd1903713d69dfa2a5d277e927c433a9628dec9c783f3e10fec5e614e1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h563653475df05f6fa11e0bd85e25736d18355ebf79f175ac31fa368c16d8fee1f68abcb5a682bffa7aa1ebd9cb3c2f8fe90618ff7449ce16a67783609873032aff38a4609553f4a2750f3c3091e1e95159e0e34acc18e5fd2928bf2650074f4304c500231d2a87775d874069760e39d17446d97cf96c97c81e5cb2eb973611de736bb562c25790570acab33ad3ca4839f269b6065c75cf920e77281e0658f5f53966c67ecc34a2f71720207a60b35d73ab94ecd36ae5cbd22bb8634e56105c7c2649ac8c09037dcc9b0640169e2b6b9dd9bc32ca09bc1eaa43c91b8874ce9ed4801209892ccb1898ad0dab762aabeb655d0e8eb811d0664c86cebbfccd88a340c1174b275095f853db806f0dccdee6ecd070385e57bf1732f85b172548be9f787deca9c5165e7be0c5302b51bb3416c4cd32c4519460f36560736a5ecf310c9c22b7df727e89931dd05a74d5ff4083152d1aae9e16dd8a80445eba7bfae3d7d745765d84129ffa89f76362c5908b96510bdd6c64dc39e56bb73f9b788f5bd11c16d8232edb7272df1ecf71cc2bbfa942d9f8c6fd5e321e958bac5abc9b8f2cfad3325690981bdf9fc73eb603ada7689482c9fde811558f77a904d12cf9eac577c936b84c2161769332d472cd89f0ea82cef84cfa1ad72634b628dc93015f2f3acf9c3a6b2906225505e8396910fa45594ef43afe4a8efed9ea7142188e02a5651a988dbc1dfaebda45ba17142996e0eb2fddc436b7e74aebfc8ee2585e67cc45098d307cfdf37e03e0d3f876e72af427d10db76e9c953387983584ea32837fcf2bc38a3c3cbe71742b3c1272fdaf12d01b61bd81128d29bbc13a69e3fa1a12bdada79a4b11eaf867abaefb53a4632f1bfac8378a4b697e04928b9b0624e82794538611c99fa22762;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'ha5a709f109e78db0cd448ca1e30e4bf375ee3ea53ce3f3817887b40de6a1cfab0f91ea41c33739930fa7fadf20081a062e4d6f63f0afa9c1dd44ac02ea4a3a879206e7564efa9d8c89066be5fd4becc9610824596f03907e86e0b67ea11c9f0aefa08909f40ada7c86bd24e36114a5e67e8d5d9e62f5f6d27547c82c4480cba3f5c961d0da1157af48a1b77a66f54b18e28e333368538512bb738127f3bf03573610122c2a8f17c131e9d94dd886b89f6d6963486492f50daf996f8d77f6533a8a23b291eae9b4dc04b95916b3410708f6c5f063653030b6cf4b8056d51e72ee9ca034bb5a25c28eb1214244e5c3bc62bf1c7ab749ef5c9753f458f59d5753a815b4710fc30191920fdb6a61a04e1eca13927082488441631f11e5548a1f71eff7720893107c31390a00466ac7a21f68844c23a2c5d89045483a561e401a81e2f7369adfc74cf7ff6f871375d51d08be1f9dc726ee89887e2b2d8433dd9bb1ebcbd7c5ece4f7ddabcda8802abfa40ee0c2bfa3340ff4bbc20324e5f151157e65f940c8c8599da3124c8b43e62fe2ab9966bdc13d9ca4c4a9865a50f1ccd7f1454be543c849e49d07672ccbb78568fab26b4d833c726666095cb186b9c10a67717ba62e2240dcee680c3ad5ba24056a960fb6708039cc8183316c67b4531f9043c76c85023a8501339006d0fe1f136667cd27b60693d14560d1d1ebe24492bb18ac0d47730e12b34fd7138fd079e009d88a4ef22bd186cae10f6e2cd8db80f69cc9723e86c56f1de69a00973a8b3f05ffe4234523ccbb5ca736c9d8ba5f823027d711c149585cb5601221f8fd827c9d64b69c4d4a2c165ef6d5624fd9118a38321d88b4e2832d655094f2a0927e7f6b3fbab49f556ad0a8595e74e7a2ff0baf20507b1b4655f474bd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h508d1f4b06547b94872e81ebdf3a2732fd048ac139aedb0be251cd10659bfbde463fe490951c307de5c3ef44468bc00b1ac6d5e220b218ac318308e4d92611dc172f5fe971592ab38aefe372990ee4c7bd094de4e9701396ce8d705f5e3087a7f5a48f402c155acbb7a3f642f5704991e2f59726c1348611c2a9dae3aca1a56e224b63cc9f1f9042c562bd404b0ac5f578ff03c9929c78d3c49cd8b478097f0a6074f1dc759ebac165838e20556b2514fb860fc5963393df1d793befa86acc4f86a461966b11baf064365d63260522c7daf6afbf47fe393b63cf8715f6df1206255eb18159fef3d535e3f396836dc75636594792a32bda236cb56ba2bcb5139d6f0b2bed9b037222f6109de7dbfed577f2b46b4cffce6cebbabb412e8b5e9c3078c4f77b040fe4923ba37749f900aa2d7f2bf8ef0c81b9148afc7e2c8ce1fb30ec865c618912286421588a0d8398f51e9fc36382cfeffef531ac5215dcfc3f693a75872a56f8698f996206eb938ac7aa4d7325b2923b52b7b77855014c76b55ea1857aca51f4a1ec0809c01d3186ffbe78f1035f65d01e49a745c8d6e1d9209d9ff2955de0459e12504e92ee059cdc027384d4321cbd509ac009dca27535876c9b3a38bf26c3a8eddb0c98e907cad043b9b2210b6242879a18731f7af554a10469497c743177c13343337570a4ec1ccadf1317d66bbcb041be919d2f9c19b87e0c262109e71ab3ffc90fc595cc0920e46b84981ed16a4c8b9449f37a165364c37c03bd138c93f548d3634f295b52aaa59da1a71c7828270be18a57115b25b8c7944d825fe7ffa1368add849dcacf14310d6e8cee1e6cdcc09cb347f5521602d3ff173791c78390ae12765a3b6a2abcfa7c6b74ca39adf81b525388cde580c2d0961fb80bcd41e5bb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h8fb8e162373b00e4d13fb90ebbd1f7d0df81797ac8b4715e03954945713ea883bbb51a884da35dc363a6a0b076829b7e98563fb16f95a71d3dfb93c994dd64ec9a67f2903dec0b8f4bc95f8399074a0bf7dcde050c377d4d055f5f6e95b5a7e982bdf0c9d33744959299062ed109746823407e7c6f626878d9d458afc5f103b7c2953c89a589ec112c17bf7a9a6343970df31da9ba7b39a52cb26139987f7108b9ace13652f354ef9ba5a6c16657e02c9421035af09288c53d22b50c8d38c7e7789e3f539bf9f85c3ac46166b2a6ffcad78f13438f21491bc9f3280af6704e306fae5ae3685a775d9b6e33a9ee90613f4a825245977321af8bf11117133587ea299c8a7cceb22aaef228e97b0f957b75c29788b8c7202f2a52f22f4010a36d75343d5208253769e0a10b843d7ed7cf38587b973878ae79732fe7ab0169ae5f1f00d44437f2dffd31803e33877dc7916f624a5949ea59fe1c6f23dc0197edf2c5f10c99bfb584996cc3be80e928aca80f79478fe2c109579c2785412c8ac63b3e412a16b8344338f3ff87fd0f52f67c08d5feec85394697580628b0b4a16e9dec6a631b2eae6b63057907e52e6ac838d7057dbf73290830859a8e8be24cad1d5962b827663523b601525bf151db21b89449299fd514bde43e6ff7ec5b7aa5b922f4fd7ac3197a8f38dd7d13452a9af9a77b09f73822cdfaccb24c4468ab2bdc8b5a27cea94aeab8e7bdbb519a950d7f705ccfc88730ac96ca3f4a5df9257cc3dd965d7431e6ee61db08233fe70154075d31523bd29b180556b1dfa1d96110d2cac9cfcacede0d4eeca275074eae59a370e4ca1c3c400521f39e3279222922a6c218ae671478ff48bf2a63c472f1c35bf6c63594feca08c0997cea2889b6b5acda1e4b476722f8c6b6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h54d44a37dd8e9274c0a8d776592623bfd79dabdea95a50294901300634434875a91566ee630bfe4c721e101aadcfe1a42b17ecfcfa5045f969d42213581fe5d66a306b9aff77e418107f2fd5a87c9083833c4cd83e46b95117fb20f3159ec40dc066f855322f4722935aeb70b06b1d7162d0b3b5c9db9bbc1607200ebc35ba9155a815e0988d391b71d254405b1f03579c4d6fc4c8a613518a18068e6472fba081c4af803d3a4d90c2890050b0b559c5a440fa8df8169c310be238411f3d83fbc54b213a9a41a64c26922ada431db16c6841bb1fd49ab86c1ba5eebae6fa2ab498a89eb567cb23871244af4c2e0dbd107fbf9255d32025a3249105215d85ab80bfd596675ff8f16621b578858fb4a5ba9b3380b21ea7b54ed6ade2ac13519dedd11a918bb5d76fb10295cd4bde5cd4e9fc7692422f8c8cd5da0efd81c9572118c55e8bef9e6334388ac890c61988e237de62d8b0ce730180a37ff8026999fe723585baa05510037a2d1d0723340053a8a7874d58650f3d19e168a8a14193e7b61d506395d57d715f1dd7ca1d52546df0aa1f50e7881ec56e87445fce5fdeb72f16a8009de4af054931e602bbca00ba8dec8bfe727db494bb247a0f3094db82747035dacf7ad16838650f2e9231483a6718b7dc69a85f66482c329bd2ded6f8f6b9a49ff9ff6a7438adc9ca16f396b4068574289c246be880105cc519e666a79edd32e9cef8c6ab7d81a229ba2242a9dbda021f89fe2a00e69eaf0b45ae4e050060bdb2fab2c01a9b6afa76901b9f9dcaadec1ad54f40648b9006b2ec497daa1592b35923734524b00151f19b10ec12c64f649a13cdbc72e58af31b09402ab592f2ea9de661ec153b9f4aa18d62406a7f1567ee14744bdddd557ec80a39b6fa9bc55903e5c6794a2e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hd79bf6a3f2208cd7a5c320f2fa0afbfe83f91383f193da74af8e9f6032f99f3eb60bc3f5ff04dfd4f675b5457140b7c6e5e65d42c23b818a776070de1d76ab4581aed3c76c3559a26ab76a71c472288e3e3612569b00c546d93c656d496dbb729c939d916e3bf12c88e5d7271836b47c43cf0e918b86518858f897b1ddc789781872bafa88424466facc5dad8a60a9550b6141e3ae74b93fa135fa2610814165c0770b7cabaf3cba6ffd1aa577a6200a5bfc2b7d8f308fc1f830b5b15f488959241807e0606e913caadbb5fd50e027045662da4d5a674d01447ad5e66df50072dc32f729e82014d3c4aed44cbfda8474e6ff9f5814f24edf94f1325929cb51b678959e3c2d6dfedb1d4c9d2aa10d1c0559e8d992f512eb7bc92141fa94cde83592223e6c33d24cd9a3adccefe53f38b33e47d672dac3c22b8ce120562e486f61b2d49bf827a2f75955dd4ffbe00d713cc7b1119a56d63f78615703989beeade6dd953f928b20b3b247ea3d1106439ca4a4aa481fbc4981cedb8663a578a1155296749e98eef7ce9a151db173418759ce54f9d191c155ca7e71d96a1e24c1ba2a8df10595d5d44043c24f10599264ba3ccadb7970d63f90d4464c2f0346c24a1b3f696c9d618c1471b63c2bd64bd541651d793db7d524a7ab959418fb47690a377992328b55f82854cf7235efd965a79f87a3a31b36508583a017c36ceaae30cc4fc68358acad6cc664ba9a8221dd8c14b0beb82f30756b3f9165a1d396c70e05b9f6ad83533ab4d08638c20c64a0caee430c0ea9b8eb9d393653e167fcf26f4a9a0ae607149ce7219451abe0675a94082055d23eb03af1e38f3a82297b358478c900db4b32a00e90955bef548d5517262ee98f23c4064a71394680a5644a3042687f4288f6a84d22;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hde59472a1afb082c9a552fa3426dcf9caeb5119b5b3e605e18999f929cefe9f61138e24b3ae793c609d5d6113e6ce7402cbf6b5c86c49bfa66748338e105b85e0a27739a41235f1123bb3f346e081b41af641a4f72b059263cd85107dcad333b40d5a04edd54ee52ab757b3b75236f146db70cacb518dae3d0b9a8bca9130d57ea6b80fdef965b328f6f09a84d80aa2d34066ad3d6c0593040ffe8bff0c6a035ff25af2827a41ebf9c8b6e2f2c21ca1322a1d3a583a8e3196751b2bec759ef8c7895d573de4e9afbe337b7c2673d1a722865c46a5614c99fd7e4486aa409752cb0203a374b3684081034fcf4ed947d2aeb7ce10a4dd16b26821cc04257b5c7da0302587904c21c8a7caadd6a02276be9da3662b2377f3b35013840d07bbd44e10c7bfccc7f9257ad8aa94b88f698969f712bc3082346c1cdc68022d9642c3e39aab52b56f7da918880c572e07649cc3ede720002f822e14e7daf84ebdde3af8ca8adbadc7f76e3d55b5071ba37b2dd23ca9f0ceb21151da3699bd17b1621cbf605b62b4742d2c0870d04665e928906a669cb6dd736b479b5caf7175b0b2ea1002280fe1a16e9da0c469403a719bc4c1545b7307b12641e55e091b1bd6d2c3b03b250832579441e9d981d5cf062528a1325ced57a4e4b5a80ea2e8dc83464f87df25e205bae3f0e033940b45a7feac979f01e62528108e5299abcee0da2e6eb1e37c39f8552cef3e1f92e198295e964e20ce0f6a092c89fb1a380f8d01c1a26844154d6e5d0273f04466c8d3be999d48b16e169357c09b424db6ed80f22ce6ec78b0404c142c7ee63b9fd7ece3a7516f0d43a66c3bd0cfc545fe0c352e3d719cd2db2d1724f05ad1b41dd4bf77ff522913e5e15be8e053b8729fdfb09f93b59d53f45bdc002ee7458;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hcec39ffe15b64380b7a5826992ebc8360072fd9d17c1f3f1038214d332e94b757b7fab661aae9904df4156e1e49c43b1dd58d1e410c5e63675c29ee43e7252342194f13402fd106f7ec33d413acaba67b49e9518e8b54da203f3c50fc6985d33a53557d77412148350616c0e8e3540fb1d26f3990eee53f6af6158635fade89d47060455763329412f7199cb188e7ea6d4afeb4e3a5eb07414c7a0d4419d96890fe810422cdeca5c8f20a8488b571fac14aa763082adfff850fa3530624560fe8b003071252686e1074bbe2f7d94ecf3c6dd8423a11a6407d0f95eaca2f4b79f876e8d26511aa67bb29402124e40115d7fd86baef67d4a4ea0df1b67094a60b35af0906fb63207836b445cc927844cc58236d3befcf6b487875c9bc62d372bab74f248f46b34bac889cfc9959b1915fc39072d4973768908213d1e8131c60029a6e68e6e1261c8e05bff5acb03c446e0ab0c40007f2b50c64301128e8ef6dcbfa31a12d0c32c91ebf4561ba44d94dcfbed8f28e10ae42bbac6435a26143cc6a16e8a22102887b47f83b72bb593139044299b41a25e41c58a0fef188cc9ac408f6a9e16903b66f2b8a2bd4abe45bc54f92d4ed8b559eaa4582fc7b62dab50a3576fa0d2d3fa1f82f86655af312f897d4b128b459a2a0cb04688e6c758077f59783cd862995e495c7bbeb228dcf2d51d2bbe883daa15a7b96e53778ddd0bcbd03c04fd129f7dd0ec0acfc764a6d990b539d5f7901259b887047fbf64e2fa527e370b83f7c07a52ce2885e92a3680ec5dd4e26899b900d45d1224838376e8ca796abfcd6be43b27a126ab41a12fa8a450bc0357a82a1a177b533106cfbdc5fe7a75b21926a3a707ecc5103ed7fe2690f9e2885ffa8353d8f29604be773258bc02ee902dfbed2dd5e20f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h81f532bd91964f2a3b6aca30df89852ed261b4bcea29ceaf7d19fc427bc0942629131057b434a9d4c37023d1b6ebfa6b12bfe2f197eca64733558b15b478ffeae142564c3018d0692ea863e7d78efa975cfbbf95288267d9e10e84e5eac4ec296ac33e19d889ddc585acd399070e628474979333cb8ff5975da6fad24f84060b8f74dd667841e5b14027ef2cf269902815646221927fe66cfd7e426c360ddd8b37a328fddff3581bdc9c6289aa0b0eb54eb4b03dd31aa04fb101074fd46bc16c9cb32418fd48f968f53b88b338b745357c1c004f4334dc22f815ffc957e3d7828b3c4af20a83387f030202a30cd097ab9f0c996237c323393c086f52458ff212f6976fb9bffca6b4d6871efc9aa933a00e5d4e0f4b03220119d4f4f60e5ffe1a1c27474606e5d1612d3646d04177ac0bdf5a40ff87eea738b96a6bb55b2d71fecade7aae86b12ac5c1194cf7462b4e5fef94d4cc1c863af1ae0bd2933e6edff0be980ef9f9750ce77f613133893b4eb04dc64bacb2e7f1f080ba658b63d68c788647f526d32ce654151888e3b5c87d3e5cc41f94baea7526f85e45c833427623bf2b64762e41d910e0cdd314a57accf179230e031403363ed940875d8e220b20700bde60a4362a4c0e010466c81fccfff6e68cae29e4c3190f8b85ec19261537698d0cccf9c75d58e57ad7b8b25fb6f419ad1e9e852417a68a326a2b248fcebb440762131a106acc1f292867b01bf96db23c328fe743d34177d4be20fcb1170a83d1c926efbed045b664fef717ceb7275b4aa3b82cc4545b4ec305ea8f08dba2a70ff0e76960a6c11b4776f2c38df385efff70e33c1a9f2aa2d8c5b528ac3459b02236c4bf441aa7481d22a4950875237af3e87c9016a109e6389e1466827686cbcaa7e6654a65ee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h356b3b5ef196102627216dcdd721c40491e6daf8c14b3bec8e97662063a7ac3e9f88f08eae88000961bc46f20e4da1656c0f1d7b3950e8a8bac613f84c51ad23f46637d535410fec7da8de1d70f7a80501cff7d3d27fcef91c290e06c5b8b9cff18c6d4eec14feb2f9ffeddce52ba24c5628e5f9cb4391d1d83dc1401b84ac11b18f8ccd58507df89b2acc669d86124c98a30a6ed745723904c23e2d330d8b52569447d62656471ad0279355019d59639aa61a6a8638e67743b02337784bb528d0bfdbe3aec9d2333a16867076e4de7cc0ab799ff2a7809ed51bf43f698c1792a9ba5861b7c2393327b75a3d03774127fc915cf43f7e5ee9f9f9bdc5a984bafb1dafed16a1a7a582529c2e134bf34adc67f77680612742af354b945535956fa812f0a625b9ac683fe3bdafe726e7ef89ae13f88d20a37666b53ae03927f1ea0808d3c9a490d53e058bc88fbb77b40adc394c0a36f7e47f8c3ad42845ad2094adab08fe9bc844a648728e0e0228f15760884fe4dbe2d74885d567364ae227bd4b69d26a24d2063aa2dc6a51b80234d167d22e28a0056ed0ccf5b6ae670da0a8931ec2299def080d189d7af7e7fb186223f1937ff24a6ac7bb64451b4b770efa37e4848809cea5aabf2a3d5a5e4f83c442482ac2eab67650c8d67e045d656b641399f8af50e31056b85a73ada1a25b178ecc4108c6248b825406dfbbe7a50e7b963f80a04a072a355dd24547f5c4649ecbfcad5d63709958023d460a8f5744c1b97f26d6bc2629699f52df157f6fd7bcee5cf6fcf2445762c686ce91035c65e36ce8e98d05e306df1422ccd0627e4ce3e4d1872d50bd8d033e36464518e3f1fbaac26dc4737e665883ee58984f525516f4491310db565beb0168741dabef82d2e2f2692afb5007a2dc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h1d0b54edcbdedc9a12a9e1e7d8138d8adbb1fed85a71eee2a30ba44b94ba43b5a0fffaaa2f7b5674e6fc759552a3648a714f9ce0204aa690ca2b6c0051a9074e29c3b2d9af421445a08d73503fb01be05429ee74f64c2761a7adf020bec05a15a2aef9e987caf5182431d8bf04d7a461acd5d4c39c79eb7b321686116ca734cbd2161812eae5607285d316a6c31101121b16332adba2eff77cc16ac657546071877af4ec7601cb3508df79ac43a48e85386a46474aaad57255ab356c3024da477ebe87a6262981dad726f6506cbdb383bb0d30dc3847282ad2fa158489f28c228acddad6cad54e5db65ec45378f29a0fd04f87701a8b860f4833beb4f102dc9b72a9a3979d993b74932f489c9e8b6c918d16f67f067419f04842f1c503ec4bc273c2054241e9c54fb5a38f262251fc0a219337193b1e45e97b9924631b705200b37dec9ed4a03ae09d9f25783d46b6cd59cc21a33b001a2c3429c18a41649d46821097ccd8fa16fde2050f265f542bd8383435f11ffd7306e91e687f1c1a0846a8c0aba70314be492e3cfce256648f9c0a6b526322f0365d151550821f5da06c218bd6c13e949ba489065c7529f0b2beaded12fceb9db7184f434b1a0767acbb7fbefe5b93ade94afbc8b30ad8afac40d8c00b8d1d750be8b84182b888df1fc697f2ddd521813d64c20f192ad5dd6948f8d4269cf74c9e298a18a666c6eac52ca2cda4bba35b0b7b4f4f81e7b030a9900538bf99a8b2eb5bbe008994aa6e46dc2a69df7069ac35057b8f1daade7f1b4bd6b47f235799bae73d65b5a22495c7b4dacc425e3d61d01f83d112a5f364d9e53f8d53f11c09f0e0e1fa060f33761ad0a5b860164b5fdaaaedacc959b2a3d2276feed7df06f1b3bc607da893b2b79116021cb01665fb31b2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h37c3eef1ba679cfdbb47779f1cc45da14498b2a61474ea81a1ca877401cb05f910e110e1a537405a8a714af920badd75d869acd00c9fdb32f9f7e33b9f7f35990e35e5e76bbbaa2bbd9e7252d6fd107f5e8fe12f2a2a1a09e60578942d3baeb70d8e2b2b7772c83a4941b3049eb1320c680ff76a958c7426067f76de4f6508879c0e0138bf0d6f8a21dc3dee14247cf86e4b1b8cf75dc3eb2f9042aa59c5e42ae20d220240a17d96902e1c4aba7c9c377106d6f12a772e7480f7ccd9feffdbea2c2cb4b046d19978db2c900ffc69b53a896694c027012c6270173270d0a5fe19dd4ece30e858a87b2f3cf03e8f490830691b6308003b9a901432055d890dd122a17987c0383f24649b852c4b1da9eb981359e9168dea72be389f91d0efee1e42b6f5adb44555522db3284ae9d7870f8a0f64c9fa98dc31752743090e8106f018115ffee145a9c14466d40b0e22722227e24307031db68fa9d783226f7e79da6d407d757268b5a7375bbe08306fae9e65dc3669d0ec4187c86f5a761634da2f6581c37990bd8175655ebf5c3188ca099755255b026a427f98ddd0bad0ce4770217e21cda73935de49a8a7375c0585c88f0c86d271af84334a08c7f30bb8065d1fc2132c97cb9c571f2356078b359d9ab6724ef0fd14b2d57a87ae4b8b7acee4dd8a23c3d4bd0225ef7ea00b5c3bc93af9b5969ea72adb2264eb06b0449a00c2a7cfb43ab4d8db9a77a75afe764a2d371962e49e062abed662597edd2d3ea88b1093821f849c7243e8d0c94346118b91b4d094392356b57ea2ba06ecafe248cce733349d0d41a9b555f10f74ae3071fc74ca81a15d6bb1d46237bd5a34961c5e0fd3e4c94eeb3226d44ecff09f9b0c178ed7ef7539d3cce262658282d862e39e2020787e9320750581;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h7454e4819154dc94b1f1b4a3f6ab4a26ba99e7cb58f531da52a68f99ef18a9bfeb017b746b9e6fdef6e0ade45cc366719a9841edf7ccc06694445a0f97dda396caab3e2d4e83e9c8b489926c72e53a3589e96870f0ab9f20e0cf40ae59bedfd5fc52a33f74bfe761c1bc72b8e17fcdfeb8633952b2c3d2bc3d6ef6423307e3802caf81f4bcdca9561c9fd358932c8a45a4618af8e1d2f20194b202d9692c415a19c90e335290acbbfcb68a9e179efe6d8c70b68a5c7c2767d7ab4343c13da71cd7187f4c7bc163ef84d01b483d0e192bcece3a130957082cb38d3dff3877029aa6b54a01e0b9243e0aade8216817054e408591cf5906aaf767693faeabdddfcc610c704b8f020e8ee5d1e09a60c28a3ce3134df22541d2dd3ab57fa3f7c2fd49d4624a8eb0886017e17a097afc6faf968e4e347dc5de9fb5079284a40b98c03dbf7c274f2d31bd076bbaa39e426fe417dea42b8091586d114315e8f006ac77349dc3b126d484d052eeae61a8ca3290fcbb1f953eeb47e92f53fd0495d40507a6f3b30dcc5c01dcb9f6ffb97cba2416617e3710fca6d079283876678494c882d46fb1fd122638decd2f6d2ad3a8b399c47ba4a93f13b1656d4a11980b18e242eecfde659d1794338f17584d41013d30d6b443506b6b4fc7d2e4e834738b0a9c4f01dbec8b39de7bf7d30a637e0331a90e3d0b0a58edb3d9beabb9da28c985506ef18b015820fc176019b62e3d5f7bd0321ac9addbbea56463eb8a8dd39183d0970d8735d3c7adfaa9be65cb7c896641ac10e5c901aad634a3134667bdf225a83b363ef3d938efe828443e1a70a43ea3f03a79c100c6281c28a7d2b2a115a5f200509969741751164e1e936b3b880c6c06e8539adaa8521e7554cf5b68e2fc3e10c3e79a7a002e6d39;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h9ca01b09af09cc3e965d957389ea2d977aacd5e3abfcf847e409fa63780bc7bfd01be95cdc897f3dd03effe618449e719d2df8ab73a45bc669aee8d84ab16555ecd1c7194012011cd764b2604790cd0a9d2ec7a5a8faab0859124ecd86f3bc3fb84b1c457a6b4b3d35cd47b57d119d9a8617104272b86ab8c6ef0457181c70d5b07f5314f64891d22204b2bb2cd506aebdc199248131026756bff002fdf2a75a7f101ec44c64880b22fc6aede5c7e9c421213c212338f3a982e39dd2384be8e29199611884350d795f5fd060495162f0c918ff066e6c100af89b3b42ca35c1b91905ad1cfad076bc1f70a695f1dcda85cd73568069281900f7a412a4999539887615614866ac81f2a644b66b0a940688b13ae9e43cd5179cb72c2ead64d66f8da70f234651d8eb85ec13d1d84258296525506a90550f863b512b98a1f731f5c6f0b2a2a57fdf85b5ebc059021d250d8691d09da935b7fcf5fd1b9b4e901e340a36e0dff90aa0b2439a79456939d81c94e6cf017e7debc20acccd0da2e588bd1ddf737f831389a4f83e97b80cd49ec160c00654e5cf5f7dfd2e46c22a03db9c7d3162967fd1400e5e5159a66b8f569eff4d17ab2ba5bb9126015a3342be07581449e72eac1ab92f0a5e92cb9b8ba40f2cfe5360af23da66aea6d0232a45d0713c53ba863e72472b0614719768b4c5f1cad896c2c8999b7cfbbe48609e981b61822dc551cd8e5370175291bd20c5c31fa6cc99a38051c772fadb6214decff2d38a5144bbe6452708ade6d571c767941d79fd38fdeb1f4c00def6555bd818458f7c6143fc9fe502a80991a406e4056ec7af70f6735f8ea834cb7374de1b67d6990da4357d5b46b05062ab8a7d6583317617094ba41914658b5398a3d02afb7f021efdebdf367c169c55;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h55f38b20acb854cc01ecfd1169af7e2ec786ca30b34c8d895e60be62617a646df6a28ad28501ed235b6443e757c3fbca2c90109fe248261c02c7db5ca95f9c0ce47b4a343fb2c3138e457f03b7f9ca7c6af1c5a727bafe3488eb67d5d4a70754ebd6ae1001286f7fb3409aa6fd8e82d19988b9254aaa5e1abac0055a53f86da67fa08bb6f14278c3b53d5d613f90eda01d9474cdb09c296806121974ff7ffb6fa44c78100bb1104e45b16a1b5d56155c65feecfbf4d96ecbe40ec335144f315c01a1de5dc7e817511b67d2677534200b9b4af7551c08b837e1a8218769c22adbd64590d877e2a49b19211897527a0385c26b1c5827d7b9fcc5593b77d846fa50bb76c190d62436cca008739850c79a89e017654e4a7c2c5d975ddc8e477fddc9866aff79fd2a6ff6cbd125fb4ff30d5bc7e234374e8bd2fb63b95e8c1c5539530e5d2a4817aa1ee602cb0d27bdf243f2b2057fb2b872e845dc6185a82ac17eb9b87c4271fc7146bcbd48901af92389b2c07ac2ecd211ddc8456e4aac21cf9967347127a9f827eef0920ac8a8349ea2e524139bd4a21afdcdfbdfb90fc92835a23a1c9adc37f000755d7dad15d158e0c900f3b6f0d7cffbab24b3130853cc2e30e8252818312f12b3329a493a67310ea80e6bb9c1022dbfcc8921839d1125018067cf3cd721024db7e06b373a52082f2341e3acef1ca85e681dac6700b1f81477aff544863af6120db6c9ee77520d637fccf6090f495e62b5081fc0a0835aebd0f62cc923dc41713ddadb6e194a3825b54312a2582ed222fdb0318b949f1d02ac6e1831bb08c3bd826246f095badd8ba28df404d6a8332385b7d3addfb277150e435c4f326f49b846514a7b66551d3a128e9a8f8ee64614fa4de5e9d8dc87de9ac635369d4e19c533;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hfb1a0ef7526d15381f1d1a97cee7932ed6d24ae0bd91d170ac67370e4ac6124e68575c0e0b82a19e301ae3ceb452e5c7838bb603c409c6c1f73996dfb29a800537fab139f22b2924c045c91ed7582161520bc55777dbb14b394966f87d5a28e541084272973d4d21e99a15620656b576af37b056aaab0f655fde2020b57865e5d81a133cd9487b5d2386fbb181f45b6e64342be80d28ce928c0b276f15ea8af5f6f56106b36bb77f9c84a6e1f62d931b562d58371be69a6badd7012c937c45721d66a70e7789a69fe127ecd00ce9ad508572935ad66139431c129f3fb88e1f41d67f7762fc6c7480b7b9dcc81986f045a8ca1145adaf77cfdafa2da599cd1ccc793007f00edeb6f7711852b0ecf90278ca664163a43738c62d20b020c6c5ecaed021dde5fa2c57ed5a769f47aa5daeb83267d425c73c1d43db099f5c4b7a378b7a17278cf5813b4b45ec954a851649de5524b5612bd70ee3ba1ef1ed3863e24e188da6a30bc5cd5be71e25280a3b76a8b71817b33745c1f794384dc1a8b383a95b628c87054520ffe978b1d1bfabeacc7be34051fb14012386a9251d8a0f6d102bddc400cddf8261a6a942bf7b72d126501129b6f52903a2373bab0237c107e14a1a8eef03eed41c57c9e221977c08a8c9391dd9bbffa2a466291e54fabbd381c94ffe5dcb8c3e9f4d951a99b1625bf38d00e674609c82718d98dd6dc83f0420ba907cc6116aca4e5e596c0a57fa1a79dc7db12c6a0ebb0ffd36fcfeaee89823da6f600d20af16a4581a7ea0f0c42cffdaf0ba45755499fbea45e9913bfa1b1c3d82680b409bba7853d9a98fa768cf0963a4bfd2892d0ec2281e20633fa7513edaa69959c7daf29fc4bfd2bbf60f8a74fcc432b7b5ec8b66246240ccf9b98ed33f1c967bb4657ae9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h36d7d1c31745086371fd4892b2d9e002355ac615fb5fdd1bd3a5e7937f7aa0072b02614bf7aa3c330191bf50c9f35bfea29ce01d5a0e6475c5a8f7c5d8a1b5c45ee47e538ef659ea4ea3283231b8e0db6418d32d633ba375ed4307dfeb33013f4e244888b2d86d3c60cd30b39f94466bc5a721f8cb0726bfbbd77eb18746f31399b55fbd51c28d66c1909ff504d3bf93d756aca4a88a797c752ade49bed1754237172762b50999d6467ccb052d052f4a4581092db7c78568a10a5b92f87402146a5620bd5bcc8ec3058d02ecb676f1a2e3c92e275b0e1bd5b96f38ba0877df8f5649d281f7575c0a5d2cdf03df4670903574af24b7c4dd9d97ec5885f5f664ec1dfadcc7581ef96de86f75e15601f34c8be249fb26c06f82ba8a8e988065e7095b49a25b829501c1cde5911c41f51cb8bbd37453bbdf88a66e77795a384ae423e939f9d656573a1bc086628170beed6b42274ab13a14adca90d8338bf582d9fdd9fa1d4a4be99c66904404c44d997ae0f8fcf9c33107b999c9ac98c2ea3b2a354ddd5a090e9a24cbcc59d41ab2e3a7f84747144e7386bf6456700f2be51741b43d9b1fce4be2a50dddb3e6f6a0d60d095375cda119ca47850d7bfe0aa2acc1c1912073d3b8d98a4a3c0ce3d471584601359e77b0c02b259d6572bf6b1fc19f2686d8ed49e21bf2d19d7edbbd63441570f5df41e07c9aec3d9d7283f056eaa5e1ef2246896079ed8559e88c8d164bfaa03a44c71841f219f23f74b765598cfba890baeb2895d8efb33520e1f348f2cae9befc19bb44cc81c4868e0634b4721ee4d48cfe4b47958d3bdc2c2c4cb6f9d6d6ba60caf5e662b16060c46d420ffc983e9e529e42565c463ddf752f343732e4f6bac23f385c40b921c8d8767e38ac6017dc132d81bbe1d1de;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h182c3521ba40e5f927eec11c3f2063523474c389d41ff121b801273d190170fd06dad7ba13dc1aafb0feb604d0d55ee046433e351f8c16787872f287266ef267e12813076782ee675b1332d62f074e4fc51d11e570855d84e5a8a58acbe46d58e312e6e036e3ee70905ac34baa88a53ec38904daf24dbf1b87b2d0f2e60cc84aa58b3eaa3669ca1a0da3a1384250d76da14259189feaeb1be873a1649a05b68d2d9b4ffeef7e1bdaecb775a91dd557d055192b86dd1e74afccf682e55785265e3eab0fc608183ac4e40b0d8765fcba659525d19fced38ac8d429a56721d3d1089d92ca3d12f907ca3e7fcdf66282f6f78022863fb7f0d4ebf57cdfd37611290b5a2ea9c7d42bdbf2acb7dd46558551c55556994f9e7a6e906920abf9773900e50f53fc81facf834b53d7fc3dfd6961baf05dc56b775d721f7e0c6667529f5c0d2805503b62b4679a4f34490266353957e04768e64dd73b639dbe7618f17c877a71f0ea538740b594c0a179e4e9f3b5a031b41e1a5ae6c2e770b8200abe47a799e1dfdced382b2e307c3024b9cdcd5b717eaa095520ae4430175d8679a65c96ad7ddba15b0aee5e4ec8eda778a29765425eff850de05e4d92975730a7060fda1ba9679c741fdea548ba52cbb206d76f764422f8a9551db528474045d2d7dddd506547841d8f8dc66f6e199e8ded40f268141bc75ef67b563c82f640d30cf40b32af9a908346e3f8541705e2efbaef239c1c6f8491d05376de331f6b53d5adf3d0b361f71511fc10ec390a98a0764ac8eac1dd555878d814dc864a72d02b8b048154801b59cea70fe4420f5202b2ee796aeaee74ab28f17684e6b89c86abf09989575debb1b0c8d73f4c6b5f3f2b482ea9e85f660788eb860b92c8eedef899b093f62e168dd0781b9f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hc161a20dd2cc128ed66d4d3b6aa605c374b08ce568616af14c56f8980fca750e23de8b6b0dcaccfb804156e4635c53d117108b0d8e2afea2d93da5bf33b4070a8616a2c48b073214d2f1458b2c703232150214340715afe87d38fc33f3b7f186a6f15b30669158feae30439e4ce54b1d8760f6ebacb0255c85865a341dc3a94df8168cb4c5e1eda32b6de00ab834bb3bf946ef3efc137422ceb76ef2d32c39a7decc72039457edb483254e041a6fffca1ca47a76872470107ec6a435afdcafefc8d31758f05fc0acf0dc033545cc51ced273ac0ad7e813ee7cd311ece28f43f66356b7c0ee32e063c8e2bd6becc54a359bf18c0804c6353c523c87218c3b9a96a463f25f9a964bd49f8566e1a25815c9b05c61c5a335224618281506443217cc4d5ae9df9e8228f100c4b724e22d48211f2bc9026b27d2795249890c70fdd583b2c6b8a28d44e356253c7914c686e48fad70a09073ebc2a6162451990190fcf789bcb344ec90b3810130b42da26174fa7641c2a90a6c75056a5475528ef3e444254c1c40dbb1c708c89a94fd24c888e13005e238e91219183376107ea3e309fc9d4d420c27225cdc9b04d8bd068ed199afc3a48a67d067efd83ac643c6563aa56683a9d89579f3e18f3cf74f7ec88300d496d53657c601dcc835df218a96e72a96e1ec3719b27f1a489f593b50643f236b050388f7da8d6c691b8ff4aecf90fea79a1af98bd55a90953438a30acec49f32f93b156c751f287f09e7e1e8826ef469ecf3e3f2c215d55888bff89e5a5c6a588daf16c9e590e268248d7e83feaa352c56713e4a565de11d11952e9ccb98b0ab7e604bf17c310b0e0aa086e276e1d837bf80205051d97e85ee5581b648373d09268a9b9507f33dbe149fd5ee9efc35c478d2c52b516633;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h8a505cc6ef95a5f8dabc84e577af5496dc0dd505dad3451520c8d475118e825133f8a07c270f636ead2f74a358b09d69d96e84f09269499ec850e4fcb1cd48fa25e8db1066b0c40b355d812e1bc892894be00d00aa1b198e6cfd27eb0c195184dc5f4151554672a3c20ddda956e2ffc90efbcb1785eab7f55c9d65b815eccd6237651808954fbe1d75f294e41cbbf87f231c2e089bf5826c935a344a996400b958ba03d8b867a83d5d504209d42c54f991db20d479ee2fc32c41cd43b3886fdc77dd7f5d52e17fadfa5e31098499f4083c486d51635629e0c2c85069ab476c95ae9575d28570046e2e2383b3a2f198e467cf2827b013c283d96b31e6ceb0a54975b1a27368ee626c3fae00e93fcda7e09acf171f0079a6b6c5374dfc6147a92c0eec196b3ef3ed076f320d96e5b836b7d39d210dd0a3f35837df3a7ef3f95838ba409b0ea899e898384f0ed4103cdb5054f91f9bfe695bb9014ac25b87d349a2a6c5d66ccb744a85159af6ce1774a376cca72b645ba0a14ab64442289975fb34434f3e2b788e37b9aa42abd59009c7d5c6d2a4db137ab4c68cf2f7dc8c0e08b355403aa1c8222f22a5ac68901709628102f4790fe66f5f6497da31bfb3816d1d286efe4458c0a2bfdadf9f89fd42f661f84c2a3fb2da2dada738365c53eef6a72f49f9e4bf339356123db4bd95e20bb2a5a68a6a9f836d1b425b665d117e34609d610fc36ef14db62bf59d4774b2857f2d0ffa838212786fe5cdb6c88f118246a0022ad53b0d67e232a33bd0db084575991f724307083932bd64d906b236682dde68ca406b9aac7c29131e5f0e5520df0da6a4fc435fc3d571aa71074ad01f9c51050b61e294875221655cc74334a25102a06442bf67dc01af88a7bf2fbea05ffbe681ed083e0f5a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hff0c835fc064a7d31c0db4a70ac07163260d9e976c775e40cd989480efce6232df868159a2ec75f1cd6c1e7dc57891e1b52299a2c8ff5eaec23e240e8738021da03c87058b5cc4939192c2101ee4116909d852c8bc9165fa37f365fd9d1ab148a79aaa0d5ea870a17ad16c569462d43312da5b4b0a344694630f486a412dab5d33b33c07335ee565656418fa03a756031be1983b909634718a8ba2ee1d7e6b3c32cc224a1e2a527df7d9adbf308c01f72f221fc580e0dffbaaf1e357e82682b985327b407aa6e7f32d13e62e410846f404ac017767ca55294d344c9a9725a69cf2754aa5084c3281397b29d3b9076ce0f9cdc491b377aece1b5d79177027eaf716cbfbba817393e7406dfb8e06584dcdd79f8195bded3e4a1fcba24ac5f60c7bc4475448d7d6e1b262ceffc7d3bedff9c4a08e216ba1370c00acb66c069985017c2374442eccf64a9ac4a4e8a7dd4cc487ccd9664c17474e066b5c9185eb8d3fd7267909a81af88d8029c0ebad9dfac4c8ed3e590104d20548ea641bdef09238eb7092e79e9aaafbe2bb027e97c0eb38cb556629085e75fa4ce5c5e1c57b48e504b0e6e7c0447f0fc791a0703b8bf89460d65bad2b4e2ca29b134ecc486c48cbc3c4c47b5527f2ecb458d3df51c004e67e53784fc58b18cf370403e82492c8338ab259c23f43f253253fbf8121baf2bf4668d45d278998cf94aec2b034e2bdc4cc63a8c83a5767869d8999ddd44987388b4b8b78188f99ef45df57b28cc4ab5aee62fa69c83adeef1ba3a3f67fc6f1eb8eec12666ac11b70efb9d8c8bc6ae4a7ce50afef9861607e7d2c5458229f53104c77c30429ef4ec6ed26ab1f7491160a8068489e98cb936199b9953fa67efddc96bb92ac0cf9c28d99323c0c7a42e4dfe615be91ba0499ab;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hb22d065283005958f30212d0723de86fcb85a6fef8f8bab8dfb2238e55df28b521b78e06236c7c3043b037049a02b72c83404e6cb6816a4c3b236d8c4620c685918f5fad4fcb26a04047d0262187d367d1d7ca1d5558458a982e0be915d55f0e090002a8c40e318829d61af02f4e75c3a830079727528a854177aec111d4dc42fa86845768300052594dc7106bdf3de1cce0d1daf01df4a51a05cb75b26de1b4fee57858c8c6a3bd3a33d3155d6c93a03cf19913b9c16ce7c603638bab21e6910e39e10ad04ebe2e6b2b0d91b80e48e52f930baf5f268d3f59f599b0c91af5bf6fe14258138b6f7dfa01298adf96f03b9576c83eb6639218fd9a5b3db49758f16ec86a9737f9d9000be6c2765ade3521846841b6b579e197adf15cfb3a3c00a68b2e976137844e60671b3065f921fcbe9f4bc210bc1db7f1facff17456c6450e3a5552aa2d29578ee8e2f0953d2570c176217c2f5588533324c89097670ecb99a6ce03dcaeb8356f51b16b3f06c985b732d22031fada24eaf5a9ec56826ecc687169c555c741c477df485b4384c44bfbf65345dc022ded6211c13ab85ef3e49781da11eebdd9528fe79dad782edde2c74ba2f49010ec2f0793adfdf54b10498189903ec45911a05ecde9c678e86568415aaa2a9640ccce9d3cde1527879bebf8ceea671501eddd1d9300dca4559fa17a1fcfa405aa2e116c853b57a23553402ea956085b3e2d6bab1075cec9589aaba0ff07b7926f3bb149057bcd35fe1aa3285ed2995fb9f1db39ea6db2b0164a1314dcee38d3955a825def91d3c01c9ceddfea7fac861f5d285de3e8477aacb2b64e25549fd3335e9cefd3c9a75392ab31e535c814db157990a9570f5b9f97a08761accefe8fde559b5c8d94cb829234af4e6328cc573184aa98;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hff60c5e032b6bd5b0142d4f5ff5ac0907ebdb8bff08884f030efd0bea88e047295f1de3913a09870c4f6c7bae9a7521b30899264b5e8a1e04791c8a9ac0607f6b2033f497a4b0cc29af5fec904b7a9d776f6f3d59690caf2986f600248314dba793d474ec7f916e750e571e0ee49cc7de16e7cde425ff6a146dafed489e58f93176f5ea88211cd8700d719d99f7c7993e41b4730f75ff4f021be11234cf6666c962f701050c4eba5a8ad4d69c5c8b8b3d28c5ba184c0eea50f8b47d64c259d1763e3514f791dfde745501a009b4bad3d9c93856d4c9555cdb4c2c30df142138e6883eb9d2031d233b2c11aa527d3f5037306902049a97c953f9d83a6f4f3916e9229019f6a676fcea330db42420e766ac50533ed3779e98199c2060bc42cdeca8bd4f1bf82e49e9305c3f5f7792de14625b395c1fc2586fd8e6839239cb892d7a03b464009241141ea8e866066fae2f9e29466c9c6dd460cf29c4e7833bbff81562420eba7018104cff546e732705b0b104d69635d18f2a57059be0968ee71787ac4740a6b533b0d451e468b5219e09c405261f7e23af62eaa1f2abc1f52ae0a6d9e1ba64c8763a39ad3b72dea62f2269302251d01f3439302bbe1d20b676f97db457957c60ac4acf072e5e1fe32be8ef85577914dab000205308fc777e7fa7ee0f3c45394621b8c2241c0d122cbed7ae05dc0e0df2b2b61672cbc5b23531084ce83b6d9e22bb37f5221eb30eae20cc220b9e5574f87d52d24ab304a3bc32744c7254500658402109c4785f6b1ef9ead0d8f1f0cc73c65ba95fa1b7cd72bbece44455942a1c960199754be33608428f21f3cdd9216304de18091c2e0ebeb0f6176be0869d7ac96d8e714c65d0cbb060650075d3c7bf49076427902048e24ae1c483e2f4393de5d6b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hd5e0770689e8fe9156020fff9d1efad7e731ac6f876cb6090606b91d597c097ec4795a47ee4ead27c60262b3c5dba1812b63d73cf70ab16468f7ccc8a06de7b5db4505342fb001bacb0e4e0b1c6b523472e33a755c023a5a5521fc96b90ca47c6ba0e7e3e25409ff1fdaf466031a4444bbe922c11d66c91382ac68fac5d81390be949ce09e2cf6d1ae505881f58943d20f713da64e0b7eaacab45bc9626f66b1e8f50e1e5467e1477cf4792617429e1aab434c40a6e8cea96e2f08ad74605f63cfdd0a8c335b5f4d8cf7234474e4e21804a614251cca6bb01e77c66fd50cb99830bb6c708385f2611fe2507786f878f9111269b6532a038014683cad01a3edbdf370324d21cc8121ee48c76b24f21208af3bedc765b07d9215a623527866684330c0e1c92999bbc60c0cd5386dab7e55671669b560bad58e2d1a30c7716c20597178f71afda576e35962f8642a03cbb7bd999250df3ded59c0f259a8b80cf345487d1ebc43fe5e26cc59ef4483b3cb1aef5620da29533e90ce5efdafc9ae2db6713104807000944ade2c957b209f45af8116fc23c0d5f2048e0fffb735d886c4cc95314672932ffa013a82342c6783bfc8f9c536f7cd2554f394b4df2e1921d0c1f06dffd074db4b71545189528a2e288bf5b604a23a4217c12bc3608e0d1976ae3df58ff5eeadfffaca82d16b1461b1df0974f4755073e4eaf734e001a81c138b0305ba5be79b12fd526e26a477c19bd48156a6d6c3af4b959b912cb44ab3cd734ec2591f8e4f076930ac95689067a1bc33433ee8e1a84e80da2a03aa7925aed859a91012b380f8c79099f02adb837b87931abece6505103b4192fbefe9ef28abba42b458417dd534baa62321a32f2447e94fbabad7a9321121bd5aa6d8638845ccd61af00a05f0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h3b805c30c1aed834fe3b0b45a23865ef5e0c2ed2e6445a4ecfcb7b949335753e2acfd0924d1f1e8af8f1294b7e86ac99557dface19e36bf38e95f7882f08deb400baf9f27be6e4b25a4a3c1f26dbfde711ec6160de588eb661877cc92243feb3273b8c50c318dbd7ed8acea4b75b6171c790ad889c26dfa0034f55086265bcf7ababe02c02336c8069a74b8889590978a4b8254cb1552e1f62b9f9b6f25cf68dff3bd49c34db43179f32e0ed8d0b4927f01ade1b22ef660cf9c0cb6f26d78f7c3be520441fdfaf6e173e56fbe6e54180091de5ac83f41a32fa87ecc670da2c74decdd2ec43cd335574b7ab4182bdd6aaf6f25af3d69e15f7709de8feee5ba98fcaf5eed5d55451ff894727d6a932304646ba124cc83a2e7f273ffed1696631e133fa9aff1118aafda1aaf7e83bae15e52b608c7467c7aa632e0fbe9749d696b422f5c1f9ce8b640288b909b9aa1000759a34c9143dc442b7013bce6a66afa877481dc6a887259613ef54179a6b8144b03a84d1c390876c140c3e9767af9e40ab0312cc15a21e9c36c196bf61b114220ee8ed55645e503309b588273d6f0695f9b377b5dfc8ddc626e6dda386a495e7dc4ad662074ebda52cbdf7839e3d7d3df894a70915a60b6df2e5a68cdeb6b321f1592251f79c4d0659562e42776f21be4e30677862453d1bcd78a127653c05ea1409804fd43bcd8a2cdbbf76fc785dc0cab224ed3f95d464bc1ec2a6ee919be59185a1b08e3d7023c98011a430d5905e3ba6f0107e779655ecac5689879a32abe944b16a7d70f084404ca326158ba1608685df8497dc96922e8d4bcf47f73793fa7261a6b4e4da9b93f303a22e042a5f76141e2d993302c9b3b2055894e00d5303dddb03683f17a48eaa9c35d9f1aacf1c67a5bbda875cf40;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hf7e74dc617947b3c9d36c131324f44cbd71e900397a958c67f6f6b5d5292b02c0008b2e383b8c7ce0ce9df622583816c8bd8dfa6235a6f466659b6a9658e70597cf94681bc66b52790ba10bda09ce698472f50fe6409874a299f635b9ad2b22c96c94935c3f09d4245f6c556ea6f8bf9690712650baf2e0de96d9bd17269206f34b81ada4101d58d163c16bcf80868575e04c25ca15114a166094adb7a8ffcfdd9389f419f950bb32093c6388349849faa0ba20659cf1d7ca06179b6c611177555ed3ef233394bbd9fd359c1978e4357eea95f6598eb0513618dd999df2fedd83e3f7bc034b252c0be973dd9407b754830828c69e82092be8f732a3bc64b441e1d9f603ec96503b4bda0f9ac4c140ce05a9851a61d0213709afb333b4a496be2a40a8d6aec70854bfecf1458b3fd44a59bfdc726608520adc5cdbf37786c34194b2c2f2fd94f25af5990e05e3a8afee7ac3f27113600a633609d088ffe026962dad80f1945fec21071142d8d9b9e33f37ca4bacbda9c3dc16c10350cb4af12d246e00fd07360e0d3c581d5f007f66cc9d1e4c7c617d2f89763e4a4e917c1990b8d26bd29bf631525db25d81387c5fc8bad4f4d31a6f02c199e64280c4d89a29006ba52cc3d9e2081a83227832e223dff02cb7749b325a9bfa88ab565af7dc67b8d57ed4d45e3efa41ee695a8a441718531b557be3d92a4fa22742a458d731d6fb4f133dabb1fcab21f435ecbcad9fbde9cbd672045011e991b539ad8aaf2db49ff5bfa467ed119ecd51613f128cb42574ee4bb05a9066a0ab2a668eedb583f0e20518762b162f929bdd2fe91433420be5afe70e202e4f61e5a615e8ae2829dd74627570cf245511888673fb84f1024a5b5fa05c3ad17b90484f6c26a39b066bdc6bc19a62515c01b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hb90ea062104cdce7b4870ba7911b3ec8c1b56e97fe59a4e069be4833e007209f4604add8bbc68372aaad1f733bf493e392f31daf3eded81f8d4b8f94beb3a34bd149912d5de6e116819542b969a294e79cadabb084abf802c855c071cbb77cc3ec8dea6f43a9de41843b8bc168f35cd311d09f73abbb73da0aae5822182093284b021b3568e92c6ae5592dcf0411519a16baab5ba24b73173081ad39781d5f48ff6eefd2069cddc5ab60a1ee30cfebfe006ba56461ca47103372c7896e6874efdee4d615e860df4ad12d2c2cf7ef2fa6ecec617e6444efcdcf0bc099f54ed18e27c5eea93d15f4231fb1411a4a724262c28e06c91c207062128d8da117e5db5a0850204b7f8cdc7b57b10b273e286e496d2f5e3806dfd6588bf8e722ac07c5cf0f981778cb02523795a2cbfeb9c5c96994595b2e328a1aee54ea9ccfe7480631851839351dd06328d428635a99044a1ff0173622a6fe439dbb2aa643e09b583fba7257fea6bef74be4b08ad15aa26a6795c2298159b711b644a69793cf43cc4444bd6d44efd9644af612613c0b779876d5ecb1463148c092e2041540bfe318a8a0265f331f705762074dab8b11b83e466344e170d76ecd217e3b53c76fde9cb93821318aaf65c2b44857b3e49db0fa50228c78f730e6b63b1cddfaa4aa759101c41727365778c5ec08ca3dc876501a0fe2171adca3554198249a39a82f9abbf37842f432cf8a3092132ff566999f07c0c624085485b95ee56484835b917dac3f4f2617a651d229e0070a660fdf0b031933497566f7119dd98d04a52757111be72c783dd4550847996125dafd8e88b93eda8f24a322604ce4ace824ccfea9e8dd25e99fa03c5422f4c236248fee4428f9f870538c1edadaf7c24acbf15a6037a15c47bf2db3cd201e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h1352e98d26f73ad69898be25e0db1b90648eb743e1aea7bf1f026e0b9ed30cd6f595ef51f407f853b8ed5a968bd8d3160cbe99ec2adbed4a7d1090dfc1fca8462b7eb225f2f3a2d2b68ad9f09d14bd9f948ee9945bf9ca65eb70ab4bc73f7dffdfec4af207cf2a760cf484840dc81bdb4c03997747e5a8bd77a73818a78c83984be64630ec365e3b9ab0a503c1cd1852b82fb830dfc124289afc17590cfbd515dd960f06c64d80116a3c83bb9f0330802fd40476f3738be1bedaec646216e29f3e2e80eb4d4ca3569264f16846793e4e794bee7ef8636a763154ef9758a37453a1f5dcabcca0c13086568c63bcf8f2028d48f8e1fd06fa13a2ac7e0c5302dbdad9cbfcc00876e08e69bc52d014a1048eb4a6f6e42bcfbd6248727297c5dfe8e7a51f45fb1cfd1eb2af58ece79adb79853cf118f7963eac27f2e84fd8bad177874bb55926b5a05845d10cf3682705e04e3bbd5524f62efed4d482474bf0d705712cd1fd177564aa82693e0d46507642da3832cb4cf9fbf7151827918607a3c7b450bc48c3d91feb35ff6c02c9032730cdde306353bcf8388f26b8c88cee97037525286e2039adb7c26c6cef0c343b5b9da41df7eec638172c3d86716537d17c3b0d5234e904adf77e54226e29a82719c90067c1c2a53c9ab43fb88ebee11f43b4ddb8cc80a0c0dcc3d35edcb70223d9448a29dc693ae3b5a2491fe84ffad9dd38562c21caf34e5d9aa6ea197c638ca6f3531849f407ae475a7cebc9a5bdc482fe125ccea112abccfafdae62a7932786f74ec29fb2ddd282c2a76f08a4a7d5d4087a4757b272d8a2f630112ec6f66b9b7adf35b57ae7d2957a5aadb68dac5b3d35a3c8a5650d4a7574b551a6733957a03a66346be5fa6144df916feaf164f4c4d12f1a96eee4fcc6a9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h32faa0581f0479130753cefbbe779824fbbb1945ec05aa9c1ed5879c68890e0eda054ea510eb99b8beeae837d2a808f4a4eed5556922423321066d02baf15109899a83ed5ac979f43d4635977b77ed15805e6ef9577ee023d5c22bdbb92781a42b06b36b3fd5cbb33a399bbfcb758c82c6cfb67408cd5e87a84c43f9998d8e01000decc33f9e243ef43422c02171a39bd076c7cfeaf46c3c5b5cec6526ddcb4b89dd55525b7785dc856d828403f73978d79346590c33c4b13452338f6168771ce0d4b05e2e28e54c509365683de0106fc8929db33523093048807d66830c19e565f8b7e82c57a7bdc67a760d58c57fb876326055a615312c408e598dea04691fcebacccc705142f3f16d8fa7551ba3f3faaa8737854152a64ff9938381adbaa3c0c119609035091f1c0d6bc136766ef479e61d43dc0e57313a2825c55d2cada5c0bab21e82fd3d58c1fceb691276eb49e24473ef1693f784ac57ddc53d958d78ddbf889a6624ca825816e4f9d505461d3cb8a6807ab5764faf63f18d8eb2716b8fac3d38ffa8a3fc64788cae6e4d8b79d47e0d53e722557a4cc3b61cdf30a40366f922656ec338094f76b6057ec175cb99b29e6e39005c6a7be67719214746df4da558eae00cc203a66a692d09a0d20a149835f18292176f21b496956c802a16aae1bc1afbc033ac742dda5fa810390596cffdedfb498329e5bef40c478b89e480d7029b6296a37a0cbc453766d64a482d4fefbe11ff929fdd0fe7e33c6e62038edfca0f9961f9b977dbc2625673871faa9387f696eddfbcdef3be021a0631b1ce919f743d74f67c9a9fd6e96352c71bb94a819bd430ce67ff0e32b9b6231a85e75366024538ce759550f9c6f4c3ff049eedba4df22519c5bec7657c57763eb39176ef837005c18d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h508c41d0dcf4664e8da1bac6ac0223b2ed5df584aec8a14c5f347ca7411ee6621a90d2644d141752a93cf7ca65319a158332e952808f7c12596bc796d6ea117bee092fd55ed8aadf768f27bd1672090cf1fab5cd20d5989a17d22831b8cb19fd0c7f1487f77e29ec1d16e31497e676c350ea065e140a6f7efb0a2d664990eb098f7025c6ffff6f3d136f494c86b918deeec49d7f74ce4bc45e68a17c2495c6361880c9cd22cc9a0cbc01d257bf587ea741ab2ffbd6a0c2d393fdb246decf47bbb3c7de71a7f7f0964e8362d19fe52a172493d9039090f6cf83684fa4742744bb84bc928a2875928aca6177d3fd067452cd5ec82460c22aed9e105a65927b1c54c16f3171fe32c771e8f31355a56f5a3f57ace99cf388d6fd0ae3870459f2e36ee321c66957de4c1e4b9192f21a4df1c802c7fa488edbe16492e1e18f7246d4e9abe924b0c159522b0850c66c276ec44c07559a7dfd1de17210c4f12b5845c1e6175894c56ceba50860834c4ef948289b98544ae8589473360a1d066c91746a09682f9fe488443f759313a6f6ce038888ccc48b046d7d2ef65b038cc27ead6acba044db4998e7150c7c45111b9bff4761002ddab8b130db3821cac64b50e6d77fc8689c871fdece67e5547b71381a3ec049973c2605a55f9e22a3ad1201034a10c24b3f80d68d3130ef184306e3163bfbdb64bd1c8f2d300ff22195407b609b430cbc9a0ed48f3397a4bc0264bfb250c56e742aa5def35f6c7da4b17106f6334356bd837396e4eb9be23b6fc66c42fa51a8ee7e546207441f8df94244acab01668a4b13f832011f31a7f91b3910ec3659ac9aa8678fd3202868b7b4ea52960d06d7f0a3c0c5802e030d3a2ac7d4d3772c4bb8164575a1276a51842050d534f902d33bf574ac24fe40;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h52e533eaf14b96b603abc36aed90e13146c02447d9bc5f3258a8371f4b280d2c32efba653b48acbd2bdf3b73d042955a9b501ef4dba5a69762880850e1bd46f33e275272ef1126013ecef5b592ff08bf55a921f2543eeff10f0eccbed5280f2589fd3123be6ebfbdf321a00f913d5aeef5f8ec37962cb9a37b1081dc07df6a709aa599dce346df6278cea0aed70543cf3976521d3416ab4212b7aa153d652c753a983b0b4be6ffcc9b55a033334d5c605a1173cd027b77d044ff2f47f650000b4628f05c3b874f7c5dc981336833e427a43ce187aa05e9fee21b656c2db8878d6021be99074e0548e19b6efd04ee7dcd5c5f57168eebd94e3fd81009cc2c351b18965818d273ec678b932a9ff8b15dbc35283d15f5e65293695beacb7d51603d437d0b526373d57d410c3c370b409f3cbf1f55375a35072ba0eb0bd8a54caec0313a46f37ec086f5e5604df1da70496e897511523ffd683ee71d13c524e7da037ff5e2e358a2517c92c6c5c963d828b83f788a1513403a218489f2a067b660ffdc2e2f075b5e006bead6b3ac2c4da39e85308d5bdecf6eb5f4c932c02539417cd773f6d62d9cf859f0c5f68d61d7a8d2b4d94dd64fc5836c8e2477e345b3f0f905ac8af9051ea8b48513f495a9aef1547cb093421640687d2997daf965eb01feba4a5293f5d52de747f3aac22cfe11843ede2327be31053dd1caf98a82ca140ead7cb1d680be3eadb7efce4fac2763cceb26722c8675a52726eb381f6be39ada357f071c23c437df2d45e5d7a9467c055d1bd677003ecd102dfbf2467afcd9fc8e00a44a4bdc89e56866213478039ffc7ffa938e5fa385485802484063b87e63581f786507f0972d6dcdc0fc8e898e7670cc9c6ec4f3cca0c315a6b01b14daba178396caa2b96b30;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h17f5dd8517f5f9f98047034df5b1316db9ade590236f67d1b3edcf914db5e7cb944a17cb893abe80c97e0b57a06c706f521d339dfb9cfbb9e689fee9491061396f35429a99f62e60e322df3651ea1cf9cbd580376c9f0ca397a1057febeaa10866bc07a06f530b676600a1ec3575f2bec0087da09aa3c0128535f32d932ff6b118881fb501f3179d4020937c0ce25042a9a39f917ea2279f9be12de2c0d0b255d613e8ecdfee34d80b685158b85d7e5789a26e84180b15d7ea3ad4ce756a273b19a951034fac4727d031cff342c9876526e69944b50ca6083d4f08ad05d874837cd00d8092292263284a80eb2ebe1c0373669af86975e66d98022cd59a01d87aedcb0dbbbd207828e97159e23cb8cf835f41f58c9f83dd4f69aee3992f43921d57892830b973008999b23ca8c5c480545cce49d62b9972a8c4a262c29af15bac0705c6bc6857026bc45cdd042c978af42787d9051c423f532206b0045d7880037ed363359642bdcf10244a6d7dfb39b6603760a4daa5516fc335cdcb724dd536b05efd144107234ca7d424762f55049ab6ff9af1f99b0b8515aa8f63ac7a3aadf168c5b8225e4950a3ca2ac32b99f33ae607c517505f618baa62bf06d67c5f0b19048ad8f5058fc6e90bc687147d9e19a1d2ebf497d3fc658b467314a95981f1dbdc938d220cae7307ccde348a1309ba6e1dea78e9f73e52cf8d26b30758175e1c2fb7db4b3490935bd12eecf9c15f3602c7d077508ea34364da014d82462a14e1a20cf63b6095cf03d2bec91b31db8adbf8a13db14218ca1cc9de7feebefd5fd6d9ee7cbdc3eb0bc9308e0c05e8145bcb7974b2eacd48f7866ee9d8fce8e7ad708e103f2f865ee8423c569d0e46fb57f523646e01a430ddffb3202d2f21868cc397dd7c55e85e8c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hf7ba53c6e1d01f15997156c4ec00c92fc64511466bc50c96b0c6f7daeb22b36e40a1cb78322a8300662dc2d7fcdf505be7b81678faf175559f3f2e29f9a78f9c56d06e5fdfe3b404740d43075b2556688a3b94dae1817e8afe505593d2d5ad46be33f600c70f988b53db72161cf2b24c7f40ce1b9f1718c60398ff80ce4cc133a9f530ebf7fa594478b12b4902a573f74e0d860044badb8aea5a312660e2e0525b8dd1c50871caf303bca97ead7f91f54516ae57910ada4da3754b9c6b00482f1c705f6e36a11387bfc9f47e3fc32be2c9e45cb3581a8b21257f554ae92a3c4c640637aa6f4910a5c10bc0fbb8a04bbaf6dab40794d70ea992a7d57e18ea0540e2b519bc0fcfba06dcda5d50ac179ee2eb6b358c4a7f8dcb66bb74e921bba6520a74e49e8cb275e1795457ec54f4060290fa2af721d0129c47bf6041e4c7388cc7d2c501f4d09ccc28feffa203579e538492d4539276325213154cb09826d4fccb7267175884efcd67ac2c9ae36d87467b31146f4c363bf8a2959e175db12e482eca69ea5132997cfaf2d93609850f0bd9435281b6c1b4bdc581902565f925f2feda8f0a5dc29e5089de2d9ffa1e7b0bd5d8a62061ae3933eb21cea8d3b961b8c59d443aa76ec68f1c9f0124a6bf9602f17e0bc716e78ab964d1c0f839b9211b25325a161be1c5f8b18743d49bbccff8cb9c3e3fff080fed141256bc9d33f72510dda13dda347d21de642d4e59b42baf002ec3f24f7aeba0e3aaec921eff42c50c424ba860b07057c81064924c8f2bf4f33563b366f831f2b3b99e113d9c5df018b7e220ee91a244624b7554329fce1e07227d8d2a760212117c265692d14c3b4381b0a3a261a0a9808b28ed23393de325ef1685ff5334038307056d5b3e322db8a64e0c719d36;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h3a9a1102581f4017c2ea449f80d6ba1169d55a2afeb9c06e9d0ea481cd18595e849eae88c9aa59121be824a3fd4c9efb5af767a4c2a96673c1ccd4ec432d25401cb1beffb11dc234e62a4955768e0a5d0391e3ce5c9f84ef6484934d0f17049e8eb545c85b5f3aba34636b150454e2809b72bbaf1e3b74937d15f3a1aa1e8665f4118d85ee4b34e05cb5777aae97e591d7cc9feb8f7837fe0e4f8e960c891b81927cb98a63fe0e0afd9d78aa6dea0f26ce8c6af40133b3a1235a6897076eb2c2d45efc12fb561968ed560090928602879ca5ead7f5c630b031bf2546d36518f80ed6ca6d2a5d88cfffd270290166fea64dc7a788909f66cf32de65fce39127bf26c744c12e31178a74b619182ee6c9af86bdf46a800a8e57f9a159c3ecefc457b9c97cb0ca5125b018f14958c8470175d93900cc388d3b2de9c8cfd75c4d9777e381461b3be597f8cea9a2387c68ae6eaec830c30bc482d6a128412b7159e55842bfc60f4e3dc25f0e26b64129b2c333f1daa9736b35eb21ae1460434a99f9430b7efe9d6039ed58d0cab6bb788caf64a78b4ccdc15baae2fe2fee158e49dc033b944b9fd667def2dc9d86eb6f30f59633378d5c26e8fff72cff3f9e841ce1f94584c4022c52a0914d2e8dbe39b0ddd19836cbc31bc8c89d8153d3bf756bd8e0b0af08a49438739f60fc4f10f559eabbcf22383a4c4078df3a8a1934530a1a742662d8e0748bcd01fd2b380c7507bd2bfa04ab8a2ccaea29e96c4570e410cedebbea5d57495dc5f98afe72fe58669adbc9336146eac25f91ed2ef6cf3892058115406df628197d284affd1698af598b36ce2f0f8c68acf75f59a8f0a77c19666649c5f5d74b4290318b1794f03efaff09bccaf0bd8b4d1494abe9862da22f9905bd1b96351e0c8b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h4198acdba91959f9915a4228a1a482b3111461c31f7f7c74bac6d11ddae78c5a8b286496636e558bc5623f08f7906a0f4904d424ee3d4bc2b0c1630b81b7defad7d8f7e685638ca712547bae0475a2950e9383b998deab4e6e83443fad64922f35664250e41dcc722da3c9d293089f95405cb2682a3fffe1aa2b8404458113f47feca41449f98cea350bf809911b55e16446d3927955f3da80ebec35662237c2029dfa1e7734357407d129977432ecae5f06e1460c41c5ffba3fb3cbbc0de03d6cf8b8bbacee455b2877ba8e634b8af1c6dde15277e5e4d119e090353a528fc7943084c7d26a0980137782bd0a63afcb209ea8c3e113a60842baae4ac63e230355675f564aea3270ed6baf098aa97463e5a42572dee3d8af21932de092abea6e6a3682bc04e5d21dc1527146eb4d96d5abd734f976622f6dadd9027f3958396587da4199a7e4888380b851f94147a6a404ca9fd0c7243f5f20fdf420dca3f48c384decc283932d0d848eb38313f749198365ddb9c6202a842b7ae982d7890e9d3454a1cb53942adc15040c8b2478a9eba63554710924893f5a3a4d8f5d8b12248aa71c268bbaba3b324543c70d4ee7e1813ba0ed1dd8de5638f4268ff322ce3ae02596cf9ac64987aa9f42682754a63f19a7238ba6c0404d208a1064bc35d6800ce2c286f30222c97a66f6a7ff49d00a05f2b1ff845ab077e233ed24463d0d789f0583f9a8859a740f24e15247b06572878128b0588975b50c588cd52ab81e4821e936bc142494476aba93c576955b040510eb08e1299a13d451aaffcb1fa7730082ceaf9afc7185b820292ae201fc5ace4805316bf42964b8c1165d6967f1051988c69e370f97681b59739f2fedeba3daef015e5a350f90f4ccd68414d7df247d17d8d40c0fc322;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h439ad27f2061bbbab5bd62340c26317d5fdecafa893d642170dad6fa5cc2416444e9072e9530c903f3188a2471ca86139ed7f18274620eabf52025028453c32ece9407f562b103ee16ec9f8c54c34e8b770c79c30badb0b95a1355b1e525f57e68ea79599634dd84b758917f3b1a540e861d84c8ce3f51b7cc905688b7e3ceef11a5bfaff74c5fe12364a7ed6d3a0bec10ca65976044479acab2273649e77b6d2da6872267e348e5037ea136b7f74d62509eb1283f9a1e480325c0c8eba2f2dc2af4a304070b222481d9306ec6118dbd3ddab5ee176ec295138e110f3114e2f89d51b2ff3fa905814dbe87c0fbc849cd88e9545e9bf8701bf69b72fc8051b6a12a96c9657621c2cd23b56c5768ce3ac52f28f396c4133572e2a42a1dbd63d88036a2d3c5154fbf979ce3a30532ae9a081287f935688f6e3212cd12a5b850777e5446f22f4573a680ea36e38813dfc8ad30312f4e7ab58e3a4bb0f5d31bbe7c8dc0e759bba728f3060ca495f7147c2d0d8fd6d9aa7b74366b170d1494b227b73006751d15eb188a0035f5d5df66c5a6bfe0c856808653831172912cf309b86f18ad19764ff60deff09871a44e36f1b12be76944073e2b446c2d625ba5b9a540ec232a765979bc3895f55e82a89d130c0171ca30f87724740e8540bca6595c14508c9256b181e0741db8f6d4e36973476533c9d49ddfc2a7471d59f4e691ab37780172a6c2a9427ba3cb53e463acc189c49e23ab2a0cc446ccbd17cdcb7c969362015d3dff4e03b2003d71c5f953fbb4c8b792430d12df72a0f5289510a0ef707489880891c6a547c49f2319f600f660916c915426d2f4f90a97a1b524021515d2dc393da780d32851d7bc92c4bfd1d111f62b86e8442d47fcbf49beb247e5d4de391f976f8004913b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h9944f1eddd849531f00171bf64f21598f48e4d60d3acad12f2b06d9eebe958407ab4a0da13934a5599cbc258403c6db4aba03f1ffd3e359ec802e055cf1a248d1b8d4fc494d6296a553852cef386af2adead2e1cde96f276a3b7fd159509c50c82d9aa50336e9ca8d88334695f4da7fb42baa3b6d7bcd4e42e8de3bfe205a0648b83dc524e1bb4902605f2645876e43ad515f2c03abe8b9d09ba831d6765dea6dc2b3cae9c2a80b0af21a6d28e4c201d10c7dd33754898631793ad98eb9f5f5a1945aae36a0c7cea5a3c3041f857df9b846cc41f0039eba5da59d3ea5239253f5ff569473bafd2d1ddac2e4a9af4d6b538682a5c38755acebb83ebc4d04b0caf613f9b56ac4a7718e4a16ecee734e4110544108754573443321f77e613dde96a559d52fea4afe03f14356a7b9a8d07d9a3aaa048c3fa9a9dda6e3ec0afd0027690d768df9051c748edfba7aa31b1f301dedaf960033b8f85d1e5607b4c67e3b64488dc925653e10e2e790125e96c51e5470e8e04b84be548fdd87c7b8a35ce4490fe6efc9c84f97d709962142afa8059c29d91c488bd7888b05728e7beba75606954417f0bf4a66cef3cae5cfa723d33a4434846dbc8df98a284795ca6345473723fb9ccf4a984d32ba96e3df57488e1c6b9a4039ed61d24db4bb4c6e5bcda81d747747f21501dbc8c52238f59b6742d30890f6da57b4af502bcf9719741e8967faf6dd2a038ec016f7e6dd43d3bea05efeb03725815f3a639c16c55dfde4ffcb11ee82f491cc14b22ffb0ab018beebbc44d0a06063aac8ca9746032b1146d7bc8a91fef644f9756feed1249274d8d8f1f6b6191d98b03562ad535f866b17f5b31a94032fc4e951ce0dba0929754e6254259d896d00b51627301d0662b57a247db6b9150c1272c00;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hc9eab4ed1af22d55f5a24913463aa9dbccefceff5dd03ef051fb9562517f670991f0f6014784905bfd008cc6934152951c63c86cdd28847fe3e302eb32fd0e263e816f65c291f9da6d5adfdfd4d4a26367eb3930cdc05a093785099b63045ed51b9b8eafd2c04b796bc34196c30a4f61307741c03e1742884429a618bbd239cb977a0ef043f048aa00dc8b10f4857459ab244e1b143c698629767c07c38579073fec27e48ec0081a36bcc413fccb2289d6d87b22ce876a8a04fadbfc7acfe5595c150382cacabb4ce6e7b2db185d8ced26649d0f1b70aec066f7c91ac83ec975fdbc56aad30b4dd5afb488411270901b7ae36cf4b9ce49efdfc8f12f42bb82c41dd3845e46c1b03e2e87caad013af78ba2a7c2cd2edaca4065eab60ab1f32dcfdd503624294ea3dc8111b7ae8aa0869a53ab50a920d060fdbf914abb92746c63ebf4f6e9e2af92956c2d826d708ce21978b64c0fe6d30ca5b92e4b0b4e3d7b0139f13504070f17f7a06ebbd0a59a8ce44b6827d505ec35955184f822031e56bc9307386f36ab3b2e1b2b2ceac839af41fbe19a635728ff37bad412d5dce1914f06f20686878cf72e2914a07b32bfff65534257327d51ac4055987a532f03adaad10b9e94f1ef3ea828d4d8b9b57c1c0e1d3bba3eff6edbb3d3a54491ff4d680b6a43b1af04930e120973041fa88a6de755cc22a14b60d382b3211eb4ad50850c8d1368b984710bd4c6aff20b23debca7a69a8cef3ab7e846f624e86db49e3be3c75538c1a45db9f97b974deeaa9fd952570a7941009e4456182c569c97e70d3c119d1417a0ceed3bb0e41c64695547a8e60de060e51298f9f0e30b16c1db592bb0356d27ec5c8752bef901456396a1fe6ce5340572f40acdf74425c86c57782c308cb70c929f27a5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hfe00cff57db48ba255a1ec4d443a163244681cb154157027273a342a7a1cbbf2aa7a14d836b32182b82eb9d3addee68b8162e1f0b5b215e48e244532d57b3ae398a8e923ec1ac9fbd6dad0b9b8421932653239f029dbc59550bec0f7e9c2ee99e7ee5bea669e5e59341faef45c23f608ee50df4e21bd598d2dec5669a48eac35d2992c328670cd9703e4906e54400970e382771899ce97cde027438e4da203a71f32a0cfcb0a22d44b5628bbfcfa0518260862b45f1faafb71157b188a9d315f4d9c58ac9171148fea6625bc92670c5b7bce68582bdba7ef479d3ddbaee32a743f6cb9801f7b7ec670f0a7635f7cde85a4d08aadf5e15041b94cf4ff04c5b5f3d3e98a9f0a32849f41f7bcd849e41d2de8f66efe2596996b2450113e2b36c1f4fccc56e19c7451fd2934ed5884bac7d209fbd2aefce263d551c779dc3e907e2438a3ec04ce225a852b3dddfce0b4c36f4d0f65f7b06ddafa6365920275cd37b9209c1f5250a6df17d3a3fd685e9a88d9d45f0978f4a0eff1337f8a24cf761b700316961169a3a50dd7e40d7101b426c2f2b91112b7f33635d451009b2f4a94cf1933dc249774ef253ebd26141e00e23563e9227ea182271cc318e3936c180333392ff637b0523f60e70de3033daf8d5a3144f0f6773e5b47e811f5a93e3dbd9e88eef761df2c7f951e530b481895a4e1e764fd7f261c70c380072c83b69d8f271bbd79e33b18284ad33aa9600c018510c70728a5808b15030083f2b779d6d910e889649bc83158d1d19b2f6a6bb8f13d7654d964cfd5502f9e71dea68baff9d61a5a6745db1b7d364ae9c76d8a25680995f363d6b4c87476f0aeced733477473ec91c71a7741f8124182b1036d55f037d5b6245e12c06b5eca3e63f7b5833af4ae00932923402325;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h7e297c5d56e6dd0a3e02bb5bf166dd588fb3049a19700369c2acbdcfbe7a3001414fc11ff87a2cc551f0a8d0ab5e0b12b0b52c6b0a5f00c8d50049560d0c3e00426e77f02d05cd6b84cf12d251bc7bd784c467b094fddb17b62bb5d33b7027712fb57f4dcef1b56fca6bfe57308c91ff33e5d4e3179e8391b9fc1f65a426c7acf8215db69a0d447d94ccd436324269d27cb8010d58865cf6f14cb6b8fef4e06e34b62e50c4b3daa388bade70f2bc8bcd1573d83f0e497ed45bf4c69019355e8b74d9682a321c4d7b866504f4de1319f88ef8d39710ef1f8815f58336685247066875fab016e1e9a47791bfe6f6738042f23d2e4355ecdf3e99665195fb5745c504c82196ff24cc43e7872e606db647e45e6f3a04ae2a3a8eb3ac1bd69b016eefe702d73d6a90864292b5dc0201655a4ccf4d30865645d35479129da1fe306e20f25f9ac1732797c9dacf6d4d16366bdf920f3d1a555673ccfdb5bc10d7c07f00a77e3b2c4e6867e75f736c82151b1915971d3a49eaa29dbee8afd4b8b85d37cd8607313641eb9aa02e3f1827445b3c99900a72cdadfb741ea63f1b5a6069f3efd266cc6b4f7c61de790c3216cfb881a4de69e0d373198a32969eeda688868dbb9259dcc83431c2d5352d55994b42a9f31572572d3f9e7e0d3dfdd3a9860eab40944929035d9602f929d7e9f866f787fa929808ac49becf7dcce87d2afb0fe1adeda0af7d4173305f62b4942c211725f51de565f56fc55d31d5ef5557314f60df2d71145a6525632aaaa039c7321fb21c9c2233a5e0a631a240135da481ec4e1343b6395269c9232a0c416e1cf6f29d7edcca5a0a0000535d0be82ada8b56161c93a0c35382aef7b00519c184751a51fb26d5429901fe7c5a5455fee765afe7f442f1bf180dfedbe5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hf7580e7b9d357f9c6e769c5eabe73d3b9af55fa836187e2795c8b412c053f8f5f8bdb9ad8e33c0443b9d2105e040aef99cd06214ea5a2b0dbaae27d7af8e31c9a46dd00accc03698921308db47bff3a9939cb246efdb0a5caec53d95659d5806825633b34b3753651eb438ee489ae16aef40fda83d183863883c973b2fa687e107975fcc83b5e422bb6dc762207d4262f0a69055ed056a824d3a6b45bc752e4dc1910621b84d54c6fd672f48c4d6bce21273194bcd6fa26be106947ec8028edd0c277d0fe18a1fac181ae1e5d70e05c5c69cc4ab41ed74d99ec070506fc51c0b06e8bd2b7dfa4c0fecf6dd889257d0db613a334f73c568a93d25c2d5052f46e75a829485dc144cfa0686b87fc56835a060d5631e323bac4672af710c812f48700cc708a4b7e9facb1617503dc2079dbd9fc713e95785bc06f25828d63ad3d347b4e8752d7441c2945f851d68e0acd6be220a945c49c22ec06ac3ca1cb9cee79c1160d3ce0155178b2978c5094420ccaaa7ef883605ae4e752d2f5239cfd71278580ceb0d98ea1148994f19336f504bf5aef3d53971aeafc9892747214b70fe732303341e3e834507c5f7ffd67049a4f06ca9a8c05cf30438e169009abaeeb44ceaa47deeb567679e489b8c0d223bab1bbf096d91d282e0d6ebd7bbc74841a14bc4cc3486c8d2ad8fa8fc90f6b5483a00db9060ffa8d564b607a04381ea02cd32095c14fec6df118519329929aea3ad5530897b2a99a885d5cd39cdd256c85714213f6574385062c379fe1162901d080ae2590c51c2189f75fba2ba0aa4a7a0d1e9c7a4395ef4baf5cb089729e570ccd8350f43232552015bbb0ca894dcd11d0a22d441dac10317cc14e1fb946fb7be99ef34ecd3209b7a03d4f781e97e561530b63c5cb349d67b95;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'ha4608b224026d619543e7835f09ebf6b5fe9c19ab53cc254121a52806526e6135346b4d3f0b6e5590f89028b55fb4ecbc0a226111dc122d431e89e6e165c7f64f492ad0ce85fc3a6491aa67cb13b963eb1001edbec79fc8ecbd2dc353f793b925e041af10d150ec5a82e341eaf84694a95f19fb1d08d299bfcb6c1e5ea53653d5745149f8a80910f670b1bfb825142a79af1329ef1595e881e3939d7026db4b8f6d6c76f135446864d624dd1cfaddb522a83733444a27bab8bde55e8b4a0a96d8ee85430339dad26e209a8a7ae08516f0f5118867179b07d156cf10da29014876885b1804da07a39a245629a874deaae0eca8fca9a3ce6c6fc02a408a1c89a9bf68778d2c820cdf539c04d685cccaaacf5773d4d0401a3e6eb474d87f3d8adec5e6df11d718ec89e5c585aacf17910b92a2e2a0008a41ba5eda792a2e33b83b04207d41430ccb004ba170e1e9bdb209f713646e79263235283c73402085951b9fb450681ca755d6227c5e94f38f9855692d2ac95211b43a457f18caa6bfaab7e3b92297037e95d80304235e9cbd86258ca1aeee7b4e1bb5a31c0a6b98e152d76331e7b711c41ff2bf31952685ced3b987329927bce3df24369f123cce43e9b749066172e48110ae425030bef2222157d8065ad7109892b33518329c7a056293535238fd1a81da475cdaf4099a0a6acd85ef32cdc2d4a847b7fa11087827a7ae86ef3f71b1b8e5037e2a533b545577e0a7240d5732d1953b0be7d75716b5c3c44f74979608e1181d51345a7fa9c5abed7e8432289c7a8e344e469f548f86b4ba1faa967bad0d15bdafe06743e70381a767813d053ff6d6402935122c252a2f70fae01cb891eb4eec494687d49a9d0dd5fc9e375c59be532a4bb2e9759f5b2884226db17982743853a;
        #1
        $finish();
    end
endmodule
