module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        input wire src32_,
        input wire src33_,
        input wire src34_,
        input wire src35_,
        input wire src36_,
        input wire src37_,
        input wire src38_,
        input wire src39_,
        input wire src40_,
        input wire src41_,
        input wire src42_,
        input wire src43_,
        input wire src44_,
        input wire src45_,
        input wire src46_,
        input wire src47_,
        input wire src48_,
        input wire src49_,
        input wire src50_,
        input wire src51_,
        input wire src52_,
        input wire src53_,
        input wire src54_,
        input wire src55_,
        input wire src56_,
        input wire src57_,
        input wire src58_,
        input wire src59_,
        input wire src60_,
        input wire src61_,
        input wire src62_,
        input wire src63_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39,
        output wire [0:0] dst40,
        output wire [0:0] dst41,
        output wire [0:0] dst42,
        output wire [0:0] dst43,
        output wire [0:0] dst44,
        output wire [0:0] dst45,
        output wire [0:0] dst46,
        output wire [0:0] dst47,
        output wire [0:0] dst48,
        output wire [0:0] dst49,
        output wire [0:0] dst50,
        output wire [0:0] dst51,
        output wire [0:0] dst52,
        output wire [0:0] dst53,
        output wire [0:0] dst54,
        output wire [0:0] dst55,
        output wire [0:0] dst56,
        output wire [0:0] dst57,
        output wire [0:0] dst58,
        output wire [0:0] dst59,
        output wire [0:0] dst60,
        output wire [0:0] dst61,
        output wire [0:0] dst62,
        output wire [0:0] dst63,
        output wire [0:0] dst64,
        output wire [0:0] dst65,
        output wire [0:0] dst66,
        output wire [0:0] dst67,
        output wire [0:0] dst68,
        output wire [0:0] dst69,
        output wire [0:0] dst70,
        output wire [0:0] dst71,
        output wire [0:0] dst72);
    reg [485:0] src0;
    reg [485:0] src1;
    reg [485:0] src2;
    reg [485:0] src3;
    reg [485:0] src4;
    reg [485:0] src5;
    reg [485:0] src6;
    reg [485:0] src7;
    reg [485:0] src8;
    reg [485:0] src9;
    reg [485:0] src10;
    reg [485:0] src11;
    reg [485:0] src12;
    reg [485:0] src13;
    reg [485:0] src14;
    reg [485:0] src15;
    reg [485:0] src16;
    reg [485:0] src17;
    reg [485:0] src18;
    reg [485:0] src19;
    reg [485:0] src20;
    reg [485:0] src21;
    reg [485:0] src22;
    reg [485:0] src23;
    reg [485:0] src24;
    reg [485:0] src25;
    reg [485:0] src26;
    reg [485:0] src27;
    reg [485:0] src28;
    reg [485:0] src29;
    reg [485:0] src30;
    reg [485:0] src31;
    reg [485:0] src32;
    reg [485:0] src33;
    reg [485:0] src34;
    reg [485:0] src35;
    reg [485:0] src36;
    reg [485:0] src37;
    reg [485:0] src38;
    reg [485:0] src39;
    reg [485:0] src40;
    reg [485:0] src41;
    reg [485:0] src42;
    reg [485:0] src43;
    reg [485:0] src44;
    reg [485:0] src45;
    reg [485:0] src46;
    reg [485:0] src47;
    reg [485:0] src48;
    reg [485:0] src49;
    reg [485:0] src50;
    reg [485:0] src51;
    reg [485:0] src52;
    reg [485:0] src53;
    reg [485:0] src54;
    reg [485:0] src55;
    reg [485:0] src56;
    reg [485:0] src57;
    reg [485:0] src58;
    reg [485:0] src59;
    reg [485:0] src60;
    reg [485:0] src61;
    reg [485:0] src62;
    reg [485:0] src63;
    compressor_CLA486_64 compressor_CLA486_64(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .src32(src32),
            .src33(src33),
            .src34(src34),
            .src35(src35),
            .src36(src36),
            .src37(src37),
            .src38(src38),
            .src39(src39),
            .src40(src40),
            .src41(src41),
            .src42(src42),
            .src43(src43),
            .src44(src44),
            .src45(src45),
            .src46(src46),
            .src47(src47),
            .src48(src48),
            .src49(src49),
            .src50(src50),
            .src51(src51),
            .src52(src52),
            .src53(src53),
            .src54(src54),
            .src55(src55),
            .src56(src56),
            .src57(src57),
            .src58(src58),
            .src59(src59),
            .src60(src60),
            .src61(src61),
            .src62(src62),
            .src63(src63),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39),
            .dst40(dst40),
            .dst41(dst41),
            .dst42(dst42),
            .dst43(dst43),
            .dst44(dst44),
            .dst45(dst45),
            .dst46(dst46),
            .dst47(dst47),
            .dst48(dst48),
            .dst49(dst49),
            .dst50(dst50),
            .dst51(dst51),
            .dst52(dst52),
            .dst53(dst53),
            .dst54(dst54),
            .dst55(dst55),
            .dst56(dst56),
            .dst57(dst57),
            .dst58(dst58),
            .dst59(dst59),
            .dst60(dst60),
            .dst61(dst61),
            .dst62(dst62),
            .dst63(dst63),
            .dst64(dst64),
            .dst65(dst65),
            .dst66(dst66),
            .dst67(dst67),
            .dst68(dst68),
            .dst69(dst69),
            .dst70(dst70),
            .dst71(dst71),
            .dst72(dst72));
    initial begin
        src0 <= 486'h0;
        src1 <= 486'h0;
        src2 <= 486'h0;
        src3 <= 486'h0;
        src4 <= 486'h0;
        src5 <= 486'h0;
        src6 <= 486'h0;
        src7 <= 486'h0;
        src8 <= 486'h0;
        src9 <= 486'h0;
        src10 <= 486'h0;
        src11 <= 486'h0;
        src12 <= 486'h0;
        src13 <= 486'h0;
        src14 <= 486'h0;
        src15 <= 486'h0;
        src16 <= 486'h0;
        src17 <= 486'h0;
        src18 <= 486'h0;
        src19 <= 486'h0;
        src20 <= 486'h0;
        src21 <= 486'h0;
        src22 <= 486'h0;
        src23 <= 486'h0;
        src24 <= 486'h0;
        src25 <= 486'h0;
        src26 <= 486'h0;
        src27 <= 486'h0;
        src28 <= 486'h0;
        src29 <= 486'h0;
        src30 <= 486'h0;
        src31 <= 486'h0;
        src32 <= 486'h0;
        src33 <= 486'h0;
        src34 <= 486'h0;
        src35 <= 486'h0;
        src36 <= 486'h0;
        src37 <= 486'h0;
        src38 <= 486'h0;
        src39 <= 486'h0;
        src40 <= 486'h0;
        src41 <= 486'h0;
        src42 <= 486'h0;
        src43 <= 486'h0;
        src44 <= 486'h0;
        src45 <= 486'h0;
        src46 <= 486'h0;
        src47 <= 486'h0;
        src48 <= 486'h0;
        src49 <= 486'h0;
        src50 <= 486'h0;
        src51 <= 486'h0;
        src52 <= 486'h0;
        src53 <= 486'h0;
        src54 <= 486'h0;
        src55 <= 486'h0;
        src56 <= 486'h0;
        src57 <= 486'h0;
        src58 <= 486'h0;
        src59 <= 486'h0;
        src60 <= 486'h0;
        src61 <= 486'h0;
        src62 <= 486'h0;
        src63 <= 486'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
        src32 <= {src32, src32_};
        src33 <= {src33, src33_};
        src34 <= {src34, src34_};
        src35 <= {src35, src35_};
        src36 <= {src36, src36_};
        src37 <= {src37, src37_};
        src38 <= {src38, src38_};
        src39 <= {src39, src39_};
        src40 <= {src40, src40_};
        src41 <= {src41, src41_};
        src42 <= {src42, src42_};
        src43 <= {src43, src43_};
        src44 <= {src44, src44_};
        src45 <= {src45, src45_};
        src46 <= {src46, src46_};
        src47 <= {src47, src47_};
        src48 <= {src48, src48_};
        src49 <= {src49, src49_};
        src50 <= {src50, src50_};
        src51 <= {src51, src51_};
        src52 <= {src52, src52_};
        src53 <= {src53, src53_};
        src54 <= {src54, src54_};
        src55 <= {src55, src55_};
        src56 <= {src56, src56_};
        src57 <= {src57, src57_};
        src58 <= {src58, src58_};
        src59 <= {src59, src59_};
        src60 <= {src60, src60_};
        src61 <= {src61, src61_};
        src62 <= {src62, src62_};
        src63 <= {src63, src63_};
    end
endmodule
module compressor_CLA486_64(
    input [485:0]src0,
    input [485:0]src1,
    input [485:0]src2,
    input [485:0]src3,
    input [485:0]src4,
    input [485:0]src5,
    input [485:0]src6,
    input [485:0]src7,
    input [485:0]src8,
    input [485:0]src9,
    input [485:0]src10,
    input [485:0]src11,
    input [485:0]src12,
    input [485:0]src13,
    input [485:0]src14,
    input [485:0]src15,
    input [485:0]src16,
    input [485:0]src17,
    input [485:0]src18,
    input [485:0]src19,
    input [485:0]src20,
    input [485:0]src21,
    input [485:0]src22,
    input [485:0]src23,
    input [485:0]src24,
    input [485:0]src25,
    input [485:0]src26,
    input [485:0]src27,
    input [485:0]src28,
    input [485:0]src29,
    input [485:0]src30,
    input [485:0]src31,
    input [485:0]src32,
    input [485:0]src33,
    input [485:0]src34,
    input [485:0]src35,
    input [485:0]src36,
    input [485:0]src37,
    input [485:0]src38,
    input [485:0]src39,
    input [485:0]src40,
    input [485:0]src41,
    input [485:0]src42,
    input [485:0]src43,
    input [485:0]src44,
    input [485:0]src45,
    input [485:0]src46,
    input [485:0]src47,
    input [485:0]src48,
    input [485:0]src49,
    input [485:0]src50,
    input [485:0]src51,
    input [485:0]src52,
    input [485:0]src53,
    input [485:0]src54,
    input [485:0]src55,
    input [485:0]src56,
    input [485:0]src57,
    input [485:0]src58,
    input [485:0]src59,
    input [485:0]src60,
    input [485:0]src61,
    input [485:0]src62,
    input [485:0]src63,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39,
    output dst40,
    output dst41,
    output dst42,
    output dst43,
    output dst44,
    output dst45,
    output dst46,
    output dst47,
    output dst48,
    output dst49,
    output dst50,
    output dst51,
    output dst52,
    output dst53,
    output dst54,
    output dst55,
    output dst56,
    output dst57,
    output dst58,
    output dst59,
    output dst60,
    output dst61,
    output dst62,
    output dst63,
    output dst64,
    output dst65,
    output dst66,
    output dst67,
    output dst68,
    output dst69,
    output dst70,
    output dst71,
    output dst72);

    wire [0:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [0:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    wire [1:0] comp_out39;
    wire [1:0] comp_out40;
    wire [1:0] comp_out41;
    wire [1:0] comp_out42;
    wire [1:0] comp_out43;
    wire [1:0] comp_out44;
    wire [1:0] comp_out45;
    wire [0:0] comp_out46;
    wire [1:0] comp_out47;
    wire [1:0] comp_out48;
    wire [1:0] comp_out49;
    wire [1:0] comp_out50;
    wire [1:0] comp_out51;
    wire [1:0] comp_out52;
    wire [1:0] comp_out53;
    wire [1:0] comp_out54;
    wire [1:0] comp_out55;
    wire [1:0] comp_out56;
    wire [1:0] comp_out57;
    wire [1:0] comp_out58;
    wire [1:0] comp_out59;
    wire [1:0] comp_out60;
    wire [1:0] comp_out61;
    wire [1:0] comp_out62;
    wire [1:0] comp_out63;
    wire [1:0] comp_out64;
    wire [1:0] comp_out65;
    wire [1:0] comp_out66;
    wire [1:0] comp_out67;
    wire [1:0] comp_out68;
    wire [1:0] comp_out69;
    wire [1:0] comp_out70;
    wire [1:0] comp_out71;
    wire [1:0] comp_out72;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39),
        .dst40(comp_out40),
        .dst41(comp_out41),
        .dst42(comp_out42),
        .dst43(comp_out43),
        .dst44(comp_out44),
        .dst45(comp_out45),
        .dst46(comp_out46),
        .dst47(comp_out47),
        .dst48(comp_out48),
        .dst49(comp_out49),
        .dst50(comp_out50),
        .dst51(comp_out51),
        .dst52(comp_out52),
        .dst53(comp_out53),
        .dst54(comp_out54),
        .dst55(comp_out55),
        .dst56(comp_out56),
        .dst57(comp_out57),
        .dst58(comp_out58),
        .dst59(comp_out59),
        .dst60(comp_out60),
        .dst61(comp_out61),
        .dst62(comp_out62),
        .dst63(comp_out63),
        .dst64(comp_out64),
        .dst65(comp_out65),
        .dst66(comp_out66),
        .dst67(comp_out67),
        .dst68(comp_out68),
        .dst69(comp_out69),
        .dst70(comp_out70),
        .dst71(comp_out71),
        .dst72(comp_out72)
    );
    LookAheadCarryUnit256 LCU256(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out72[0], comp_out71[0], comp_out70[0], comp_out69[0], comp_out68[0], comp_out67[0], comp_out66[0], comp_out65[0], comp_out64[0], comp_out63[0], comp_out62[0], comp_out61[0], comp_out60[0], comp_out59[0], comp_out58[0], comp_out57[0], comp_out56[0], comp_out55[0], comp_out54[0], comp_out53[0], comp_out52[0], comp_out51[0], comp_out50[0], comp_out49[0], comp_out48[0], comp_out47[0], comp_out46[0], comp_out45[0], comp_out44[0], comp_out43[0], comp_out42[0], comp_out41[0], comp_out40[0], comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out72[1], comp_out71[1], comp_out70[1], comp_out69[1], comp_out68[1], comp_out67[1], comp_out66[1], comp_out65[1], comp_out64[1], comp_out63[1], comp_out62[1], comp_out61[1], comp_out60[1], comp_out59[1], comp_out58[1], comp_out57[1], comp_out56[1], comp_out55[1], comp_out54[1], comp_out53[1], comp_out52[1], comp_out51[1], comp_out50[1], comp_out49[1], comp_out48[1], comp_out47[1], 1'h0, comp_out45[1], comp_out44[1], comp_out43[1], comp_out42[1], comp_out41[1], comp_out40[1], comp_out39[1], comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], 1'h0, comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], 1'h0}),
        .dst({dst72, dst71, dst70, dst69, dst68, dst67, dst66, dst65, dst64, dst63, dst62, dst61, dst60, dst59, dst58, dst57, dst56, dst55, dst54, dst53, dst52, dst51, dst50, dst49, dst48, dst47, dst46, dst45, dst44, dst43, dst42, dst41, dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [485:0] src0,
      input wire [485:0] src1,
      input wire [485:0] src2,
      input wire [485:0] src3,
      input wire [485:0] src4,
      input wire [485:0] src5,
      input wire [485:0] src6,
      input wire [485:0] src7,
      input wire [485:0] src8,
      input wire [485:0] src9,
      input wire [485:0] src10,
      input wire [485:0] src11,
      input wire [485:0] src12,
      input wire [485:0] src13,
      input wire [485:0] src14,
      input wire [485:0] src15,
      input wire [485:0] src16,
      input wire [485:0] src17,
      input wire [485:0] src18,
      input wire [485:0] src19,
      input wire [485:0] src20,
      input wire [485:0] src21,
      input wire [485:0] src22,
      input wire [485:0] src23,
      input wire [485:0] src24,
      input wire [485:0] src25,
      input wire [485:0] src26,
      input wire [485:0] src27,
      input wire [485:0] src28,
      input wire [485:0] src29,
      input wire [485:0] src30,
      input wire [485:0] src31,
      input wire [485:0] src32,
      input wire [485:0] src33,
      input wire [485:0] src34,
      input wire [485:0] src35,
      input wire [485:0] src36,
      input wire [485:0] src37,
      input wire [485:0] src38,
      input wire [485:0] src39,
      input wire [485:0] src40,
      input wire [485:0] src41,
      input wire [485:0] src42,
      input wire [485:0] src43,
      input wire [485:0] src44,
      input wire [485:0] src45,
      input wire [485:0] src46,
      input wire [485:0] src47,
      input wire [485:0] src48,
      input wire [485:0] src49,
      input wire [485:0] src50,
      input wire [485:0] src51,
      input wire [485:0] src52,
      input wire [485:0] src53,
      input wire [485:0] src54,
      input wire [485:0] src55,
      input wire [485:0] src56,
      input wire [485:0] src57,
      input wire [485:0] src58,
      input wire [485:0] src59,
      input wire [485:0] src60,
      input wire [485:0] src61,
      input wire [485:0] src62,
      input wire [485:0] src63,
      output wire [0:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [0:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38,
      output wire [1:0] dst39,
      output wire [1:0] dst40,
      output wire [1:0] dst41,
      output wire [1:0] dst42,
      output wire [1:0] dst43,
      output wire [1:0] dst44,
      output wire [1:0] dst45,
      output wire [0:0] dst46,
      output wire [1:0] dst47,
      output wire [1:0] dst48,
      output wire [1:0] dst49,
      output wire [1:0] dst50,
      output wire [1:0] dst51,
      output wire [1:0] dst52,
      output wire [1:0] dst53,
      output wire [1:0] dst54,
      output wire [1:0] dst55,
      output wire [1:0] dst56,
      output wire [1:0] dst57,
      output wire [1:0] dst58,
      output wire [1:0] dst59,
      output wire [1:0] dst60,
      output wire [1:0] dst61,
      output wire [1:0] dst62,
      output wire [1:0] dst63,
      output wire [1:0] dst64,
      output wire [1:0] dst65,
      output wire [1:0] dst66,
      output wire [1:0] dst67,
      output wire [1:0] dst68,
      output wire [1:0] dst69,
      output wire [1:0] dst70,
      output wire [1:0] dst71,
      output wire [1:0] dst72);

   wire [485:0] stage0_0;
   wire [485:0] stage0_1;
   wire [485:0] stage0_2;
   wire [485:0] stage0_3;
   wire [485:0] stage0_4;
   wire [485:0] stage0_5;
   wire [485:0] stage0_6;
   wire [485:0] stage0_7;
   wire [485:0] stage0_8;
   wire [485:0] stage0_9;
   wire [485:0] stage0_10;
   wire [485:0] stage0_11;
   wire [485:0] stage0_12;
   wire [485:0] stage0_13;
   wire [485:0] stage0_14;
   wire [485:0] stage0_15;
   wire [485:0] stage0_16;
   wire [485:0] stage0_17;
   wire [485:0] stage0_18;
   wire [485:0] stage0_19;
   wire [485:0] stage0_20;
   wire [485:0] stage0_21;
   wire [485:0] stage0_22;
   wire [485:0] stage0_23;
   wire [485:0] stage0_24;
   wire [485:0] stage0_25;
   wire [485:0] stage0_26;
   wire [485:0] stage0_27;
   wire [485:0] stage0_28;
   wire [485:0] stage0_29;
   wire [485:0] stage0_30;
   wire [485:0] stage0_31;
   wire [485:0] stage0_32;
   wire [485:0] stage0_33;
   wire [485:0] stage0_34;
   wire [485:0] stage0_35;
   wire [485:0] stage0_36;
   wire [485:0] stage0_37;
   wire [485:0] stage0_38;
   wire [485:0] stage0_39;
   wire [485:0] stage0_40;
   wire [485:0] stage0_41;
   wire [485:0] stage0_42;
   wire [485:0] stage0_43;
   wire [485:0] stage0_44;
   wire [485:0] stage0_45;
   wire [485:0] stage0_46;
   wire [485:0] stage0_47;
   wire [485:0] stage0_48;
   wire [485:0] stage0_49;
   wire [485:0] stage0_50;
   wire [485:0] stage0_51;
   wire [485:0] stage0_52;
   wire [485:0] stage0_53;
   wire [485:0] stage0_54;
   wire [485:0] stage0_55;
   wire [485:0] stage0_56;
   wire [485:0] stage0_57;
   wire [485:0] stage0_58;
   wire [485:0] stage0_59;
   wire [485:0] stage0_60;
   wire [485:0] stage0_61;
   wire [485:0] stage0_62;
   wire [485:0] stage0_63;
   wire [124:0] stage1_0;
   wire [175:0] stage1_1;
   wire [157:0] stage1_2;
   wire [214:0] stage1_3;
   wire [227:0] stage1_4;
   wire [197:0] stage1_5;
   wire [213:0] stage1_6;
   wire [220:0] stage1_7;
   wire [205:0] stage1_8;
   wire [213:0] stage1_9;
   wire [284:0] stage1_10;
   wire [276:0] stage1_11;
   wire [188:0] stage1_12;
   wire [304:0] stage1_13;
   wire [218:0] stage1_14;
   wire [170:0] stage1_15;
   wire [221:0] stage1_16;
   wire [228:0] stage1_17;
   wire [208:0] stage1_18;
   wire [275:0] stage1_19;
   wire [267:0] stage1_20;
   wire [189:0] stage1_21;
   wire [170:0] stage1_22;
   wire [286:0] stage1_23;
   wire [213:0] stage1_24;
   wire [183:0] stage1_25;
   wire [250:0] stage1_26;
   wire [205:0] stage1_27;
   wire [223:0] stage1_28;
   wire [228:0] stage1_29;
   wire [191:0] stage1_30;
   wire [217:0] stage1_31;
   wire [216:0] stage1_32;
   wire [258:0] stage1_33;
   wire [189:0] stage1_34;
   wire [216:0] stage1_35;
   wire [201:0] stage1_36;
   wire [307:0] stage1_37;
   wire [264:0] stage1_38;
   wire [212:0] stage1_39;
   wire [303:0] stage1_40;
   wire [170:0] stage1_41;
   wire [173:0] stage1_42;
   wire [253:0] stage1_43;
   wire [255:0] stage1_44;
   wire [211:0] stage1_45;
   wire [297:0] stage1_46;
   wire [235:0] stage1_47;
   wire [197:0] stage1_48;
   wire [172:0] stage1_49;
   wire [189:0] stage1_50;
   wire [274:0] stage1_51;
   wire [198:0] stage1_52;
   wire [168:0] stage1_53;
   wire [230:0] stage1_54;
   wire [266:0] stage1_55;
   wire [186:0] stage1_56;
   wire [188:0] stage1_57;
   wire [219:0] stage1_58;
   wire [205:0] stage1_59;
   wire [214:0] stage1_60;
   wire [218:0] stage1_61;
   wire [192:0] stage1_62;
   wire [307:0] stage1_63;
   wire [123:0] stage1_64;
   wire [53:0] stage1_65;
   wire [37:0] stage2_0;
   wire [53:0] stage2_1;
   wire [62:0] stage2_2;
   wire [113:0] stage2_3;
   wire [111:0] stage2_4;
   wire [151:0] stage2_5;
   wire [91:0] stage2_6;
   wire [72:0] stage2_7;
   wire [159:0] stage2_8;
   wire [142:0] stage2_9;
   wire [163:0] stage2_10;
   wire [138:0] stage2_11;
   wire [106:0] stage2_12;
   wire [77:0] stage2_13;
   wire [107:0] stage2_14;
   wire [140:0] stage2_15;
   wire [82:0] stage2_16;
   wire [86:0] stage2_17;
   wire [118:0] stage2_18;
   wire [112:0] stage2_19;
   wire [92:0] stage2_20;
   wire [127:0] stage2_21;
   wire [107:0] stage2_22;
   wire [75:0] stage2_23;
   wire [101:0] stage2_24;
   wire [95:0] stage2_25;
   wire [84:0] stage2_26;
   wire [105:0] stage2_27;
   wire [91:0] stage2_28;
   wire [86:0] stage2_29;
   wire [116:0] stage2_30;
   wire [98:0] stage2_31;
   wire [105:0] stage2_32;
   wire [75:0] stage2_33;
   wire [131:0] stage2_34;
   wire [132:0] stage2_35;
   wire [74:0] stage2_36;
   wire [89:0] stage2_37;
   wire [139:0] stage2_38;
   wire [136:0] stage2_39;
   wire [112:0] stage2_40;
   wire [105:0] stage2_41;
   wire [85:0] stage2_42;
   wire [78:0] stage2_43;
   wire [118:0] stage2_44;
   wire [117:0] stage2_45;
   wire [87:0] stage2_46;
   wire [103:0] stage2_47;
   wire [129:0] stage2_48;
   wire [95:0] stage2_49;
   wire [85:0] stage2_50;
   wire [87:0] stage2_51;
   wire [104:0] stage2_52;
   wire [114:0] stage2_53;
   wire [99:0] stage2_54;
   wire [105:0] stage2_55;
   wire [114:0] stage2_56;
   wire [65:0] stage2_57;
   wire [85:0] stage2_58;
   wire [109:0] stage2_59;
   wire [84:0] stage2_60;
   wire [74:0] stage2_61;
   wire [104:0] stage2_62;
   wire [98:0] stage2_63;
   wire [141:0] stage2_64;
   wire [55:0] stage2_65;
   wire [41:0] stage2_66;
   wire [20:0] stage3_0;
   wire [21:0] stage3_1;
   wire [42:0] stage3_2;
   wire [28:0] stage3_3;
   wire [111:0] stage3_4;
   wire [52:0] stage3_5;
   wire [77:0] stage3_6;
   wire [50:0] stage3_7;
   wire [34:0] stage3_8;
   wire [53:0] stage3_9;
   wire [99:0] stage3_10;
   wire [57:0] stage3_11;
   wire [67:0] stage3_12;
   wire [56:0] stage3_13;
   wire [31:0] stage3_14;
   wire [47:0] stage3_15;
   wire [50:0] stage3_16;
   wire [35:0] stage3_17;
   wire [59:0] stage3_18;
   wire [47:0] stage3_19;
   wire [82:0] stage3_20;
   wire [38:0] stage3_21;
   wire [72:0] stage3_22;
   wire [42:0] stage3_23;
   wire [28:0] stage3_24;
   wire [32:0] stage3_25;
   wire [48:0] stage3_26;
   wire [48:0] stage3_27;
   wire [56:0] stage3_28;
   wire [47:0] stage3_29;
   wire [41:0] stage3_30;
   wire [37:0] stage3_31;
   wire [53:0] stage3_32;
   wire [45:0] stage3_33;
   wire [41:0] stage3_34;
   wire [56:0] stage3_35;
   wire [45:0] stage3_36;
   wire [52:0] stage3_37;
   wire [59:0] stage3_38;
   wire [57:0] stage3_39;
   wire [51:0] stage3_40;
   wire [42:0] stage3_41;
   wire [49:0] stage3_42;
   wire [45:0] stage3_43;
   wire [40:0] stage3_44;
   wire [43:0] stage3_45;
   wire [57:0] stage3_46;
   wire [43:0] stage3_47;
   wire [41:0] stage3_48;
   wire [41:0] stage3_49;
   wire [46:0] stage3_50;
   wire [62:0] stage3_51;
   wire [62:0] stage3_52;
   wire [74:0] stage3_53;
   wire [38:0] stage3_54;
   wire [66:0] stage3_55;
   wire [31:0] stage3_56;
   wire [53:0] stage3_57;
   wire [61:0] stage3_58;
   wire [49:0] stage3_59;
   wire [41:0] stage3_60;
   wire [52:0] stage3_61;
   wire [33:0] stage3_62;
   wire [47:0] stage3_63;
   wire [50:0] stage3_64;
   wire [37:0] stage3_65;
   wire [37:0] stage3_66;
   wire [13:0] stage3_67;
   wire [5:0] stage3_68;
   wire [8:0] stage4_0;
   wire [6:0] stage4_1;
   wire [10:0] stage4_2;
   wire [16:0] stage4_3;
   wire [30:0] stage4_4;
   wire [35:0] stage4_5;
   wire [23:0] stage4_6;
   wire [38:0] stage4_7;
   wire [27:0] stage4_8;
   wire [13:0] stage4_9;
   wire [41:0] stage4_10;
   wire [28:0] stage4_11;
   wire [23:0] stage4_12;
   wire [31:0] stage4_13;
   wire [29:0] stage4_14;
   wire [14:0] stage4_15;
   wire [26:0] stage4_16;
   wire [17:0] stage4_17;
   wire [20:0] stage4_18;
   wire [28:0] stage4_19;
   wire [33:0] stage4_20;
   wire [36:0] stage4_21;
   wire [17:0] stage4_22;
   wire [20:0] stage4_23;
   wire [21:0] stage4_24;
   wire [20:0] stage4_25;
   wire [18:0] stage4_26;
   wire [26:0] stage4_27;
   wire [18:0] stage4_28;
   wire [21:0] stage4_29;
   wire [32:0] stage4_30;
   wire [14:0] stage4_31;
   wire [29:0] stage4_32;
   wire [28:0] stage4_33;
   wire [18:0] stage4_34;
   wire [35:0] stage4_35;
   wire [35:0] stage4_36;
   wire [17:0] stage4_37;
   wire [19:0] stage4_38;
   wire [23:0] stage4_39;
   wire [27:0] stage4_40;
   wire [19:0] stage4_41;
   wire [37:0] stage4_42;
   wire [13:0] stage4_43;
   wire [24:0] stage4_44;
   wire [28:0] stage4_45;
   wire [16:0] stage4_46;
   wire [20:0] stage4_47;
   wire [22:0] stage4_48;
   wire [12:0] stage4_49;
   wire [21:0] stage4_50;
   wire [35:0] stage4_51;
   wire [18:0] stage4_52;
   wire [43:0] stage4_53;
   wire [25:0] stage4_54;
   wire [38:0] stage4_55;
   wire [13:0] stage4_56;
   wire [25:0] stage4_57;
   wire [23:0] stage4_58;
   wire [20:0] stage4_59;
   wire [21:0] stage4_60;
   wire [31:0] stage4_61;
   wire [16:0] stage4_62;
   wire [13:0] stage4_63;
   wire [33:0] stage4_64;
   wire [35:0] stage4_65;
   wire [10:0] stage4_66;
   wire [10:0] stage4_67;
   wire [13:0] stage4_68;
   wire [1:0] stage4_69;
   wire [4:0] stage5_0;
   wire [1:0] stage5_1;
   wire [4:0] stage5_2;
   wire [7:0] stage5_3;
   wire [10:0] stage5_4;
   wire [15:0] stage5_5;
   wire [9:0] stage5_6;
   wire [10:0] stage5_7;
   wire [18:0] stage5_8;
   wire [10:0] stage5_9;
   wire [20:0] stage5_10;
   wire [13:0] stage5_11;
   wire [10:0] stage5_12;
   wire [14:0] stage5_13;
   wire [15:0] stage5_14;
   wire [11:0] stage5_15;
   wire [7:0] stage5_16;
   wire [6:0] stage5_17;
   wire [11:0] stage5_18;
   wire [15:0] stage5_19;
   wire [13:0] stage5_20;
   wire [10:0] stage5_21;
   wire [13:0] stage5_22;
   wire [9:0] stage5_23;
   wire [8:0] stage5_24;
   wire [9:0] stage5_25;
   wire [14:0] stage5_26;
   wire [5:0] stage5_27;
   wire [9:0] stage5_28;
   wire [14:0] stage5_29;
   wire [8:0] stage5_30;
   wire [9:0] stage5_31;
   wire [19:0] stage5_32;
   wire [11:0] stage5_33;
   wire [13:0] stage5_34;
   wire [13:0] stage5_35;
   wire [12:0] stage5_36;
   wire [10:0] stage5_37;
   wire [9:0] stage5_38;
   wire [9:0] stage5_39;
   wire [10:0] stage5_40;
   wire [8:0] stage5_41;
   wire [18:0] stage5_42;
   wire [10:0] stage5_43;
   wire [12:0] stage5_44;
   wire [14:0] stage5_45;
   wire [11:0] stage5_46;
   wire [11:0] stage5_47;
   wire [13:0] stage5_48;
   wire [5:0] stage5_49;
   wire [11:0] stage5_50;
   wire [18:0] stage5_51;
   wire [9:0] stage5_52;
   wire [12:0] stage5_53;
   wire [16:0] stage5_54;
   wire [21:0] stage5_55;
   wire [8:0] stage5_56;
   wire [13:0] stage5_57;
   wire [15:0] stage5_58;
   wire [7:0] stage5_59;
   wire [14:0] stage5_60;
   wire [15:0] stage5_61;
   wire [11:0] stage5_62;
   wire [8:0] stage5_63;
   wire [14:0] stage5_64;
   wire [17:0] stage5_65;
   wire [7:0] stage5_66;
   wire [10:0] stage5_67;
   wire [13:0] stage5_68;
   wire [2:0] stage5_69;
   wire [0:0] stage5_70;
   wire [4:0] stage6_0;
   wire [1:0] stage6_1;
   wire [4:0] stage6_2;
   wire [1:0] stage6_3;
   wire [5:0] stage6_4;
   wire [3:0] stage6_5;
   wire [7:0] stage6_6;
   wire [4:0] stage6_7;
   wire [5:0] stage6_8;
   wire [9:0] stage6_9;
   wire [4:0] stage6_10;
   wire [6:0] stage6_11;
   wire [6:0] stage6_12;
   wire [9:0] stage6_13;
   wire [6:0] stage6_14;
   wire [5:0] stage6_15;
   wire [4:0] stage6_16;
   wire [4:0] stage6_17;
   wire [5:0] stage6_18;
   wire [4:0] stage6_19;
   wire [5:0] stage6_20;
   wire [5:0] stage6_21;
   wire [5:0] stage6_22;
   wire [6:0] stage6_23;
   wire [6:0] stage6_24;
   wire [2:0] stage6_25;
   wire [7:0] stage6_26;
   wire [4:0] stage6_27;
   wire [5:0] stage6_28;
   wire [5:0] stage6_29;
   wire [4:0] stage6_30;
   wire [5:0] stage6_31;
   wire [5:0] stage6_32;
   wire [5:0] stage6_33;
   wire [8:0] stage6_34;
   wire [4:0] stage6_35;
   wire [5:0] stage6_36;
   wire [5:0] stage6_37;
   wire [4:0] stage6_38;
   wire [3:0] stage6_39;
   wire [5:0] stage6_40;
   wire [7:0] stage6_41;
   wire [6:0] stage6_42;
   wire [6:0] stage6_43;
   wire [4:0] stage6_44;
   wire [8:0] stage6_45;
   wire [4:0] stage6_46;
   wire [6:0] stage6_47;
   wire [4:0] stage6_48;
   wire [5:0] stage6_49;
   wire [2:0] stage6_50;
   wire [7:0] stage6_51;
   wire [6:0] stage6_52;
   wire [4:0] stage6_53;
   wire [5:0] stage6_54;
   wire [9:0] stage6_55;
   wire [9:0] stage6_56;
   wire [6:0] stage6_57;
   wire [5:0] stage6_58;
   wire [4:0] stage6_59;
   wire [4:0] stage6_60;
   wire [8:0] stage6_61;
   wire [5:0] stage6_62;
   wire [4:0] stage6_63;
   wire [8:0] stage6_64;
   wire [4:0] stage6_65;
   wire [4:0] stage6_66;
   wire [4:0] stage6_67;
   wire [16:0] stage6_68;
   wire [4:0] stage6_69;
   wire [0:0] stage6_70;
   wire [4:0] stage7_0;
   wire [1:0] stage7_1;
   wire [4:0] stage7_2;
   wire [1:0] stage7_3;
   wire [0:0] stage7_4;
   wire [1:0] stage7_5;
   wire [2:0] stage7_6;
   wire [2:0] stage7_7;
   wire [4:0] stage7_8;
   wire [5:0] stage7_9;
   wire [1:0] stage7_10;
   wire [3:0] stage7_11;
   wire [1:0] stage7_12;
   wire [5:0] stage7_13;
   wire [2:0] stage7_14;
   wire [5:0] stage7_15;
   wire [2:0] stage7_16;
   wire [1:0] stage7_17;
   wire [1:0] stage7_18;
   wire [6:0] stage7_19;
   wire [2:0] stage7_20;
   wire [5:0] stage7_21;
   wire [6:0] stage7_22;
   wire [0:0] stage7_23;
   wire [3:0] stage7_24;
   wire [1:0] stage7_25;
   wire [5:0] stage7_26;
   wire [4:0] stage7_27;
   wire [0:0] stage7_28;
   wire [4:0] stage7_29;
   wire [6:0] stage7_30;
   wire [1:0] stage7_31;
   wire [5:0] stage7_32;
   wire [0:0] stage7_33;
   wire [5:0] stage7_34;
   wire [5:0] stage7_35;
   wire [0:0] stage7_36;
   wire [1:0] stage7_37;
   wire [6:0] stage7_38;
   wire [0:0] stage7_39;
   wire [6:0] stage7_40;
   wire [4:0] stage7_41;
   wire [2:0] stage7_42;
   wire [3:0] stage7_43;
   wire [1:0] stage7_44;
   wire [4:0] stage7_45;
   wire [2:0] stage7_46;
   wire [7:0] stage7_47;
   wire [0:0] stage7_48;
   wire [1:0] stage7_49;
   wire [2:0] stage7_50;
   wire [3:0] stage7_51;
   wire [3:0] stage7_52;
   wire [5:0] stage7_53;
   wire [0:0] stage7_54;
   wire [6:0] stage7_55;
   wire [6:0] stage7_56;
   wire [1:0] stage7_57;
   wire [1:0] stage7_58;
   wire [6:0] stage7_59;
   wire [5:0] stage7_60;
   wire [1:0] stage7_61;
   wire [1:0] stage7_62;
   wire [2:0] stage7_63;
   wire [3:0] stage7_64;
   wire [2:0] stage7_65;
   wire [5:0] stage7_66;
   wire [0:0] stage7_67;
   wire [4:0] stage7_68;
   wire [4:0] stage7_69;
   wire [2:0] stage7_70;
   wire [1:0] stage7_71;
   wire [0:0] stage8_0;
   wire [1:0] stage8_1;
   wire [1:0] stage8_2;
   wire [1:0] stage8_3;
   wire [1:0] stage8_4;
   wire [1:0] stage8_5;
   wire [0:0] stage8_6;
   wire [1:0] stage8_7;
   wire [1:0] stage8_8;
   wire [1:0] stage8_9;
   wire [1:0] stage8_10;
   wire [1:0] stage8_11;
   wire [1:0] stage8_12;
   wire [1:0] stage8_13;
   wire [1:0] stage8_14;
   wire [1:0] stage8_15;
   wire [1:0] stage8_16;
   wire [1:0] stage8_17;
   wire [1:0] stage8_18;
   wire [1:0] stage8_19;
   wire [1:0] stage8_20;
   wire [1:0] stage8_21;
   wire [1:0] stage8_22;
   wire [1:0] stage8_23;
   wire [1:0] stage8_24;
   wire [1:0] stage8_25;
   wire [1:0] stage8_26;
   wire [1:0] stage8_27;
   wire [1:0] stage8_28;
   wire [1:0] stage8_29;
   wire [1:0] stage8_30;
   wire [1:0] stage8_31;
   wire [1:0] stage8_32;
   wire [1:0] stage8_33;
   wire [1:0] stage8_34;
   wire [1:0] stage8_35;
   wire [1:0] stage8_36;
   wire [1:0] stage8_37;
   wire [1:0] stage8_38;
   wire [1:0] stage8_39;
   wire [1:0] stage8_40;
   wire [1:0] stage8_41;
   wire [1:0] stage8_42;
   wire [1:0] stage8_43;
   wire [1:0] stage8_44;
   wire [1:0] stage8_45;
   wire [0:0] stage8_46;
   wire [1:0] stage8_47;
   wire [1:0] stage8_48;
   wire [1:0] stage8_49;
   wire [1:0] stage8_50;
   wire [1:0] stage8_51;
   wire [1:0] stage8_52;
   wire [1:0] stage8_53;
   wire [1:0] stage8_54;
   wire [1:0] stage8_55;
   wire [1:0] stage8_56;
   wire [1:0] stage8_57;
   wire [1:0] stage8_58;
   wire [1:0] stage8_59;
   wire [1:0] stage8_60;
   wire [1:0] stage8_61;
   wire [1:0] stage8_62;
   wire [1:0] stage8_63;
   wire [1:0] stage8_64;
   wire [1:0] stage8_65;
   wire [1:0] stage8_66;
   wire [1:0] stage8_67;
   wire [1:0] stage8_68;
   wire [1:0] stage8_69;
   wire [1:0] stage8_70;
   wire [1:0] stage8_71;
   wire [1:0] stage8_72;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign stage0_32 = src32;
   assign stage0_33 = src33;
   assign stage0_34 = src34;
   assign stage0_35 = src35;
   assign stage0_36 = src36;
   assign stage0_37 = src37;
   assign stage0_38 = src38;
   assign stage0_39 = src39;
   assign stage0_40 = src40;
   assign stage0_41 = src41;
   assign stage0_42 = src42;
   assign stage0_43 = src43;
   assign stage0_44 = src44;
   assign stage0_45 = src45;
   assign stage0_46 = src46;
   assign stage0_47 = src47;
   assign stage0_48 = src48;
   assign stage0_49 = src49;
   assign stage0_50 = src50;
   assign stage0_51 = src51;
   assign stage0_52 = src52;
   assign stage0_53 = src53;
   assign stage0_54 = src54;
   assign stage0_55 = src55;
   assign stage0_56 = src56;
   assign stage0_57 = src57;
   assign stage0_58 = src58;
   assign stage0_59 = src59;
   assign stage0_60 = src60;
   assign stage0_61 = src61;
   assign stage0_62 = src62;
   assign stage0_63 = src63;
   assign dst0 = stage8_0;
   assign dst1 = stage8_1;
   assign dst2 = stage8_2;
   assign dst3 = stage8_3;
   assign dst4 = stage8_4;
   assign dst5 = stage8_5;
   assign dst6 = stage8_6;
   assign dst7 = stage8_7;
   assign dst8 = stage8_8;
   assign dst9 = stage8_9;
   assign dst10 = stage8_10;
   assign dst11 = stage8_11;
   assign dst12 = stage8_12;
   assign dst13 = stage8_13;
   assign dst14 = stage8_14;
   assign dst15 = stage8_15;
   assign dst16 = stage8_16;
   assign dst17 = stage8_17;
   assign dst18 = stage8_18;
   assign dst19 = stage8_19;
   assign dst20 = stage8_20;
   assign dst21 = stage8_21;
   assign dst22 = stage8_22;
   assign dst23 = stage8_23;
   assign dst24 = stage8_24;
   assign dst25 = stage8_25;
   assign dst26 = stage8_26;
   assign dst27 = stage8_27;
   assign dst28 = stage8_28;
   assign dst29 = stage8_29;
   assign dst30 = stage8_30;
   assign dst31 = stage8_31;
   assign dst32 = stage8_32;
   assign dst33 = stage8_33;
   assign dst34 = stage8_34;
   assign dst35 = stage8_35;
   assign dst36 = stage8_36;
   assign dst37 = stage8_37;
   assign dst38 = stage8_38;
   assign dst39 = stage8_39;
   assign dst40 = stage8_40;
   assign dst41 = stage8_41;
   assign dst42 = stage8_42;
   assign dst43 = stage8_43;
   assign dst44 = stage8_44;
   assign dst45 = stage8_45;
   assign dst46 = stage8_46;
   assign dst47 = stage8_47;
   assign dst48 = stage8_48;
   assign dst49 = stage8_49;
   assign dst50 = stage8_50;
   assign dst51 = stage8_51;
   assign dst52 = stage8_52;
   assign dst53 = stage8_53;
   assign dst54 = stage8_54;
   assign dst55 = stage8_55;
   assign dst56 = stage8_56;
   assign dst57 = stage8_57;
   assign dst58 = stage8_58;
   assign dst59 = stage8_59;
   assign dst60 = stage8_60;
   assign dst61 = stage8_61;
   assign dst62 = stage8_62;
   assign dst63 = stage8_63;
   assign dst64 = stage8_64;
   assign dst65 = stage8_65;
   assign dst66 = stage8_66;
   assign dst67 = stage8_67;
   assign dst68 = stage8_68;
   assign dst69 = stage8_69;
   assign dst70 = stage8_70;
   assign dst71 = stage8_71;
   assign dst72 = stage8_72;

   gpc117_4 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5], stage0_0[6]},
      {stage0_1[0]},
      {stage0_2[0]},
      {stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc117_4 gpc1 (
      {stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13]},
      {stage0_1[1]},
      {stage0_2[1]},
      {stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc117_4 gpc2 (
      {stage0_0[14], stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_1[2]},
      {stage0_2[2]},
      {stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc117_4 gpc3 (
      {stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27]},
      {stage0_1[3]},
      {stage0_2[3]},
      {stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc117_4 gpc4 (
      {stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[4]},
      {stage0_2[4]},
      {stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc117_4 gpc5 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41]},
      {stage0_1[5]},
      {stage0_2[5]},
      {stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc117_4 gpc6 (
      {stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48]},
      {stage0_1[6]},
      {stage0_2[6]},
      {stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc117_4 gpc7 (
      {stage0_0[49], stage0_0[50], stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54], stage0_0[55]},
      {stage0_1[7]},
      {stage0_2[7]},
      {stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc117_4 gpc8 (
      {stage0_0[56], stage0_0[57], stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_1[8]},
      {stage0_2[8]},
      {stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc117_4 gpc9 (
      {stage0_0[63], stage0_0[64], stage0_0[65], stage0_0[66], stage0_0[67], stage0_0[68], stage0_0[69]},
      {stage0_1[9]},
      {stage0_2[9]},
      {stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc117_4 gpc10 (
      {stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74], stage0_0[75], stage0_0[76]},
      {stage0_1[10]},
      {stage0_2[10]},
      {stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc117_4 gpc11 (
      {stage0_0[77], stage0_0[78], stage0_0[79], stage0_0[80], stage0_0[81], stage0_0[82], stage0_0[83]},
      {stage0_1[11]},
      {stage0_2[11]},
      {stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc117_4 gpc12 (
      {stage0_0[84], stage0_0[85], stage0_0[86], stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90]},
      {stage0_1[12]},
      {stage0_2[12]},
      {stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc1163_5 gpc13 (
      {stage0_0[91], stage0_0[92], stage0_0[93]},
      {stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18]},
      {stage0_2[13]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc1163_5 gpc14 (
      {stage0_0[94], stage0_0[95], stage0_0[96]},
      {stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24]},
      {stage0_2[14]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc1163_5 gpc15 (
      {stage0_0[97], stage0_0[98], stage0_0[99]},
      {stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30]},
      {stage0_2[15]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc1163_5 gpc16 (
      {stage0_0[100], stage0_0[101], stage0_0[102]},
      {stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36]},
      {stage0_2[16]},
      {stage0_3[3]},
      {stage1_4[3],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc1163_5 gpc17 (
      {stage0_0[103], stage0_0[104], stage0_0[105]},
      {stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42]},
      {stage0_2[17]},
      {stage0_3[4]},
      {stage1_4[4],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc1163_5 gpc18 (
      {stage0_0[106], stage0_0[107], stage0_0[108]},
      {stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48]},
      {stage0_2[18]},
      {stage0_3[5]},
      {stage1_4[5],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc1163_5 gpc19 (
      {stage0_0[109], stage0_0[110], stage0_0[111]},
      {stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53], stage0_1[54]},
      {stage0_2[19]},
      {stage0_3[6]},
      {stage1_4[6],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc1163_5 gpc20 (
      {stage0_0[112], stage0_0[113], stage0_0[114]},
      {stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59], stage0_1[60]},
      {stage0_2[20]},
      {stage0_3[7]},
      {stage1_4[7],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc1163_5 gpc21 (
      {stage0_0[115], stage0_0[116], stage0_0[117]},
      {stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65], stage0_1[66]},
      {stage0_2[21]},
      {stage0_3[8]},
      {stage1_4[8],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc1163_5 gpc22 (
      {stage0_0[118], stage0_0[119], stage0_0[120]},
      {stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71], stage0_1[72]},
      {stage0_2[22]},
      {stage0_3[9]},
      {stage1_4[9],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc1163_5 gpc23 (
      {stage0_0[121], stage0_0[122], stage0_0[123]},
      {stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77], stage0_1[78]},
      {stage0_2[23]},
      {stage0_3[10]},
      {stage1_4[10],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc1163_5 gpc24 (
      {stage0_0[124], stage0_0[125], stage0_0[126]},
      {stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83], stage0_1[84]},
      {stage0_2[24]},
      {stage0_3[11]},
      {stage1_4[11],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc1163_5 gpc25 (
      {stage0_0[127], stage0_0[128], stage0_0[129]},
      {stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89], stage0_1[90]},
      {stage0_2[25]},
      {stage0_3[12]},
      {stage1_4[12],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc1163_5 gpc26 (
      {stage0_0[130], stage0_0[131], stage0_0[132]},
      {stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95], stage0_1[96]},
      {stage0_2[26]},
      {stage0_3[13]},
      {stage1_4[13],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc1163_5 gpc27 (
      {stage0_0[133], stage0_0[134], stage0_0[135]},
      {stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101], stage0_1[102]},
      {stage0_2[27]},
      {stage0_3[14]},
      {stage1_4[14],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc1163_5 gpc28 (
      {stage0_0[136], stage0_0[137], stage0_0[138]},
      {stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107], stage0_1[108]},
      {stage0_2[28]},
      {stage0_3[15]},
      {stage1_4[15],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc1163_5 gpc29 (
      {stage0_0[139], stage0_0[140], stage0_0[141]},
      {stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113], stage0_1[114]},
      {stage0_2[29]},
      {stage0_3[16]},
      {stage1_4[16],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc1163_5 gpc30 (
      {stage0_0[142], stage0_0[143], stage0_0[144]},
      {stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119], stage0_1[120]},
      {stage0_2[30]},
      {stage0_3[17]},
      {stage1_4[17],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc1163_5 gpc31 (
      {stage0_0[145], stage0_0[146], stage0_0[147]},
      {stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125], stage0_1[126]},
      {stage0_2[31]},
      {stage0_3[18]},
      {stage1_4[18],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc1163_5 gpc32 (
      {stage0_0[148], stage0_0[149], stage0_0[150]},
      {stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131], stage0_1[132]},
      {stage0_2[32]},
      {stage0_3[19]},
      {stage1_4[19],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc1163_5 gpc33 (
      {stage0_0[151], stage0_0[152], stage0_0[153]},
      {stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137], stage0_1[138]},
      {stage0_2[33]},
      {stage0_3[20]},
      {stage1_4[20],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc1163_5 gpc34 (
      {stage0_0[154], stage0_0[155], stage0_0[156]},
      {stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143], stage0_1[144]},
      {stage0_2[34]},
      {stage0_3[21]},
      {stage1_4[21],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc1163_5 gpc35 (
      {stage0_0[157], stage0_0[158], stage0_0[159]},
      {stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149], stage0_1[150]},
      {stage0_2[35]},
      {stage0_3[22]},
      {stage1_4[22],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc1163_5 gpc36 (
      {stage0_0[160], stage0_0[161], stage0_0[162]},
      {stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155], stage0_1[156]},
      {stage0_2[36]},
      {stage0_3[23]},
      {stage1_4[23],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc1163_5 gpc37 (
      {stage0_0[163], stage0_0[164], stage0_0[165]},
      {stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161], stage0_1[162]},
      {stage0_2[37]},
      {stage0_3[24]},
      {stage1_4[24],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc1163_5 gpc38 (
      {stage0_0[166], stage0_0[167], stage0_0[168]},
      {stage0_1[163], stage0_1[164], stage0_1[165], stage0_1[166], stage0_1[167], stage0_1[168]},
      {stage0_2[38]},
      {stage0_3[25]},
      {stage1_4[25],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc1163_5 gpc39 (
      {stage0_0[169], stage0_0[170], stage0_0[171]},
      {stage0_1[169], stage0_1[170], stage0_1[171], stage0_1[172], stage0_1[173], stage0_1[174]},
      {stage0_2[39]},
      {stage0_3[26]},
      {stage1_4[26],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc1163_5 gpc40 (
      {stage0_0[172], stage0_0[173], stage0_0[174]},
      {stage0_1[175], stage0_1[176], stage0_1[177], stage0_1[178], stage0_1[179], stage0_1[180]},
      {stage0_2[40]},
      {stage0_3[27]},
      {stage1_4[27],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc1163_5 gpc41 (
      {stage0_0[175], stage0_0[176], stage0_0[177]},
      {stage0_1[181], stage0_1[182], stage0_1[183], stage0_1[184], stage0_1[185], stage0_1[186]},
      {stage0_2[41]},
      {stage0_3[28]},
      {stage1_4[28],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc606_5 gpc42 (
      {stage0_0[178], stage0_0[179], stage0_0[180], stage0_0[181], stage0_0[182], stage0_0[183]},
      {stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47]},
      {stage1_4[29],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc606_5 gpc43 (
      {stage0_0[184], stage0_0[185], stage0_0[186], stage0_0[187], stage0_0[188], stage0_0[189]},
      {stage0_2[48], stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53]},
      {stage1_4[30],stage1_3[43],stage1_2[43],stage1_1[43],stage1_0[43]}
   );
   gpc606_5 gpc44 (
      {stage0_0[190], stage0_0[191], stage0_0[192], stage0_0[193], stage0_0[194], stage0_0[195]},
      {stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59]},
      {stage1_4[31],stage1_3[44],stage1_2[44],stage1_1[44],stage1_0[44]}
   );
   gpc606_5 gpc45 (
      {stage0_0[196], stage0_0[197], stage0_0[198], stage0_0[199], stage0_0[200], stage0_0[201]},
      {stage0_2[60], stage0_2[61], stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65]},
      {stage1_4[32],stage1_3[45],stage1_2[45],stage1_1[45],stage1_0[45]}
   );
   gpc606_5 gpc46 (
      {stage0_0[202], stage0_0[203], stage0_0[204], stage0_0[205], stage0_0[206], stage0_0[207]},
      {stage0_2[66], stage0_2[67], stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71]},
      {stage1_4[33],stage1_3[46],stage1_2[46],stage1_1[46],stage1_0[46]}
   );
   gpc606_5 gpc47 (
      {stage0_0[208], stage0_0[209], stage0_0[210], stage0_0[211], stage0_0[212], stage0_0[213]},
      {stage0_2[72], stage0_2[73], stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77]},
      {stage1_4[34],stage1_3[47],stage1_2[47],stage1_1[47],stage1_0[47]}
   );
   gpc606_5 gpc48 (
      {stage0_0[214], stage0_0[215], stage0_0[216], stage0_0[217], stage0_0[218], stage0_0[219]},
      {stage0_2[78], stage0_2[79], stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83]},
      {stage1_4[35],stage1_3[48],stage1_2[48],stage1_1[48],stage1_0[48]}
   );
   gpc606_5 gpc49 (
      {stage0_0[220], stage0_0[221], stage0_0[222], stage0_0[223], stage0_0[224], stage0_0[225]},
      {stage0_2[84], stage0_2[85], stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89]},
      {stage1_4[36],stage1_3[49],stage1_2[49],stage1_1[49],stage1_0[49]}
   );
   gpc606_5 gpc50 (
      {stage0_0[226], stage0_0[227], stage0_0[228], stage0_0[229], stage0_0[230], stage0_0[231]},
      {stage0_2[90], stage0_2[91], stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95]},
      {stage1_4[37],stage1_3[50],stage1_2[50],stage1_1[50],stage1_0[50]}
   );
   gpc606_5 gpc51 (
      {stage0_0[232], stage0_0[233], stage0_0[234], stage0_0[235], stage0_0[236], stage0_0[237]},
      {stage0_2[96], stage0_2[97], stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101]},
      {stage1_4[38],stage1_3[51],stage1_2[51],stage1_1[51],stage1_0[51]}
   );
   gpc606_5 gpc52 (
      {stage0_0[238], stage0_0[239], stage0_0[240], stage0_0[241], stage0_0[242], stage0_0[243]},
      {stage0_2[102], stage0_2[103], stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107]},
      {stage1_4[39],stage1_3[52],stage1_2[52],stage1_1[52],stage1_0[52]}
   );
   gpc606_5 gpc53 (
      {stage0_0[244], stage0_0[245], stage0_0[246], stage0_0[247], stage0_0[248], stage0_0[249]},
      {stage0_2[108], stage0_2[109], stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113]},
      {stage1_4[40],stage1_3[53],stage1_2[53],stage1_1[53],stage1_0[53]}
   );
   gpc606_5 gpc54 (
      {stage0_0[250], stage0_0[251], stage0_0[252], stage0_0[253], stage0_0[254], stage0_0[255]},
      {stage0_2[114], stage0_2[115], stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119]},
      {stage1_4[41],stage1_3[54],stage1_2[54],stage1_1[54],stage1_0[54]}
   );
   gpc606_5 gpc55 (
      {stage0_0[256], stage0_0[257], stage0_0[258], stage0_0[259], stage0_0[260], stage0_0[261]},
      {stage0_2[120], stage0_2[121], stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125]},
      {stage1_4[42],stage1_3[55],stage1_2[55],stage1_1[55],stage1_0[55]}
   );
   gpc606_5 gpc56 (
      {stage0_0[262], stage0_0[263], stage0_0[264], stage0_0[265], stage0_0[266], stage0_0[267]},
      {stage0_2[126], stage0_2[127], stage0_2[128], stage0_2[129], stage0_2[130], stage0_2[131]},
      {stage1_4[43],stage1_3[56],stage1_2[56],stage1_1[56],stage1_0[56]}
   );
   gpc606_5 gpc57 (
      {stage0_0[268], stage0_0[269], stage0_0[270], stage0_0[271], stage0_0[272], stage0_0[273]},
      {stage0_2[132], stage0_2[133], stage0_2[134], stage0_2[135], stage0_2[136], stage0_2[137]},
      {stage1_4[44],stage1_3[57],stage1_2[57],stage1_1[57],stage1_0[57]}
   );
   gpc606_5 gpc58 (
      {stage0_0[274], stage0_0[275], stage0_0[276], stage0_0[277], stage0_0[278], stage0_0[279]},
      {stage0_2[138], stage0_2[139], stage0_2[140], stage0_2[141], stage0_2[142], stage0_2[143]},
      {stage1_4[45],stage1_3[58],stage1_2[58],stage1_1[58],stage1_0[58]}
   );
   gpc606_5 gpc59 (
      {stage0_0[280], stage0_0[281], stage0_0[282], stage0_0[283], stage0_0[284], stage0_0[285]},
      {stage0_2[144], stage0_2[145], stage0_2[146], stage0_2[147], stage0_2[148], stage0_2[149]},
      {stage1_4[46],stage1_3[59],stage1_2[59],stage1_1[59],stage1_0[59]}
   );
   gpc606_5 gpc60 (
      {stage0_0[286], stage0_0[287], stage0_0[288], stage0_0[289], stage0_0[290], stage0_0[291]},
      {stage0_2[150], stage0_2[151], stage0_2[152], stage0_2[153], stage0_2[154], stage0_2[155]},
      {stage1_4[47],stage1_3[60],stage1_2[60],stage1_1[60],stage1_0[60]}
   );
   gpc606_5 gpc61 (
      {stage0_0[292], stage0_0[293], stage0_0[294], stage0_0[295], stage0_0[296], stage0_0[297]},
      {stage0_2[156], stage0_2[157], stage0_2[158], stage0_2[159], stage0_2[160], stage0_2[161]},
      {stage1_4[48],stage1_3[61],stage1_2[61],stage1_1[61],stage1_0[61]}
   );
   gpc606_5 gpc62 (
      {stage0_0[298], stage0_0[299], stage0_0[300], stage0_0[301], stage0_0[302], stage0_0[303]},
      {stage0_2[162], stage0_2[163], stage0_2[164], stage0_2[165], stage0_2[166], stage0_2[167]},
      {stage1_4[49],stage1_3[62],stage1_2[62],stage1_1[62],stage1_0[62]}
   );
   gpc606_5 gpc63 (
      {stage0_0[304], stage0_0[305], stage0_0[306], stage0_0[307], stage0_0[308], stage0_0[309]},
      {stage0_2[168], stage0_2[169], stage0_2[170], stage0_2[171], stage0_2[172], stage0_2[173]},
      {stage1_4[50],stage1_3[63],stage1_2[63],stage1_1[63],stage1_0[63]}
   );
   gpc606_5 gpc64 (
      {stage0_0[310], stage0_0[311], stage0_0[312], stage0_0[313], stage0_0[314], stage0_0[315]},
      {stage0_2[174], stage0_2[175], stage0_2[176], stage0_2[177], stage0_2[178], stage0_2[179]},
      {stage1_4[51],stage1_3[64],stage1_2[64],stage1_1[64],stage1_0[64]}
   );
   gpc606_5 gpc65 (
      {stage0_0[316], stage0_0[317], stage0_0[318], stage0_0[319], stage0_0[320], stage0_0[321]},
      {stage0_2[180], stage0_2[181], stage0_2[182], stage0_2[183], stage0_2[184], stage0_2[185]},
      {stage1_4[52],stage1_3[65],stage1_2[65],stage1_1[65],stage1_0[65]}
   );
   gpc606_5 gpc66 (
      {stage0_0[322], stage0_0[323], stage0_0[324], stage0_0[325], stage0_0[326], stage0_0[327]},
      {stage0_2[186], stage0_2[187], stage0_2[188], stage0_2[189], stage0_2[190], stage0_2[191]},
      {stage1_4[53],stage1_3[66],stage1_2[66],stage1_1[66],stage1_0[66]}
   );
   gpc606_5 gpc67 (
      {stage0_0[328], stage0_0[329], stage0_0[330], stage0_0[331], stage0_0[332], stage0_0[333]},
      {stage0_2[192], stage0_2[193], stage0_2[194], stage0_2[195], stage0_2[196], stage0_2[197]},
      {stage1_4[54],stage1_3[67],stage1_2[67],stage1_1[67],stage1_0[67]}
   );
   gpc606_5 gpc68 (
      {stage0_0[334], stage0_0[335], stage0_0[336], stage0_0[337], stage0_0[338], stage0_0[339]},
      {stage0_2[198], stage0_2[199], stage0_2[200], stage0_2[201], stage0_2[202], stage0_2[203]},
      {stage1_4[55],stage1_3[68],stage1_2[68],stage1_1[68],stage1_0[68]}
   );
   gpc606_5 gpc69 (
      {stage0_0[340], stage0_0[341], stage0_0[342], stage0_0[343], stage0_0[344], stage0_0[345]},
      {stage0_2[204], stage0_2[205], stage0_2[206], stage0_2[207], stage0_2[208], stage0_2[209]},
      {stage1_4[56],stage1_3[69],stage1_2[69],stage1_1[69],stage1_0[69]}
   );
   gpc606_5 gpc70 (
      {stage0_0[346], stage0_0[347], stage0_0[348], stage0_0[349], stage0_0[350], stage0_0[351]},
      {stage0_2[210], stage0_2[211], stage0_2[212], stage0_2[213], stage0_2[214], stage0_2[215]},
      {stage1_4[57],stage1_3[70],stage1_2[70],stage1_1[70],stage1_0[70]}
   );
   gpc606_5 gpc71 (
      {stage0_0[352], stage0_0[353], stage0_0[354], stage0_0[355], stage0_0[356], stage0_0[357]},
      {stage0_2[216], stage0_2[217], stage0_2[218], stage0_2[219], stage0_2[220], stage0_2[221]},
      {stage1_4[58],stage1_3[71],stage1_2[71],stage1_1[71],stage1_0[71]}
   );
   gpc606_5 gpc72 (
      {stage0_0[358], stage0_0[359], stage0_0[360], stage0_0[361], stage0_0[362], stage0_0[363]},
      {stage0_2[222], stage0_2[223], stage0_2[224], stage0_2[225], stage0_2[226], stage0_2[227]},
      {stage1_4[59],stage1_3[72],stage1_2[72],stage1_1[72],stage1_0[72]}
   );
   gpc606_5 gpc73 (
      {stage0_0[364], stage0_0[365], stage0_0[366], stage0_0[367], stage0_0[368], stage0_0[369]},
      {stage0_2[228], stage0_2[229], stage0_2[230], stage0_2[231], stage0_2[232], stage0_2[233]},
      {stage1_4[60],stage1_3[73],stage1_2[73],stage1_1[73],stage1_0[73]}
   );
   gpc606_5 gpc74 (
      {stage0_0[370], stage0_0[371], stage0_0[372], stage0_0[373], stage0_0[374], stage0_0[375]},
      {stage0_2[234], stage0_2[235], stage0_2[236], stage0_2[237], stage0_2[238], stage0_2[239]},
      {stage1_4[61],stage1_3[74],stage1_2[74],stage1_1[74],stage1_0[74]}
   );
   gpc606_5 gpc75 (
      {stage0_0[376], stage0_0[377], stage0_0[378], stage0_0[379], stage0_0[380], stage0_0[381]},
      {stage0_2[240], stage0_2[241], stage0_2[242], stage0_2[243], stage0_2[244], stage0_2[245]},
      {stage1_4[62],stage1_3[75],stage1_2[75],stage1_1[75],stage1_0[75]}
   );
   gpc606_5 gpc76 (
      {stage0_0[382], stage0_0[383], stage0_0[384], stage0_0[385], stage0_0[386], stage0_0[387]},
      {stage0_2[246], stage0_2[247], stage0_2[248], stage0_2[249], stage0_2[250], stage0_2[251]},
      {stage1_4[63],stage1_3[76],stage1_2[76],stage1_1[76],stage1_0[76]}
   );
   gpc606_5 gpc77 (
      {stage0_0[388], stage0_0[389], stage0_0[390], stage0_0[391], stage0_0[392], stage0_0[393]},
      {stage0_2[252], stage0_2[253], stage0_2[254], stage0_2[255], stage0_2[256], stage0_2[257]},
      {stage1_4[64],stage1_3[77],stage1_2[77],stage1_1[77],stage1_0[77]}
   );
   gpc606_5 gpc78 (
      {stage0_0[394], stage0_0[395], stage0_0[396], stage0_0[397], stage0_0[398], stage0_0[399]},
      {stage0_2[258], stage0_2[259], stage0_2[260], stage0_2[261], stage0_2[262], stage0_2[263]},
      {stage1_4[65],stage1_3[78],stage1_2[78],stage1_1[78],stage1_0[78]}
   );
   gpc606_5 gpc79 (
      {stage0_0[400], stage0_0[401], stage0_0[402], stage0_0[403], stage0_0[404], stage0_0[405]},
      {stage0_2[264], stage0_2[265], stage0_2[266], stage0_2[267], stage0_2[268], stage0_2[269]},
      {stage1_4[66],stage1_3[79],stage1_2[79],stage1_1[79],stage1_0[79]}
   );
   gpc606_5 gpc80 (
      {stage0_0[406], stage0_0[407], stage0_0[408], stage0_0[409], stage0_0[410], stage0_0[411]},
      {stage0_2[270], stage0_2[271], stage0_2[272], stage0_2[273], stage0_2[274], stage0_2[275]},
      {stage1_4[67],stage1_3[80],stage1_2[80],stage1_1[80],stage1_0[80]}
   );
   gpc606_5 gpc81 (
      {stage0_0[412], stage0_0[413], stage0_0[414], stage0_0[415], stage0_0[416], stage0_0[417]},
      {stage0_2[276], stage0_2[277], stage0_2[278], stage0_2[279], stage0_2[280], stage0_2[281]},
      {stage1_4[68],stage1_3[81],stage1_2[81],stage1_1[81],stage1_0[81]}
   );
   gpc606_5 gpc82 (
      {stage0_0[418], stage0_0[419], stage0_0[420], stage0_0[421], stage0_0[422], stage0_0[423]},
      {stage0_2[282], stage0_2[283], stage0_2[284], stage0_2[285], stage0_2[286], stage0_2[287]},
      {stage1_4[69],stage1_3[82],stage1_2[82],stage1_1[82],stage1_0[82]}
   );
   gpc606_5 gpc83 (
      {stage0_0[424], stage0_0[425], stage0_0[426], stage0_0[427], stage0_0[428], stage0_0[429]},
      {stage0_2[288], stage0_2[289], stage0_2[290], stage0_2[291], stage0_2[292], stage0_2[293]},
      {stage1_4[70],stage1_3[83],stage1_2[83],stage1_1[83],stage1_0[83]}
   );
   gpc606_5 gpc84 (
      {stage0_0[430], stage0_0[431], stage0_0[432], stage0_0[433], stage0_0[434], stage0_0[435]},
      {stage0_2[294], stage0_2[295], stage0_2[296], stage0_2[297], stage0_2[298], stage0_2[299]},
      {stage1_4[71],stage1_3[84],stage1_2[84],stage1_1[84],stage1_0[84]}
   );
   gpc606_5 gpc85 (
      {stage0_0[436], stage0_0[437], stage0_0[438], stage0_0[439], stage0_0[440], stage0_0[441]},
      {stage0_2[300], stage0_2[301], stage0_2[302], stage0_2[303], stage0_2[304], stage0_2[305]},
      {stage1_4[72],stage1_3[85],stage1_2[85],stage1_1[85],stage1_0[85]}
   );
   gpc606_5 gpc86 (
      {stage0_0[442], stage0_0[443], stage0_0[444], stage0_0[445], stage0_0[446], stage0_0[447]},
      {stage0_2[306], stage0_2[307], stage0_2[308], stage0_2[309], stage0_2[310], stage0_2[311]},
      {stage1_4[73],stage1_3[86],stage1_2[86],stage1_1[86],stage1_0[86]}
   );
   gpc606_5 gpc87 (
      {stage0_1[187], stage0_1[188], stage0_1[189], stage0_1[190], stage0_1[191], stage0_1[192]},
      {stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32], stage0_3[33], stage0_3[34]},
      {stage1_5[0],stage1_4[74],stage1_3[87],stage1_2[87],stage1_1[87]}
   );
   gpc606_5 gpc88 (
      {stage0_1[193], stage0_1[194], stage0_1[195], stage0_1[196], stage0_1[197], stage0_1[198]},
      {stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39], stage0_3[40]},
      {stage1_5[1],stage1_4[75],stage1_3[88],stage1_2[88],stage1_1[88]}
   );
   gpc606_5 gpc89 (
      {stage0_1[199], stage0_1[200], stage0_1[201], stage0_1[202], stage0_1[203], stage0_1[204]},
      {stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46]},
      {stage1_5[2],stage1_4[76],stage1_3[89],stage1_2[89],stage1_1[89]}
   );
   gpc606_5 gpc90 (
      {stage0_1[205], stage0_1[206], stage0_1[207], stage0_1[208], stage0_1[209], stage0_1[210]},
      {stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50], stage0_3[51], stage0_3[52]},
      {stage1_5[3],stage1_4[77],stage1_3[90],stage1_2[90],stage1_1[90]}
   );
   gpc606_5 gpc91 (
      {stage0_1[211], stage0_1[212], stage0_1[213], stage0_1[214], stage0_1[215], stage0_1[216]},
      {stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56], stage0_3[57], stage0_3[58]},
      {stage1_5[4],stage1_4[78],stage1_3[91],stage1_2[91],stage1_1[91]}
   );
   gpc606_5 gpc92 (
      {stage0_1[217], stage0_1[218], stage0_1[219], stage0_1[220], stage0_1[221], stage0_1[222]},
      {stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62], stage0_3[63], stage0_3[64]},
      {stage1_5[5],stage1_4[79],stage1_3[92],stage1_2[92],stage1_1[92]}
   );
   gpc606_5 gpc93 (
      {stage0_1[223], stage0_1[224], stage0_1[225], stage0_1[226], stage0_1[227], stage0_1[228]},
      {stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68], stage0_3[69], stage0_3[70]},
      {stage1_5[6],stage1_4[80],stage1_3[93],stage1_2[93],stage1_1[93]}
   );
   gpc606_5 gpc94 (
      {stage0_1[229], stage0_1[230], stage0_1[231], stage0_1[232], stage0_1[233], stage0_1[234]},
      {stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74], stage0_3[75], stage0_3[76]},
      {stage1_5[7],stage1_4[81],stage1_3[94],stage1_2[94],stage1_1[94]}
   );
   gpc606_5 gpc95 (
      {stage0_1[235], stage0_1[236], stage0_1[237], stage0_1[238], stage0_1[239], stage0_1[240]},
      {stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80], stage0_3[81], stage0_3[82]},
      {stage1_5[8],stage1_4[82],stage1_3[95],stage1_2[95],stage1_1[95]}
   );
   gpc606_5 gpc96 (
      {stage0_1[241], stage0_1[242], stage0_1[243], stage0_1[244], stage0_1[245], stage0_1[246]},
      {stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86], stage0_3[87], stage0_3[88]},
      {stage1_5[9],stage1_4[83],stage1_3[96],stage1_2[96],stage1_1[96]}
   );
   gpc606_5 gpc97 (
      {stage0_1[247], stage0_1[248], stage0_1[249], stage0_1[250], stage0_1[251], stage0_1[252]},
      {stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92], stage0_3[93], stage0_3[94]},
      {stage1_5[10],stage1_4[84],stage1_3[97],stage1_2[97],stage1_1[97]}
   );
   gpc606_5 gpc98 (
      {stage0_1[253], stage0_1[254], stage0_1[255], stage0_1[256], stage0_1[257], stage0_1[258]},
      {stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98], stage0_3[99], stage0_3[100]},
      {stage1_5[11],stage1_4[85],stage1_3[98],stage1_2[98],stage1_1[98]}
   );
   gpc606_5 gpc99 (
      {stage0_1[259], stage0_1[260], stage0_1[261], stage0_1[262], stage0_1[263], stage0_1[264]},
      {stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104], stage0_3[105], stage0_3[106]},
      {stage1_5[12],stage1_4[86],stage1_3[99],stage1_2[99],stage1_1[99]}
   );
   gpc606_5 gpc100 (
      {stage0_1[265], stage0_1[266], stage0_1[267], stage0_1[268], stage0_1[269], stage0_1[270]},
      {stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110], stage0_3[111], stage0_3[112]},
      {stage1_5[13],stage1_4[87],stage1_3[100],stage1_2[100],stage1_1[100]}
   );
   gpc606_5 gpc101 (
      {stage0_1[271], stage0_1[272], stage0_1[273], stage0_1[274], stage0_1[275], stage0_1[276]},
      {stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116], stage0_3[117], stage0_3[118]},
      {stage1_5[14],stage1_4[88],stage1_3[101],stage1_2[101],stage1_1[101]}
   );
   gpc606_5 gpc102 (
      {stage0_1[277], stage0_1[278], stage0_1[279], stage0_1[280], stage0_1[281], stage0_1[282]},
      {stage0_3[119], stage0_3[120], stage0_3[121], stage0_3[122], stage0_3[123], stage0_3[124]},
      {stage1_5[15],stage1_4[89],stage1_3[102],stage1_2[102],stage1_1[102]}
   );
   gpc606_5 gpc103 (
      {stage0_1[283], stage0_1[284], stage0_1[285], stage0_1[286], stage0_1[287], stage0_1[288]},
      {stage0_3[125], stage0_3[126], stage0_3[127], stage0_3[128], stage0_3[129], stage0_3[130]},
      {stage1_5[16],stage1_4[90],stage1_3[103],stage1_2[103],stage1_1[103]}
   );
   gpc606_5 gpc104 (
      {stage0_1[289], stage0_1[290], stage0_1[291], stage0_1[292], stage0_1[293], stage0_1[294]},
      {stage0_3[131], stage0_3[132], stage0_3[133], stage0_3[134], stage0_3[135], stage0_3[136]},
      {stage1_5[17],stage1_4[91],stage1_3[104],stage1_2[104],stage1_1[104]}
   );
   gpc606_5 gpc105 (
      {stage0_1[295], stage0_1[296], stage0_1[297], stage0_1[298], stage0_1[299], stage0_1[300]},
      {stage0_3[137], stage0_3[138], stage0_3[139], stage0_3[140], stage0_3[141], stage0_3[142]},
      {stage1_5[18],stage1_4[92],stage1_3[105],stage1_2[105],stage1_1[105]}
   );
   gpc606_5 gpc106 (
      {stage0_1[301], stage0_1[302], stage0_1[303], stage0_1[304], stage0_1[305], stage0_1[306]},
      {stage0_3[143], stage0_3[144], stage0_3[145], stage0_3[146], stage0_3[147], stage0_3[148]},
      {stage1_5[19],stage1_4[93],stage1_3[106],stage1_2[106],stage1_1[106]}
   );
   gpc606_5 gpc107 (
      {stage0_1[307], stage0_1[308], stage0_1[309], stage0_1[310], stage0_1[311], stage0_1[312]},
      {stage0_3[149], stage0_3[150], stage0_3[151], stage0_3[152], stage0_3[153], stage0_3[154]},
      {stage1_5[20],stage1_4[94],stage1_3[107],stage1_2[107],stage1_1[107]}
   );
   gpc606_5 gpc108 (
      {stage0_1[313], stage0_1[314], stage0_1[315], stage0_1[316], stage0_1[317], stage0_1[318]},
      {stage0_3[155], stage0_3[156], stage0_3[157], stage0_3[158], stage0_3[159], stage0_3[160]},
      {stage1_5[21],stage1_4[95],stage1_3[108],stage1_2[108],stage1_1[108]}
   );
   gpc606_5 gpc109 (
      {stage0_1[319], stage0_1[320], stage0_1[321], stage0_1[322], stage0_1[323], stage0_1[324]},
      {stage0_3[161], stage0_3[162], stage0_3[163], stage0_3[164], stage0_3[165], stage0_3[166]},
      {stage1_5[22],stage1_4[96],stage1_3[109],stage1_2[109],stage1_1[109]}
   );
   gpc606_5 gpc110 (
      {stage0_1[325], stage0_1[326], stage0_1[327], stage0_1[328], stage0_1[329], stage0_1[330]},
      {stage0_3[167], stage0_3[168], stage0_3[169], stage0_3[170], stage0_3[171], stage0_3[172]},
      {stage1_5[23],stage1_4[97],stage1_3[110],stage1_2[110],stage1_1[110]}
   );
   gpc606_5 gpc111 (
      {stage0_1[331], stage0_1[332], stage0_1[333], stage0_1[334], stage0_1[335], stage0_1[336]},
      {stage0_3[173], stage0_3[174], stage0_3[175], stage0_3[176], stage0_3[177], stage0_3[178]},
      {stage1_5[24],stage1_4[98],stage1_3[111],stage1_2[111],stage1_1[111]}
   );
   gpc606_5 gpc112 (
      {stage0_1[337], stage0_1[338], stage0_1[339], stage0_1[340], stage0_1[341], stage0_1[342]},
      {stage0_3[179], stage0_3[180], stage0_3[181], stage0_3[182], stage0_3[183], stage0_3[184]},
      {stage1_5[25],stage1_4[99],stage1_3[112],stage1_2[112],stage1_1[112]}
   );
   gpc606_5 gpc113 (
      {stage0_1[343], stage0_1[344], stage0_1[345], stage0_1[346], stage0_1[347], stage0_1[348]},
      {stage0_3[185], stage0_3[186], stage0_3[187], stage0_3[188], stage0_3[189], stage0_3[190]},
      {stage1_5[26],stage1_4[100],stage1_3[113],stage1_2[113],stage1_1[113]}
   );
   gpc606_5 gpc114 (
      {stage0_1[349], stage0_1[350], stage0_1[351], stage0_1[352], stage0_1[353], stage0_1[354]},
      {stage0_3[191], stage0_3[192], stage0_3[193], stage0_3[194], stage0_3[195], stage0_3[196]},
      {stage1_5[27],stage1_4[101],stage1_3[114],stage1_2[114],stage1_1[114]}
   );
   gpc606_5 gpc115 (
      {stage0_1[355], stage0_1[356], stage0_1[357], stage0_1[358], stage0_1[359], stage0_1[360]},
      {stage0_3[197], stage0_3[198], stage0_3[199], stage0_3[200], stage0_3[201], stage0_3[202]},
      {stage1_5[28],stage1_4[102],stage1_3[115],stage1_2[115],stage1_1[115]}
   );
   gpc606_5 gpc116 (
      {stage0_1[361], stage0_1[362], stage0_1[363], stage0_1[364], stage0_1[365], stage0_1[366]},
      {stage0_3[203], stage0_3[204], stage0_3[205], stage0_3[206], stage0_3[207], stage0_3[208]},
      {stage1_5[29],stage1_4[103],stage1_3[116],stage1_2[116],stage1_1[116]}
   );
   gpc606_5 gpc117 (
      {stage0_1[367], stage0_1[368], stage0_1[369], stage0_1[370], stage0_1[371], stage0_1[372]},
      {stage0_3[209], stage0_3[210], stage0_3[211], stage0_3[212], stage0_3[213], stage0_3[214]},
      {stage1_5[30],stage1_4[104],stage1_3[117],stage1_2[117],stage1_1[117]}
   );
   gpc606_5 gpc118 (
      {stage0_1[373], stage0_1[374], stage0_1[375], stage0_1[376], stage0_1[377], stage0_1[378]},
      {stage0_3[215], stage0_3[216], stage0_3[217], stage0_3[218], stage0_3[219], stage0_3[220]},
      {stage1_5[31],stage1_4[105],stage1_3[118],stage1_2[118],stage1_1[118]}
   );
   gpc606_5 gpc119 (
      {stage0_1[379], stage0_1[380], stage0_1[381], stage0_1[382], stage0_1[383], stage0_1[384]},
      {stage0_3[221], stage0_3[222], stage0_3[223], stage0_3[224], stage0_3[225], stage0_3[226]},
      {stage1_5[32],stage1_4[106],stage1_3[119],stage1_2[119],stage1_1[119]}
   );
   gpc606_5 gpc120 (
      {stage0_1[385], stage0_1[386], stage0_1[387], stage0_1[388], stage0_1[389], stage0_1[390]},
      {stage0_3[227], stage0_3[228], stage0_3[229], stage0_3[230], stage0_3[231], stage0_3[232]},
      {stage1_5[33],stage1_4[107],stage1_3[120],stage1_2[120],stage1_1[120]}
   );
   gpc606_5 gpc121 (
      {stage0_1[391], stage0_1[392], stage0_1[393], stage0_1[394], stage0_1[395], stage0_1[396]},
      {stage0_3[233], stage0_3[234], stage0_3[235], stage0_3[236], stage0_3[237], stage0_3[238]},
      {stage1_5[34],stage1_4[108],stage1_3[121],stage1_2[121],stage1_1[121]}
   );
   gpc606_5 gpc122 (
      {stage0_1[397], stage0_1[398], stage0_1[399], stage0_1[400], stage0_1[401], stage0_1[402]},
      {stage0_3[239], stage0_3[240], stage0_3[241], stage0_3[242], stage0_3[243], stage0_3[244]},
      {stage1_5[35],stage1_4[109],stage1_3[122],stage1_2[122],stage1_1[122]}
   );
   gpc606_5 gpc123 (
      {stage0_1[403], stage0_1[404], stage0_1[405], stage0_1[406], stage0_1[407], stage0_1[408]},
      {stage0_3[245], stage0_3[246], stage0_3[247], stage0_3[248], stage0_3[249], stage0_3[250]},
      {stage1_5[36],stage1_4[110],stage1_3[123],stage1_2[123],stage1_1[123]}
   );
   gpc606_5 gpc124 (
      {stage0_1[409], stage0_1[410], stage0_1[411], stage0_1[412], stage0_1[413], stage0_1[414]},
      {stage0_3[251], stage0_3[252], stage0_3[253], stage0_3[254], stage0_3[255], stage0_3[256]},
      {stage1_5[37],stage1_4[111],stage1_3[124],stage1_2[124],stage1_1[124]}
   );
   gpc606_5 gpc125 (
      {stage0_1[415], stage0_1[416], stage0_1[417], stage0_1[418], stage0_1[419], stage0_1[420]},
      {stage0_3[257], stage0_3[258], stage0_3[259], stage0_3[260], stage0_3[261], stage0_3[262]},
      {stage1_5[38],stage1_4[112],stage1_3[125],stage1_2[125],stage1_1[125]}
   );
   gpc606_5 gpc126 (
      {stage0_1[421], stage0_1[422], stage0_1[423], stage0_1[424], stage0_1[425], stage0_1[426]},
      {stage0_3[263], stage0_3[264], stage0_3[265], stage0_3[266], stage0_3[267], stage0_3[268]},
      {stage1_5[39],stage1_4[113],stage1_3[126],stage1_2[126],stage1_1[126]}
   );
   gpc606_5 gpc127 (
      {stage0_1[427], stage0_1[428], stage0_1[429], stage0_1[430], stage0_1[431], stage0_1[432]},
      {stage0_3[269], stage0_3[270], stage0_3[271], stage0_3[272], stage0_3[273], stage0_3[274]},
      {stage1_5[40],stage1_4[114],stage1_3[127],stage1_2[127],stage1_1[127]}
   );
   gpc606_5 gpc128 (
      {stage0_1[433], stage0_1[434], stage0_1[435], stage0_1[436], stage0_1[437], stage0_1[438]},
      {stage0_3[275], stage0_3[276], stage0_3[277], stage0_3[278], stage0_3[279], stage0_3[280]},
      {stage1_5[41],stage1_4[115],stage1_3[128],stage1_2[128],stage1_1[128]}
   );
   gpc606_5 gpc129 (
      {stage0_2[312], stage0_2[313], stage0_2[314], stage0_2[315], stage0_2[316], stage0_2[317]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[42],stage1_4[116],stage1_3[129],stage1_2[129]}
   );
   gpc606_5 gpc130 (
      {stage0_2[318], stage0_2[319], stage0_2[320], stage0_2[321], stage0_2[322], stage0_2[323]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[43],stage1_4[117],stage1_3[130],stage1_2[130]}
   );
   gpc606_5 gpc131 (
      {stage0_2[324], stage0_2[325], stage0_2[326], stage0_2[327], stage0_2[328], stage0_2[329]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[44],stage1_4[118],stage1_3[131],stage1_2[131]}
   );
   gpc606_5 gpc132 (
      {stage0_2[330], stage0_2[331], stage0_2[332], stage0_2[333], stage0_2[334], stage0_2[335]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[45],stage1_4[119],stage1_3[132],stage1_2[132]}
   );
   gpc606_5 gpc133 (
      {stage0_2[336], stage0_2[337], stage0_2[338], stage0_2[339], stage0_2[340], stage0_2[341]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[46],stage1_4[120],stage1_3[133],stage1_2[133]}
   );
   gpc606_5 gpc134 (
      {stage0_2[342], stage0_2[343], stage0_2[344], stage0_2[345], stage0_2[346], stage0_2[347]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[47],stage1_4[121],stage1_3[134],stage1_2[134]}
   );
   gpc606_5 gpc135 (
      {stage0_2[348], stage0_2[349], stage0_2[350], stage0_2[351], stage0_2[352], stage0_2[353]},
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage1_6[6],stage1_5[48],stage1_4[122],stage1_3[135],stage1_2[135]}
   );
   gpc606_5 gpc136 (
      {stage0_2[354], stage0_2[355], stage0_2[356], stage0_2[357], stage0_2[358], stage0_2[359]},
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage1_6[7],stage1_5[49],stage1_4[123],stage1_3[136],stage1_2[136]}
   );
   gpc606_5 gpc137 (
      {stage0_2[360], stage0_2[361], stage0_2[362], stage0_2[363], stage0_2[364], stage0_2[365]},
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage1_6[8],stage1_5[50],stage1_4[124],stage1_3[137],stage1_2[137]}
   );
   gpc606_5 gpc138 (
      {stage0_2[366], stage0_2[367], stage0_2[368], stage0_2[369], stage0_2[370], stage0_2[371]},
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage1_6[9],stage1_5[51],stage1_4[125],stage1_3[138],stage1_2[138]}
   );
   gpc606_5 gpc139 (
      {stage0_2[372], stage0_2[373], stage0_2[374], stage0_2[375], stage0_2[376], stage0_2[377]},
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage1_6[10],stage1_5[52],stage1_4[126],stage1_3[139],stage1_2[139]}
   );
   gpc606_5 gpc140 (
      {stage0_2[378], stage0_2[379], stage0_2[380], stage0_2[381], stage0_2[382], stage0_2[383]},
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage1_6[11],stage1_5[53],stage1_4[127],stage1_3[140],stage1_2[140]}
   );
   gpc606_5 gpc141 (
      {stage0_2[384], stage0_2[385], stage0_2[386], stage0_2[387], stage0_2[388], stage0_2[389]},
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage1_6[12],stage1_5[54],stage1_4[128],stage1_3[141],stage1_2[141]}
   );
   gpc606_5 gpc142 (
      {stage0_2[390], stage0_2[391], stage0_2[392], stage0_2[393], stage0_2[394], stage0_2[395]},
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage1_6[13],stage1_5[55],stage1_4[129],stage1_3[142],stage1_2[142]}
   );
   gpc606_5 gpc143 (
      {stage0_2[396], stage0_2[397], stage0_2[398], stage0_2[399], stage0_2[400], stage0_2[401]},
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage1_6[14],stage1_5[56],stage1_4[130],stage1_3[143],stage1_2[143]}
   );
   gpc606_5 gpc144 (
      {stage0_2[402], stage0_2[403], stage0_2[404], stage0_2[405], stage0_2[406], stage0_2[407]},
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage1_6[15],stage1_5[57],stage1_4[131],stage1_3[144],stage1_2[144]}
   );
   gpc606_5 gpc145 (
      {stage0_2[408], stage0_2[409], stage0_2[410], stage0_2[411], stage0_2[412], stage0_2[413]},
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage1_6[16],stage1_5[58],stage1_4[132],stage1_3[145],stage1_2[145]}
   );
   gpc606_5 gpc146 (
      {stage0_2[414], stage0_2[415], stage0_2[416], stage0_2[417], stage0_2[418], stage0_2[419]},
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage1_6[17],stage1_5[59],stage1_4[133],stage1_3[146],stage1_2[146]}
   );
   gpc606_5 gpc147 (
      {stage0_2[420], stage0_2[421], stage0_2[422], stage0_2[423], stage0_2[424], stage0_2[425]},
      {stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113]},
      {stage1_6[18],stage1_5[60],stage1_4[134],stage1_3[147],stage1_2[147]}
   );
   gpc606_5 gpc148 (
      {stage0_2[426], stage0_2[427], stage0_2[428], stage0_2[429], stage0_2[430], stage0_2[431]},
      {stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119]},
      {stage1_6[19],stage1_5[61],stage1_4[135],stage1_3[148],stage1_2[148]}
   );
   gpc606_5 gpc149 (
      {stage0_2[432], stage0_2[433], stage0_2[434], stage0_2[435], stage0_2[436], stage0_2[437]},
      {stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125]},
      {stage1_6[20],stage1_5[62],stage1_4[136],stage1_3[149],stage1_2[149]}
   );
   gpc606_5 gpc150 (
      {stage0_2[438], stage0_2[439], stage0_2[440], stage0_2[441], stage0_2[442], stage0_2[443]},
      {stage0_4[126], stage0_4[127], stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131]},
      {stage1_6[21],stage1_5[63],stage1_4[137],stage1_3[150],stage1_2[150]}
   );
   gpc606_5 gpc151 (
      {stage0_2[444], stage0_2[445], stage0_2[446], stage0_2[447], stage0_2[448], stage0_2[449]},
      {stage0_4[132], stage0_4[133], stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137]},
      {stage1_6[22],stage1_5[64],stage1_4[138],stage1_3[151],stage1_2[151]}
   );
   gpc606_5 gpc152 (
      {stage0_2[450], stage0_2[451], stage0_2[452], stage0_2[453], stage0_2[454], stage0_2[455]},
      {stage0_4[138], stage0_4[139], stage0_4[140], stage0_4[141], stage0_4[142], stage0_4[143]},
      {stage1_6[23],stage1_5[65],stage1_4[139],stage1_3[152],stage1_2[152]}
   );
   gpc606_5 gpc153 (
      {stage0_2[456], stage0_2[457], stage0_2[458], stage0_2[459], stage0_2[460], stage0_2[461]},
      {stage0_4[144], stage0_4[145], stage0_4[146], stage0_4[147], stage0_4[148], stage0_4[149]},
      {stage1_6[24],stage1_5[66],stage1_4[140],stage1_3[153],stage1_2[153]}
   );
   gpc606_5 gpc154 (
      {stage0_2[462], stage0_2[463], stage0_2[464], stage0_2[465], stage0_2[466], stage0_2[467]},
      {stage0_4[150], stage0_4[151], stage0_4[152], stage0_4[153], stage0_4[154], stage0_4[155]},
      {stage1_6[25],stage1_5[67],stage1_4[141],stage1_3[154],stage1_2[154]}
   );
   gpc606_5 gpc155 (
      {stage0_2[468], stage0_2[469], stage0_2[470], stage0_2[471], stage0_2[472], stage0_2[473]},
      {stage0_4[156], stage0_4[157], stage0_4[158], stage0_4[159], stage0_4[160], stage0_4[161]},
      {stage1_6[26],stage1_5[68],stage1_4[142],stage1_3[155],stage1_2[155]}
   );
   gpc606_5 gpc156 (
      {stage0_2[474], stage0_2[475], stage0_2[476], stage0_2[477], stage0_2[478], stage0_2[479]},
      {stage0_4[162], stage0_4[163], stage0_4[164], stage0_4[165], stage0_4[166], stage0_4[167]},
      {stage1_6[27],stage1_5[69],stage1_4[143],stage1_3[156],stage1_2[156]}
   );
   gpc606_5 gpc157 (
      {stage0_2[480], stage0_2[481], stage0_2[482], stage0_2[483], stage0_2[484], stage0_2[485]},
      {stage0_4[168], stage0_4[169], stage0_4[170], stage0_4[171], stage0_4[172], stage0_4[173]},
      {stage1_6[28],stage1_5[70],stage1_4[144],stage1_3[157],stage1_2[157]}
   );
   gpc615_5 gpc158 (
      {stage0_3[281], stage0_3[282], stage0_3[283], stage0_3[284], stage0_3[285]},
      {stage0_4[174]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[29],stage1_5[71],stage1_4[145],stage1_3[158]}
   );
   gpc615_5 gpc159 (
      {stage0_3[286], stage0_3[287], stage0_3[288], stage0_3[289], stage0_3[290]},
      {stage0_4[175]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[30],stage1_5[72],stage1_4[146],stage1_3[159]}
   );
   gpc615_5 gpc160 (
      {stage0_3[291], stage0_3[292], stage0_3[293], stage0_3[294], stage0_3[295]},
      {stage0_4[176]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[31],stage1_5[73],stage1_4[147],stage1_3[160]}
   );
   gpc615_5 gpc161 (
      {stage0_3[296], stage0_3[297], stage0_3[298], stage0_3[299], stage0_3[300]},
      {stage0_4[177]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[32],stage1_5[74],stage1_4[148],stage1_3[161]}
   );
   gpc615_5 gpc162 (
      {stage0_3[301], stage0_3[302], stage0_3[303], stage0_3[304], stage0_3[305]},
      {stage0_4[178]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[33],stage1_5[75],stage1_4[149],stage1_3[162]}
   );
   gpc615_5 gpc163 (
      {stage0_3[306], stage0_3[307], stage0_3[308], stage0_3[309], stage0_3[310]},
      {stage0_4[179]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[34],stage1_5[76],stage1_4[150],stage1_3[163]}
   );
   gpc615_5 gpc164 (
      {stage0_3[311], stage0_3[312], stage0_3[313], stage0_3[314], stage0_3[315]},
      {stage0_4[180]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[35],stage1_5[77],stage1_4[151],stage1_3[164]}
   );
   gpc615_5 gpc165 (
      {stage0_3[316], stage0_3[317], stage0_3[318], stage0_3[319], stage0_3[320]},
      {stage0_4[181]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage1_7[7],stage1_6[36],stage1_5[78],stage1_4[152],stage1_3[165]}
   );
   gpc615_5 gpc166 (
      {stage0_3[321], stage0_3[322], stage0_3[323], stage0_3[324], stage0_3[325]},
      {stage0_4[182]},
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage1_7[8],stage1_6[37],stage1_5[79],stage1_4[153],stage1_3[166]}
   );
   gpc615_5 gpc167 (
      {stage0_3[326], stage0_3[327], stage0_3[328], stage0_3[329], stage0_3[330]},
      {stage0_4[183]},
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage1_7[9],stage1_6[38],stage1_5[80],stage1_4[154],stage1_3[167]}
   );
   gpc615_5 gpc168 (
      {stage0_3[331], stage0_3[332], stage0_3[333], stage0_3[334], stage0_3[335]},
      {stage0_4[184]},
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage1_7[10],stage1_6[39],stage1_5[81],stage1_4[155],stage1_3[168]}
   );
   gpc615_5 gpc169 (
      {stage0_3[336], stage0_3[337], stage0_3[338], stage0_3[339], stage0_3[340]},
      {stage0_4[185]},
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage1_7[11],stage1_6[40],stage1_5[82],stage1_4[156],stage1_3[169]}
   );
   gpc615_5 gpc170 (
      {stage0_3[341], stage0_3[342], stage0_3[343], stage0_3[344], stage0_3[345]},
      {stage0_4[186]},
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage1_7[12],stage1_6[41],stage1_5[83],stage1_4[157],stage1_3[170]}
   );
   gpc615_5 gpc171 (
      {stage0_3[346], stage0_3[347], stage0_3[348], stage0_3[349], stage0_3[350]},
      {stage0_4[187]},
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage1_7[13],stage1_6[42],stage1_5[84],stage1_4[158],stage1_3[171]}
   );
   gpc615_5 gpc172 (
      {stage0_3[351], stage0_3[352], stage0_3[353], stage0_3[354], stage0_3[355]},
      {stage0_4[188]},
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage1_7[14],stage1_6[43],stage1_5[85],stage1_4[159],stage1_3[172]}
   );
   gpc615_5 gpc173 (
      {stage0_3[356], stage0_3[357], stage0_3[358], stage0_3[359], stage0_3[360]},
      {stage0_4[189]},
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage1_7[15],stage1_6[44],stage1_5[86],stage1_4[160],stage1_3[173]}
   );
   gpc615_5 gpc174 (
      {stage0_3[361], stage0_3[362], stage0_3[363], stage0_3[364], stage0_3[365]},
      {stage0_4[190]},
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage1_7[16],stage1_6[45],stage1_5[87],stage1_4[161],stage1_3[174]}
   );
   gpc615_5 gpc175 (
      {stage0_3[366], stage0_3[367], stage0_3[368], stage0_3[369], stage0_3[370]},
      {stage0_4[191]},
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage1_7[17],stage1_6[46],stage1_5[88],stage1_4[162],stage1_3[175]}
   );
   gpc615_5 gpc176 (
      {stage0_3[371], stage0_3[372], stage0_3[373], stage0_3[374], stage0_3[375]},
      {stage0_4[192]},
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage1_7[18],stage1_6[47],stage1_5[89],stage1_4[163],stage1_3[176]}
   );
   gpc615_5 gpc177 (
      {stage0_3[376], stage0_3[377], stage0_3[378], stage0_3[379], stage0_3[380]},
      {stage0_4[193]},
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage1_7[19],stage1_6[48],stage1_5[90],stage1_4[164],stage1_3[177]}
   );
   gpc615_5 gpc178 (
      {stage0_3[381], stage0_3[382], stage0_3[383], stage0_3[384], stage0_3[385]},
      {stage0_4[194]},
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage1_7[20],stage1_6[49],stage1_5[91],stage1_4[165],stage1_3[178]}
   );
   gpc615_5 gpc179 (
      {stage0_3[386], stage0_3[387], stage0_3[388], stage0_3[389], stage0_3[390]},
      {stage0_4[195]},
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage1_7[21],stage1_6[50],stage1_5[92],stage1_4[166],stage1_3[179]}
   );
   gpc615_5 gpc180 (
      {stage0_3[391], stage0_3[392], stage0_3[393], stage0_3[394], stage0_3[395]},
      {stage0_4[196]},
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage1_7[22],stage1_6[51],stage1_5[93],stage1_4[167],stage1_3[180]}
   );
   gpc615_5 gpc181 (
      {stage0_3[396], stage0_3[397], stage0_3[398], stage0_3[399], stage0_3[400]},
      {stage0_4[197]},
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage1_7[23],stage1_6[52],stage1_5[94],stage1_4[168],stage1_3[181]}
   );
   gpc615_5 gpc182 (
      {stage0_3[401], stage0_3[402], stage0_3[403], stage0_3[404], stage0_3[405]},
      {stage0_4[198]},
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage1_7[24],stage1_6[53],stage1_5[95],stage1_4[169],stage1_3[182]}
   );
   gpc615_5 gpc183 (
      {stage0_3[406], stage0_3[407], stage0_3[408], stage0_3[409], stage0_3[410]},
      {stage0_4[199]},
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155]},
      {stage1_7[25],stage1_6[54],stage1_5[96],stage1_4[170],stage1_3[183]}
   );
   gpc615_5 gpc184 (
      {stage0_3[411], stage0_3[412], stage0_3[413], stage0_3[414], stage0_3[415]},
      {stage0_4[200]},
      {stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161]},
      {stage1_7[26],stage1_6[55],stage1_5[97],stage1_4[171],stage1_3[184]}
   );
   gpc615_5 gpc185 (
      {stage0_3[416], stage0_3[417], stage0_3[418], stage0_3[419], stage0_3[420]},
      {stage0_4[201]},
      {stage0_5[162], stage0_5[163], stage0_5[164], stage0_5[165], stage0_5[166], stage0_5[167]},
      {stage1_7[27],stage1_6[56],stage1_5[98],stage1_4[172],stage1_3[185]}
   );
   gpc615_5 gpc186 (
      {stage0_3[421], stage0_3[422], stage0_3[423], stage0_3[424], stage0_3[425]},
      {stage0_4[202]},
      {stage0_5[168], stage0_5[169], stage0_5[170], stage0_5[171], stage0_5[172], stage0_5[173]},
      {stage1_7[28],stage1_6[57],stage1_5[99],stage1_4[173],stage1_3[186]}
   );
   gpc615_5 gpc187 (
      {stage0_3[426], stage0_3[427], stage0_3[428], stage0_3[429], stage0_3[430]},
      {stage0_4[203]},
      {stage0_5[174], stage0_5[175], stage0_5[176], stage0_5[177], stage0_5[178], stage0_5[179]},
      {stage1_7[29],stage1_6[58],stage1_5[100],stage1_4[174],stage1_3[187]}
   );
   gpc615_5 gpc188 (
      {stage0_3[431], stage0_3[432], stage0_3[433], stage0_3[434], stage0_3[435]},
      {stage0_4[204]},
      {stage0_5[180], stage0_5[181], stage0_5[182], stage0_5[183], stage0_5[184], stage0_5[185]},
      {stage1_7[30],stage1_6[59],stage1_5[101],stage1_4[175],stage1_3[188]}
   );
   gpc615_5 gpc189 (
      {stage0_3[436], stage0_3[437], stage0_3[438], stage0_3[439], stage0_3[440]},
      {stage0_4[205]},
      {stage0_5[186], stage0_5[187], stage0_5[188], stage0_5[189], stage0_5[190], stage0_5[191]},
      {stage1_7[31],stage1_6[60],stage1_5[102],stage1_4[176],stage1_3[189]}
   );
   gpc615_5 gpc190 (
      {stage0_3[441], stage0_3[442], stage0_3[443], stage0_3[444], stage0_3[445]},
      {stage0_4[206]},
      {stage0_5[192], stage0_5[193], stage0_5[194], stage0_5[195], stage0_5[196], stage0_5[197]},
      {stage1_7[32],stage1_6[61],stage1_5[103],stage1_4[177],stage1_3[190]}
   );
   gpc615_5 gpc191 (
      {stage0_3[446], stage0_3[447], stage0_3[448], stage0_3[449], stage0_3[450]},
      {stage0_4[207]},
      {stage0_5[198], stage0_5[199], stage0_5[200], stage0_5[201], stage0_5[202], stage0_5[203]},
      {stage1_7[33],stage1_6[62],stage1_5[104],stage1_4[178],stage1_3[191]}
   );
   gpc615_5 gpc192 (
      {stage0_3[451], stage0_3[452], stage0_3[453], stage0_3[454], stage0_3[455]},
      {stage0_4[208]},
      {stage0_5[204], stage0_5[205], stage0_5[206], stage0_5[207], stage0_5[208], stage0_5[209]},
      {stage1_7[34],stage1_6[63],stage1_5[105],stage1_4[179],stage1_3[192]}
   );
   gpc615_5 gpc193 (
      {stage0_3[456], stage0_3[457], stage0_3[458], stage0_3[459], stage0_3[460]},
      {stage0_4[209]},
      {stage0_5[210], stage0_5[211], stage0_5[212], stage0_5[213], stage0_5[214], stage0_5[215]},
      {stage1_7[35],stage1_6[64],stage1_5[106],stage1_4[180],stage1_3[193]}
   );
   gpc615_5 gpc194 (
      {stage0_3[461], stage0_3[462], stage0_3[463], stage0_3[464], stage0_3[465]},
      {stage0_4[210]},
      {stage0_5[216], stage0_5[217], stage0_5[218], stage0_5[219], stage0_5[220], stage0_5[221]},
      {stage1_7[36],stage1_6[65],stage1_5[107],stage1_4[181],stage1_3[194]}
   );
   gpc606_5 gpc195 (
      {stage0_4[211], stage0_4[212], stage0_4[213], stage0_4[214], stage0_4[215], stage0_4[216]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[37],stage1_6[66],stage1_5[108],stage1_4[182]}
   );
   gpc606_5 gpc196 (
      {stage0_4[217], stage0_4[218], stage0_4[219], stage0_4[220], stage0_4[221], stage0_4[222]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[38],stage1_6[67],stage1_5[109],stage1_4[183]}
   );
   gpc606_5 gpc197 (
      {stage0_4[223], stage0_4[224], stage0_4[225], stage0_4[226], stage0_4[227], stage0_4[228]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[39],stage1_6[68],stage1_5[110],stage1_4[184]}
   );
   gpc606_5 gpc198 (
      {stage0_4[229], stage0_4[230], stage0_4[231], stage0_4[232], stage0_4[233], stage0_4[234]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[40],stage1_6[69],stage1_5[111],stage1_4[185]}
   );
   gpc606_5 gpc199 (
      {stage0_4[235], stage0_4[236], stage0_4[237], stage0_4[238], stage0_4[239], stage0_4[240]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[41],stage1_6[70],stage1_5[112],stage1_4[186]}
   );
   gpc606_5 gpc200 (
      {stage0_4[241], stage0_4[242], stage0_4[243], stage0_4[244], stage0_4[245], stage0_4[246]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[42],stage1_6[71],stage1_5[113],stage1_4[187]}
   );
   gpc606_5 gpc201 (
      {stage0_4[247], stage0_4[248], stage0_4[249], stage0_4[250], stage0_4[251], stage0_4[252]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[43],stage1_6[72],stage1_5[114],stage1_4[188]}
   );
   gpc606_5 gpc202 (
      {stage0_4[253], stage0_4[254], stage0_4[255], stage0_4[256], stage0_4[257], stage0_4[258]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[44],stage1_6[73],stage1_5[115],stage1_4[189]}
   );
   gpc606_5 gpc203 (
      {stage0_4[259], stage0_4[260], stage0_4[261], stage0_4[262], stage0_4[263], stage0_4[264]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[45],stage1_6[74],stage1_5[116],stage1_4[190]}
   );
   gpc606_5 gpc204 (
      {stage0_4[265], stage0_4[266], stage0_4[267], stage0_4[268], stage0_4[269], stage0_4[270]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[46],stage1_6[75],stage1_5[117],stage1_4[191]}
   );
   gpc606_5 gpc205 (
      {stage0_4[271], stage0_4[272], stage0_4[273], stage0_4[274], stage0_4[275], stage0_4[276]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[47],stage1_6[76],stage1_5[118],stage1_4[192]}
   );
   gpc606_5 gpc206 (
      {stage0_4[277], stage0_4[278], stage0_4[279], stage0_4[280], stage0_4[281], stage0_4[282]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[48],stage1_6[77],stage1_5[119],stage1_4[193]}
   );
   gpc606_5 gpc207 (
      {stage0_4[283], stage0_4[284], stage0_4[285], stage0_4[286], stage0_4[287], stage0_4[288]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[49],stage1_6[78],stage1_5[120],stage1_4[194]}
   );
   gpc606_5 gpc208 (
      {stage0_4[289], stage0_4[290], stage0_4[291], stage0_4[292], stage0_4[293], stage0_4[294]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[50],stage1_6[79],stage1_5[121],stage1_4[195]}
   );
   gpc606_5 gpc209 (
      {stage0_4[295], stage0_4[296], stage0_4[297], stage0_4[298], stage0_4[299], stage0_4[300]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[51],stage1_6[80],stage1_5[122],stage1_4[196]}
   );
   gpc606_5 gpc210 (
      {stage0_4[301], stage0_4[302], stage0_4[303], stage0_4[304], stage0_4[305], stage0_4[306]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[52],stage1_6[81],stage1_5[123],stage1_4[197]}
   );
   gpc606_5 gpc211 (
      {stage0_4[307], stage0_4[308], stage0_4[309], stage0_4[310], stage0_4[311], stage0_4[312]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[53],stage1_6[82],stage1_5[124],stage1_4[198]}
   );
   gpc606_5 gpc212 (
      {stage0_4[313], stage0_4[314], stage0_4[315], stage0_4[316], stage0_4[317], stage0_4[318]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[54],stage1_6[83],stage1_5[125],stage1_4[199]}
   );
   gpc606_5 gpc213 (
      {stage0_4[319], stage0_4[320], stage0_4[321], stage0_4[322], stage0_4[323], stage0_4[324]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[55],stage1_6[84],stage1_5[126],stage1_4[200]}
   );
   gpc606_5 gpc214 (
      {stage0_4[325], stage0_4[326], stage0_4[327], stage0_4[328], stage0_4[329], stage0_4[330]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[56],stage1_6[85],stage1_5[127],stage1_4[201]}
   );
   gpc606_5 gpc215 (
      {stage0_4[331], stage0_4[332], stage0_4[333], stage0_4[334], stage0_4[335], stage0_4[336]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[57],stage1_6[86],stage1_5[128],stage1_4[202]}
   );
   gpc606_5 gpc216 (
      {stage0_4[337], stage0_4[338], stage0_4[339], stage0_4[340], stage0_4[341], stage0_4[342]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[21],stage1_7[58],stage1_6[87],stage1_5[129],stage1_4[203]}
   );
   gpc606_5 gpc217 (
      {stage0_4[343], stage0_4[344], stage0_4[345], stage0_4[346], stage0_4[347], stage0_4[348]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[22],stage1_7[59],stage1_6[88],stage1_5[130],stage1_4[204]}
   );
   gpc606_5 gpc218 (
      {stage0_4[349], stage0_4[350], stage0_4[351], stage0_4[352], stage0_4[353], stage0_4[354]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[23],stage1_7[60],stage1_6[89],stage1_5[131],stage1_4[205]}
   );
   gpc606_5 gpc219 (
      {stage0_4[355], stage0_4[356], stage0_4[357], stage0_4[358], stage0_4[359], stage0_4[360]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[24],stage1_7[61],stage1_6[90],stage1_5[132],stage1_4[206]}
   );
   gpc606_5 gpc220 (
      {stage0_4[361], stage0_4[362], stage0_4[363], stage0_4[364], stage0_4[365], stage0_4[366]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[25],stage1_7[62],stage1_6[91],stage1_5[133],stage1_4[207]}
   );
   gpc606_5 gpc221 (
      {stage0_4[367], stage0_4[368], stage0_4[369], stage0_4[370], stage0_4[371], stage0_4[372]},
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage1_8[26],stage1_7[63],stage1_6[92],stage1_5[134],stage1_4[208]}
   );
   gpc606_5 gpc222 (
      {stage0_4[373], stage0_4[374], stage0_4[375], stage0_4[376], stage0_4[377], stage0_4[378]},
      {stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167]},
      {stage1_8[27],stage1_7[64],stage1_6[93],stage1_5[135],stage1_4[209]}
   );
   gpc606_5 gpc223 (
      {stage0_4[379], stage0_4[380], stage0_4[381], stage0_4[382], stage0_4[383], stage0_4[384]},
      {stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173]},
      {stage1_8[28],stage1_7[65],stage1_6[94],stage1_5[136],stage1_4[210]}
   );
   gpc606_5 gpc224 (
      {stage0_4[385], stage0_4[386], stage0_4[387], stage0_4[388], stage0_4[389], stage0_4[390]},
      {stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179]},
      {stage1_8[29],stage1_7[66],stage1_6[95],stage1_5[137],stage1_4[211]}
   );
   gpc606_5 gpc225 (
      {stage0_4[391], stage0_4[392], stage0_4[393], stage0_4[394], stage0_4[395], stage0_4[396]},
      {stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184], stage0_6[185]},
      {stage1_8[30],stage1_7[67],stage1_6[96],stage1_5[138],stage1_4[212]}
   );
   gpc606_5 gpc226 (
      {stage0_4[397], stage0_4[398], stage0_4[399], stage0_4[400], stage0_4[401], stage0_4[402]},
      {stage0_6[186], stage0_6[187], stage0_6[188], stage0_6[189], stage0_6[190], stage0_6[191]},
      {stage1_8[31],stage1_7[68],stage1_6[97],stage1_5[139],stage1_4[213]}
   );
   gpc606_5 gpc227 (
      {stage0_4[403], stage0_4[404], stage0_4[405], stage0_4[406], stage0_4[407], stage0_4[408]},
      {stage0_6[192], stage0_6[193], stage0_6[194], stage0_6[195], stage0_6[196], stage0_6[197]},
      {stage1_8[32],stage1_7[69],stage1_6[98],stage1_5[140],stage1_4[214]}
   );
   gpc606_5 gpc228 (
      {stage0_4[409], stage0_4[410], stage0_4[411], stage0_4[412], stage0_4[413], stage0_4[414]},
      {stage0_6[198], stage0_6[199], stage0_6[200], stage0_6[201], stage0_6[202], stage0_6[203]},
      {stage1_8[33],stage1_7[70],stage1_6[99],stage1_5[141],stage1_4[215]}
   );
   gpc606_5 gpc229 (
      {stage0_4[415], stage0_4[416], stage0_4[417], stage0_4[418], stage0_4[419], stage0_4[420]},
      {stage0_6[204], stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208], stage0_6[209]},
      {stage1_8[34],stage1_7[71],stage1_6[100],stage1_5[142],stage1_4[216]}
   );
   gpc606_5 gpc230 (
      {stage0_4[421], stage0_4[422], stage0_4[423], stage0_4[424], stage0_4[425], stage0_4[426]},
      {stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214], stage0_6[215]},
      {stage1_8[35],stage1_7[72],stage1_6[101],stage1_5[143],stage1_4[217]}
   );
   gpc606_5 gpc231 (
      {stage0_4[427], stage0_4[428], stage0_4[429], stage0_4[430], stage0_4[431], stage0_4[432]},
      {stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219], stage0_6[220], stage0_6[221]},
      {stage1_8[36],stage1_7[73],stage1_6[102],stage1_5[144],stage1_4[218]}
   );
   gpc606_5 gpc232 (
      {stage0_4[433], stage0_4[434], stage0_4[435], stage0_4[436], stage0_4[437], stage0_4[438]},
      {stage0_6[222], stage0_6[223], stage0_6[224], stage0_6[225], stage0_6[226], stage0_6[227]},
      {stage1_8[37],stage1_7[74],stage1_6[103],stage1_5[145],stage1_4[219]}
   );
   gpc606_5 gpc233 (
      {stage0_4[439], stage0_4[440], stage0_4[441], stage0_4[442], stage0_4[443], stage0_4[444]},
      {stage0_6[228], stage0_6[229], stage0_6[230], stage0_6[231], stage0_6[232], stage0_6[233]},
      {stage1_8[38],stage1_7[75],stage1_6[104],stage1_5[146],stage1_4[220]}
   );
   gpc606_5 gpc234 (
      {stage0_4[445], stage0_4[446], stage0_4[447], stage0_4[448], stage0_4[449], stage0_4[450]},
      {stage0_6[234], stage0_6[235], stage0_6[236], stage0_6[237], stage0_6[238], stage0_6[239]},
      {stage1_8[39],stage1_7[76],stage1_6[105],stage1_5[147],stage1_4[221]}
   );
   gpc606_5 gpc235 (
      {stage0_4[451], stage0_4[452], stage0_4[453], stage0_4[454], stage0_4[455], stage0_4[456]},
      {stage0_6[240], stage0_6[241], stage0_6[242], stage0_6[243], stage0_6[244], stage0_6[245]},
      {stage1_8[40],stage1_7[77],stage1_6[106],stage1_5[148],stage1_4[222]}
   );
   gpc606_5 gpc236 (
      {stage0_4[457], stage0_4[458], stage0_4[459], stage0_4[460], stage0_4[461], stage0_4[462]},
      {stage0_6[246], stage0_6[247], stage0_6[248], stage0_6[249], stage0_6[250], stage0_6[251]},
      {stage1_8[41],stage1_7[78],stage1_6[107],stage1_5[149],stage1_4[223]}
   );
   gpc606_5 gpc237 (
      {stage0_4[463], stage0_4[464], stage0_4[465], stage0_4[466], stage0_4[467], stage0_4[468]},
      {stage0_6[252], stage0_6[253], stage0_6[254], stage0_6[255], stage0_6[256], stage0_6[257]},
      {stage1_8[42],stage1_7[79],stage1_6[108],stage1_5[150],stage1_4[224]}
   );
   gpc606_5 gpc238 (
      {stage0_4[469], stage0_4[470], stage0_4[471], stage0_4[472], stage0_4[473], stage0_4[474]},
      {stage0_6[258], stage0_6[259], stage0_6[260], stage0_6[261], stage0_6[262], stage0_6[263]},
      {stage1_8[43],stage1_7[80],stage1_6[109],stage1_5[151],stage1_4[225]}
   );
   gpc606_5 gpc239 (
      {stage0_4[475], stage0_4[476], stage0_4[477], stage0_4[478], stage0_4[479], stage0_4[480]},
      {stage0_6[264], stage0_6[265], stage0_6[266], stage0_6[267], stage0_6[268], stage0_6[269]},
      {stage1_8[44],stage1_7[81],stage1_6[110],stage1_5[152],stage1_4[226]}
   );
   gpc606_5 gpc240 (
      {stage0_4[481], stage0_4[482], stage0_4[483], stage0_4[484], stage0_4[485], 1'b0},
      {stage0_6[270], stage0_6[271], stage0_6[272], stage0_6[273], stage0_6[274], stage0_6[275]},
      {stage1_8[45],stage1_7[82],stage1_6[111],stage1_5[153],stage1_4[227]}
   );
   gpc606_5 gpc241 (
      {stage0_5[222], stage0_5[223], stage0_5[224], stage0_5[225], stage0_5[226], stage0_5[227]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[46],stage1_7[83],stage1_6[112],stage1_5[154]}
   );
   gpc606_5 gpc242 (
      {stage0_5[228], stage0_5[229], stage0_5[230], stage0_5[231], stage0_5[232], stage0_5[233]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[47],stage1_7[84],stage1_6[113],stage1_5[155]}
   );
   gpc606_5 gpc243 (
      {stage0_5[234], stage0_5[235], stage0_5[236], stage0_5[237], stage0_5[238], stage0_5[239]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[48],stage1_7[85],stage1_6[114],stage1_5[156]}
   );
   gpc606_5 gpc244 (
      {stage0_5[240], stage0_5[241], stage0_5[242], stage0_5[243], stage0_5[244], stage0_5[245]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[49],stage1_7[86],stage1_6[115],stage1_5[157]}
   );
   gpc606_5 gpc245 (
      {stage0_5[246], stage0_5[247], stage0_5[248], stage0_5[249], stage0_5[250], stage0_5[251]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[50],stage1_7[87],stage1_6[116],stage1_5[158]}
   );
   gpc606_5 gpc246 (
      {stage0_5[252], stage0_5[253], stage0_5[254], stage0_5[255], stage0_5[256], stage0_5[257]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[51],stage1_7[88],stage1_6[117],stage1_5[159]}
   );
   gpc606_5 gpc247 (
      {stage0_5[258], stage0_5[259], stage0_5[260], stage0_5[261], stage0_5[262], stage0_5[263]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[52],stage1_7[89],stage1_6[118],stage1_5[160]}
   );
   gpc606_5 gpc248 (
      {stage0_5[264], stage0_5[265], stage0_5[266], stage0_5[267], stage0_5[268], stage0_5[269]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[53],stage1_7[90],stage1_6[119],stage1_5[161]}
   );
   gpc606_5 gpc249 (
      {stage0_5[270], stage0_5[271], stage0_5[272], stage0_5[273], stage0_5[274], stage0_5[275]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[54],stage1_7[91],stage1_6[120],stage1_5[162]}
   );
   gpc606_5 gpc250 (
      {stage0_5[276], stage0_5[277], stage0_5[278], stage0_5[279], stage0_5[280], stage0_5[281]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[55],stage1_7[92],stage1_6[121],stage1_5[163]}
   );
   gpc606_5 gpc251 (
      {stage0_5[282], stage0_5[283], stage0_5[284], stage0_5[285], stage0_5[286], stage0_5[287]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[56],stage1_7[93],stage1_6[122],stage1_5[164]}
   );
   gpc606_5 gpc252 (
      {stage0_5[288], stage0_5[289], stage0_5[290], stage0_5[291], stage0_5[292], stage0_5[293]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[57],stage1_7[94],stage1_6[123],stage1_5[165]}
   );
   gpc606_5 gpc253 (
      {stage0_5[294], stage0_5[295], stage0_5[296], stage0_5[297], stage0_5[298], stage0_5[299]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[58],stage1_7[95],stage1_6[124],stage1_5[166]}
   );
   gpc606_5 gpc254 (
      {stage0_5[300], stage0_5[301], stage0_5[302], stage0_5[303], stage0_5[304], stage0_5[305]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[59],stage1_7[96],stage1_6[125],stage1_5[167]}
   );
   gpc606_5 gpc255 (
      {stage0_5[306], stage0_5[307], stage0_5[308], stage0_5[309], stage0_5[310], stage0_5[311]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[60],stage1_7[97],stage1_6[126],stage1_5[168]}
   );
   gpc606_5 gpc256 (
      {stage0_5[312], stage0_5[313], stage0_5[314], stage0_5[315], stage0_5[316], stage0_5[317]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[61],stage1_7[98],stage1_6[127],stage1_5[169]}
   );
   gpc606_5 gpc257 (
      {stage0_5[318], stage0_5[319], stage0_5[320], stage0_5[321], stage0_5[322], stage0_5[323]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[62],stage1_7[99],stage1_6[128],stage1_5[170]}
   );
   gpc606_5 gpc258 (
      {stage0_5[324], stage0_5[325], stage0_5[326], stage0_5[327], stage0_5[328], stage0_5[329]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[63],stage1_7[100],stage1_6[129],stage1_5[171]}
   );
   gpc606_5 gpc259 (
      {stage0_5[330], stage0_5[331], stage0_5[332], stage0_5[333], stage0_5[334], stage0_5[335]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[64],stage1_7[101],stage1_6[130],stage1_5[172]}
   );
   gpc606_5 gpc260 (
      {stage0_5[336], stage0_5[337], stage0_5[338], stage0_5[339], stage0_5[340], stage0_5[341]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[65],stage1_7[102],stage1_6[131],stage1_5[173]}
   );
   gpc606_5 gpc261 (
      {stage0_5[342], stage0_5[343], stage0_5[344], stage0_5[345], stage0_5[346], stage0_5[347]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[66],stage1_7[103],stage1_6[132],stage1_5[174]}
   );
   gpc606_5 gpc262 (
      {stage0_5[348], stage0_5[349], stage0_5[350], stage0_5[351], stage0_5[352], stage0_5[353]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[67],stage1_7[104],stage1_6[133],stage1_5[175]}
   );
   gpc606_5 gpc263 (
      {stage0_5[354], stage0_5[355], stage0_5[356], stage0_5[357], stage0_5[358], stage0_5[359]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[68],stage1_7[105],stage1_6[134],stage1_5[176]}
   );
   gpc606_5 gpc264 (
      {stage0_5[360], stage0_5[361], stage0_5[362], stage0_5[363], stage0_5[364], stage0_5[365]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[69],stage1_7[106],stage1_6[135],stage1_5[177]}
   );
   gpc606_5 gpc265 (
      {stage0_5[366], stage0_5[367], stage0_5[368], stage0_5[369], stage0_5[370], stage0_5[371]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[70],stage1_7[107],stage1_6[136],stage1_5[178]}
   );
   gpc606_5 gpc266 (
      {stage0_5[372], stage0_5[373], stage0_5[374], stage0_5[375], stage0_5[376], stage0_5[377]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[71],stage1_7[108],stage1_6[137],stage1_5[179]}
   );
   gpc606_5 gpc267 (
      {stage0_5[378], stage0_5[379], stage0_5[380], stage0_5[381], stage0_5[382], stage0_5[383]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[72],stage1_7[109],stage1_6[138],stage1_5[180]}
   );
   gpc606_5 gpc268 (
      {stage0_5[384], stage0_5[385], stage0_5[386], stage0_5[387], stage0_5[388], stage0_5[389]},
      {stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167]},
      {stage1_9[27],stage1_8[73],stage1_7[110],stage1_6[139],stage1_5[181]}
   );
   gpc606_5 gpc269 (
      {stage0_5[390], stage0_5[391], stage0_5[392], stage0_5[393], stage0_5[394], stage0_5[395]},
      {stage0_7[168], stage0_7[169], stage0_7[170], stage0_7[171], stage0_7[172], stage0_7[173]},
      {stage1_9[28],stage1_8[74],stage1_7[111],stage1_6[140],stage1_5[182]}
   );
   gpc606_5 gpc270 (
      {stage0_5[396], stage0_5[397], stage0_5[398], stage0_5[399], stage0_5[400], stage0_5[401]},
      {stage0_7[174], stage0_7[175], stage0_7[176], stage0_7[177], stage0_7[178], stage0_7[179]},
      {stage1_9[29],stage1_8[75],stage1_7[112],stage1_6[141],stage1_5[183]}
   );
   gpc606_5 gpc271 (
      {stage0_5[402], stage0_5[403], stage0_5[404], stage0_5[405], stage0_5[406], stage0_5[407]},
      {stage0_7[180], stage0_7[181], stage0_7[182], stage0_7[183], stage0_7[184], stage0_7[185]},
      {stage1_9[30],stage1_8[76],stage1_7[113],stage1_6[142],stage1_5[184]}
   );
   gpc606_5 gpc272 (
      {stage0_5[408], stage0_5[409], stage0_5[410], stage0_5[411], stage0_5[412], stage0_5[413]},
      {stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189], stage0_7[190], stage0_7[191]},
      {stage1_9[31],stage1_8[77],stage1_7[114],stage1_6[143],stage1_5[185]}
   );
   gpc606_5 gpc273 (
      {stage0_5[414], stage0_5[415], stage0_5[416], stage0_5[417], stage0_5[418], stage0_5[419]},
      {stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195], stage0_7[196], stage0_7[197]},
      {stage1_9[32],stage1_8[78],stage1_7[115],stage1_6[144],stage1_5[186]}
   );
   gpc606_5 gpc274 (
      {stage0_5[420], stage0_5[421], stage0_5[422], stage0_5[423], stage0_5[424], stage0_5[425]},
      {stage0_7[198], stage0_7[199], stage0_7[200], stage0_7[201], stage0_7[202], stage0_7[203]},
      {stage1_9[33],stage1_8[79],stage1_7[116],stage1_6[145],stage1_5[187]}
   );
   gpc606_5 gpc275 (
      {stage0_5[426], stage0_5[427], stage0_5[428], stage0_5[429], stage0_5[430], stage0_5[431]},
      {stage0_7[204], stage0_7[205], stage0_7[206], stage0_7[207], stage0_7[208], stage0_7[209]},
      {stage1_9[34],stage1_8[80],stage1_7[117],stage1_6[146],stage1_5[188]}
   );
   gpc606_5 gpc276 (
      {stage0_5[432], stage0_5[433], stage0_5[434], stage0_5[435], stage0_5[436], stage0_5[437]},
      {stage0_7[210], stage0_7[211], stage0_7[212], stage0_7[213], stage0_7[214], stage0_7[215]},
      {stage1_9[35],stage1_8[81],stage1_7[118],stage1_6[147],stage1_5[189]}
   );
   gpc606_5 gpc277 (
      {stage0_5[438], stage0_5[439], stage0_5[440], stage0_5[441], stage0_5[442], stage0_5[443]},
      {stage0_7[216], stage0_7[217], stage0_7[218], stage0_7[219], stage0_7[220], stage0_7[221]},
      {stage1_9[36],stage1_8[82],stage1_7[119],stage1_6[148],stage1_5[190]}
   );
   gpc606_5 gpc278 (
      {stage0_5[444], stage0_5[445], stage0_5[446], stage0_5[447], stage0_5[448], stage0_5[449]},
      {stage0_7[222], stage0_7[223], stage0_7[224], stage0_7[225], stage0_7[226], stage0_7[227]},
      {stage1_9[37],stage1_8[83],stage1_7[120],stage1_6[149],stage1_5[191]}
   );
   gpc606_5 gpc279 (
      {stage0_5[450], stage0_5[451], stage0_5[452], stage0_5[453], stage0_5[454], stage0_5[455]},
      {stage0_7[228], stage0_7[229], stage0_7[230], stage0_7[231], stage0_7[232], stage0_7[233]},
      {stage1_9[38],stage1_8[84],stage1_7[121],stage1_6[150],stage1_5[192]}
   );
   gpc606_5 gpc280 (
      {stage0_5[456], stage0_5[457], stage0_5[458], stage0_5[459], stage0_5[460], stage0_5[461]},
      {stage0_7[234], stage0_7[235], stage0_7[236], stage0_7[237], stage0_7[238], stage0_7[239]},
      {stage1_9[39],stage1_8[85],stage1_7[122],stage1_6[151],stage1_5[193]}
   );
   gpc606_5 gpc281 (
      {stage0_5[462], stage0_5[463], stage0_5[464], stage0_5[465], stage0_5[466], stage0_5[467]},
      {stage0_7[240], stage0_7[241], stage0_7[242], stage0_7[243], stage0_7[244], stage0_7[245]},
      {stage1_9[40],stage1_8[86],stage1_7[123],stage1_6[152],stage1_5[194]}
   );
   gpc606_5 gpc282 (
      {stage0_5[468], stage0_5[469], stage0_5[470], stage0_5[471], stage0_5[472], stage0_5[473]},
      {stage0_7[246], stage0_7[247], stage0_7[248], stage0_7[249], stage0_7[250], stage0_7[251]},
      {stage1_9[41],stage1_8[87],stage1_7[124],stage1_6[153],stage1_5[195]}
   );
   gpc606_5 gpc283 (
      {stage0_5[474], stage0_5[475], stage0_5[476], stage0_5[477], stage0_5[478], stage0_5[479]},
      {stage0_7[252], stage0_7[253], stage0_7[254], stage0_7[255], stage0_7[256], stage0_7[257]},
      {stage1_9[42],stage1_8[88],stage1_7[125],stage1_6[154],stage1_5[196]}
   );
   gpc606_5 gpc284 (
      {stage0_5[480], stage0_5[481], stage0_5[482], stage0_5[483], stage0_5[484], stage0_5[485]},
      {stage0_7[258], stage0_7[259], stage0_7[260], stage0_7[261], stage0_7[262], stage0_7[263]},
      {stage1_9[43],stage1_8[89],stage1_7[126],stage1_6[155],stage1_5[197]}
   );
   gpc615_5 gpc285 (
      {stage0_6[276], stage0_6[277], stage0_6[278], stage0_6[279], stage0_6[280]},
      {stage0_7[264]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[44],stage1_8[90],stage1_7[127],stage1_6[156]}
   );
   gpc615_5 gpc286 (
      {stage0_6[281], stage0_6[282], stage0_6[283], stage0_6[284], stage0_6[285]},
      {stage0_7[265]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[45],stage1_8[91],stage1_7[128],stage1_6[157]}
   );
   gpc615_5 gpc287 (
      {stage0_6[286], stage0_6[287], stage0_6[288], stage0_6[289], stage0_6[290]},
      {stage0_7[266]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[46],stage1_8[92],stage1_7[129],stage1_6[158]}
   );
   gpc615_5 gpc288 (
      {stage0_6[291], stage0_6[292], stage0_6[293], stage0_6[294], stage0_6[295]},
      {stage0_7[267]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[47],stage1_8[93],stage1_7[130],stage1_6[159]}
   );
   gpc615_5 gpc289 (
      {stage0_6[296], stage0_6[297], stage0_6[298], stage0_6[299], stage0_6[300]},
      {stage0_7[268]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[48],stage1_8[94],stage1_7[131],stage1_6[160]}
   );
   gpc615_5 gpc290 (
      {stage0_6[301], stage0_6[302], stage0_6[303], stage0_6[304], stage0_6[305]},
      {stage0_7[269]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[49],stage1_8[95],stage1_7[132],stage1_6[161]}
   );
   gpc615_5 gpc291 (
      {stage0_6[306], stage0_6[307], stage0_6[308], stage0_6[309], stage0_6[310]},
      {stage0_7[270]},
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage1_10[6],stage1_9[50],stage1_8[96],stage1_7[133],stage1_6[162]}
   );
   gpc615_5 gpc292 (
      {stage0_6[311], stage0_6[312], stage0_6[313], stage0_6[314], stage0_6[315]},
      {stage0_7[271]},
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage1_10[7],stage1_9[51],stage1_8[97],stage1_7[134],stage1_6[163]}
   );
   gpc615_5 gpc293 (
      {stage0_6[316], stage0_6[317], stage0_6[318], stage0_6[319], stage0_6[320]},
      {stage0_7[272]},
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage1_10[8],stage1_9[52],stage1_8[98],stage1_7[135],stage1_6[164]}
   );
   gpc615_5 gpc294 (
      {stage0_6[321], stage0_6[322], stage0_6[323], stage0_6[324], stage0_6[325]},
      {stage0_7[273]},
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage1_10[9],stage1_9[53],stage1_8[99],stage1_7[136],stage1_6[165]}
   );
   gpc615_5 gpc295 (
      {stage0_6[326], stage0_6[327], stage0_6[328], stage0_6[329], stage0_6[330]},
      {stage0_7[274]},
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage1_10[10],stage1_9[54],stage1_8[100],stage1_7[137],stage1_6[166]}
   );
   gpc615_5 gpc296 (
      {stage0_6[331], stage0_6[332], stage0_6[333], stage0_6[334], stage0_6[335]},
      {stage0_7[275]},
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage1_10[11],stage1_9[55],stage1_8[101],stage1_7[138],stage1_6[167]}
   );
   gpc615_5 gpc297 (
      {stage0_6[336], stage0_6[337], stage0_6[338], stage0_6[339], stage0_6[340]},
      {stage0_7[276]},
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77]},
      {stage1_10[12],stage1_9[56],stage1_8[102],stage1_7[139],stage1_6[168]}
   );
   gpc615_5 gpc298 (
      {stage0_6[341], stage0_6[342], stage0_6[343], stage0_6[344], stage0_6[345]},
      {stage0_7[277]},
      {stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83]},
      {stage1_10[13],stage1_9[57],stage1_8[103],stage1_7[140],stage1_6[169]}
   );
   gpc615_5 gpc299 (
      {stage0_6[346], stage0_6[347], stage0_6[348], stage0_6[349], stage0_6[350]},
      {stage0_7[278]},
      {stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89]},
      {stage1_10[14],stage1_9[58],stage1_8[104],stage1_7[141],stage1_6[170]}
   );
   gpc615_5 gpc300 (
      {stage0_6[351], stage0_6[352], stage0_6[353], stage0_6[354], stage0_6[355]},
      {stage0_7[279]},
      {stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95]},
      {stage1_10[15],stage1_9[59],stage1_8[105],stage1_7[142],stage1_6[171]}
   );
   gpc615_5 gpc301 (
      {stage0_6[356], stage0_6[357], stage0_6[358], stage0_6[359], stage0_6[360]},
      {stage0_7[280]},
      {stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101]},
      {stage1_10[16],stage1_9[60],stage1_8[106],stage1_7[143],stage1_6[172]}
   );
   gpc615_5 gpc302 (
      {stage0_6[361], stage0_6[362], stage0_6[363], stage0_6[364], stage0_6[365]},
      {stage0_7[281]},
      {stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107]},
      {stage1_10[17],stage1_9[61],stage1_8[107],stage1_7[144],stage1_6[173]}
   );
   gpc615_5 gpc303 (
      {stage0_6[366], stage0_6[367], stage0_6[368], stage0_6[369], stage0_6[370]},
      {stage0_7[282]},
      {stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113]},
      {stage1_10[18],stage1_9[62],stage1_8[108],stage1_7[145],stage1_6[174]}
   );
   gpc615_5 gpc304 (
      {stage0_6[371], stage0_6[372], stage0_6[373], stage0_6[374], stage0_6[375]},
      {stage0_7[283]},
      {stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119]},
      {stage1_10[19],stage1_9[63],stage1_8[109],stage1_7[146],stage1_6[175]}
   );
   gpc615_5 gpc305 (
      {stage0_6[376], stage0_6[377], stage0_6[378], stage0_6[379], stage0_6[380]},
      {stage0_7[284]},
      {stage0_8[120], stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125]},
      {stage1_10[20],stage1_9[64],stage1_8[110],stage1_7[147],stage1_6[176]}
   );
   gpc615_5 gpc306 (
      {stage0_6[381], stage0_6[382], stage0_6[383], stage0_6[384], stage0_6[385]},
      {stage0_7[285]},
      {stage0_8[126], stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131]},
      {stage1_10[21],stage1_9[65],stage1_8[111],stage1_7[148],stage1_6[177]}
   );
   gpc615_5 gpc307 (
      {stage0_6[386], stage0_6[387], stage0_6[388], stage0_6[389], stage0_6[390]},
      {stage0_7[286]},
      {stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137]},
      {stage1_10[22],stage1_9[66],stage1_8[112],stage1_7[149],stage1_6[178]}
   );
   gpc615_5 gpc308 (
      {stage0_6[391], stage0_6[392], stage0_6[393], stage0_6[394], stage0_6[395]},
      {stage0_7[287]},
      {stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143]},
      {stage1_10[23],stage1_9[67],stage1_8[113],stage1_7[150],stage1_6[179]}
   );
   gpc615_5 gpc309 (
      {stage0_6[396], stage0_6[397], stage0_6[398], stage0_6[399], stage0_6[400]},
      {stage0_7[288]},
      {stage0_8[144], stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149]},
      {stage1_10[24],stage1_9[68],stage1_8[114],stage1_7[151],stage1_6[180]}
   );
   gpc615_5 gpc310 (
      {stage0_6[401], stage0_6[402], stage0_6[403], stage0_6[404], stage0_6[405]},
      {stage0_7[289]},
      {stage0_8[150], stage0_8[151], stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155]},
      {stage1_10[25],stage1_9[69],stage1_8[115],stage1_7[152],stage1_6[181]}
   );
   gpc615_5 gpc311 (
      {stage0_6[406], stage0_6[407], stage0_6[408], stage0_6[409], stage0_6[410]},
      {stage0_7[290]},
      {stage0_8[156], stage0_8[157], stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161]},
      {stage1_10[26],stage1_9[70],stage1_8[116],stage1_7[153],stage1_6[182]}
   );
   gpc615_5 gpc312 (
      {stage0_6[411], stage0_6[412], stage0_6[413], stage0_6[414], stage0_6[415]},
      {stage0_7[291]},
      {stage0_8[162], stage0_8[163], stage0_8[164], stage0_8[165], stage0_8[166], stage0_8[167]},
      {stage1_10[27],stage1_9[71],stage1_8[117],stage1_7[154],stage1_6[183]}
   );
   gpc615_5 gpc313 (
      {stage0_6[416], stage0_6[417], stage0_6[418], stage0_6[419], stage0_6[420]},
      {stage0_7[292]},
      {stage0_8[168], stage0_8[169], stage0_8[170], stage0_8[171], stage0_8[172], stage0_8[173]},
      {stage1_10[28],stage1_9[72],stage1_8[118],stage1_7[155],stage1_6[184]}
   );
   gpc615_5 gpc314 (
      {stage0_6[421], stage0_6[422], stage0_6[423], stage0_6[424], stage0_6[425]},
      {stage0_7[293]},
      {stage0_8[174], stage0_8[175], stage0_8[176], stage0_8[177], stage0_8[178], stage0_8[179]},
      {stage1_10[29],stage1_9[73],stage1_8[119],stage1_7[156],stage1_6[185]}
   );
   gpc615_5 gpc315 (
      {stage0_6[426], stage0_6[427], stage0_6[428], stage0_6[429], stage0_6[430]},
      {stage0_7[294]},
      {stage0_8[180], stage0_8[181], stage0_8[182], stage0_8[183], stage0_8[184], stage0_8[185]},
      {stage1_10[30],stage1_9[74],stage1_8[120],stage1_7[157],stage1_6[186]}
   );
   gpc615_5 gpc316 (
      {stage0_6[431], stage0_6[432], stage0_6[433], stage0_6[434], stage0_6[435]},
      {stage0_7[295]},
      {stage0_8[186], stage0_8[187], stage0_8[188], stage0_8[189], stage0_8[190], stage0_8[191]},
      {stage1_10[31],stage1_9[75],stage1_8[121],stage1_7[158],stage1_6[187]}
   );
   gpc615_5 gpc317 (
      {stage0_6[436], stage0_6[437], stage0_6[438], stage0_6[439], stage0_6[440]},
      {stage0_7[296]},
      {stage0_8[192], stage0_8[193], stage0_8[194], stage0_8[195], stage0_8[196], stage0_8[197]},
      {stage1_10[32],stage1_9[76],stage1_8[122],stage1_7[159],stage1_6[188]}
   );
   gpc615_5 gpc318 (
      {stage0_6[441], stage0_6[442], stage0_6[443], stage0_6[444], stage0_6[445]},
      {stage0_7[297]},
      {stage0_8[198], stage0_8[199], stage0_8[200], stage0_8[201], stage0_8[202], stage0_8[203]},
      {stage1_10[33],stage1_9[77],stage1_8[123],stage1_7[160],stage1_6[189]}
   );
   gpc615_5 gpc319 (
      {stage0_6[446], stage0_6[447], stage0_6[448], stage0_6[449], stage0_6[450]},
      {stage0_7[298]},
      {stage0_8[204], stage0_8[205], stage0_8[206], stage0_8[207], stage0_8[208], stage0_8[209]},
      {stage1_10[34],stage1_9[78],stage1_8[124],stage1_7[161],stage1_6[190]}
   );
   gpc615_5 gpc320 (
      {stage0_6[451], stage0_6[452], stage0_6[453], stage0_6[454], stage0_6[455]},
      {stage0_7[299]},
      {stage0_8[210], stage0_8[211], stage0_8[212], stage0_8[213], stage0_8[214], stage0_8[215]},
      {stage1_10[35],stage1_9[79],stage1_8[125],stage1_7[162],stage1_6[191]}
   );
   gpc615_5 gpc321 (
      {stage0_6[456], stage0_6[457], stage0_6[458], stage0_6[459], stage0_6[460]},
      {stage0_7[300]},
      {stage0_8[216], stage0_8[217], stage0_8[218], stage0_8[219], stage0_8[220], stage0_8[221]},
      {stage1_10[36],stage1_9[80],stage1_8[126],stage1_7[163],stage1_6[192]}
   );
   gpc615_5 gpc322 (
      {stage0_6[461], stage0_6[462], stage0_6[463], stage0_6[464], stage0_6[465]},
      {stage0_7[301]},
      {stage0_8[222], stage0_8[223], stage0_8[224], stage0_8[225], stage0_8[226], stage0_8[227]},
      {stage1_10[37],stage1_9[81],stage1_8[127],stage1_7[164],stage1_6[193]}
   );
   gpc615_5 gpc323 (
      {stage0_7[302], stage0_7[303], stage0_7[304], stage0_7[305], stage0_7[306]},
      {stage0_8[228]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[38],stage1_9[82],stage1_8[128],stage1_7[165]}
   );
   gpc615_5 gpc324 (
      {stage0_7[307], stage0_7[308], stage0_7[309], stage0_7[310], stage0_7[311]},
      {stage0_8[229]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[39],stage1_9[83],stage1_8[129],stage1_7[166]}
   );
   gpc615_5 gpc325 (
      {stage0_7[312], stage0_7[313], stage0_7[314], stage0_7[315], stage0_7[316]},
      {stage0_8[230]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[40],stage1_9[84],stage1_8[130],stage1_7[167]}
   );
   gpc615_5 gpc326 (
      {stage0_7[317], stage0_7[318], stage0_7[319], stage0_7[320], stage0_7[321]},
      {stage0_8[231]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[41],stage1_9[85],stage1_8[131],stage1_7[168]}
   );
   gpc615_5 gpc327 (
      {stage0_7[322], stage0_7[323], stage0_7[324], stage0_7[325], stage0_7[326]},
      {stage0_8[232]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[42],stage1_9[86],stage1_8[132],stage1_7[169]}
   );
   gpc615_5 gpc328 (
      {stage0_7[327], stage0_7[328], stage0_7[329], stage0_7[330], stage0_7[331]},
      {stage0_8[233]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[43],stage1_9[87],stage1_8[133],stage1_7[170]}
   );
   gpc615_5 gpc329 (
      {stage0_7[332], stage0_7[333], stage0_7[334], stage0_7[335], stage0_7[336]},
      {stage0_8[234]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[44],stage1_9[88],stage1_8[134],stage1_7[171]}
   );
   gpc615_5 gpc330 (
      {stage0_7[337], stage0_7[338], stage0_7[339], stage0_7[340], stage0_7[341]},
      {stage0_8[235]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[45],stage1_9[89],stage1_8[135],stage1_7[172]}
   );
   gpc615_5 gpc331 (
      {stage0_7[342], stage0_7[343], stage0_7[344], stage0_7[345], stage0_7[346]},
      {stage0_8[236]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[46],stage1_9[90],stage1_8[136],stage1_7[173]}
   );
   gpc615_5 gpc332 (
      {stage0_7[347], stage0_7[348], stage0_7[349], stage0_7[350], stage0_7[351]},
      {stage0_8[237]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[47],stage1_9[91],stage1_8[137],stage1_7[174]}
   );
   gpc615_5 gpc333 (
      {stage0_7[352], stage0_7[353], stage0_7[354], stage0_7[355], stage0_7[356]},
      {stage0_8[238]},
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage1_11[10],stage1_10[48],stage1_9[92],stage1_8[138],stage1_7[175]}
   );
   gpc615_5 gpc334 (
      {stage0_7[357], stage0_7[358], stage0_7[359], stage0_7[360], stage0_7[361]},
      {stage0_8[239]},
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage1_11[11],stage1_10[49],stage1_9[93],stage1_8[139],stage1_7[176]}
   );
   gpc615_5 gpc335 (
      {stage0_7[362], stage0_7[363], stage0_7[364], stage0_7[365], stage0_7[366]},
      {stage0_8[240]},
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage1_11[12],stage1_10[50],stage1_9[94],stage1_8[140],stage1_7[177]}
   );
   gpc615_5 gpc336 (
      {stage0_7[367], stage0_7[368], stage0_7[369], stage0_7[370], stage0_7[371]},
      {stage0_8[241]},
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage1_11[13],stage1_10[51],stage1_9[95],stage1_8[141],stage1_7[178]}
   );
   gpc615_5 gpc337 (
      {stage0_7[372], stage0_7[373], stage0_7[374], stage0_7[375], stage0_7[376]},
      {stage0_8[242]},
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage1_11[14],stage1_10[52],stage1_9[96],stage1_8[142],stage1_7[179]}
   );
   gpc615_5 gpc338 (
      {stage0_7[377], stage0_7[378], stage0_7[379], stage0_7[380], stage0_7[381]},
      {stage0_8[243]},
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage1_11[15],stage1_10[53],stage1_9[97],stage1_8[143],stage1_7[180]}
   );
   gpc615_5 gpc339 (
      {stage0_7[382], stage0_7[383], stage0_7[384], stage0_7[385], stage0_7[386]},
      {stage0_8[244]},
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage1_11[16],stage1_10[54],stage1_9[98],stage1_8[144],stage1_7[181]}
   );
   gpc615_5 gpc340 (
      {stage0_7[387], stage0_7[388], stage0_7[389], stage0_7[390], stage0_7[391]},
      {stage0_8[245]},
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage1_11[17],stage1_10[55],stage1_9[99],stage1_8[145],stage1_7[182]}
   );
   gpc615_5 gpc341 (
      {stage0_7[392], stage0_7[393], stage0_7[394], stage0_7[395], stage0_7[396]},
      {stage0_8[246]},
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage1_11[18],stage1_10[56],stage1_9[100],stage1_8[146],stage1_7[183]}
   );
   gpc615_5 gpc342 (
      {stage0_7[397], stage0_7[398], stage0_7[399], stage0_7[400], stage0_7[401]},
      {stage0_8[247]},
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage1_11[19],stage1_10[57],stage1_9[101],stage1_8[147],stage1_7[184]}
   );
   gpc615_5 gpc343 (
      {stage0_7[402], stage0_7[403], stage0_7[404], stage0_7[405], stage0_7[406]},
      {stage0_8[248]},
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage1_11[20],stage1_10[58],stage1_9[102],stage1_8[148],stage1_7[185]}
   );
   gpc615_5 gpc344 (
      {stage0_7[407], stage0_7[408], stage0_7[409], stage0_7[410], stage0_7[411]},
      {stage0_8[249]},
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage1_11[21],stage1_10[59],stage1_9[103],stage1_8[149],stage1_7[186]}
   );
   gpc615_5 gpc345 (
      {stage0_7[412], stage0_7[413], stage0_7[414], stage0_7[415], stage0_7[416]},
      {stage0_8[250]},
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage1_11[22],stage1_10[60],stage1_9[104],stage1_8[150],stage1_7[187]}
   );
   gpc615_5 gpc346 (
      {stage0_7[417], stage0_7[418], stage0_7[419], stage0_7[420], stage0_7[421]},
      {stage0_8[251]},
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage1_11[23],stage1_10[61],stage1_9[105],stage1_8[151],stage1_7[188]}
   );
   gpc615_5 gpc347 (
      {stage0_7[422], stage0_7[423], stage0_7[424], stage0_7[425], stage0_7[426]},
      {stage0_8[252]},
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149]},
      {stage1_11[24],stage1_10[62],stage1_9[106],stage1_8[152],stage1_7[189]}
   );
   gpc615_5 gpc348 (
      {stage0_7[427], stage0_7[428], stage0_7[429], stage0_7[430], stage0_7[431]},
      {stage0_8[253]},
      {stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage1_11[25],stage1_10[63],stage1_9[107],stage1_8[153],stage1_7[190]}
   );
   gpc615_5 gpc349 (
      {stage0_7[432], stage0_7[433], stage0_7[434], stage0_7[435], stage0_7[436]},
      {stage0_8[254]},
      {stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160], stage0_9[161]},
      {stage1_11[26],stage1_10[64],stage1_9[108],stage1_8[154],stage1_7[191]}
   );
   gpc615_5 gpc350 (
      {stage0_7[437], stage0_7[438], stage0_7[439], stage0_7[440], stage0_7[441]},
      {stage0_8[255]},
      {stage0_9[162], stage0_9[163], stage0_9[164], stage0_9[165], stage0_9[166], stage0_9[167]},
      {stage1_11[27],stage1_10[65],stage1_9[109],stage1_8[155],stage1_7[192]}
   );
   gpc615_5 gpc351 (
      {stage0_7[442], stage0_7[443], stage0_7[444], stage0_7[445], stage0_7[446]},
      {stage0_8[256]},
      {stage0_9[168], stage0_9[169], stage0_9[170], stage0_9[171], stage0_9[172], stage0_9[173]},
      {stage1_11[28],stage1_10[66],stage1_9[110],stage1_8[156],stage1_7[193]}
   );
   gpc615_5 gpc352 (
      {stage0_7[447], stage0_7[448], stage0_7[449], stage0_7[450], stage0_7[451]},
      {stage0_8[257]},
      {stage0_9[174], stage0_9[175], stage0_9[176], stage0_9[177], stage0_9[178], stage0_9[179]},
      {stage1_11[29],stage1_10[67],stage1_9[111],stage1_8[157],stage1_7[194]}
   );
   gpc615_5 gpc353 (
      {stage0_7[452], stage0_7[453], stage0_7[454], stage0_7[455], stage0_7[456]},
      {stage0_8[258]},
      {stage0_9[180], stage0_9[181], stage0_9[182], stage0_9[183], stage0_9[184], stage0_9[185]},
      {stage1_11[30],stage1_10[68],stage1_9[112],stage1_8[158],stage1_7[195]}
   );
   gpc615_5 gpc354 (
      {stage0_7[457], stage0_7[458], stage0_7[459], stage0_7[460], stage0_7[461]},
      {stage0_8[259]},
      {stage0_9[186], stage0_9[187], stage0_9[188], stage0_9[189], stage0_9[190], stage0_9[191]},
      {stage1_11[31],stage1_10[69],stage1_9[113],stage1_8[159],stage1_7[196]}
   );
   gpc606_5 gpc355 (
      {stage0_8[260], stage0_8[261], stage0_8[262], stage0_8[263], stage0_8[264], stage0_8[265]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[32],stage1_10[70],stage1_9[114],stage1_8[160]}
   );
   gpc606_5 gpc356 (
      {stage0_8[266], stage0_8[267], stage0_8[268], stage0_8[269], stage0_8[270], stage0_8[271]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[33],stage1_10[71],stage1_9[115],stage1_8[161]}
   );
   gpc606_5 gpc357 (
      {stage0_8[272], stage0_8[273], stage0_8[274], stage0_8[275], stage0_8[276], stage0_8[277]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[34],stage1_10[72],stage1_9[116],stage1_8[162]}
   );
   gpc606_5 gpc358 (
      {stage0_8[278], stage0_8[279], stage0_8[280], stage0_8[281], stage0_8[282], stage0_8[283]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[35],stage1_10[73],stage1_9[117],stage1_8[163]}
   );
   gpc606_5 gpc359 (
      {stage0_8[284], stage0_8[285], stage0_8[286], stage0_8[287], stage0_8[288], stage0_8[289]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[36],stage1_10[74],stage1_9[118],stage1_8[164]}
   );
   gpc606_5 gpc360 (
      {stage0_8[290], stage0_8[291], stage0_8[292], stage0_8[293], stage0_8[294], stage0_8[295]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[37],stage1_10[75],stage1_9[119],stage1_8[165]}
   );
   gpc606_5 gpc361 (
      {stage0_8[296], stage0_8[297], stage0_8[298], stage0_8[299], stage0_8[300], stage0_8[301]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[38],stage1_10[76],stage1_9[120],stage1_8[166]}
   );
   gpc606_5 gpc362 (
      {stage0_8[302], stage0_8[303], stage0_8[304], stage0_8[305], stage0_8[306], stage0_8[307]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[39],stage1_10[77],stage1_9[121],stage1_8[167]}
   );
   gpc606_5 gpc363 (
      {stage0_8[308], stage0_8[309], stage0_8[310], stage0_8[311], stage0_8[312], stage0_8[313]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[40],stage1_10[78],stage1_9[122],stage1_8[168]}
   );
   gpc606_5 gpc364 (
      {stage0_8[314], stage0_8[315], stage0_8[316], stage0_8[317], stage0_8[318], stage0_8[319]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[41],stage1_10[79],stage1_9[123],stage1_8[169]}
   );
   gpc606_5 gpc365 (
      {stage0_8[320], stage0_8[321], stage0_8[322], stage0_8[323], stage0_8[324], stage0_8[325]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[42],stage1_10[80],stage1_9[124],stage1_8[170]}
   );
   gpc606_5 gpc366 (
      {stage0_8[326], stage0_8[327], stage0_8[328], stage0_8[329], stage0_8[330], stage0_8[331]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[43],stage1_10[81],stage1_9[125],stage1_8[171]}
   );
   gpc606_5 gpc367 (
      {stage0_8[332], stage0_8[333], stage0_8[334], stage0_8[335], stage0_8[336], stage0_8[337]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[44],stage1_10[82],stage1_9[126],stage1_8[172]}
   );
   gpc606_5 gpc368 (
      {stage0_8[338], stage0_8[339], stage0_8[340], stage0_8[341], stage0_8[342], stage0_8[343]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[45],stage1_10[83],stage1_9[127],stage1_8[173]}
   );
   gpc606_5 gpc369 (
      {stage0_8[344], stage0_8[345], stage0_8[346], stage0_8[347], stage0_8[348], stage0_8[349]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[46],stage1_10[84],stage1_9[128],stage1_8[174]}
   );
   gpc606_5 gpc370 (
      {stage0_8[350], stage0_8[351], stage0_8[352], stage0_8[353], stage0_8[354], stage0_8[355]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[47],stage1_10[85],stage1_9[129],stage1_8[175]}
   );
   gpc606_5 gpc371 (
      {stage0_8[356], stage0_8[357], stage0_8[358], stage0_8[359], stage0_8[360], stage0_8[361]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[48],stage1_10[86],stage1_9[130],stage1_8[176]}
   );
   gpc606_5 gpc372 (
      {stage0_8[362], stage0_8[363], stage0_8[364], stage0_8[365], stage0_8[366], stage0_8[367]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[49],stage1_10[87],stage1_9[131],stage1_8[177]}
   );
   gpc606_5 gpc373 (
      {stage0_8[368], stage0_8[369], stage0_8[370], stage0_8[371], stage0_8[372], stage0_8[373]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[50],stage1_10[88],stage1_9[132],stage1_8[178]}
   );
   gpc606_5 gpc374 (
      {stage0_8[374], stage0_8[375], stage0_8[376], stage0_8[377], stage0_8[378], stage0_8[379]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[51],stage1_10[89],stage1_9[133],stage1_8[179]}
   );
   gpc606_5 gpc375 (
      {stage0_8[380], stage0_8[381], stage0_8[382], stage0_8[383], stage0_8[384], stage0_8[385]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[52],stage1_10[90],stage1_9[134],stage1_8[180]}
   );
   gpc606_5 gpc376 (
      {stage0_8[386], stage0_8[387], stage0_8[388], stage0_8[389], stage0_8[390], stage0_8[391]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[53],stage1_10[91],stage1_9[135],stage1_8[181]}
   );
   gpc606_5 gpc377 (
      {stage0_8[392], stage0_8[393], stage0_8[394], stage0_8[395], stage0_8[396], stage0_8[397]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[54],stage1_10[92],stage1_9[136],stage1_8[182]}
   );
   gpc606_5 gpc378 (
      {stage0_8[398], stage0_8[399], stage0_8[400], stage0_8[401], stage0_8[402], stage0_8[403]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[55],stage1_10[93],stage1_9[137],stage1_8[183]}
   );
   gpc606_5 gpc379 (
      {stage0_8[404], stage0_8[405], stage0_8[406], stage0_8[407], stage0_8[408], stage0_8[409]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[56],stage1_10[94],stage1_9[138],stage1_8[184]}
   );
   gpc606_5 gpc380 (
      {stage0_8[410], stage0_8[411], stage0_8[412], stage0_8[413], stage0_8[414], stage0_8[415]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[57],stage1_10[95],stage1_9[139],stage1_8[185]}
   );
   gpc606_5 gpc381 (
      {stage0_8[416], stage0_8[417], stage0_8[418], stage0_8[419], stage0_8[420], stage0_8[421]},
      {stage0_10[156], stage0_10[157], stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161]},
      {stage1_12[26],stage1_11[58],stage1_10[96],stage1_9[140],stage1_8[186]}
   );
   gpc606_5 gpc382 (
      {stage0_8[422], stage0_8[423], stage0_8[424], stage0_8[425], stage0_8[426], stage0_8[427]},
      {stage0_10[162], stage0_10[163], stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167]},
      {stage1_12[27],stage1_11[59],stage1_10[97],stage1_9[141],stage1_8[187]}
   );
   gpc606_5 gpc383 (
      {stage0_8[428], stage0_8[429], stage0_8[430], stage0_8[431], stage0_8[432], stage0_8[433]},
      {stage0_10[168], stage0_10[169], stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173]},
      {stage1_12[28],stage1_11[60],stage1_10[98],stage1_9[142],stage1_8[188]}
   );
   gpc606_5 gpc384 (
      {stage0_8[434], stage0_8[435], stage0_8[436], stage0_8[437], stage0_8[438], stage0_8[439]},
      {stage0_10[174], stage0_10[175], stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179]},
      {stage1_12[29],stage1_11[61],stage1_10[99],stage1_9[143],stage1_8[189]}
   );
   gpc606_5 gpc385 (
      {stage0_8[440], stage0_8[441], stage0_8[442], stage0_8[443], stage0_8[444], stage0_8[445]},
      {stage0_10[180], stage0_10[181], stage0_10[182], stage0_10[183], stage0_10[184], stage0_10[185]},
      {stage1_12[30],stage1_11[62],stage1_10[100],stage1_9[144],stage1_8[190]}
   );
   gpc606_5 gpc386 (
      {stage0_8[446], stage0_8[447], stage0_8[448], stage0_8[449], stage0_8[450], stage0_8[451]},
      {stage0_10[186], stage0_10[187], stage0_10[188], stage0_10[189], stage0_10[190], stage0_10[191]},
      {stage1_12[31],stage1_11[63],stage1_10[101],stage1_9[145],stage1_8[191]}
   );
   gpc606_5 gpc387 (
      {stage0_8[452], stage0_8[453], stage0_8[454], stage0_8[455], stage0_8[456], stage0_8[457]},
      {stage0_10[192], stage0_10[193], stage0_10[194], stage0_10[195], stage0_10[196], stage0_10[197]},
      {stage1_12[32],stage1_11[64],stage1_10[102],stage1_9[146],stage1_8[192]}
   );
   gpc606_5 gpc388 (
      {stage0_8[458], stage0_8[459], stage0_8[460], stage0_8[461], stage0_8[462], stage0_8[463]},
      {stage0_10[198], stage0_10[199], stage0_10[200], stage0_10[201], stage0_10[202], stage0_10[203]},
      {stage1_12[33],stage1_11[65],stage1_10[103],stage1_9[147],stage1_8[193]}
   );
   gpc606_5 gpc389 (
      {stage0_8[464], stage0_8[465], stage0_8[466], stage0_8[467], stage0_8[468], stage0_8[469]},
      {stage0_10[204], stage0_10[205], stage0_10[206], stage0_10[207], stage0_10[208], stage0_10[209]},
      {stage1_12[34],stage1_11[66],stage1_10[104],stage1_9[148],stage1_8[194]}
   );
   gpc606_5 gpc390 (
      {stage0_8[470], stage0_8[471], stage0_8[472], stage0_8[473], stage0_8[474], stage0_8[475]},
      {stage0_10[210], stage0_10[211], stage0_10[212], stage0_10[213], stage0_10[214], stage0_10[215]},
      {stage1_12[35],stage1_11[67],stage1_10[105],stage1_9[149],stage1_8[195]}
   );
   gpc606_5 gpc391 (
      {stage0_9[192], stage0_9[193], stage0_9[194], stage0_9[195], stage0_9[196], stage0_9[197]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[36],stage1_11[68],stage1_10[106],stage1_9[150]}
   );
   gpc606_5 gpc392 (
      {stage0_9[198], stage0_9[199], stage0_9[200], stage0_9[201], stage0_9[202], stage0_9[203]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[37],stage1_11[69],stage1_10[107],stage1_9[151]}
   );
   gpc606_5 gpc393 (
      {stage0_9[204], stage0_9[205], stage0_9[206], stage0_9[207], stage0_9[208], stage0_9[209]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[38],stage1_11[70],stage1_10[108],stage1_9[152]}
   );
   gpc606_5 gpc394 (
      {stage0_9[210], stage0_9[211], stage0_9[212], stage0_9[213], stage0_9[214], stage0_9[215]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[39],stage1_11[71],stage1_10[109],stage1_9[153]}
   );
   gpc606_5 gpc395 (
      {stage0_9[216], stage0_9[217], stage0_9[218], stage0_9[219], stage0_9[220], stage0_9[221]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[40],stage1_11[72],stage1_10[110],stage1_9[154]}
   );
   gpc606_5 gpc396 (
      {stage0_9[222], stage0_9[223], stage0_9[224], stage0_9[225], stage0_9[226], stage0_9[227]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[41],stage1_11[73],stage1_10[111],stage1_9[155]}
   );
   gpc606_5 gpc397 (
      {stage0_9[228], stage0_9[229], stage0_9[230], stage0_9[231], stage0_9[232], stage0_9[233]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[42],stage1_11[74],stage1_10[112],stage1_9[156]}
   );
   gpc606_5 gpc398 (
      {stage0_9[234], stage0_9[235], stage0_9[236], stage0_9[237], stage0_9[238], stage0_9[239]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[43],stage1_11[75],stage1_10[113],stage1_9[157]}
   );
   gpc606_5 gpc399 (
      {stage0_9[240], stage0_9[241], stage0_9[242], stage0_9[243], stage0_9[244], stage0_9[245]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[44],stage1_11[76],stage1_10[114],stage1_9[158]}
   );
   gpc606_5 gpc400 (
      {stage0_9[246], stage0_9[247], stage0_9[248], stage0_9[249], stage0_9[250], stage0_9[251]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[45],stage1_11[77],stage1_10[115],stage1_9[159]}
   );
   gpc606_5 gpc401 (
      {stage0_9[252], stage0_9[253], stage0_9[254], stage0_9[255], stage0_9[256], stage0_9[257]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[46],stage1_11[78],stage1_10[116],stage1_9[160]}
   );
   gpc606_5 gpc402 (
      {stage0_9[258], stage0_9[259], stage0_9[260], stage0_9[261], stage0_9[262], stage0_9[263]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[47],stage1_11[79],stage1_10[117],stage1_9[161]}
   );
   gpc606_5 gpc403 (
      {stage0_9[264], stage0_9[265], stage0_9[266], stage0_9[267], stage0_9[268], stage0_9[269]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[48],stage1_11[80],stage1_10[118],stage1_9[162]}
   );
   gpc606_5 gpc404 (
      {stage0_9[270], stage0_9[271], stage0_9[272], stage0_9[273], stage0_9[274], stage0_9[275]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[49],stage1_11[81],stage1_10[119],stage1_9[163]}
   );
   gpc606_5 gpc405 (
      {stage0_9[276], stage0_9[277], stage0_9[278], stage0_9[279], stage0_9[280], stage0_9[281]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[50],stage1_11[82],stage1_10[120],stage1_9[164]}
   );
   gpc606_5 gpc406 (
      {stage0_9[282], stage0_9[283], stage0_9[284], stage0_9[285], stage0_9[286], stage0_9[287]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[51],stage1_11[83],stage1_10[121],stage1_9[165]}
   );
   gpc606_5 gpc407 (
      {stage0_9[288], stage0_9[289], stage0_9[290], stage0_9[291], stage0_9[292], stage0_9[293]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[52],stage1_11[84],stage1_10[122],stage1_9[166]}
   );
   gpc606_5 gpc408 (
      {stage0_9[294], stage0_9[295], stage0_9[296], stage0_9[297], stage0_9[298], stage0_9[299]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[53],stage1_11[85],stage1_10[123],stage1_9[167]}
   );
   gpc606_5 gpc409 (
      {stage0_9[300], stage0_9[301], stage0_9[302], stage0_9[303], stage0_9[304], stage0_9[305]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[54],stage1_11[86],stage1_10[124],stage1_9[168]}
   );
   gpc606_5 gpc410 (
      {stage0_9[306], stage0_9[307], stage0_9[308], stage0_9[309], stage0_9[310], stage0_9[311]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[55],stage1_11[87],stage1_10[125],stage1_9[169]}
   );
   gpc606_5 gpc411 (
      {stage0_9[312], stage0_9[313], stage0_9[314], stage0_9[315], stage0_9[316], stage0_9[317]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[56],stage1_11[88],stage1_10[126],stage1_9[170]}
   );
   gpc606_5 gpc412 (
      {stage0_9[318], stage0_9[319], stage0_9[320], stage0_9[321], stage0_9[322], stage0_9[323]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[57],stage1_11[89],stage1_10[127],stage1_9[171]}
   );
   gpc606_5 gpc413 (
      {stage0_9[324], stage0_9[325], stage0_9[326], stage0_9[327], stage0_9[328], stage0_9[329]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[58],stage1_11[90],stage1_10[128],stage1_9[172]}
   );
   gpc606_5 gpc414 (
      {stage0_9[330], stage0_9[331], stage0_9[332], stage0_9[333], stage0_9[334], stage0_9[335]},
      {stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage1_13[23],stage1_12[59],stage1_11[91],stage1_10[129],stage1_9[173]}
   );
   gpc606_5 gpc415 (
      {stage0_9[336], stage0_9[337], stage0_9[338], stage0_9[339], stage0_9[340], stage0_9[341]},
      {stage0_11[144], stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage1_13[24],stage1_12[60],stage1_11[92],stage1_10[130],stage1_9[174]}
   );
   gpc606_5 gpc416 (
      {stage0_9[342], stage0_9[343], stage0_9[344], stage0_9[345], stage0_9[346], stage0_9[347]},
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154], stage0_11[155]},
      {stage1_13[25],stage1_12[61],stage1_11[93],stage1_10[131],stage1_9[175]}
   );
   gpc606_5 gpc417 (
      {stage0_9[348], stage0_9[349], stage0_9[350], stage0_9[351], stage0_9[352], stage0_9[353]},
      {stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159], stage0_11[160], stage0_11[161]},
      {stage1_13[26],stage1_12[62],stage1_11[94],stage1_10[132],stage1_9[176]}
   );
   gpc606_5 gpc418 (
      {stage0_9[354], stage0_9[355], stage0_9[356], stage0_9[357], stage0_9[358], stage0_9[359]},
      {stage0_11[162], stage0_11[163], stage0_11[164], stage0_11[165], stage0_11[166], stage0_11[167]},
      {stage1_13[27],stage1_12[63],stage1_11[95],stage1_10[133],stage1_9[177]}
   );
   gpc606_5 gpc419 (
      {stage0_9[360], stage0_9[361], stage0_9[362], stage0_9[363], stage0_9[364], stage0_9[365]},
      {stage0_11[168], stage0_11[169], stage0_11[170], stage0_11[171], stage0_11[172], stage0_11[173]},
      {stage1_13[28],stage1_12[64],stage1_11[96],stage1_10[134],stage1_9[178]}
   );
   gpc606_5 gpc420 (
      {stage0_9[366], stage0_9[367], stage0_9[368], stage0_9[369], stage0_9[370], stage0_9[371]},
      {stage0_11[174], stage0_11[175], stage0_11[176], stage0_11[177], stage0_11[178], stage0_11[179]},
      {stage1_13[29],stage1_12[65],stage1_11[97],stage1_10[135],stage1_9[179]}
   );
   gpc606_5 gpc421 (
      {stage0_9[372], stage0_9[373], stage0_9[374], stage0_9[375], stage0_9[376], stage0_9[377]},
      {stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183], stage0_11[184], stage0_11[185]},
      {stage1_13[30],stage1_12[66],stage1_11[98],stage1_10[136],stage1_9[180]}
   );
   gpc606_5 gpc422 (
      {stage0_9[378], stage0_9[379], stage0_9[380], stage0_9[381], stage0_9[382], stage0_9[383]},
      {stage0_11[186], stage0_11[187], stage0_11[188], stage0_11[189], stage0_11[190], stage0_11[191]},
      {stage1_13[31],stage1_12[67],stage1_11[99],stage1_10[137],stage1_9[181]}
   );
   gpc606_5 gpc423 (
      {stage0_9[384], stage0_9[385], stage0_9[386], stage0_9[387], stage0_9[388], stage0_9[389]},
      {stage0_11[192], stage0_11[193], stage0_11[194], stage0_11[195], stage0_11[196], stage0_11[197]},
      {stage1_13[32],stage1_12[68],stage1_11[100],stage1_10[138],stage1_9[182]}
   );
   gpc606_5 gpc424 (
      {stage0_9[390], stage0_9[391], stage0_9[392], stage0_9[393], stage0_9[394], stage0_9[395]},
      {stage0_11[198], stage0_11[199], stage0_11[200], stage0_11[201], stage0_11[202], stage0_11[203]},
      {stage1_13[33],stage1_12[69],stage1_11[101],stage1_10[139],stage1_9[183]}
   );
   gpc606_5 gpc425 (
      {stage0_9[396], stage0_9[397], stage0_9[398], stage0_9[399], stage0_9[400], stage0_9[401]},
      {stage0_11[204], stage0_11[205], stage0_11[206], stage0_11[207], stage0_11[208], stage0_11[209]},
      {stage1_13[34],stage1_12[70],stage1_11[102],stage1_10[140],stage1_9[184]}
   );
   gpc606_5 gpc426 (
      {stage0_9[402], stage0_9[403], stage0_9[404], stage0_9[405], stage0_9[406], stage0_9[407]},
      {stage0_11[210], stage0_11[211], stage0_11[212], stage0_11[213], stage0_11[214], stage0_11[215]},
      {stage1_13[35],stage1_12[71],stage1_11[103],stage1_10[141],stage1_9[185]}
   );
   gpc606_5 gpc427 (
      {stage0_9[408], stage0_9[409], stage0_9[410], stage0_9[411], stage0_9[412], stage0_9[413]},
      {stage0_11[216], stage0_11[217], stage0_11[218], stage0_11[219], stage0_11[220], stage0_11[221]},
      {stage1_13[36],stage1_12[72],stage1_11[104],stage1_10[142],stage1_9[186]}
   );
   gpc606_5 gpc428 (
      {stage0_9[414], stage0_9[415], stage0_9[416], stage0_9[417], stage0_9[418], stage0_9[419]},
      {stage0_11[222], stage0_11[223], stage0_11[224], stage0_11[225], stage0_11[226], stage0_11[227]},
      {stage1_13[37],stage1_12[73],stage1_11[105],stage1_10[143],stage1_9[187]}
   );
   gpc606_5 gpc429 (
      {stage0_9[420], stage0_9[421], stage0_9[422], stage0_9[423], stage0_9[424], stage0_9[425]},
      {stage0_11[228], stage0_11[229], stage0_11[230], stage0_11[231], stage0_11[232], stage0_11[233]},
      {stage1_13[38],stage1_12[74],stage1_11[106],stage1_10[144],stage1_9[188]}
   );
   gpc606_5 gpc430 (
      {stage0_9[426], stage0_9[427], stage0_9[428], stage0_9[429], stage0_9[430], stage0_9[431]},
      {stage0_11[234], stage0_11[235], stage0_11[236], stage0_11[237], stage0_11[238], stage0_11[239]},
      {stage1_13[39],stage1_12[75],stage1_11[107],stage1_10[145],stage1_9[189]}
   );
   gpc606_5 gpc431 (
      {stage0_9[432], stage0_9[433], stage0_9[434], stage0_9[435], stage0_9[436], stage0_9[437]},
      {stage0_11[240], stage0_11[241], stage0_11[242], stage0_11[243], stage0_11[244], stage0_11[245]},
      {stage1_13[40],stage1_12[76],stage1_11[108],stage1_10[146],stage1_9[190]}
   );
   gpc606_5 gpc432 (
      {stage0_9[438], stage0_9[439], stage0_9[440], stage0_9[441], stage0_9[442], stage0_9[443]},
      {stage0_11[246], stage0_11[247], stage0_11[248], stage0_11[249], stage0_11[250], stage0_11[251]},
      {stage1_13[41],stage1_12[77],stage1_11[109],stage1_10[147],stage1_9[191]}
   );
   gpc606_5 gpc433 (
      {stage0_9[444], stage0_9[445], stage0_9[446], stage0_9[447], stage0_9[448], stage0_9[449]},
      {stage0_11[252], stage0_11[253], stage0_11[254], stage0_11[255], stage0_11[256], stage0_11[257]},
      {stage1_13[42],stage1_12[78],stage1_11[110],stage1_10[148],stage1_9[192]}
   );
   gpc606_5 gpc434 (
      {stage0_9[450], stage0_9[451], stage0_9[452], stage0_9[453], stage0_9[454], stage0_9[455]},
      {stage0_11[258], stage0_11[259], stage0_11[260], stage0_11[261], stage0_11[262], stage0_11[263]},
      {stage1_13[43],stage1_12[79],stage1_11[111],stage1_10[149],stage1_9[193]}
   );
   gpc606_5 gpc435 (
      {stage0_9[456], stage0_9[457], stage0_9[458], stage0_9[459], stage0_9[460], stage0_9[461]},
      {stage0_11[264], stage0_11[265], stage0_11[266], stage0_11[267], stage0_11[268], stage0_11[269]},
      {stage1_13[44],stage1_12[80],stage1_11[112],stage1_10[150],stage1_9[194]}
   );
   gpc606_5 gpc436 (
      {stage0_9[462], stage0_9[463], stage0_9[464], stage0_9[465], stage0_9[466], stage0_9[467]},
      {stage0_11[270], stage0_11[271], stage0_11[272], stage0_11[273], stage0_11[274], stage0_11[275]},
      {stage1_13[45],stage1_12[81],stage1_11[113],stage1_10[151],stage1_9[195]}
   );
   gpc2135_5 gpc437 (
      {stage0_10[216], stage0_10[217], stage0_10[218], stage0_10[219], stage0_10[220]},
      {stage0_11[276], stage0_11[277], stage0_11[278]},
      {stage0_12[0]},
      {stage0_13[0], stage0_13[1]},
      {stage1_14[0],stage1_13[46],stage1_12[82],stage1_11[114],stage1_10[152]}
   );
   gpc2135_5 gpc438 (
      {stage0_10[221], stage0_10[222], stage0_10[223], stage0_10[224], stage0_10[225]},
      {stage0_11[279], stage0_11[280], stage0_11[281]},
      {stage0_12[1]},
      {stage0_13[2], stage0_13[3]},
      {stage1_14[1],stage1_13[47],stage1_12[83],stage1_11[115],stage1_10[153]}
   );
   gpc2135_5 gpc439 (
      {stage0_10[226], stage0_10[227], stage0_10[228], stage0_10[229], stage0_10[230]},
      {stage0_11[282], stage0_11[283], stage0_11[284]},
      {stage0_12[2]},
      {stage0_13[4], stage0_13[5]},
      {stage1_14[2],stage1_13[48],stage1_12[84],stage1_11[116],stage1_10[154]}
   );
   gpc2135_5 gpc440 (
      {stage0_10[231], stage0_10[232], stage0_10[233], stage0_10[234], stage0_10[235]},
      {stage0_11[285], stage0_11[286], stage0_11[287]},
      {stage0_12[3]},
      {stage0_13[6], stage0_13[7]},
      {stage1_14[3],stage1_13[49],stage1_12[85],stage1_11[117],stage1_10[155]}
   );
   gpc606_5 gpc441 (
      {stage0_10[236], stage0_10[237], stage0_10[238], stage0_10[239], stage0_10[240], stage0_10[241]},
      {stage0_12[4], stage0_12[5], stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9]},
      {stage1_14[4],stage1_13[50],stage1_12[86],stage1_11[118],stage1_10[156]}
   );
   gpc606_5 gpc442 (
      {stage0_10[242], stage0_10[243], stage0_10[244], stage0_10[245], stage0_10[246], stage0_10[247]},
      {stage0_12[10], stage0_12[11], stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15]},
      {stage1_14[5],stage1_13[51],stage1_12[87],stage1_11[119],stage1_10[157]}
   );
   gpc606_5 gpc443 (
      {stage0_10[248], stage0_10[249], stage0_10[250], stage0_10[251], stage0_10[252], stage0_10[253]},
      {stage0_12[16], stage0_12[17], stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21]},
      {stage1_14[6],stage1_13[52],stage1_12[88],stage1_11[120],stage1_10[158]}
   );
   gpc606_5 gpc444 (
      {stage0_10[254], stage0_10[255], stage0_10[256], stage0_10[257], stage0_10[258], stage0_10[259]},
      {stage0_12[22], stage0_12[23], stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27]},
      {stage1_14[7],stage1_13[53],stage1_12[89],stage1_11[121],stage1_10[159]}
   );
   gpc606_5 gpc445 (
      {stage0_10[260], stage0_10[261], stage0_10[262], stage0_10[263], stage0_10[264], stage0_10[265]},
      {stage0_12[28], stage0_12[29], stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33]},
      {stage1_14[8],stage1_13[54],stage1_12[90],stage1_11[122],stage1_10[160]}
   );
   gpc606_5 gpc446 (
      {stage0_10[266], stage0_10[267], stage0_10[268], stage0_10[269], stage0_10[270], stage0_10[271]},
      {stage0_12[34], stage0_12[35], stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39]},
      {stage1_14[9],stage1_13[55],stage1_12[91],stage1_11[123],stage1_10[161]}
   );
   gpc606_5 gpc447 (
      {stage0_10[272], stage0_10[273], stage0_10[274], stage0_10[275], stage0_10[276], stage0_10[277]},
      {stage0_12[40], stage0_12[41], stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45]},
      {stage1_14[10],stage1_13[56],stage1_12[92],stage1_11[124],stage1_10[162]}
   );
   gpc606_5 gpc448 (
      {stage0_10[278], stage0_10[279], stage0_10[280], stage0_10[281], stage0_10[282], stage0_10[283]},
      {stage0_12[46], stage0_12[47], stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51]},
      {stage1_14[11],stage1_13[57],stage1_12[93],stage1_11[125],stage1_10[163]}
   );
   gpc606_5 gpc449 (
      {stage0_10[284], stage0_10[285], stage0_10[286], stage0_10[287], stage0_10[288], stage0_10[289]},
      {stage0_12[52], stage0_12[53], stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57]},
      {stage1_14[12],stage1_13[58],stage1_12[94],stage1_11[126],stage1_10[164]}
   );
   gpc606_5 gpc450 (
      {stage0_10[290], stage0_10[291], stage0_10[292], stage0_10[293], stage0_10[294], stage0_10[295]},
      {stage0_12[58], stage0_12[59], stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63]},
      {stage1_14[13],stage1_13[59],stage1_12[95],stage1_11[127],stage1_10[165]}
   );
   gpc606_5 gpc451 (
      {stage0_10[296], stage0_10[297], stage0_10[298], stage0_10[299], stage0_10[300], stage0_10[301]},
      {stage0_12[64], stage0_12[65], stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69]},
      {stage1_14[14],stage1_13[60],stage1_12[96],stage1_11[128],stage1_10[166]}
   );
   gpc606_5 gpc452 (
      {stage0_10[302], stage0_10[303], stage0_10[304], stage0_10[305], stage0_10[306], stage0_10[307]},
      {stage0_12[70], stage0_12[71], stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75]},
      {stage1_14[15],stage1_13[61],stage1_12[97],stage1_11[129],stage1_10[167]}
   );
   gpc606_5 gpc453 (
      {stage0_10[308], stage0_10[309], stage0_10[310], stage0_10[311], stage0_10[312], stage0_10[313]},
      {stage0_12[76], stage0_12[77], stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81]},
      {stage1_14[16],stage1_13[62],stage1_12[98],stage1_11[130],stage1_10[168]}
   );
   gpc615_5 gpc454 (
      {stage0_10[314], stage0_10[315], stage0_10[316], stage0_10[317], stage0_10[318]},
      {stage0_11[288]},
      {stage0_12[82], stage0_12[83], stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87]},
      {stage1_14[17],stage1_13[63],stage1_12[99],stage1_11[131],stage1_10[169]}
   );
   gpc615_5 gpc455 (
      {stage0_10[319], stage0_10[320], stage0_10[321], stage0_10[322], stage0_10[323]},
      {stage0_11[289]},
      {stage0_12[88], stage0_12[89], stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93]},
      {stage1_14[18],stage1_13[64],stage1_12[100],stage1_11[132],stage1_10[170]}
   );
   gpc615_5 gpc456 (
      {stage0_10[324], stage0_10[325], stage0_10[326], stage0_10[327], stage0_10[328]},
      {stage0_11[290]},
      {stage0_12[94], stage0_12[95], stage0_12[96], stage0_12[97], stage0_12[98], stage0_12[99]},
      {stage1_14[19],stage1_13[65],stage1_12[101],stage1_11[133],stage1_10[171]}
   );
   gpc615_5 gpc457 (
      {stage0_10[329], stage0_10[330], stage0_10[331], stage0_10[332], stage0_10[333]},
      {stage0_11[291]},
      {stage0_12[100], stage0_12[101], stage0_12[102], stage0_12[103], stage0_12[104], stage0_12[105]},
      {stage1_14[20],stage1_13[66],stage1_12[102],stage1_11[134],stage1_10[172]}
   );
   gpc615_5 gpc458 (
      {stage0_10[334], stage0_10[335], stage0_10[336], stage0_10[337], stage0_10[338]},
      {stage0_11[292]},
      {stage0_12[106], stage0_12[107], stage0_12[108], stage0_12[109], stage0_12[110], stage0_12[111]},
      {stage1_14[21],stage1_13[67],stage1_12[103],stage1_11[135],stage1_10[173]}
   );
   gpc615_5 gpc459 (
      {stage0_10[339], stage0_10[340], stage0_10[341], stage0_10[342], stage0_10[343]},
      {stage0_11[293]},
      {stage0_12[112], stage0_12[113], stage0_12[114], stage0_12[115], stage0_12[116], stage0_12[117]},
      {stage1_14[22],stage1_13[68],stage1_12[104],stage1_11[136],stage1_10[174]}
   );
   gpc615_5 gpc460 (
      {stage0_10[344], stage0_10[345], stage0_10[346], stage0_10[347], stage0_10[348]},
      {stage0_11[294]},
      {stage0_12[118], stage0_12[119], stage0_12[120], stage0_12[121], stage0_12[122], stage0_12[123]},
      {stage1_14[23],stage1_13[69],stage1_12[105],stage1_11[137],stage1_10[175]}
   );
   gpc615_5 gpc461 (
      {stage0_10[349], stage0_10[350], stage0_10[351], stage0_10[352], stage0_10[353]},
      {stage0_11[295]},
      {stage0_12[124], stage0_12[125], stage0_12[126], stage0_12[127], stage0_12[128], stage0_12[129]},
      {stage1_14[24],stage1_13[70],stage1_12[106],stage1_11[138],stage1_10[176]}
   );
   gpc615_5 gpc462 (
      {stage0_10[354], stage0_10[355], stage0_10[356], stage0_10[357], stage0_10[358]},
      {stage0_11[296]},
      {stage0_12[130], stage0_12[131], stage0_12[132], stage0_12[133], stage0_12[134], stage0_12[135]},
      {stage1_14[25],stage1_13[71],stage1_12[107],stage1_11[139],stage1_10[177]}
   );
   gpc615_5 gpc463 (
      {stage0_10[359], stage0_10[360], stage0_10[361], stage0_10[362], stage0_10[363]},
      {stage0_11[297]},
      {stage0_12[136], stage0_12[137], stage0_12[138], stage0_12[139], stage0_12[140], stage0_12[141]},
      {stage1_14[26],stage1_13[72],stage1_12[108],stage1_11[140],stage1_10[178]}
   );
   gpc615_5 gpc464 (
      {stage0_10[364], stage0_10[365], stage0_10[366], stage0_10[367], stage0_10[368]},
      {stage0_11[298]},
      {stage0_12[142], stage0_12[143], stage0_12[144], stage0_12[145], stage0_12[146], stage0_12[147]},
      {stage1_14[27],stage1_13[73],stage1_12[109],stage1_11[141],stage1_10[179]}
   );
   gpc615_5 gpc465 (
      {stage0_10[369], stage0_10[370], stage0_10[371], stage0_10[372], stage0_10[373]},
      {stage0_11[299]},
      {stage0_12[148], stage0_12[149], stage0_12[150], stage0_12[151], stage0_12[152], stage0_12[153]},
      {stage1_14[28],stage1_13[74],stage1_12[110],stage1_11[142],stage1_10[180]}
   );
   gpc615_5 gpc466 (
      {stage0_10[374], stage0_10[375], stage0_10[376], stage0_10[377], stage0_10[378]},
      {stage0_11[300]},
      {stage0_12[154], stage0_12[155], stage0_12[156], stage0_12[157], stage0_12[158], stage0_12[159]},
      {stage1_14[29],stage1_13[75],stage1_12[111],stage1_11[143],stage1_10[181]}
   );
   gpc615_5 gpc467 (
      {stage0_10[379], stage0_10[380], stage0_10[381], stage0_10[382], stage0_10[383]},
      {stage0_11[301]},
      {stage0_12[160], stage0_12[161], stage0_12[162], stage0_12[163], stage0_12[164], stage0_12[165]},
      {stage1_14[30],stage1_13[76],stage1_12[112],stage1_11[144],stage1_10[182]}
   );
   gpc615_5 gpc468 (
      {stage0_11[302], stage0_11[303], stage0_11[304], stage0_11[305], stage0_11[306]},
      {stage0_12[166]},
      {stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11], stage0_13[12], stage0_13[13]},
      {stage1_15[0],stage1_14[31],stage1_13[77],stage1_12[113],stage1_11[145]}
   );
   gpc615_5 gpc469 (
      {stage0_11[307], stage0_11[308], stage0_11[309], stage0_11[310], stage0_11[311]},
      {stage0_12[167]},
      {stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17], stage0_13[18], stage0_13[19]},
      {stage1_15[1],stage1_14[32],stage1_13[78],stage1_12[114],stage1_11[146]}
   );
   gpc615_5 gpc470 (
      {stage0_11[312], stage0_11[313], stage0_11[314], stage0_11[315], stage0_11[316]},
      {stage0_12[168]},
      {stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23], stage0_13[24], stage0_13[25]},
      {stage1_15[2],stage1_14[33],stage1_13[79],stage1_12[115],stage1_11[147]}
   );
   gpc615_5 gpc471 (
      {stage0_11[317], stage0_11[318], stage0_11[319], stage0_11[320], stage0_11[321]},
      {stage0_12[169]},
      {stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29], stage0_13[30], stage0_13[31]},
      {stage1_15[3],stage1_14[34],stage1_13[80],stage1_12[116],stage1_11[148]}
   );
   gpc615_5 gpc472 (
      {stage0_11[322], stage0_11[323], stage0_11[324], stage0_11[325], stage0_11[326]},
      {stage0_12[170]},
      {stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35], stage0_13[36], stage0_13[37]},
      {stage1_15[4],stage1_14[35],stage1_13[81],stage1_12[117],stage1_11[149]}
   );
   gpc615_5 gpc473 (
      {stage0_11[327], stage0_11[328], stage0_11[329], stage0_11[330], stage0_11[331]},
      {stage0_12[171]},
      {stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41], stage0_13[42], stage0_13[43]},
      {stage1_15[5],stage1_14[36],stage1_13[82],stage1_12[118],stage1_11[150]}
   );
   gpc615_5 gpc474 (
      {stage0_11[332], stage0_11[333], stage0_11[334], stage0_11[335], stage0_11[336]},
      {stage0_12[172]},
      {stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47], stage0_13[48], stage0_13[49]},
      {stage1_15[6],stage1_14[37],stage1_13[83],stage1_12[119],stage1_11[151]}
   );
   gpc615_5 gpc475 (
      {stage0_11[337], stage0_11[338], stage0_11[339], stage0_11[340], stage0_11[341]},
      {stage0_12[173]},
      {stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53], stage0_13[54], stage0_13[55]},
      {stage1_15[7],stage1_14[38],stage1_13[84],stage1_12[120],stage1_11[152]}
   );
   gpc615_5 gpc476 (
      {stage0_11[342], stage0_11[343], stage0_11[344], stage0_11[345], stage0_11[346]},
      {stage0_12[174]},
      {stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59], stage0_13[60], stage0_13[61]},
      {stage1_15[8],stage1_14[39],stage1_13[85],stage1_12[121],stage1_11[153]}
   );
   gpc615_5 gpc477 (
      {stage0_11[347], stage0_11[348], stage0_11[349], stage0_11[350], stage0_11[351]},
      {stage0_12[175]},
      {stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65], stage0_13[66], stage0_13[67]},
      {stage1_15[9],stage1_14[40],stage1_13[86],stage1_12[122],stage1_11[154]}
   );
   gpc615_5 gpc478 (
      {stage0_11[352], stage0_11[353], stage0_11[354], stage0_11[355], stage0_11[356]},
      {stage0_12[176]},
      {stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71], stage0_13[72], stage0_13[73]},
      {stage1_15[10],stage1_14[41],stage1_13[87],stage1_12[123],stage1_11[155]}
   );
   gpc615_5 gpc479 (
      {stage0_11[357], stage0_11[358], stage0_11[359], stage0_11[360], stage0_11[361]},
      {stage0_12[177]},
      {stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77], stage0_13[78], stage0_13[79]},
      {stage1_15[11],stage1_14[42],stage1_13[88],stage1_12[124],stage1_11[156]}
   );
   gpc615_5 gpc480 (
      {stage0_11[362], stage0_11[363], stage0_11[364], stage0_11[365], stage0_11[366]},
      {stage0_12[178]},
      {stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83], stage0_13[84], stage0_13[85]},
      {stage1_15[12],stage1_14[43],stage1_13[89],stage1_12[125],stage1_11[157]}
   );
   gpc615_5 gpc481 (
      {stage0_12[179], stage0_12[180], stage0_12[181], stage0_12[182], stage0_12[183]},
      {stage0_13[86]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[13],stage1_14[44],stage1_13[90],stage1_12[126]}
   );
   gpc615_5 gpc482 (
      {stage0_12[184], stage0_12[185], stage0_12[186], stage0_12[187], stage0_12[188]},
      {stage0_13[87]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[14],stage1_14[45],stage1_13[91],stage1_12[127]}
   );
   gpc615_5 gpc483 (
      {stage0_12[189], stage0_12[190], stage0_12[191], stage0_12[192], stage0_12[193]},
      {stage0_13[88]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[15],stage1_14[46],stage1_13[92],stage1_12[128]}
   );
   gpc615_5 gpc484 (
      {stage0_12[194], stage0_12[195], stage0_12[196], stage0_12[197], stage0_12[198]},
      {stage0_13[89]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[16],stage1_14[47],stage1_13[93],stage1_12[129]}
   );
   gpc615_5 gpc485 (
      {stage0_12[199], stage0_12[200], stage0_12[201], stage0_12[202], stage0_12[203]},
      {stage0_13[90]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[17],stage1_14[48],stage1_13[94],stage1_12[130]}
   );
   gpc615_5 gpc486 (
      {stage0_12[204], stage0_12[205], stage0_12[206], stage0_12[207], stage0_12[208]},
      {stage0_13[91]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[18],stage1_14[49],stage1_13[95],stage1_12[131]}
   );
   gpc615_5 gpc487 (
      {stage0_12[209], stage0_12[210], stage0_12[211], stage0_12[212], stage0_12[213]},
      {stage0_13[92]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[19],stage1_14[50],stage1_13[96],stage1_12[132]}
   );
   gpc615_5 gpc488 (
      {stage0_12[214], stage0_12[215], stage0_12[216], stage0_12[217], stage0_12[218]},
      {stage0_13[93]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[20],stage1_14[51],stage1_13[97],stage1_12[133]}
   );
   gpc615_5 gpc489 (
      {stage0_12[219], stage0_12[220], stage0_12[221], stage0_12[222], stage0_12[223]},
      {stage0_13[94]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[21],stage1_14[52],stage1_13[98],stage1_12[134]}
   );
   gpc615_5 gpc490 (
      {stage0_12[224], stage0_12[225], stage0_12[226], stage0_12[227], stage0_12[228]},
      {stage0_13[95]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[22],stage1_14[53],stage1_13[99],stage1_12[135]}
   );
   gpc615_5 gpc491 (
      {stage0_12[229], stage0_12[230], stage0_12[231], stage0_12[232], stage0_12[233]},
      {stage0_13[96]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[23],stage1_14[54],stage1_13[100],stage1_12[136]}
   );
   gpc615_5 gpc492 (
      {stage0_12[234], stage0_12[235], stage0_12[236], stage0_12[237], stage0_12[238]},
      {stage0_13[97]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[24],stage1_14[55],stage1_13[101],stage1_12[137]}
   );
   gpc615_5 gpc493 (
      {stage0_12[239], stage0_12[240], stage0_12[241], stage0_12[242], stage0_12[243]},
      {stage0_13[98]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[25],stage1_14[56],stage1_13[102],stage1_12[138]}
   );
   gpc615_5 gpc494 (
      {stage0_12[244], stage0_12[245], stage0_12[246], stage0_12[247], stage0_12[248]},
      {stage0_13[99]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[26],stage1_14[57],stage1_13[103],stage1_12[139]}
   );
   gpc615_5 gpc495 (
      {stage0_12[249], stage0_12[250], stage0_12[251], stage0_12[252], stage0_12[253]},
      {stage0_13[100]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[27],stage1_14[58],stage1_13[104],stage1_12[140]}
   );
   gpc615_5 gpc496 (
      {stage0_12[254], stage0_12[255], stage0_12[256], stage0_12[257], stage0_12[258]},
      {stage0_13[101]},
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage1_16[15],stage1_15[28],stage1_14[59],stage1_13[105],stage1_12[141]}
   );
   gpc615_5 gpc497 (
      {stage0_12[259], stage0_12[260], stage0_12[261], stage0_12[262], stage0_12[263]},
      {stage0_13[102]},
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage1_16[16],stage1_15[29],stage1_14[60],stage1_13[106],stage1_12[142]}
   );
   gpc615_5 gpc498 (
      {stage0_12[264], stage0_12[265], stage0_12[266], stage0_12[267], stage0_12[268]},
      {stage0_13[103]},
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage1_16[17],stage1_15[30],stage1_14[61],stage1_13[107],stage1_12[143]}
   );
   gpc615_5 gpc499 (
      {stage0_12[269], stage0_12[270], stage0_12[271], stage0_12[272], stage0_12[273]},
      {stage0_13[104]},
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113]},
      {stage1_16[18],stage1_15[31],stage1_14[62],stage1_13[108],stage1_12[144]}
   );
   gpc615_5 gpc500 (
      {stage0_12[274], stage0_12[275], stage0_12[276], stage0_12[277], stage0_12[278]},
      {stage0_13[105]},
      {stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119]},
      {stage1_16[19],stage1_15[32],stage1_14[63],stage1_13[109],stage1_12[145]}
   );
   gpc615_5 gpc501 (
      {stage0_12[279], stage0_12[280], stage0_12[281], stage0_12[282], stage0_12[283]},
      {stage0_13[106]},
      {stage0_14[120], stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125]},
      {stage1_16[20],stage1_15[33],stage1_14[64],stage1_13[110],stage1_12[146]}
   );
   gpc615_5 gpc502 (
      {stage0_12[284], stage0_12[285], stage0_12[286], stage0_12[287], stage0_12[288]},
      {stage0_13[107]},
      {stage0_14[126], stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131]},
      {stage1_16[21],stage1_15[34],stage1_14[65],stage1_13[111],stage1_12[147]}
   );
   gpc615_5 gpc503 (
      {stage0_12[289], stage0_12[290], stage0_12[291], stage0_12[292], stage0_12[293]},
      {stage0_13[108]},
      {stage0_14[132], stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137]},
      {stage1_16[22],stage1_15[35],stage1_14[66],stage1_13[112],stage1_12[148]}
   );
   gpc615_5 gpc504 (
      {stage0_12[294], stage0_12[295], stage0_12[296], stage0_12[297], stage0_12[298]},
      {stage0_13[109]},
      {stage0_14[138], stage0_14[139], stage0_14[140], stage0_14[141], stage0_14[142], stage0_14[143]},
      {stage1_16[23],stage1_15[36],stage1_14[67],stage1_13[113],stage1_12[149]}
   );
   gpc615_5 gpc505 (
      {stage0_12[299], stage0_12[300], stage0_12[301], stage0_12[302], stage0_12[303]},
      {stage0_13[110]},
      {stage0_14[144], stage0_14[145], stage0_14[146], stage0_14[147], stage0_14[148], stage0_14[149]},
      {stage1_16[24],stage1_15[37],stage1_14[68],stage1_13[114],stage1_12[150]}
   );
   gpc615_5 gpc506 (
      {stage0_12[304], stage0_12[305], stage0_12[306], stage0_12[307], stage0_12[308]},
      {stage0_13[111]},
      {stage0_14[150], stage0_14[151], stage0_14[152], stage0_14[153], stage0_14[154], stage0_14[155]},
      {stage1_16[25],stage1_15[38],stage1_14[69],stage1_13[115],stage1_12[151]}
   );
   gpc615_5 gpc507 (
      {stage0_12[309], stage0_12[310], stage0_12[311], stage0_12[312], stage0_12[313]},
      {stage0_13[112]},
      {stage0_14[156], stage0_14[157], stage0_14[158], stage0_14[159], stage0_14[160], stage0_14[161]},
      {stage1_16[26],stage1_15[39],stage1_14[70],stage1_13[116],stage1_12[152]}
   );
   gpc615_5 gpc508 (
      {stage0_12[314], stage0_12[315], stage0_12[316], stage0_12[317], stage0_12[318]},
      {stage0_13[113]},
      {stage0_14[162], stage0_14[163], stage0_14[164], stage0_14[165], stage0_14[166], stage0_14[167]},
      {stage1_16[27],stage1_15[40],stage1_14[71],stage1_13[117],stage1_12[153]}
   );
   gpc615_5 gpc509 (
      {stage0_12[319], stage0_12[320], stage0_12[321], stage0_12[322], stage0_12[323]},
      {stage0_13[114]},
      {stage0_14[168], stage0_14[169], stage0_14[170], stage0_14[171], stage0_14[172], stage0_14[173]},
      {stage1_16[28],stage1_15[41],stage1_14[72],stage1_13[118],stage1_12[154]}
   );
   gpc615_5 gpc510 (
      {stage0_12[324], stage0_12[325], stage0_12[326], stage0_12[327], stage0_12[328]},
      {stage0_13[115]},
      {stage0_14[174], stage0_14[175], stage0_14[176], stage0_14[177], stage0_14[178], stage0_14[179]},
      {stage1_16[29],stage1_15[42],stage1_14[73],stage1_13[119],stage1_12[155]}
   );
   gpc615_5 gpc511 (
      {stage0_12[329], stage0_12[330], stage0_12[331], stage0_12[332], stage0_12[333]},
      {stage0_13[116]},
      {stage0_14[180], stage0_14[181], stage0_14[182], stage0_14[183], stage0_14[184], stage0_14[185]},
      {stage1_16[30],stage1_15[43],stage1_14[74],stage1_13[120],stage1_12[156]}
   );
   gpc615_5 gpc512 (
      {stage0_12[334], stage0_12[335], stage0_12[336], stage0_12[337], stage0_12[338]},
      {stage0_13[117]},
      {stage0_14[186], stage0_14[187], stage0_14[188], stage0_14[189], stage0_14[190], stage0_14[191]},
      {stage1_16[31],stage1_15[44],stage1_14[75],stage1_13[121],stage1_12[157]}
   );
   gpc615_5 gpc513 (
      {stage0_12[339], stage0_12[340], stage0_12[341], stage0_12[342], stage0_12[343]},
      {stage0_13[118]},
      {stage0_14[192], stage0_14[193], stage0_14[194], stage0_14[195], stage0_14[196], stage0_14[197]},
      {stage1_16[32],stage1_15[45],stage1_14[76],stage1_13[122],stage1_12[158]}
   );
   gpc615_5 gpc514 (
      {stage0_12[344], stage0_12[345], stage0_12[346], stage0_12[347], stage0_12[348]},
      {stage0_13[119]},
      {stage0_14[198], stage0_14[199], stage0_14[200], stage0_14[201], stage0_14[202], stage0_14[203]},
      {stage1_16[33],stage1_15[46],stage1_14[77],stage1_13[123],stage1_12[159]}
   );
   gpc615_5 gpc515 (
      {stage0_12[349], stage0_12[350], stage0_12[351], stage0_12[352], stage0_12[353]},
      {stage0_13[120]},
      {stage0_14[204], stage0_14[205], stage0_14[206], stage0_14[207], stage0_14[208], stage0_14[209]},
      {stage1_16[34],stage1_15[47],stage1_14[78],stage1_13[124],stage1_12[160]}
   );
   gpc615_5 gpc516 (
      {stage0_12[354], stage0_12[355], stage0_12[356], stage0_12[357], stage0_12[358]},
      {stage0_13[121]},
      {stage0_14[210], stage0_14[211], stage0_14[212], stage0_14[213], stage0_14[214], stage0_14[215]},
      {stage1_16[35],stage1_15[48],stage1_14[79],stage1_13[125],stage1_12[161]}
   );
   gpc615_5 gpc517 (
      {stage0_12[359], stage0_12[360], stage0_12[361], stage0_12[362], stage0_12[363]},
      {stage0_13[122]},
      {stage0_14[216], stage0_14[217], stage0_14[218], stage0_14[219], stage0_14[220], stage0_14[221]},
      {stage1_16[36],stage1_15[49],stage1_14[80],stage1_13[126],stage1_12[162]}
   );
   gpc615_5 gpc518 (
      {stage0_12[364], stage0_12[365], stage0_12[366], stage0_12[367], stage0_12[368]},
      {stage0_13[123]},
      {stage0_14[222], stage0_14[223], stage0_14[224], stage0_14[225], stage0_14[226], stage0_14[227]},
      {stage1_16[37],stage1_15[50],stage1_14[81],stage1_13[127],stage1_12[163]}
   );
   gpc615_5 gpc519 (
      {stage0_12[369], stage0_12[370], stage0_12[371], stage0_12[372], stage0_12[373]},
      {stage0_13[124]},
      {stage0_14[228], stage0_14[229], stage0_14[230], stage0_14[231], stage0_14[232], stage0_14[233]},
      {stage1_16[38],stage1_15[51],stage1_14[82],stage1_13[128],stage1_12[164]}
   );
   gpc615_5 gpc520 (
      {stage0_12[374], stage0_12[375], stage0_12[376], stage0_12[377], stage0_12[378]},
      {stage0_13[125]},
      {stage0_14[234], stage0_14[235], stage0_14[236], stage0_14[237], stage0_14[238], stage0_14[239]},
      {stage1_16[39],stage1_15[52],stage1_14[83],stage1_13[129],stage1_12[165]}
   );
   gpc615_5 gpc521 (
      {stage0_12[379], stage0_12[380], stage0_12[381], stage0_12[382], stage0_12[383]},
      {stage0_13[126]},
      {stage0_14[240], stage0_14[241], stage0_14[242], stage0_14[243], stage0_14[244], stage0_14[245]},
      {stage1_16[40],stage1_15[53],stage1_14[84],stage1_13[130],stage1_12[166]}
   );
   gpc615_5 gpc522 (
      {stage0_12[384], stage0_12[385], stage0_12[386], stage0_12[387], stage0_12[388]},
      {stage0_13[127]},
      {stage0_14[246], stage0_14[247], stage0_14[248], stage0_14[249], stage0_14[250], stage0_14[251]},
      {stage1_16[41],stage1_15[54],stage1_14[85],stage1_13[131],stage1_12[167]}
   );
   gpc615_5 gpc523 (
      {stage0_12[389], stage0_12[390], stage0_12[391], stage0_12[392], stage0_12[393]},
      {stage0_13[128]},
      {stage0_14[252], stage0_14[253], stage0_14[254], stage0_14[255], stage0_14[256], stage0_14[257]},
      {stage1_16[42],stage1_15[55],stage1_14[86],stage1_13[132],stage1_12[168]}
   );
   gpc615_5 gpc524 (
      {stage0_12[394], stage0_12[395], stage0_12[396], stage0_12[397], stage0_12[398]},
      {stage0_13[129]},
      {stage0_14[258], stage0_14[259], stage0_14[260], stage0_14[261], stage0_14[262], stage0_14[263]},
      {stage1_16[43],stage1_15[56],stage1_14[87],stage1_13[133],stage1_12[169]}
   );
   gpc615_5 gpc525 (
      {stage0_12[399], stage0_12[400], stage0_12[401], stage0_12[402], stage0_12[403]},
      {stage0_13[130]},
      {stage0_14[264], stage0_14[265], stage0_14[266], stage0_14[267], stage0_14[268], stage0_14[269]},
      {stage1_16[44],stage1_15[57],stage1_14[88],stage1_13[134],stage1_12[170]}
   );
   gpc615_5 gpc526 (
      {stage0_12[404], stage0_12[405], stage0_12[406], stage0_12[407], stage0_12[408]},
      {stage0_13[131]},
      {stage0_14[270], stage0_14[271], stage0_14[272], stage0_14[273], stage0_14[274], stage0_14[275]},
      {stage1_16[45],stage1_15[58],stage1_14[89],stage1_13[135],stage1_12[171]}
   );
   gpc615_5 gpc527 (
      {stage0_12[409], stage0_12[410], stage0_12[411], stage0_12[412], stage0_12[413]},
      {stage0_13[132]},
      {stage0_14[276], stage0_14[277], stage0_14[278], stage0_14[279], stage0_14[280], stage0_14[281]},
      {stage1_16[46],stage1_15[59],stage1_14[90],stage1_13[136],stage1_12[172]}
   );
   gpc615_5 gpc528 (
      {stage0_12[414], stage0_12[415], stage0_12[416], stage0_12[417], stage0_12[418]},
      {stage0_13[133]},
      {stage0_14[282], stage0_14[283], stage0_14[284], stage0_14[285], stage0_14[286], stage0_14[287]},
      {stage1_16[47],stage1_15[60],stage1_14[91],stage1_13[137],stage1_12[173]}
   );
   gpc615_5 gpc529 (
      {stage0_12[419], stage0_12[420], stage0_12[421], stage0_12[422], stage0_12[423]},
      {stage0_13[134]},
      {stage0_14[288], stage0_14[289], stage0_14[290], stage0_14[291], stage0_14[292], stage0_14[293]},
      {stage1_16[48],stage1_15[61],stage1_14[92],stage1_13[138],stage1_12[174]}
   );
   gpc615_5 gpc530 (
      {stage0_12[424], stage0_12[425], stage0_12[426], stage0_12[427], stage0_12[428]},
      {stage0_13[135]},
      {stage0_14[294], stage0_14[295], stage0_14[296], stage0_14[297], stage0_14[298], stage0_14[299]},
      {stage1_16[49],stage1_15[62],stage1_14[93],stage1_13[139],stage1_12[175]}
   );
   gpc615_5 gpc531 (
      {stage0_12[429], stage0_12[430], stage0_12[431], stage0_12[432], stage0_12[433]},
      {stage0_13[136]},
      {stage0_14[300], stage0_14[301], stage0_14[302], stage0_14[303], stage0_14[304], stage0_14[305]},
      {stage1_16[50],stage1_15[63],stage1_14[94],stage1_13[140],stage1_12[176]}
   );
   gpc615_5 gpc532 (
      {stage0_12[434], stage0_12[435], stage0_12[436], stage0_12[437], stage0_12[438]},
      {stage0_13[137]},
      {stage0_14[306], stage0_14[307], stage0_14[308], stage0_14[309], stage0_14[310], stage0_14[311]},
      {stage1_16[51],stage1_15[64],stage1_14[95],stage1_13[141],stage1_12[177]}
   );
   gpc615_5 gpc533 (
      {stage0_12[439], stage0_12[440], stage0_12[441], stage0_12[442], stage0_12[443]},
      {stage0_13[138]},
      {stage0_14[312], stage0_14[313], stage0_14[314], stage0_14[315], stage0_14[316], stage0_14[317]},
      {stage1_16[52],stage1_15[65],stage1_14[96],stage1_13[142],stage1_12[178]}
   );
   gpc615_5 gpc534 (
      {stage0_12[444], stage0_12[445], stage0_12[446], stage0_12[447], stage0_12[448]},
      {stage0_13[139]},
      {stage0_14[318], stage0_14[319], stage0_14[320], stage0_14[321], stage0_14[322], stage0_14[323]},
      {stage1_16[53],stage1_15[66],stage1_14[97],stage1_13[143],stage1_12[179]}
   );
   gpc615_5 gpc535 (
      {stage0_12[449], stage0_12[450], stage0_12[451], stage0_12[452], stage0_12[453]},
      {stage0_13[140]},
      {stage0_14[324], stage0_14[325], stage0_14[326], stage0_14[327], stage0_14[328], stage0_14[329]},
      {stage1_16[54],stage1_15[67],stage1_14[98],stage1_13[144],stage1_12[180]}
   );
   gpc615_5 gpc536 (
      {stage0_12[454], stage0_12[455], stage0_12[456], stage0_12[457], stage0_12[458]},
      {stage0_13[141]},
      {stage0_14[330], stage0_14[331], stage0_14[332], stage0_14[333], stage0_14[334], stage0_14[335]},
      {stage1_16[55],stage1_15[68],stage1_14[99],stage1_13[145],stage1_12[181]}
   );
   gpc615_5 gpc537 (
      {stage0_12[459], stage0_12[460], stage0_12[461], stage0_12[462], stage0_12[463]},
      {stage0_13[142]},
      {stage0_14[336], stage0_14[337], stage0_14[338], stage0_14[339], stage0_14[340], stage0_14[341]},
      {stage1_16[56],stage1_15[69],stage1_14[100],stage1_13[146],stage1_12[182]}
   );
   gpc615_5 gpc538 (
      {stage0_12[464], stage0_12[465], stage0_12[466], stage0_12[467], stage0_12[468]},
      {stage0_13[143]},
      {stage0_14[342], stage0_14[343], stage0_14[344], stage0_14[345], stage0_14[346], stage0_14[347]},
      {stage1_16[57],stage1_15[70],stage1_14[101],stage1_13[147],stage1_12[183]}
   );
   gpc615_5 gpc539 (
      {stage0_12[469], stage0_12[470], stage0_12[471], stage0_12[472], stage0_12[473]},
      {stage0_13[144]},
      {stage0_14[348], stage0_14[349], stage0_14[350], stage0_14[351], stage0_14[352], stage0_14[353]},
      {stage1_16[58],stage1_15[71],stage1_14[102],stage1_13[148],stage1_12[184]}
   );
   gpc615_5 gpc540 (
      {stage0_12[474], stage0_12[475], stage0_12[476], stage0_12[477], stage0_12[478]},
      {stage0_13[145]},
      {stage0_14[354], stage0_14[355], stage0_14[356], stage0_14[357], stage0_14[358], stage0_14[359]},
      {stage1_16[59],stage1_15[72],stage1_14[103],stage1_13[149],stage1_12[185]}
   );
   gpc615_5 gpc541 (
      {stage0_12[479], stage0_12[480], stage0_12[481], stage0_12[482], stage0_12[483]},
      {stage0_13[146]},
      {stage0_14[360], stage0_14[361], stage0_14[362], stage0_14[363], stage0_14[364], stage0_14[365]},
      {stage1_16[60],stage1_15[73],stage1_14[104],stage1_13[150],stage1_12[186]}
   );
   gpc606_5 gpc542 (
      {stage0_13[147], stage0_13[148], stage0_13[149], stage0_13[150], stage0_13[151], stage0_13[152]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[61],stage1_15[74],stage1_14[105],stage1_13[151]}
   );
   gpc606_5 gpc543 (
      {stage0_13[153], stage0_13[154], stage0_13[155], stage0_13[156], stage0_13[157], stage0_13[158]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[62],stage1_15[75],stage1_14[106],stage1_13[152]}
   );
   gpc606_5 gpc544 (
      {stage0_13[159], stage0_13[160], stage0_13[161], stage0_13[162], stage0_13[163], stage0_13[164]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[63],stage1_15[76],stage1_14[107],stage1_13[153]}
   );
   gpc606_5 gpc545 (
      {stage0_13[165], stage0_13[166], stage0_13[167], stage0_13[168], stage0_13[169], stage0_13[170]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[64],stage1_15[77],stage1_14[108],stage1_13[154]}
   );
   gpc606_5 gpc546 (
      {stage0_13[171], stage0_13[172], stage0_13[173], stage0_13[174], stage0_13[175], stage0_13[176]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[65],stage1_15[78],stage1_14[109],stage1_13[155]}
   );
   gpc606_5 gpc547 (
      {stage0_13[177], stage0_13[178], stage0_13[179], stage0_13[180], stage0_13[181], stage0_13[182]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[66],stage1_15[79],stage1_14[110],stage1_13[156]}
   );
   gpc606_5 gpc548 (
      {stage0_13[183], stage0_13[184], stage0_13[185], stage0_13[186], stage0_13[187], stage0_13[188]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[67],stage1_15[80],stage1_14[111],stage1_13[157]}
   );
   gpc606_5 gpc549 (
      {stage0_13[189], stage0_13[190], stage0_13[191], stage0_13[192], stage0_13[193], stage0_13[194]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[68],stage1_15[81],stage1_14[112],stage1_13[158]}
   );
   gpc606_5 gpc550 (
      {stage0_13[195], stage0_13[196], stage0_13[197], stage0_13[198], stage0_13[199], stage0_13[200]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[69],stage1_15[82],stage1_14[113],stage1_13[159]}
   );
   gpc615_5 gpc551 (
      {stage0_13[201], stage0_13[202], stage0_13[203], stage0_13[204], stage0_13[205]},
      {stage0_14[366]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[70],stage1_15[83],stage1_14[114],stage1_13[160]}
   );
   gpc615_5 gpc552 (
      {stage0_13[206], stage0_13[207], stage0_13[208], stage0_13[209], stage0_13[210]},
      {stage0_14[367]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[71],stage1_15[84],stage1_14[115],stage1_13[161]}
   );
   gpc615_5 gpc553 (
      {stage0_13[211], stage0_13[212], stage0_13[213], stage0_13[214], stage0_13[215]},
      {stage0_14[368]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[72],stage1_15[85],stage1_14[116],stage1_13[162]}
   );
   gpc615_5 gpc554 (
      {stage0_13[216], stage0_13[217], stage0_13[218], stage0_13[219], stage0_13[220]},
      {stage0_14[369]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[73],stage1_15[86],stage1_14[117],stage1_13[163]}
   );
   gpc615_5 gpc555 (
      {stage0_13[221], stage0_13[222], stage0_13[223], stage0_13[224], stage0_13[225]},
      {stage0_14[370]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[74],stage1_15[87],stage1_14[118],stage1_13[164]}
   );
   gpc615_5 gpc556 (
      {stage0_13[226], stage0_13[227], stage0_13[228], stage0_13[229], stage0_13[230]},
      {stage0_14[371]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[75],stage1_15[88],stage1_14[119],stage1_13[165]}
   );
   gpc615_5 gpc557 (
      {stage0_13[231], stage0_13[232], stage0_13[233], stage0_13[234], stage0_13[235]},
      {stage0_14[372]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[76],stage1_15[89],stage1_14[120],stage1_13[166]}
   );
   gpc615_5 gpc558 (
      {stage0_13[236], stage0_13[237], stage0_13[238], stage0_13[239], stage0_13[240]},
      {stage0_14[373]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[77],stage1_15[90],stage1_14[121],stage1_13[167]}
   );
   gpc615_5 gpc559 (
      {stage0_13[241], stage0_13[242], stage0_13[243], stage0_13[244], stage0_13[245]},
      {stage0_14[374]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[78],stage1_15[91],stage1_14[122],stage1_13[168]}
   );
   gpc615_5 gpc560 (
      {stage0_13[246], stage0_13[247], stage0_13[248], stage0_13[249], stage0_13[250]},
      {stage0_14[375]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[79],stage1_15[92],stage1_14[123],stage1_13[169]}
   );
   gpc615_5 gpc561 (
      {stage0_13[251], stage0_13[252], stage0_13[253], stage0_13[254], stage0_13[255]},
      {stage0_14[376]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[80],stage1_15[93],stage1_14[124],stage1_13[170]}
   );
   gpc615_5 gpc562 (
      {stage0_13[256], stage0_13[257], stage0_13[258], stage0_13[259], stage0_13[260]},
      {stage0_14[377]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[81],stage1_15[94],stage1_14[125],stage1_13[171]}
   );
   gpc615_5 gpc563 (
      {stage0_13[261], stage0_13[262], stage0_13[263], stage0_13[264], stage0_13[265]},
      {stage0_14[378]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[82],stage1_15[95],stage1_14[126],stage1_13[172]}
   );
   gpc615_5 gpc564 (
      {stage0_13[266], stage0_13[267], stage0_13[268], stage0_13[269], stage0_13[270]},
      {stage0_14[379]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[83],stage1_15[96],stage1_14[127],stage1_13[173]}
   );
   gpc615_5 gpc565 (
      {stage0_13[271], stage0_13[272], stage0_13[273], stage0_13[274], stage0_13[275]},
      {stage0_14[380]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[84],stage1_15[97],stage1_14[128],stage1_13[174]}
   );
   gpc615_5 gpc566 (
      {stage0_13[276], stage0_13[277], stage0_13[278], stage0_13[279], stage0_13[280]},
      {stage0_14[381]},
      {stage0_15[144], stage0_15[145], stage0_15[146], stage0_15[147], stage0_15[148], stage0_15[149]},
      {stage1_17[24],stage1_16[85],stage1_15[98],stage1_14[129],stage1_13[175]}
   );
   gpc615_5 gpc567 (
      {stage0_13[281], stage0_13[282], stage0_13[283], stage0_13[284], stage0_13[285]},
      {stage0_14[382]},
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155]},
      {stage1_17[25],stage1_16[86],stage1_15[99],stage1_14[130],stage1_13[176]}
   );
   gpc615_5 gpc568 (
      {stage0_13[286], stage0_13[287], stage0_13[288], stage0_13[289], stage0_13[290]},
      {stage0_14[383]},
      {stage0_15[156], stage0_15[157], stage0_15[158], stage0_15[159], stage0_15[160], stage0_15[161]},
      {stage1_17[26],stage1_16[87],stage1_15[100],stage1_14[131],stage1_13[177]}
   );
   gpc615_5 gpc569 (
      {stage0_13[291], stage0_13[292], stage0_13[293], stage0_13[294], stage0_13[295]},
      {stage0_14[384]},
      {stage0_15[162], stage0_15[163], stage0_15[164], stage0_15[165], stage0_15[166], stage0_15[167]},
      {stage1_17[27],stage1_16[88],stage1_15[101],stage1_14[132],stage1_13[178]}
   );
   gpc615_5 gpc570 (
      {stage0_13[296], stage0_13[297], stage0_13[298], stage0_13[299], stage0_13[300]},
      {stage0_14[385]},
      {stage0_15[168], stage0_15[169], stage0_15[170], stage0_15[171], stage0_15[172], stage0_15[173]},
      {stage1_17[28],stage1_16[89],stage1_15[102],stage1_14[133],stage1_13[179]}
   );
   gpc615_5 gpc571 (
      {stage0_13[301], stage0_13[302], stage0_13[303], stage0_13[304], stage0_13[305]},
      {stage0_14[386]},
      {stage0_15[174], stage0_15[175], stage0_15[176], stage0_15[177], stage0_15[178], stage0_15[179]},
      {stage1_17[29],stage1_16[90],stage1_15[103],stage1_14[134],stage1_13[180]}
   );
   gpc615_5 gpc572 (
      {stage0_13[306], stage0_13[307], stage0_13[308], stage0_13[309], stage0_13[310]},
      {stage0_14[387]},
      {stage0_15[180], stage0_15[181], stage0_15[182], stage0_15[183], stage0_15[184], stage0_15[185]},
      {stage1_17[30],stage1_16[91],stage1_15[104],stage1_14[135],stage1_13[181]}
   );
   gpc615_5 gpc573 (
      {stage0_13[311], stage0_13[312], stage0_13[313], stage0_13[314], stage0_13[315]},
      {stage0_14[388]},
      {stage0_15[186], stage0_15[187], stage0_15[188], stage0_15[189], stage0_15[190], stage0_15[191]},
      {stage1_17[31],stage1_16[92],stage1_15[105],stage1_14[136],stage1_13[182]}
   );
   gpc615_5 gpc574 (
      {stage0_13[316], stage0_13[317], stage0_13[318], stage0_13[319], stage0_13[320]},
      {stage0_14[389]},
      {stage0_15[192], stage0_15[193], stage0_15[194], stage0_15[195], stage0_15[196], stage0_15[197]},
      {stage1_17[32],stage1_16[93],stage1_15[106],stage1_14[137],stage1_13[183]}
   );
   gpc615_5 gpc575 (
      {stage0_13[321], stage0_13[322], stage0_13[323], stage0_13[324], stage0_13[325]},
      {stage0_14[390]},
      {stage0_15[198], stage0_15[199], stage0_15[200], stage0_15[201], stage0_15[202], stage0_15[203]},
      {stage1_17[33],stage1_16[94],stage1_15[107],stage1_14[138],stage1_13[184]}
   );
   gpc615_5 gpc576 (
      {stage0_13[326], stage0_13[327], stage0_13[328], stage0_13[329], stage0_13[330]},
      {stage0_14[391]},
      {stage0_15[204], stage0_15[205], stage0_15[206], stage0_15[207], stage0_15[208], stage0_15[209]},
      {stage1_17[34],stage1_16[95],stage1_15[108],stage1_14[139],stage1_13[185]}
   );
   gpc615_5 gpc577 (
      {stage0_13[331], stage0_13[332], stage0_13[333], stage0_13[334], stage0_13[335]},
      {stage0_14[392]},
      {stage0_15[210], stage0_15[211], stage0_15[212], stage0_15[213], stage0_15[214], stage0_15[215]},
      {stage1_17[35],stage1_16[96],stage1_15[109],stage1_14[140],stage1_13[186]}
   );
   gpc615_5 gpc578 (
      {stage0_13[336], stage0_13[337], stage0_13[338], stage0_13[339], stage0_13[340]},
      {stage0_14[393]},
      {stage0_15[216], stage0_15[217], stage0_15[218], stage0_15[219], stage0_15[220], stage0_15[221]},
      {stage1_17[36],stage1_16[97],stage1_15[110],stage1_14[141],stage1_13[187]}
   );
   gpc615_5 gpc579 (
      {stage0_13[341], stage0_13[342], stage0_13[343], stage0_13[344], stage0_13[345]},
      {stage0_14[394]},
      {stage0_15[222], stage0_15[223], stage0_15[224], stage0_15[225], stage0_15[226], stage0_15[227]},
      {stage1_17[37],stage1_16[98],stage1_15[111],stage1_14[142],stage1_13[188]}
   );
   gpc615_5 gpc580 (
      {stage0_13[346], stage0_13[347], stage0_13[348], stage0_13[349], stage0_13[350]},
      {stage0_14[395]},
      {stage0_15[228], stage0_15[229], stage0_15[230], stage0_15[231], stage0_15[232], stage0_15[233]},
      {stage1_17[38],stage1_16[99],stage1_15[112],stage1_14[143],stage1_13[189]}
   );
   gpc615_5 gpc581 (
      {stage0_13[351], stage0_13[352], stage0_13[353], stage0_13[354], stage0_13[355]},
      {stage0_14[396]},
      {stage0_15[234], stage0_15[235], stage0_15[236], stage0_15[237], stage0_15[238], stage0_15[239]},
      {stage1_17[39],stage1_16[100],stage1_15[113],stage1_14[144],stage1_13[190]}
   );
   gpc615_5 gpc582 (
      {stage0_13[356], stage0_13[357], stage0_13[358], stage0_13[359], stage0_13[360]},
      {stage0_14[397]},
      {stage0_15[240], stage0_15[241], stage0_15[242], stage0_15[243], stage0_15[244], stage0_15[245]},
      {stage1_17[40],stage1_16[101],stage1_15[114],stage1_14[145],stage1_13[191]}
   );
   gpc615_5 gpc583 (
      {stage0_13[361], stage0_13[362], stage0_13[363], stage0_13[364], stage0_13[365]},
      {stage0_14[398]},
      {stage0_15[246], stage0_15[247], stage0_15[248], stage0_15[249], stage0_15[250], stage0_15[251]},
      {stage1_17[41],stage1_16[102],stage1_15[115],stage1_14[146],stage1_13[192]}
   );
   gpc615_5 gpc584 (
      {stage0_13[366], stage0_13[367], stage0_13[368], stage0_13[369], stage0_13[370]},
      {stage0_14[399]},
      {stage0_15[252], stage0_15[253], stage0_15[254], stage0_15[255], stage0_15[256], stage0_15[257]},
      {stage1_17[42],stage1_16[103],stage1_15[116],stage1_14[147],stage1_13[193]}
   );
   gpc615_5 gpc585 (
      {stage0_13[371], stage0_13[372], stage0_13[373], stage0_13[374], stage0_13[375]},
      {stage0_14[400]},
      {stage0_15[258], stage0_15[259], stage0_15[260], stage0_15[261], stage0_15[262], stage0_15[263]},
      {stage1_17[43],stage1_16[104],stage1_15[117],stage1_14[148],stage1_13[194]}
   );
   gpc606_5 gpc586 (
      {stage0_14[401], stage0_14[402], stage0_14[403], stage0_14[404], stage0_14[405], stage0_14[406]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[44],stage1_16[105],stage1_15[118],stage1_14[149]}
   );
   gpc606_5 gpc587 (
      {stage0_14[407], stage0_14[408], stage0_14[409], stage0_14[410], stage0_14[411], stage0_14[412]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[45],stage1_16[106],stage1_15[119],stage1_14[150]}
   );
   gpc606_5 gpc588 (
      {stage0_14[413], stage0_14[414], stage0_14[415], stage0_14[416], stage0_14[417], stage0_14[418]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[46],stage1_16[107],stage1_15[120],stage1_14[151]}
   );
   gpc615_5 gpc589 (
      {stage0_15[264], stage0_15[265], stage0_15[266], stage0_15[267], stage0_15[268]},
      {stage0_16[18]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[3],stage1_17[47],stage1_16[108],stage1_15[121]}
   );
   gpc615_5 gpc590 (
      {stage0_15[269], stage0_15[270], stage0_15[271], stage0_15[272], stage0_15[273]},
      {stage0_16[19]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[4],stage1_17[48],stage1_16[109],stage1_15[122]}
   );
   gpc615_5 gpc591 (
      {stage0_15[274], stage0_15[275], stage0_15[276], stage0_15[277], stage0_15[278]},
      {stage0_16[20]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[5],stage1_17[49],stage1_16[110],stage1_15[123]}
   );
   gpc615_5 gpc592 (
      {stage0_15[279], stage0_15[280], stage0_15[281], stage0_15[282], stage0_15[283]},
      {stage0_16[21]},
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage1_19[3],stage1_18[6],stage1_17[50],stage1_16[111],stage1_15[124]}
   );
   gpc615_5 gpc593 (
      {stage0_15[284], stage0_15[285], stage0_15[286], stage0_15[287], stage0_15[288]},
      {stage0_16[22]},
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage1_19[4],stage1_18[7],stage1_17[51],stage1_16[112],stage1_15[125]}
   );
   gpc615_5 gpc594 (
      {stage0_15[289], stage0_15[290], stage0_15[291], stage0_15[292], stage0_15[293]},
      {stage0_16[23]},
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage1_19[5],stage1_18[8],stage1_17[52],stage1_16[113],stage1_15[126]}
   );
   gpc615_5 gpc595 (
      {stage0_15[294], stage0_15[295], stage0_15[296], stage0_15[297], stage0_15[298]},
      {stage0_16[24]},
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage1_19[6],stage1_18[9],stage1_17[53],stage1_16[114],stage1_15[127]}
   );
   gpc615_5 gpc596 (
      {stage0_15[299], stage0_15[300], stage0_15[301], stage0_15[302], stage0_15[303]},
      {stage0_16[25]},
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage1_19[7],stage1_18[10],stage1_17[54],stage1_16[115],stage1_15[128]}
   );
   gpc615_5 gpc597 (
      {stage0_15[304], stage0_15[305], stage0_15[306], stage0_15[307], stage0_15[308]},
      {stage0_16[26]},
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage1_19[8],stage1_18[11],stage1_17[55],stage1_16[116],stage1_15[129]}
   );
   gpc615_5 gpc598 (
      {stage0_15[309], stage0_15[310], stage0_15[311], stage0_15[312], stage0_15[313]},
      {stage0_16[27]},
      {stage0_17[54], stage0_17[55], stage0_17[56], stage0_17[57], stage0_17[58], stage0_17[59]},
      {stage1_19[9],stage1_18[12],stage1_17[56],stage1_16[117],stage1_15[130]}
   );
   gpc615_5 gpc599 (
      {stage0_15[314], stage0_15[315], stage0_15[316], stage0_15[317], stage0_15[318]},
      {stage0_16[28]},
      {stage0_17[60], stage0_17[61], stage0_17[62], stage0_17[63], stage0_17[64], stage0_17[65]},
      {stage1_19[10],stage1_18[13],stage1_17[57],stage1_16[118],stage1_15[131]}
   );
   gpc615_5 gpc600 (
      {stage0_15[319], stage0_15[320], stage0_15[321], stage0_15[322], stage0_15[323]},
      {stage0_16[29]},
      {stage0_17[66], stage0_17[67], stage0_17[68], stage0_17[69], stage0_17[70], stage0_17[71]},
      {stage1_19[11],stage1_18[14],stage1_17[58],stage1_16[119],stage1_15[132]}
   );
   gpc615_5 gpc601 (
      {stage0_15[324], stage0_15[325], stage0_15[326], stage0_15[327], stage0_15[328]},
      {stage0_16[30]},
      {stage0_17[72], stage0_17[73], stage0_17[74], stage0_17[75], stage0_17[76], stage0_17[77]},
      {stage1_19[12],stage1_18[15],stage1_17[59],stage1_16[120],stage1_15[133]}
   );
   gpc615_5 gpc602 (
      {stage0_15[329], stage0_15[330], stage0_15[331], stage0_15[332], stage0_15[333]},
      {stage0_16[31]},
      {stage0_17[78], stage0_17[79], stage0_17[80], stage0_17[81], stage0_17[82], stage0_17[83]},
      {stage1_19[13],stage1_18[16],stage1_17[60],stage1_16[121],stage1_15[134]}
   );
   gpc615_5 gpc603 (
      {stage0_15[334], stage0_15[335], stage0_15[336], stage0_15[337], stage0_15[338]},
      {stage0_16[32]},
      {stage0_17[84], stage0_17[85], stage0_17[86], stage0_17[87], stage0_17[88], stage0_17[89]},
      {stage1_19[14],stage1_18[17],stage1_17[61],stage1_16[122],stage1_15[135]}
   );
   gpc615_5 gpc604 (
      {stage0_15[339], stage0_15[340], stage0_15[341], stage0_15[342], stage0_15[343]},
      {stage0_16[33]},
      {stage0_17[90], stage0_17[91], stage0_17[92], stage0_17[93], stage0_17[94], stage0_17[95]},
      {stage1_19[15],stage1_18[18],stage1_17[62],stage1_16[123],stage1_15[136]}
   );
   gpc615_5 gpc605 (
      {stage0_15[344], stage0_15[345], stage0_15[346], stage0_15[347], stage0_15[348]},
      {stage0_16[34]},
      {stage0_17[96], stage0_17[97], stage0_17[98], stage0_17[99], stage0_17[100], stage0_17[101]},
      {stage1_19[16],stage1_18[19],stage1_17[63],stage1_16[124],stage1_15[137]}
   );
   gpc615_5 gpc606 (
      {stage0_15[349], stage0_15[350], stage0_15[351], stage0_15[352], stage0_15[353]},
      {stage0_16[35]},
      {stage0_17[102], stage0_17[103], stage0_17[104], stage0_17[105], stage0_17[106], stage0_17[107]},
      {stage1_19[17],stage1_18[20],stage1_17[64],stage1_16[125],stage1_15[138]}
   );
   gpc615_5 gpc607 (
      {stage0_15[354], stage0_15[355], stage0_15[356], stage0_15[357], stage0_15[358]},
      {stage0_16[36]},
      {stage0_17[108], stage0_17[109], stage0_17[110], stage0_17[111], stage0_17[112], stage0_17[113]},
      {stage1_19[18],stage1_18[21],stage1_17[65],stage1_16[126],stage1_15[139]}
   );
   gpc615_5 gpc608 (
      {stage0_15[359], stage0_15[360], stage0_15[361], stage0_15[362], stage0_15[363]},
      {stage0_16[37]},
      {stage0_17[114], stage0_17[115], stage0_17[116], stage0_17[117], stage0_17[118], stage0_17[119]},
      {stage1_19[19],stage1_18[22],stage1_17[66],stage1_16[127],stage1_15[140]}
   );
   gpc615_5 gpc609 (
      {stage0_15[364], stage0_15[365], stage0_15[366], stage0_15[367], stage0_15[368]},
      {stage0_16[38]},
      {stage0_17[120], stage0_17[121], stage0_17[122], stage0_17[123], stage0_17[124], stage0_17[125]},
      {stage1_19[20],stage1_18[23],stage1_17[67],stage1_16[128],stage1_15[141]}
   );
   gpc615_5 gpc610 (
      {stage0_15[369], stage0_15[370], stage0_15[371], stage0_15[372], stage0_15[373]},
      {stage0_16[39]},
      {stage0_17[126], stage0_17[127], stage0_17[128], stage0_17[129], stage0_17[130], stage0_17[131]},
      {stage1_19[21],stage1_18[24],stage1_17[68],stage1_16[129],stage1_15[142]}
   );
   gpc615_5 gpc611 (
      {stage0_15[374], stage0_15[375], stage0_15[376], stage0_15[377], stage0_15[378]},
      {stage0_16[40]},
      {stage0_17[132], stage0_17[133], stage0_17[134], stage0_17[135], stage0_17[136], stage0_17[137]},
      {stage1_19[22],stage1_18[25],stage1_17[69],stage1_16[130],stage1_15[143]}
   );
   gpc615_5 gpc612 (
      {stage0_15[379], stage0_15[380], stage0_15[381], stage0_15[382], stage0_15[383]},
      {stage0_16[41]},
      {stage0_17[138], stage0_17[139], stage0_17[140], stage0_17[141], stage0_17[142], stage0_17[143]},
      {stage1_19[23],stage1_18[26],stage1_17[70],stage1_16[131],stage1_15[144]}
   );
   gpc615_5 gpc613 (
      {stage0_15[384], stage0_15[385], stage0_15[386], stage0_15[387], stage0_15[388]},
      {stage0_16[42]},
      {stage0_17[144], stage0_17[145], stage0_17[146], stage0_17[147], stage0_17[148], stage0_17[149]},
      {stage1_19[24],stage1_18[27],stage1_17[71],stage1_16[132],stage1_15[145]}
   );
   gpc615_5 gpc614 (
      {stage0_15[389], stage0_15[390], stage0_15[391], stage0_15[392], stage0_15[393]},
      {stage0_16[43]},
      {stage0_17[150], stage0_17[151], stage0_17[152], stage0_17[153], stage0_17[154], stage0_17[155]},
      {stage1_19[25],stage1_18[28],stage1_17[72],stage1_16[133],stage1_15[146]}
   );
   gpc615_5 gpc615 (
      {stage0_15[394], stage0_15[395], stage0_15[396], stage0_15[397], stage0_15[398]},
      {stage0_16[44]},
      {stage0_17[156], stage0_17[157], stage0_17[158], stage0_17[159], stage0_17[160], stage0_17[161]},
      {stage1_19[26],stage1_18[29],stage1_17[73],stage1_16[134],stage1_15[147]}
   );
   gpc615_5 gpc616 (
      {stage0_15[399], stage0_15[400], stage0_15[401], stage0_15[402], stage0_15[403]},
      {stage0_16[45]},
      {stage0_17[162], stage0_17[163], stage0_17[164], stage0_17[165], stage0_17[166], stage0_17[167]},
      {stage1_19[27],stage1_18[30],stage1_17[74],stage1_16[135],stage1_15[148]}
   );
   gpc615_5 gpc617 (
      {stage0_15[404], stage0_15[405], stage0_15[406], stage0_15[407], stage0_15[408]},
      {stage0_16[46]},
      {stage0_17[168], stage0_17[169], stage0_17[170], stage0_17[171], stage0_17[172], stage0_17[173]},
      {stage1_19[28],stage1_18[31],stage1_17[75],stage1_16[136],stage1_15[149]}
   );
   gpc615_5 gpc618 (
      {stage0_15[409], stage0_15[410], stage0_15[411], stage0_15[412], stage0_15[413]},
      {stage0_16[47]},
      {stage0_17[174], stage0_17[175], stage0_17[176], stage0_17[177], stage0_17[178], stage0_17[179]},
      {stage1_19[29],stage1_18[32],stage1_17[76],stage1_16[137],stage1_15[150]}
   );
   gpc615_5 gpc619 (
      {stage0_15[414], stage0_15[415], stage0_15[416], stage0_15[417], stage0_15[418]},
      {stage0_16[48]},
      {stage0_17[180], stage0_17[181], stage0_17[182], stage0_17[183], stage0_17[184], stage0_17[185]},
      {stage1_19[30],stage1_18[33],stage1_17[77],stage1_16[138],stage1_15[151]}
   );
   gpc615_5 gpc620 (
      {stage0_15[419], stage0_15[420], stage0_15[421], stage0_15[422], stage0_15[423]},
      {stage0_16[49]},
      {stage0_17[186], stage0_17[187], stage0_17[188], stage0_17[189], stage0_17[190], stage0_17[191]},
      {stage1_19[31],stage1_18[34],stage1_17[78],stage1_16[139],stage1_15[152]}
   );
   gpc615_5 gpc621 (
      {stage0_15[424], stage0_15[425], stage0_15[426], stage0_15[427], stage0_15[428]},
      {stage0_16[50]},
      {stage0_17[192], stage0_17[193], stage0_17[194], stage0_17[195], stage0_17[196], stage0_17[197]},
      {stage1_19[32],stage1_18[35],stage1_17[79],stage1_16[140],stage1_15[153]}
   );
   gpc615_5 gpc622 (
      {stage0_15[429], stage0_15[430], stage0_15[431], stage0_15[432], stage0_15[433]},
      {stage0_16[51]},
      {stage0_17[198], stage0_17[199], stage0_17[200], stage0_17[201], stage0_17[202], stage0_17[203]},
      {stage1_19[33],stage1_18[36],stage1_17[80],stage1_16[141],stage1_15[154]}
   );
   gpc615_5 gpc623 (
      {stage0_15[434], stage0_15[435], stage0_15[436], stage0_15[437], stage0_15[438]},
      {stage0_16[52]},
      {stage0_17[204], stage0_17[205], stage0_17[206], stage0_17[207], stage0_17[208], stage0_17[209]},
      {stage1_19[34],stage1_18[37],stage1_17[81],stage1_16[142],stage1_15[155]}
   );
   gpc615_5 gpc624 (
      {stage0_15[439], stage0_15[440], stage0_15[441], stage0_15[442], stage0_15[443]},
      {stage0_16[53]},
      {stage0_17[210], stage0_17[211], stage0_17[212], stage0_17[213], stage0_17[214], stage0_17[215]},
      {stage1_19[35],stage1_18[38],stage1_17[82],stage1_16[143],stage1_15[156]}
   );
   gpc615_5 gpc625 (
      {stage0_15[444], stage0_15[445], stage0_15[446], stage0_15[447], stage0_15[448]},
      {stage0_16[54]},
      {stage0_17[216], stage0_17[217], stage0_17[218], stage0_17[219], stage0_17[220], stage0_17[221]},
      {stage1_19[36],stage1_18[39],stage1_17[83],stage1_16[144],stage1_15[157]}
   );
   gpc615_5 gpc626 (
      {stage0_15[449], stage0_15[450], stage0_15[451], stage0_15[452], stage0_15[453]},
      {stage0_16[55]},
      {stage0_17[222], stage0_17[223], stage0_17[224], stage0_17[225], stage0_17[226], stage0_17[227]},
      {stage1_19[37],stage1_18[40],stage1_17[84],stage1_16[145],stage1_15[158]}
   );
   gpc615_5 gpc627 (
      {stage0_15[454], stage0_15[455], stage0_15[456], stage0_15[457], stage0_15[458]},
      {stage0_16[56]},
      {stage0_17[228], stage0_17[229], stage0_17[230], stage0_17[231], stage0_17[232], stage0_17[233]},
      {stage1_19[38],stage1_18[41],stage1_17[85],stage1_16[146],stage1_15[159]}
   );
   gpc615_5 gpc628 (
      {stage0_15[459], stage0_15[460], stage0_15[461], stage0_15[462], stage0_15[463]},
      {stage0_16[57]},
      {stage0_17[234], stage0_17[235], stage0_17[236], stage0_17[237], stage0_17[238], stage0_17[239]},
      {stage1_19[39],stage1_18[42],stage1_17[86],stage1_16[147],stage1_15[160]}
   );
   gpc615_5 gpc629 (
      {stage0_15[464], stage0_15[465], stage0_15[466], stage0_15[467], stage0_15[468]},
      {stage0_16[58]},
      {stage0_17[240], stage0_17[241], stage0_17[242], stage0_17[243], stage0_17[244], stage0_17[245]},
      {stage1_19[40],stage1_18[43],stage1_17[87],stage1_16[148],stage1_15[161]}
   );
   gpc615_5 gpc630 (
      {stage0_15[469], stage0_15[470], stage0_15[471], stage0_15[472], stage0_15[473]},
      {stage0_16[59]},
      {stage0_17[246], stage0_17[247], stage0_17[248], stage0_17[249], stage0_17[250], stage0_17[251]},
      {stage1_19[41],stage1_18[44],stage1_17[88],stage1_16[149],stage1_15[162]}
   );
   gpc615_5 gpc631 (
      {stage0_15[474], stage0_15[475], stage0_15[476], stage0_15[477], stage0_15[478]},
      {stage0_16[60]},
      {stage0_17[252], stage0_17[253], stage0_17[254], stage0_17[255], stage0_17[256], stage0_17[257]},
      {stage1_19[42],stage1_18[45],stage1_17[89],stage1_16[150],stage1_15[163]}
   );
   gpc606_5 gpc632 (
      {stage0_16[61], stage0_16[62], stage0_16[63], stage0_16[64], stage0_16[65], stage0_16[66]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[43],stage1_18[46],stage1_17[90],stage1_16[151]}
   );
   gpc606_5 gpc633 (
      {stage0_16[67], stage0_16[68], stage0_16[69], stage0_16[70], stage0_16[71], stage0_16[72]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[44],stage1_18[47],stage1_17[91],stage1_16[152]}
   );
   gpc606_5 gpc634 (
      {stage0_16[73], stage0_16[74], stage0_16[75], stage0_16[76], stage0_16[77], stage0_16[78]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[45],stage1_18[48],stage1_17[92],stage1_16[153]}
   );
   gpc606_5 gpc635 (
      {stage0_16[79], stage0_16[80], stage0_16[81], stage0_16[82], stage0_16[83], stage0_16[84]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[46],stage1_18[49],stage1_17[93],stage1_16[154]}
   );
   gpc606_5 gpc636 (
      {stage0_16[85], stage0_16[86], stage0_16[87], stage0_16[88], stage0_16[89], stage0_16[90]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage1_20[4],stage1_19[47],stage1_18[50],stage1_17[94],stage1_16[155]}
   );
   gpc606_5 gpc637 (
      {stage0_16[91], stage0_16[92], stage0_16[93], stage0_16[94], stage0_16[95], stage0_16[96]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage1_20[5],stage1_19[48],stage1_18[51],stage1_17[95],stage1_16[156]}
   );
   gpc606_5 gpc638 (
      {stage0_16[97], stage0_16[98], stage0_16[99], stage0_16[100], stage0_16[101], stage0_16[102]},
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage1_20[6],stage1_19[49],stage1_18[52],stage1_17[96],stage1_16[157]}
   );
   gpc606_5 gpc639 (
      {stage0_16[103], stage0_16[104], stage0_16[105], stage0_16[106], stage0_16[107], stage0_16[108]},
      {stage0_18[42], stage0_18[43], stage0_18[44], stage0_18[45], stage0_18[46], stage0_18[47]},
      {stage1_20[7],stage1_19[50],stage1_18[53],stage1_17[97],stage1_16[158]}
   );
   gpc606_5 gpc640 (
      {stage0_16[109], stage0_16[110], stage0_16[111], stage0_16[112], stage0_16[113], stage0_16[114]},
      {stage0_18[48], stage0_18[49], stage0_18[50], stage0_18[51], stage0_18[52], stage0_18[53]},
      {stage1_20[8],stage1_19[51],stage1_18[54],stage1_17[98],stage1_16[159]}
   );
   gpc606_5 gpc641 (
      {stage0_16[115], stage0_16[116], stage0_16[117], stage0_16[118], stage0_16[119], stage0_16[120]},
      {stage0_18[54], stage0_18[55], stage0_18[56], stage0_18[57], stage0_18[58], stage0_18[59]},
      {stage1_20[9],stage1_19[52],stage1_18[55],stage1_17[99],stage1_16[160]}
   );
   gpc606_5 gpc642 (
      {stage0_16[121], stage0_16[122], stage0_16[123], stage0_16[124], stage0_16[125], stage0_16[126]},
      {stage0_18[60], stage0_18[61], stage0_18[62], stage0_18[63], stage0_18[64], stage0_18[65]},
      {stage1_20[10],stage1_19[53],stage1_18[56],stage1_17[100],stage1_16[161]}
   );
   gpc606_5 gpc643 (
      {stage0_16[127], stage0_16[128], stage0_16[129], stage0_16[130], stage0_16[131], stage0_16[132]},
      {stage0_18[66], stage0_18[67], stage0_18[68], stage0_18[69], stage0_18[70], stage0_18[71]},
      {stage1_20[11],stage1_19[54],stage1_18[57],stage1_17[101],stage1_16[162]}
   );
   gpc606_5 gpc644 (
      {stage0_16[133], stage0_16[134], stage0_16[135], stage0_16[136], stage0_16[137], stage0_16[138]},
      {stage0_18[72], stage0_18[73], stage0_18[74], stage0_18[75], stage0_18[76], stage0_18[77]},
      {stage1_20[12],stage1_19[55],stage1_18[58],stage1_17[102],stage1_16[163]}
   );
   gpc606_5 gpc645 (
      {stage0_16[139], stage0_16[140], stage0_16[141], stage0_16[142], stage0_16[143], stage0_16[144]},
      {stage0_18[78], stage0_18[79], stage0_18[80], stage0_18[81], stage0_18[82], stage0_18[83]},
      {stage1_20[13],stage1_19[56],stage1_18[59],stage1_17[103],stage1_16[164]}
   );
   gpc606_5 gpc646 (
      {stage0_16[145], stage0_16[146], stage0_16[147], stage0_16[148], stage0_16[149], stage0_16[150]},
      {stage0_18[84], stage0_18[85], stage0_18[86], stage0_18[87], stage0_18[88], stage0_18[89]},
      {stage1_20[14],stage1_19[57],stage1_18[60],stage1_17[104],stage1_16[165]}
   );
   gpc606_5 gpc647 (
      {stage0_16[151], stage0_16[152], stage0_16[153], stage0_16[154], stage0_16[155], stage0_16[156]},
      {stage0_18[90], stage0_18[91], stage0_18[92], stage0_18[93], stage0_18[94], stage0_18[95]},
      {stage1_20[15],stage1_19[58],stage1_18[61],stage1_17[105],stage1_16[166]}
   );
   gpc606_5 gpc648 (
      {stage0_16[157], stage0_16[158], stage0_16[159], stage0_16[160], stage0_16[161], stage0_16[162]},
      {stage0_18[96], stage0_18[97], stage0_18[98], stage0_18[99], stage0_18[100], stage0_18[101]},
      {stage1_20[16],stage1_19[59],stage1_18[62],stage1_17[106],stage1_16[167]}
   );
   gpc606_5 gpc649 (
      {stage0_16[163], stage0_16[164], stage0_16[165], stage0_16[166], stage0_16[167], stage0_16[168]},
      {stage0_18[102], stage0_18[103], stage0_18[104], stage0_18[105], stage0_18[106], stage0_18[107]},
      {stage1_20[17],stage1_19[60],stage1_18[63],stage1_17[107],stage1_16[168]}
   );
   gpc606_5 gpc650 (
      {stage0_16[169], stage0_16[170], stage0_16[171], stage0_16[172], stage0_16[173], stage0_16[174]},
      {stage0_18[108], stage0_18[109], stage0_18[110], stage0_18[111], stage0_18[112], stage0_18[113]},
      {stage1_20[18],stage1_19[61],stage1_18[64],stage1_17[108],stage1_16[169]}
   );
   gpc606_5 gpc651 (
      {stage0_16[175], stage0_16[176], stage0_16[177], stage0_16[178], stage0_16[179], stage0_16[180]},
      {stage0_18[114], stage0_18[115], stage0_18[116], stage0_18[117], stage0_18[118], stage0_18[119]},
      {stage1_20[19],stage1_19[62],stage1_18[65],stage1_17[109],stage1_16[170]}
   );
   gpc606_5 gpc652 (
      {stage0_16[181], stage0_16[182], stage0_16[183], stage0_16[184], stage0_16[185], stage0_16[186]},
      {stage0_18[120], stage0_18[121], stage0_18[122], stage0_18[123], stage0_18[124], stage0_18[125]},
      {stage1_20[20],stage1_19[63],stage1_18[66],stage1_17[110],stage1_16[171]}
   );
   gpc606_5 gpc653 (
      {stage0_16[187], stage0_16[188], stage0_16[189], stage0_16[190], stage0_16[191], stage0_16[192]},
      {stage0_18[126], stage0_18[127], stage0_18[128], stage0_18[129], stage0_18[130], stage0_18[131]},
      {stage1_20[21],stage1_19[64],stage1_18[67],stage1_17[111],stage1_16[172]}
   );
   gpc606_5 gpc654 (
      {stage0_16[193], stage0_16[194], stage0_16[195], stage0_16[196], stage0_16[197], stage0_16[198]},
      {stage0_18[132], stage0_18[133], stage0_18[134], stage0_18[135], stage0_18[136], stage0_18[137]},
      {stage1_20[22],stage1_19[65],stage1_18[68],stage1_17[112],stage1_16[173]}
   );
   gpc606_5 gpc655 (
      {stage0_16[199], stage0_16[200], stage0_16[201], stage0_16[202], stage0_16[203], stage0_16[204]},
      {stage0_18[138], stage0_18[139], stage0_18[140], stage0_18[141], stage0_18[142], stage0_18[143]},
      {stage1_20[23],stage1_19[66],stage1_18[69],stage1_17[113],stage1_16[174]}
   );
   gpc606_5 gpc656 (
      {stage0_16[205], stage0_16[206], stage0_16[207], stage0_16[208], stage0_16[209], stage0_16[210]},
      {stage0_18[144], stage0_18[145], stage0_18[146], stage0_18[147], stage0_18[148], stage0_18[149]},
      {stage1_20[24],stage1_19[67],stage1_18[70],stage1_17[114],stage1_16[175]}
   );
   gpc606_5 gpc657 (
      {stage0_16[211], stage0_16[212], stage0_16[213], stage0_16[214], stage0_16[215], stage0_16[216]},
      {stage0_18[150], stage0_18[151], stage0_18[152], stage0_18[153], stage0_18[154], stage0_18[155]},
      {stage1_20[25],stage1_19[68],stage1_18[71],stage1_17[115],stage1_16[176]}
   );
   gpc606_5 gpc658 (
      {stage0_16[217], stage0_16[218], stage0_16[219], stage0_16[220], stage0_16[221], stage0_16[222]},
      {stage0_18[156], stage0_18[157], stage0_18[158], stage0_18[159], stage0_18[160], stage0_18[161]},
      {stage1_20[26],stage1_19[69],stage1_18[72],stage1_17[116],stage1_16[177]}
   );
   gpc606_5 gpc659 (
      {stage0_16[223], stage0_16[224], stage0_16[225], stage0_16[226], stage0_16[227], stage0_16[228]},
      {stage0_18[162], stage0_18[163], stage0_18[164], stage0_18[165], stage0_18[166], stage0_18[167]},
      {stage1_20[27],stage1_19[70],stage1_18[73],stage1_17[117],stage1_16[178]}
   );
   gpc606_5 gpc660 (
      {stage0_16[229], stage0_16[230], stage0_16[231], stage0_16[232], stage0_16[233], stage0_16[234]},
      {stage0_18[168], stage0_18[169], stage0_18[170], stage0_18[171], stage0_18[172], stage0_18[173]},
      {stage1_20[28],stage1_19[71],stage1_18[74],stage1_17[118],stage1_16[179]}
   );
   gpc606_5 gpc661 (
      {stage0_16[235], stage0_16[236], stage0_16[237], stage0_16[238], stage0_16[239], stage0_16[240]},
      {stage0_18[174], stage0_18[175], stage0_18[176], stage0_18[177], stage0_18[178], stage0_18[179]},
      {stage1_20[29],stage1_19[72],stage1_18[75],stage1_17[119],stage1_16[180]}
   );
   gpc606_5 gpc662 (
      {stage0_16[241], stage0_16[242], stage0_16[243], stage0_16[244], stage0_16[245], stage0_16[246]},
      {stage0_18[180], stage0_18[181], stage0_18[182], stage0_18[183], stage0_18[184], stage0_18[185]},
      {stage1_20[30],stage1_19[73],stage1_18[76],stage1_17[120],stage1_16[181]}
   );
   gpc606_5 gpc663 (
      {stage0_16[247], stage0_16[248], stage0_16[249], stage0_16[250], stage0_16[251], stage0_16[252]},
      {stage0_18[186], stage0_18[187], stage0_18[188], stage0_18[189], stage0_18[190], stage0_18[191]},
      {stage1_20[31],stage1_19[74],stage1_18[77],stage1_17[121],stage1_16[182]}
   );
   gpc606_5 gpc664 (
      {stage0_16[253], stage0_16[254], stage0_16[255], stage0_16[256], stage0_16[257], stage0_16[258]},
      {stage0_18[192], stage0_18[193], stage0_18[194], stage0_18[195], stage0_18[196], stage0_18[197]},
      {stage1_20[32],stage1_19[75],stage1_18[78],stage1_17[122],stage1_16[183]}
   );
   gpc606_5 gpc665 (
      {stage0_16[259], stage0_16[260], stage0_16[261], stage0_16[262], stage0_16[263], stage0_16[264]},
      {stage0_18[198], stage0_18[199], stage0_18[200], stage0_18[201], stage0_18[202], stage0_18[203]},
      {stage1_20[33],stage1_19[76],stage1_18[79],stage1_17[123],stage1_16[184]}
   );
   gpc606_5 gpc666 (
      {stage0_16[265], stage0_16[266], stage0_16[267], stage0_16[268], stage0_16[269], stage0_16[270]},
      {stage0_18[204], stage0_18[205], stage0_18[206], stage0_18[207], stage0_18[208], stage0_18[209]},
      {stage1_20[34],stage1_19[77],stage1_18[80],stage1_17[124],stage1_16[185]}
   );
   gpc606_5 gpc667 (
      {stage0_16[271], stage0_16[272], stage0_16[273], stage0_16[274], stage0_16[275], stage0_16[276]},
      {stage0_18[210], stage0_18[211], stage0_18[212], stage0_18[213], stage0_18[214], stage0_18[215]},
      {stage1_20[35],stage1_19[78],stage1_18[81],stage1_17[125],stage1_16[186]}
   );
   gpc606_5 gpc668 (
      {stage0_16[277], stage0_16[278], stage0_16[279], stage0_16[280], stage0_16[281], stage0_16[282]},
      {stage0_18[216], stage0_18[217], stage0_18[218], stage0_18[219], stage0_18[220], stage0_18[221]},
      {stage1_20[36],stage1_19[79],stage1_18[82],stage1_17[126],stage1_16[187]}
   );
   gpc606_5 gpc669 (
      {stage0_16[283], stage0_16[284], stage0_16[285], stage0_16[286], stage0_16[287], stage0_16[288]},
      {stage0_18[222], stage0_18[223], stage0_18[224], stage0_18[225], stage0_18[226], stage0_18[227]},
      {stage1_20[37],stage1_19[80],stage1_18[83],stage1_17[127],stage1_16[188]}
   );
   gpc606_5 gpc670 (
      {stage0_16[289], stage0_16[290], stage0_16[291], stage0_16[292], stage0_16[293], stage0_16[294]},
      {stage0_18[228], stage0_18[229], stage0_18[230], stage0_18[231], stage0_18[232], stage0_18[233]},
      {stage1_20[38],stage1_19[81],stage1_18[84],stage1_17[128],stage1_16[189]}
   );
   gpc606_5 gpc671 (
      {stage0_16[295], stage0_16[296], stage0_16[297], stage0_16[298], stage0_16[299], stage0_16[300]},
      {stage0_18[234], stage0_18[235], stage0_18[236], stage0_18[237], stage0_18[238], stage0_18[239]},
      {stage1_20[39],stage1_19[82],stage1_18[85],stage1_17[129],stage1_16[190]}
   );
   gpc606_5 gpc672 (
      {stage0_16[301], stage0_16[302], stage0_16[303], stage0_16[304], stage0_16[305], stage0_16[306]},
      {stage0_18[240], stage0_18[241], stage0_18[242], stage0_18[243], stage0_18[244], stage0_18[245]},
      {stage1_20[40],stage1_19[83],stage1_18[86],stage1_17[130],stage1_16[191]}
   );
   gpc606_5 gpc673 (
      {stage0_16[307], stage0_16[308], stage0_16[309], stage0_16[310], stage0_16[311], stage0_16[312]},
      {stage0_18[246], stage0_18[247], stage0_18[248], stage0_18[249], stage0_18[250], stage0_18[251]},
      {stage1_20[41],stage1_19[84],stage1_18[87],stage1_17[131],stage1_16[192]}
   );
   gpc606_5 gpc674 (
      {stage0_16[313], stage0_16[314], stage0_16[315], stage0_16[316], stage0_16[317], stage0_16[318]},
      {stage0_18[252], stage0_18[253], stage0_18[254], stage0_18[255], stage0_18[256], stage0_18[257]},
      {stage1_20[42],stage1_19[85],stage1_18[88],stage1_17[132],stage1_16[193]}
   );
   gpc606_5 gpc675 (
      {stage0_16[319], stage0_16[320], stage0_16[321], stage0_16[322], stage0_16[323], stage0_16[324]},
      {stage0_18[258], stage0_18[259], stage0_18[260], stage0_18[261], stage0_18[262], stage0_18[263]},
      {stage1_20[43],stage1_19[86],stage1_18[89],stage1_17[133],stage1_16[194]}
   );
   gpc606_5 gpc676 (
      {stage0_16[325], stage0_16[326], stage0_16[327], stage0_16[328], stage0_16[329], stage0_16[330]},
      {stage0_18[264], stage0_18[265], stage0_18[266], stage0_18[267], stage0_18[268], stage0_18[269]},
      {stage1_20[44],stage1_19[87],stage1_18[90],stage1_17[134],stage1_16[195]}
   );
   gpc606_5 gpc677 (
      {stage0_16[331], stage0_16[332], stage0_16[333], stage0_16[334], stage0_16[335], stage0_16[336]},
      {stage0_18[270], stage0_18[271], stage0_18[272], stage0_18[273], stage0_18[274], stage0_18[275]},
      {stage1_20[45],stage1_19[88],stage1_18[91],stage1_17[135],stage1_16[196]}
   );
   gpc606_5 gpc678 (
      {stage0_16[337], stage0_16[338], stage0_16[339], stage0_16[340], stage0_16[341], stage0_16[342]},
      {stage0_18[276], stage0_18[277], stage0_18[278], stage0_18[279], stage0_18[280], stage0_18[281]},
      {stage1_20[46],stage1_19[89],stage1_18[92],stage1_17[136],stage1_16[197]}
   );
   gpc606_5 gpc679 (
      {stage0_16[343], stage0_16[344], stage0_16[345], stage0_16[346], stage0_16[347], stage0_16[348]},
      {stage0_18[282], stage0_18[283], stage0_18[284], stage0_18[285], stage0_18[286], stage0_18[287]},
      {stage1_20[47],stage1_19[90],stage1_18[93],stage1_17[137],stage1_16[198]}
   );
   gpc606_5 gpc680 (
      {stage0_16[349], stage0_16[350], stage0_16[351], stage0_16[352], stage0_16[353], stage0_16[354]},
      {stage0_18[288], stage0_18[289], stage0_18[290], stage0_18[291], stage0_18[292], stage0_18[293]},
      {stage1_20[48],stage1_19[91],stage1_18[94],stage1_17[138],stage1_16[199]}
   );
   gpc606_5 gpc681 (
      {stage0_16[355], stage0_16[356], stage0_16[357], stage0_16[358], stage0_16[359], stage0_16[360]},
      {stage0_18[294], stage0_18[295], stage0_18[296], stage0_18[297], stage0_18[298], stage0_18[299]},
      {stage1_20[49],stage1_19[92],stage1_18[95],stage1_17[139],stage1_16[200]}
   );
   gpc606_5 gpc682 (
      {stage0_16[361], stage0_16[362], stage0_16[363], stage0_16[364], stage0_16[365], stage0_16[366]},
      {stage0_18[300], stage0_18[301], stage0_18[302], stage0_18[303], stage0_18[304], stage0_18[305]},
      {stage1_20[50],stage1_19[93],stage1_18[96],stage1_17[140],stage1_16[201]}
   );
   gpc606_5 gpc683 (
      {stage0_16[367], stage0_16[368], stage0_16[369], stage0_16[370], stage0_16[371], stage0_16[372]},
      {stage0_18[306], stage0_18[307], stage0_18[308], stage0_18[309], stage0_18[310], stage0_18[311]},
      {stage1_20[51],stage1_19[94],stage1_18[97],stage1_17[141],stage1_16[202]}
   );
   gpc606_5 gpc684 (
      {stage0_16[373], stage0_16[374], stage0_16[375], stage0_16[376], stage0_16[377], stage0_16[378]},
      {stage0_18[312], stage0_18[313], stage0_18[314], stage0_18[315], stage0_18[316], stage0_18[317]},
      {stage1_20[52],stage1_19[95],stage1_18[98],stage1_17[142],stage1_16[203]}
   );
   gpc606_5 gpc685 (
      {stage0_16[379], stage0_16[380], stage0_16[381], stage0_16[382], stage0_16[383], stage0_16[384]},
      {stage0_18[318], stage0_18[319], stage0_18[320], stage0_18[321], stage0_18[322], stage0_18[323]},
      {stage1_20[53],stage1_19[96],stage1_18[99],stage1_17[143],stage1_16[204]}
   );
   gpc606_5 gpc686 (
      {stage0_16[385], stage0_16[386], stage0_16[387], stage0_16[388], stage0_16[389], stage0_16[390]},
      {stage0_18[324], stage0_18[325], stage0_18[326], stage0_18[327], stage0_18[328], stage0_18[329]},
      {stage1_20[54],stage1_19[97],stage1_18[100],stage1_17[144],stage1_16[205]}
   );
   gpc606_5 gpc687 (
      {stage0_16[391], stage0_16[392], stage0_16[393], stage0_16[394], stage0_16[395], stage0_16[396]},
      {stage0_18[330], stage0_18[331], stage0_18[332], stage0_18[333], stage0_18[334], stage0_18[335]},
      {stage1_20[55],stage1_19[98],stage1_18[101],stage1_17[145],stage1_16[206]}
   );
   gpc606_5 gpc688 (
      {stage0_16[397], stage0_16[398], stage0_16[399], stage0_16[400], stage0_16[401], stage0_16[402]},
      {stage0_18[336], stage0_18[337], stage0_18[338], stage0_18[339], stage0_18[340], stage0_18[341]},
      {stage1_20[56],stage1_19[99],stage1_18[102],stage1_17[146],stage1_16[207]}
   );
   gpc606_5 gpc689 (
      {stage0_16[403], stage0_16[404], stage0_16[405], stage0_16[406], stage0_16[407], stage0_16[408]},
      {stage0_18[342], stage0_18[343], stage0_18[344], stage0_18[345], stage0_18[346], stage0_18[347]},
      {stage1_20[57],stage1_19[100],stage1_18[103],stage1_17[147],stage1_16[208]}
   );
   gpc606_5 gpc690 (
      {stage0_16[409], stage0_16[410], stage0_16[411], stage0_16[412], stage0_16[413], stage0_16[414]},
      {stage0_18[348], stage0_18[349], stage0_18[350], stage0_18[351], stage0_18[352], stage0_18[353]},
      {stage1_20[58],stage1_19[101],stage1_18[104],stage1_17[148],stage1_16[209]}
   );
   gpc606_5 gpc691 (
      {stage0_16[415], stage0_16[416], stage0_16[417], stage0_16[418], stage0_16[419], stage0_16[420]},
      {stage0_18[354], stage0_18[355], stage0_18[356], stage0_18[357], stage0_18[358], stage0_18[359]},
      {stage1_20[59],stage1_19[102],stage1_18[105],stage1_17[149],stage1_16[210]}
   );
   gpc606_5 gpc692 (
      {stage0_16[421], stage0_16[422], stage0_16[423], stage0_16[424], stage0_16[425], stage0_16[426]},
      {stage0_18[360], stage0_18[361], stage0_18[362], stage0_18[363], stage0_18[364], stage0_18[365]},
      {stage1_20[60],stage1_19[103],stage1_18[106],stage1_17[150],stage1_16[211]}
   );
   gpc606_5 gpc693 (
      {stage0_16[427], stage0_16[428], stage0_16[429], stage0_16[430], stage0_16[431], stage0_16[432]},
      {stage0_18[366], stage0_18[367], stage0_18[368], stage0_18[369], stage0_18[370], stage0_18[371]},
      {stage1_20[61],stage1_19[104],stage1_18[107],stage1_17[151],stage1_16[212]}
   );
   gpc606_5 gpc694 (
      {stage0_16[433], stage0_16[434], stage0_16[435], stage0_16[436], stage0_16[437], stage0_16[438]},
      {stage0_18[372], stage0_18[373], stage0_18[374], stage0_18[375], stage0_18[376], stage0_18[377]},
      {stage1_20[62],stage1_19[105],stage1_18[108],stage1_17[152],stage1_16[213]}
   );
   gpc606_5 gpc695 (
      {stage0_16[439], stage0_16[440], stage0_16[441], stage0_16[442], stage0_16[443], stage0_16[444]},
      {stage0_18[378], stage0_18[379], stage0_18[380], stage0_18[381], stage0_18[382], stage0_18[383]},
      {stage1_20[63],stage1_19[106],stage1_18[109],stage1_17[153],stage1_16[214]}
   );
   gpc606_5 gpc696 (
      {stage0_16[445], stage0_16[446], stage0_16[447], stage0_16[448], stage0_16[449], stage0_16[450]},
      {stage0_18[384], stage0_18[385], stage0_18[386], stage0_18[387], stage0_18[388], stage0_18[389]},
      {stage1_20[64],stage1_19[107],stage1_18[110],stage1_17[154],stage1_16[215]}
   );
   gpc606_5 gpc697 (
      {stage0_16[451], stage0_16[452], stage0_16[453], stage0_16[454], stage0_16[455], stage0_16[456]},
      {stage0_18[390], stage0_18[391], stage0_18[392], stage0_18[393], stage0_18[394], stage0_18[395]},
      {stage1_20[65],stage1_19[108],stage1_18[111],stage1_17[155],stage1_16[216]}
   );
   gpc606_5 gpc698 (
      {stage0_16[457], stage0_16[458], stage0_16[459], stage0_16[460], stage0_16[461], stage0_16[462]},
      {stage0_18[396], stage0_18[397], stage0_18[398], stage0_18[399], stage0_18[400], stage0_18[401]},
      {stage1_20[66],stage1_19[109],stage1_18[112],stage1_17[156],stage1_16[217]}
   );
   gpc606_5 gpc699 (
      {stage0_16[463], stage0_16[464], stage0_16[465], stage0_16[466], stage0_16[467], stage0_16[468]},
      {stage0_18[402], stage0_18[403], stage0_18[404], stage0_18[405], stage0_18[406], stage0_18[407]},
      {stage1_20[67],stage1_19[110],stage1_18[113],stage1_17[157],stage1_16[218]}
   );
   gpc606_5 gpc700 (
      {stage0_16[469], stage0_16[470], stage0_16[471], stage0_16[472], stage0_16[473], stage0_16[474]},
      {stage0_18[408], stage0_18[409], stage0_18[410], stage0_18[411], stage0_18[412], stage0_18[413]},
      {stage1_20[68],stage1_19[111],stage1_18[114],stage1_17[158],stage1_16[219]}
   );
   gpc606_5 gpc701 (
      {stage0_16[475], stage0_16[476], stage0_16[477], stage0_16[478], stage0_16[479], stage0_16[480]},
      {stage0_18[414], stage0_18[415], stage0_18[416], stage0_18[417], stage0_18[418], stage0_18[419]},
      {stage1_20[69],stage1_19[112],stage1_18[115],stage1_17[159],stage1_16[220]}
   );
   gpc606_5 gpc702 (
      {stage0_16[481], stage0_16[482], stage0_16[483], stage0_16[484], stage0_16[485], 1'b0},
      {stage0_18[420], stage0_18[421], stage0_18[422], stage0_18[423], stage0_18[424], stage0_18[425]},
      {stage1_20[70],stage1_19[113],stage1_18[116],stage1_17[160],stage1_16[221]}
   );
   gpc606_5 gpc703 (
      {stage0_17[258], stage0_17[259], stage0_17[260], stage0_17[261], stage0_17[262], stage0_17[263]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[71],stage1_19[114],stage1_18[117],stage1_17[161]}
   );
   gpc606_5 gpc704 (
      {stage0_17[264], stage0_17[265], stage0_17[266], stage0_17[267], stage0_17[268], stage0_17[269]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[72],stage1_19[115],stage1_18[118],stage1_17[162]}
   );
   gpc606_5 gpc705 (
      {stage0_17[270], stage0_17[271], stage0_17[272], stage0_17[273], stage0_17[274], stage0_17[275]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[73],stage1_19[116],stage1_18[119],stage1_17[163]}
   );
   gpc606_5 gpc706 (
      {stage0_17[276], stage0_17[277], stage0_17[278], stage0_17[279], stage0_17[280], stage0_17[281]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[74],stage1_19[117],stage1_18[120],stage1_17[164]}
   );
   gpc606_5 gpc707 (
      {stage0_17[282], stage0_17[283], stage0_17[284], stage0_17[285], stage0_17[286], stage0_17[287]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[75],stage1_19[118],stage1_18[121],stage1_17[165]}
   );
   gpc606_5 gpc708 (
      {stage0_17[288], stage0_17[289], stage0_17[290], stage0_17[291], stage0_17[292], stage0_17[293]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[76],stage1_19[119],stage1_18[122],stage1_17[166]}
   );
   gpc606_5 gpc709 (
      {stage0_17[294], stage0_17[295], stage0_17[296], stage0_17[297], stage0_17[298], stage0_17[299]},
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage1_21[6],stage1_20[77],stage1_19[120],stage1_18[123],stage1_17[167]}
   );
   gpc606_5 gpc710 (
      {stage0_17[300], stage0_17[301], stage0_17[302], stage0_17[303], stage0_17[304], stage0_17[305]},
      {stage0_19[42], stage0_19[43], stage0_19[44], stage0_19[45], stage0_19[46], stage0_19[47]},
      {stage1_21[7],stage1_20[78],stage1_19[121],stage1_18[124],stage1_17[168]}
   );
   gpc606_5 gpc711 (
      {stage0_17[306], stage0_17[307], stage0_17[308], stage0_17[309], stage0_17[310], stage0_17[311]},
      {stage0_19[48], stage0_19[49], stage0_19[50], stage0_19[51], stage0_19[52], stage0_19[53]},
      {stage1_21[8],stage1_20[79],stage1_19[122],stage1_18[125],stage1_17[169]}
   );
   gpc606_5 gpc712 (
      {stage0_17[312], stage0_17[313], stage0_17[314], stage0_17[315], stage0_17[316], stage0_17[317]},
      {stage0_19[54], stage0_19[55], stage0_19[56], stage0_19[57], stage0_19[58], stage0_19[59]},
      {stage1_21[9],stage1_20[80],stage1_19[123],stage1_18[126],stage1_17[170]}
   );
   gpc606_5 gpc713 (
      {stage0_17[318], stage0_17[319], stage0_17[320], stage0_17[321], stage0_17[322], stage0_17[323]},
      {stage0_19[60], stage0_19[61], stage0_19[62], stage0_19[63], stage0_19[64], stage0_19[65]},
      {stage1_21[10],stage1_20[81],stage1_19[124],stage1_18[127],stage1_17[171]}
   );
   gpc606_5 gpc714 (
      {stage0_17[324], stage0_17[325], stage0_17[326], stage0_17[327], stage0_17[328], stage0_17[329]},
      {stage0_19[66], stage0_19[67], stage0_19[68], stage0_19[69], stage0_19[70], stage0_19[71]},
      {stage1_21[11],stage1_20[82],stage1_19[125],stage1_18[128],stage1_17[172]}
   );
   gpc606_5 gpc715 (
      {stage0_17[330], stage0_17[331], stage0_17[332], stage0_17[333], stage0_17[334], stage0_17[335]},
      {stage0_19[72], stage0_19[73], stage0_19[74], stage0_19[75], stage0_19[76], stage0_19[77]},
      {stage1_21[12],stage1_20[83],stage1_19[126],stage1_18[129],stage1_17[173]}
   );
   gpc606_5 gpc716 (
      {stage0_17[336], stage0_17[337], stage0_17[338], stage0_17[339], stage0_17[340], stage0_17[341]},
      {stage0_19[78], stage0_19[79], stage0_19[80], stage0_19[81], stage0_19[82], stage0_19[83]},
      {stage1_21[13],stage1_20[84],stage1_19[127],stage1_18[130],stage1_17[174]}
   );
   gpc606_5 gpc717 (
      {stage0_17[342], stage0_17[343], stage0_17[344], stage0_17[345], stage0_17[346], stage0_17[347]},
      {stage0_19[84], stage0_19[85], stage0_19[86], stage0_19[87], stage0_19[88], stage0_19[89]},
      {stage1_21[14],stage1_20[85],stage1_19[128],stage1_18[131],stage1_17[175]}
   );
   gpc606_5 gpc718 (
      {stage0_17[348], stage0_17[349], stage0_17[350], stage0_17[351], stage0_17[352], stage0_17[353]},
      {stage0_19[90], stage0_19[91], stage0_19[92], stage0_19[93], stage0_19[94], stage0_19[95]},
      {stage1_21[15],stage1_20[86],stage1_19[129],stage1_18[132],stage1_17[176]}
   );
   gpc606_5 gpc719 (
      {stage0_17[354], stage0_17[355], stage0_17[356], stage0_17[357], stage0_17[358], stage0_17[359]},
      {stage0_19[96], stage0_19[97], stage0_19[98], stage0_19[99], stage0_19[100], stage0_19[101]},
      {stage1_21[16],stage1_20[87],stage1_19[130],stage1_18[133],stage1_17[177]}
   );
   gpc606_5 gpc720 (
      {stage0_17[360], stage0_17[361], stage0_17[362], stage0_17[363], stage0_17[364], stage0_17[365]},
      {stage0_19[102], stage0_19[103], stage0_19[104], stage0_19[105], stage0_19[106], stage0_19[107]},
      {stage1_21[17],stage1_20[88],stage1_19[131],stage1_18[134],stage1_17[178]}
   );
   gpc606_5 gpc721 (
      {stage0_17[366], stage0_17[367], stage0_17[368], stage0_17[369], stage0_17[370], stage0_17[371]},
      {stage0_19[108], stage0_19[109], stage0_19[110], stage0_19[111], stage0_19[112], stage0_19[113]},
      {stage1_21[18],stage1_20[89],stage1_19[132],stage1_18[135],stage1_17[179]}
   );
   gpc606_5 gpc722 (
      {stage0_17[372], stage0_17[373], stage0_17[374], stage0_17[375], stage0_17[376], stage0_17[377]},
      {stage0_19[114], stage0_19[115], stage0_19[116], stage0_19[117], stage0_19[118], stage0_19[119]},
      {stage1_21[19],stage1_20[90],stage1_19[133],stage1_18[136],stage1_17[180]}
   );
   gpc606_5 gpc723 (
      {stage0_17[378], stage0_17[379], stage0_17[380], stage0_17[381], stage0_17[382], stage0_17[383]},
      {stage0_19[120], stage0_19[121], stage0_19[122], stage0_19[123], stage0_19[124], stage0_19[125]},
      {stage1_21[20],stage1_20[91],stage1_19[134],stage1_18[137],stage1_17[181]}
   );
   gpc606_5 gpc724 (
      {stage0_17[384], stage0_17[385], stage0_17[386], stage0_17[387], stage0_17[388], stage0_17[389]},
      {stage0_19[126], stage0_19[127], stage0_19[128], stage0_19[129], stage0_19[130], stage0_19[131]},
      {stage1_21[21],stage1_20[92],stage1_19[135],stage1_18[138],stage1_17[182]}
   );
   gpc606_5 gpc725 (
      {stage0_17[390], stage0_17[391], stage0_17[392], stage0_17[393], stage0_17[394], stage0_17[395]},
      {stage0_19[132], stage0_19[133], stage0_19[134], stage0_19[135], stage0_19[136], stage0_19[137]},
      {stage1_21[22],stage1_20[93],stage1_19[136],stage1_18[139],stage1_17[183]}
   );
   gpc606_5 gpc726 (
      {stage0_17[396], stage0_17[397], stage0_17[398], stage0_17[399], stage0_17[400], stage0_17[401]},
      {stage0_19[138], stage0_19[139], stage0_19[140], stage0_19[141], stage0_19[142], stage0_19[143]},
      {stage1_21[23],stage1_20[94],stage1_19[137],stage1_18[140],stage1_17[184]}
   );
   gpc606_5 gpc727 (
      {stage0_17[402], stage0_17[403], stage0_17[404], stage0_17[405], stage0_17[406], stage0_17[407]},
      {stage0_19[144], stage0_19[145], stage0_19[146], stage0_19[147], stage0_19[148], stage0_19[149]},
      {stage1_21[24],stage1_20[95],stage1_19[138],stage1_18[141],stage1_17[185]}
   );
   gpc606_5 gpc728 (
      {stage0_17[408], stage0_17[409], stage0_17[410], stage0_17[411], stage0_17[412], stage0_17[413]},
      {stage0_19[150], stage0_19[151], stage0_19[152], stage0_19[153], stage0_19[154], stage0_19[155]},
      {stage1_21[25],stage1_20[96],stage1_19[139],stage1_18[142],stage1_17[186]}
   );
   gpc606_5 gpc729 (
      {stage0_17[414], stage0_17[415], stage0_17[416], stage0_17[417], stage0_17[418], stage0_17[419]},
      {stage0_19[156], stage0_19[157], stage0_19[158], stage0_19[159], stage0_19[160], stage0_19[161]},
      {stage1_21[26],stage1_20[97],stage1_19[140],stage1_18[143],stage1_17[187]}
   );
   gpc606_5 gpc730 (
      {stage0_17[420], stage0_17[421], stage0_17[422], stage0_17[423], stage0_17[424], stage0_17[425]},
      {stage0_19[162], stage0_19[163], stage0_19[164], stage0_19[165], stage0_19[166], stage0_19[167]},
      {stage1_21[27],stage1_20[98],stage1_19[141],stage1_18[144],stage1_17[188]}
   );
   gpc606_5 gpc731 (
      {stage0_17[426], stage0_17[427], stage0_17[428], stage0_17[429], stage0_17[430], stage0_17[431]},
      {stage0_19[168], stage0_19[169], stage0_19[170], stage0_19[171], stage0_19[172], stage0_19[173]},
      {stage1_21[28],stage1_20[99],stage1_19[142],stage1_18[145],stage1_17[189]}
   );
   gpc606_5 gpc732 (
      {stage0_17[432], stage0_17[433], stage0_17[434], stage0_17[435], stage0_17[436], stage0_17[437]},
      {stage0_19[174], stage0_19[175], stage0_19[176], stage0_19[177], stage0_19[178], stage0_19[179]},
      {stage1_21[29],stage1_20[100],stage1_19[143],stage1_18[146],stage1_17[190]}
   );
   gpc606_5 gpc733 (
      {stage0_17[438], stage0_17[439], stage0_17[440], stage0_17[441], stage0_17[442], stage0_17[443]},
      {stage0_19[180], stage0_19[181], stage0_19[182], stage0_19[183], stage0_19[184], stage0_19[185]},
      {stage1_21[30],stage1_20[101],stage1_19[144],stage1_18[147],stage1_17[191]}
   );
   gpc606_5 gpc734 (
      {stage0_17[444], stage0_17[445], stage0_17[446], stage0_17[447], stage0_17[448], stage0_17[449]},
      {stage0_19[186], stage0_19[187], stage0_19[188], stage0_19[189], stage0_19[190], stage0_19[191]},
      {stage1_21[31],stage1_20[102],stage1_19[145],stage1_18[148],stage1_17[192]}
   );
   gpc615_5 gpc735 (
      {stage0_19[192], stage0_19[193], stage0_19[194], stage0_19[195], stage0_19[196]},
      {stage0_20[0]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[0],stage1_21[32],stage1_20[103],stage1_19[146]}
   );
   gpc615_5 gpc736 (
      {stage0_19[197], stage0_19[198], stage0_19[199], stage0_19[200], stage0_19[201]},
      {stage0_20[1]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[1],stage1_21[33],stage1_20[104],stage1_19[147]}
   );
   gpc615_5 gpc737 (
      {stage0_19[202], stage0_19[203], stage0_19[204], stage0_19[205], stage0_19[206]},
      {stage0_20[2]},
      {stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17]},
      {stage1_23[2],stage1_22[2],stage1_21[34],stage1_20[105],stage1_19[148]}
   );
   gpc615_5 gpc738 (
      {stage0_19[207], stage0_19[208], stage0_19[209], stage0_19[210], stage0_19[211]},
      {stage0_20[3]},
      {stage0_21[18], stage0_21[19], stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23]},
      {stage1_23[3],stage1_22[3],stage1_21[35],stage1_20[106],stage1_19[149]}
   );
   gpc615_5 gpc739 (
      {stage0_19[212], stage0_19[213], stage0_19[214], stage0_19[215], stage0_19[216]},
      {stage0_20[4]},
      {stage0_21[24], stage0_21[25], stage0_21[26], stage0_21[27], stage0_21[28], stage0_21[29]},
      {stage1_23[4],stage1_22[4],stage1_21[36],stage1_20[107],stage1_19[150]}
   );
   gpc615_5 gpc740 (
      {stage0_19[217], stage0_19[218], stage0_19[219], stage0_19[220], stage0_19[221]},
      {stage0_20[5]},
      {stage0_21[30], stage0_21[31], stage0_21[32], stage0_21[33], stage0_21[34], stage0_21[35]},
      {stage1_23[5],stage1_22[5],stage1_21[37],stage1_20[108],stage1_19[151]}
   );
   gpc615_5 gpc741 (
      {stage0_19[222], stage0_19[223], stage0_19[224], stage0_19[225], stage0_19[226]},
      {stage0_20[6]},
      {stage0_21[36], stage0_21[37], stage0_21[38], stage0_21[39], stage0_21[40], stage0_21[41]},
      {stage1_23[6],stage1_22[6],stage1_21[38],stage1_20[109],stage1_19[152]}
   );
   gpc615_5 gpc742 (
      {stage0_19[227], stage0_19[228], stage0_19[229], stage0_19[230], stage0_19[231]},
      {stage0_20[7]},
      {stage0_21[42], stage0_21[43], stage0_21[44], stage0_21[45], stage0_21[46], stage0_21[47]},
      {stage1_23[7],stage1_22[7],stage1_21[39],stage1_20[110],stage1_19[153]}
   );
   gpc615_5 gpc743 (
      {stage0_19[232], stage0_19[233], stage0_19[234], stage0_19[235], stage0_19[236]},
      {stage0_20[8]},
      {stage0_21[48], stage0_21[49], stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53]},
      {stage1_23[8],stage1_22[8],stage1_21[40],stage1_20[111],stage1_19[154]}
   );
   gpc615_5 gpc744 (
      {stage0_19[237], stage0_19[238], stage0_19[239], stage0_19[240], stage0_19[241]},
      {stage0_20[9]},
      {stage0_21[54], stage0_21[55], stage0_21[56], stage0_21[57], stage0_21[58], stage0_21[59]},
      {stage1_23[9],stage1_22[9],stage1_21[41],stage1_20[112],stage1_19[155]}
   );
   gpc615_5 gpc745 (
      {stage0_19[242], stage0_19[243], stage0_19[244], stage0_19[245], stage0_19[246]},
      {stage0_20[10]},
      {stage0_21[60], stage0_21[61], stage0_21[62], stage0_21[63], stage0_21[64], stage0_21[65]},
      {stage1_23[10],stage1_22[10],stage1_21[42],stage1_20[113],stage1_19[156]}
   );
   gpc615_5 gpc746 (
      {stage0_19[247], stage0_19[248], stage0_19[249], stage0_19[250], stage0_19[251]},
      {stage0_20[11]},
      {stage0_21[66], stage0_21[67], stage0_21[68], stage0_21[69], stage0_21[70], stage0_21[71]},
      {stage1_23[11],stage1_22[11],stage1_21[43],stage1_20[114],stage1_19[157]}
   );
   gpc615_5 gpc747 (
      {stage0_19[252], stage0_19[253], stage0_19[254], stage0_19[255], stage0_19[256]},
      {stage0_20[12]},
      {stage0_21[72], stage0_21[73], stage0_21[74], stage0_21[75], stage0_21[76], stage0_21[77]},
      {stage1_23[12],stage1_22[12],stage1_21[44],stage1_20[115],stage1_19[158]}
   );
   gpc615_5 gpc748 (
      {stage0_19[257], stage0_19[258], stage0_19[259], stage0_19[260], stage0_19[261]},
      {stage0_20[13]},
      {stage0_21[78], stage0_21[79], stage0_21[80], stage0_21[81], stage0_21[82], stage0_21[83]},
      {stage1_23[13],stage1_22[13],stage1_21[45],stage1_20[116],stage1_19[159]}
   );
   gpc615_5 gpc749 (
      {stage0_19[262], stage0_19[263], stage0_19[264], stage0_19[265], stage0_19[266]},
      {stage0_20[14]},
      {stage0_21[84], stage0_21[85], stage0_21[86], stage0_21[87], stage0_21[88], stage0_21[89]},
      {stage1_23[14],stage1_22[14],stage1_21[46],stage1_20[117],stage1_19[160]}
   );
   gpc615_5 gpc750 (
      {stage0_19[267], stage0_19[268], stage0_19[269], stage0_19[270], stage0_19[271]},
      {stage0_20[15]},
      {stage0_21[90], stage0_21[91], stage0_21[92], stage0_21[93], stage0_21[94], stage0_21[95]},
      {stage1_23[15],stage1_22[15],stage1_21[47],stage1_20[118],stage1_19[161]}
   );
   gpc615_5 gpc751 (
      {stage0_19[272], stage0_19[273], stage0_19[274], stage0_19[275], stage0_19[276]},
      {stage0_20[16]},
      {stage0_21[96], stage0_21[97], stage0_21[98], stage0_21[99], stage0_21[100], stage0_21[101]},
      {stage1_23[16],stage1_22[16],stage1_21[48],stage1_20[119],stage1_19[162]}
   );
   gpc615_5 gpc752 (
      {stage0_19[277], stage0_19[278], stage0_19[279], stage0_19[280], stage0_19[281]},
      {stage0_20[17]},
      {stage0_21[102], stage0_21[103], stage0_21[104], stage0_21[105], stage0_21[106], stage0_21[107]},
      {stage1_23[17],stage1_22[17],stage1_21[49],stage1_20[120],stage1_19[163]}
   );
   gpc615_5 gpc753 (
      {stage0_19[282], stage0_19[283], stage0_19[284], stage0_19[285], stage0_19[286]},
      {stage0_20[18]},
      {stage0_21[108], stage0_21[109], stage0_21[110], stage0_21[111], stage0_21[112], stage0_21[113]},
      {stage1_23[18],stage1_22[18],stage1_21[50],stage1_20[121],stage1_19[164]}
   );
   gpc615_5 gpc754 (
      {stage0_19[287], stage0_19[288], stage0_19[289], stage0_19[290], stage0_19[291]},
      {stage0_20[19]},
      {stage0_21[114], stage0_21[115], stage0_21[116], stage0_21[117], stage0_21[118], stage0_21[119]},
      {stage1_23[19],stage1_22[19],stage1_21[51],stage1_20[122],stage1_19[165]}
   );
   gpc615_5 gpc755 (
      {stage0_19[292], stage0_19[293], stage0_19[294], stage0_19[295], stage0_19[296]},
      {stage0_20[20]},
      {stage0_21[120], stage0_21[121], stage0_21[122], stage0_21[123], stage0_21[124], stage0_21[125]},
      {stage1_23[20],stage1_22[20],stage1_21[52],stage1_20[123],stage1_19[166]}
   );
   gpc615_5 gpc756 (
      {stage0_19[297], stage0_19[298], stage0_19[299], stage0_19[300], stage0_19[301]},
      {stage0_20[21]},
      {stage0_21[126], stage0_21[127], stage0_21[128], stage0_21[129], stage0_21[130], stage0_21[131]},
      {stage1_23[21],stage1_22[21],stage1_21[53],stage1_20[124],stage1_19[167]}
   );
   gpc615_5 gpc757 (
      {stage0_19[302], stage0_19[303], stage0_19[304], stage0_19[305], stage0_19[306]},
      {stage0_20[22]},
      {stage0_21[132], stage0_21[133], stage0_21[134], stage0_21[135], stage0_21[136], stage0_21[137]},
      {stage1_23[22],stage1_22[22],stage1_21[54],stage1_20[125],stage1_19[168]}
   );
   gpc615_5 gpc758 (
      {stage0_19[307], stage0_19[308], stage0_19[309], stage0_19[310], stage0_19[311]},
      {stage0_20[23]},
      {stage0_21[138], stage0_21[139], stage0_21[140], stage0_21[141], stage0_21[142], stage0_21[143]},
      {stage1_23[23],stage1_22[23],stage1_21[55],stage1_20[126],stage1_19[169]}
   );
   gpc615_5 gpc759 (
      {stage0_19[312], stage0_19[313], stage0_19[314], stage0_19[315], stage0_19[316]},
      {stage0_20[24]},
      {stage0_21[144], stage0_21[145], stage0_21[146], stage0_21[147], stage0_21[148], stage0_21[149]},
      {stage1_23[24],stage1_22[24],stage1_21[56],stage1_20[127],stage1_19[170]}
   );
   gpc615_5 gpc760 (
      {stage0_19[317], stage0_19[318], stage0_19[319], stage0_19[320], stage0_19[321]},
      {stage0_20[25]},
      {stage0_21[150], stage0_21[151], stage0_21[152], stage0_21[153], stage0_21[154], stage0_21[155]},
      {stage1_23[25],stage1_22[25],stage1_21[57],stage1_20[128],stage1_19[171]}
   );
   gpc615_5 gpc761 (
      {stage0_19[322], stage0_19[323], stage0_19[324], stage0_19[325], stage0_19[326]},
      {stage0_20[26]},
      {stage0_21[156], stage0_21[157], stage0_21[158], stage0_21[159], stage0_21[160], stage0_21[161]},
      {stage1_23[26],stage1_22[26],stage1_21[58],stage1_20[129],stage1_19[172]}
   );
   gpc615_5 gpc762 (
      {stage0_19[327], stage0_19[328], stage0_19[329], stage0_19[330], stage0_19[331]},
      {stage0_20[27]},
      {stage0_21[162], stage0_21[163], stage0_21[164], stage0_21[165], stage0_21[166], stage0_21[167]},
      {stage1_23[27],stage1_22[27],stage1_21[59],stage1_20[130],stage1_19[173]}
   );
   gpc615_5 gpc763 (
      {stage0_19[332], stage0_19[333], stage0_19[334], stage0_19[335], stage0_19[336]},
      {stage0_20[28]},
      {stage0_21[168], stage0_21[169], stage0_21[170], stage0_21[171], stage0_21[172], stage0_21[173]},
      {stage1_23[28],stage1_22[28],stage1_21[60],stage1_20[131],stage1_19[174]}
   );
   gpc615_5 gpc764 (
      {stage0_19[337], stage0_19[338], stage0_19[339], stage0_19[340], stage0_19[341]},
      {stage0_20[29]},
      {stage0_21[174], stage0_21[175], stage0_21[176], stage0_21[177], stage0_21[178], stage0_21[179]},
      {stage1_23[29],stage1_22[29],stage1_21[61],stage1_20[132],stage1_19[175]}
   );
   gpc615_5 gpc765 (
      {stage0_19[342], stage0_19[343], stage0_19[344], stage0_19[345], stage0_19[346]},
      {stage0_20[30]},
      {stage0_21[180], stage0_21[181], stage0_21[182], stage0_21[183], stage0_21[184], stage0_21[185]},
      {stage1_23[30],stage1_22[30],stage1_21[62],stage1_20[133],stage1_19[176]}
   );
   gpc615_5 gpc766 (
      {stage0_19[347], stage0_19[348], stage0_19[349], stage0_19[350], stage0_19[351]},
      {stage0_20[31]},
      {stage0_21[186], stage0_21[187], stage0_21[188], stage0_21[189], stage0_21[190], stage0_21[191]},
      {stage1_23[31],stage1_22[31],stage1_21[63],stage1_20[134],stage1_19[177]}
   );
   gpc615_5 gpc767 (
      {stage0_19[352], stage0_19[353], stage0_19[354], stage0_19[355], stage0_19[356]},
      {stage0_20[32]},
      {stage0_21[192], stage0_21[193], stage0_21[194], stage0_21[195], stage0_21[196], stage0_21[197]},
      {stage1_23[32],stage1_22[32],stage1_21[64],stage1_20[135],stage1_19[178]}
   );
   gpc615_5 gpc768 (
      {stage0_19[357], stage0_19[358], stage0_19[359], stage0_19[360], stage0_19[361]},
      {stage0_20[33]},
      {stage0_21[198], stage0_21[199], stage0_21[200], stage0_21[201], stage0_21[202], stage0_21[203]},
      {stage1_23[33],stage1_22[33],stage1_21[65],stage1_20[136],stage1_19[179]}
   );
   gpc615_5 gpc769 (
      {stage0_19[362], stage0_19[363], stage0_19[364], stage0_19[365], stage0_19[366]},
      {stage0_20[34]},
      {stage0_21[204], stage0_21[205], stage0_21[206], stage0_21[207], stage0_21[208], stage0_21[209]},
      {stage1_23[34],stage1_22[34],stage1_21[66],stage1_20[137],stage1_19[180]}
   );
   gpc615_5 gpc770 (
      {stage0_19[367], stage0_19[368], stage0_19[369], stage0_19[370], stage0_19[371]},
      {stage0_20[35]},
      {stage0_21[210], stage0_21[211], stage0_21[212], stage0_21[213], stage0_21[214], stage0_21[215]},
      {stage1_23[35],stage1_22[35],stage1_21[67],stage1_20[138],stage1_19[181]}
   );
   gpc615_5 gpc771 (
      {stage0_19[372], stage0_19[373], stage0_19[374], stage0_19[375], stage0_19[376]},
      {stage0_20[36]},
      {stage0_21[216], stage0_21[217], stage0_21[218], stage0_21[219], stage0_21[220], stage0_21[221]},
      {stage1_23[36],stage1_22[36],stage1_21[68],stage1_20[139],stage1_19[182]}
   );
   gpc615_5 gpc772 (
      {stage0_19[377], stage0_19[378], stage0_19[379], stage0_19[380], stage0_19[381]},
      {stage0_20[37]},
      {stage0_21[222], stage0_21[223], stage0_21[224], stage0_21[225], stage0_21[226], stage0_21[227]},
      {stage1_23[37],stage1_22[37],stage1_21[69],stage1_20[140],stage1_19[183]}
   );
   gpc615_5 gpc773 (
      {stage0_19[382], stage0_19[383], stage0_19[384], stage0_19[385], stage0_19[386]},
      {stage0_20[38]},
      {stage0_21[228], stage0_21[229], stage0_21[230], stage0_21[231], stage0_21[232], stage0_21[233]},
      {stage1_23[38],stage1_22[38],stage1_21[70],stage1_20[141],stage1_19[184]}
   );
   gpc615_5 gpc774 (
      {stage0_19[387], stage0_19[388], stage0_19[389], stage0_19[390], stage0_19[391]},
      {stage0_20[39]},
      {stage0_21[234], stage0_21[235], stage0_21[236], stage0_21[237], stage0_21[238], stage0_21[239]},
      {stage1_23[39],stage1_22[39],stage1_21[71],stage1_20[142],stage1_19[185]}
   );
   gpc615_5 gpc775 (
      {stage0_19[392], stage0_19[393], stage0_19[394], stage0_19[395], stage0_19[396]},
      {stage0_20[40]},
      {stage0_21[240], stage0_21[241], stage0_21[242], stage0_21[243], stage0_21[244], stage0_21[245]},
      {stage1_23[40],stage1_22[40],stage1_21[72],stage1_20[143],stage1_19[186]}
   );
   gpc1343_5 gpc776 (
      {stage0_20[41], stage0_20[42], stage0_20[43]},
      {stage0_21[246], stage0_21[247], stage0_21[248], stage0_21[249]},
      {stage0_22[0], stage0_22[1], stage0_22[2]},
      {stage0_23[0]},
      {stage1_24[0],stage1_23[41],stage1_22[41],stage1_21[73],stage1_20[144]}
   );
   gpc1163_5 gpc777 (
      {stage0_20[44], stage0_20[45], stage0_20[46]},
      {stage0_21[250], stage0_21[251], stage0_21[252], stage0_21[253], stage0_21[254], stage0_21[255]},
      {stage0_22[3]},
      {stage0_23[1]},
      {stage1_24[1],stage1_23[42],stage1_22[42],stage1_21[74],stage1_20[145]}
   );
   gpc1163_5 gpc778 (
      {stage0_20[47], stage0_20[48], stage0_20[49]},
      {stage0_21[256], stage0_21[257], stage0_21[258], stage0_21[259], stage0_21[260], stage0_21[261]},
      {stage0_22[4]},
      {stage0_23[2]},
      {stage1_24[2],stage1_23[43],stage1_22[43],stage1_21[75],stage1_20[146]}
   );
   gpc1163_5 gpc779 (
      {stage0_20[50], stage0_20[51], stage0_20[52]},
      {stage0_21[262], stage0_21[263], stage0_21[264], stage0_21[265], stage0_21[266], stage0_21[267]},
      {stage0_22[5]},
      {stage0_23[3]},
      {stage1_24[3],stage1_23[44],stage1_22[44],stage1_21[76],stage1_20[147]}
   );
   gpc1163_5 gpc780 (
      {stage0_20[53], stage0_20[54], stage0_20[55]},
      {stage0_21[268], stage0_21[269], stage0_21[270], stage0_21[271], stage0_21[272], stage0_21[273]},
      {stage0_22[6]},
      {stage0_23[4]},
      {stage1_24[4],stage1_23[45],stage1_22[45],stage1_21[77],stage1_20[148]}
   );
   gpc1163_5 gpc781 (
      {stage0_20[56], stage0_20[57], stage0_20[58]},
      {stage0_21[274], stage0_21[275], stage0_21[276], stage0_21[277], stage0_21[278], stage0_21[279]},
      {stage0_22[7]},
      {stage0_23[5]},
      {stage1_24[5],stage1_23[46],stage1_22[46],stage1_21[78],stage1_20[149]}
   );
   gpc1163_5 gpc782 (
      {stage0_20[59], stage0_20[60], stage0_20[61]},
      {stage0_21[280], stage0_21[281], stage0_21[282], stage0_21[283], stage0_21[284], stage0_21[285]},
      {stage0_22[8]},
      {stage0_23[6]},
      {stage1_24[6],stage1_23[47],stage1_22[47],stage1_21[79],stage1_20[150]}
   );
   gpc606_5 gpc783 (
      {stage0_20[62], stage0_20[63], stage0_20[64], stage0_20[65], stage0_20[66], stage0_20[67]},
      {stage0_22[9], stage0_22[10], stage0_22[11], stage0_22[12], stage0_22[13], stage0_22[14]},
      {stage1_24[7],stage1_23[48],stage1_22[48],stage1_21[80],stage1_20[151]}
   );
   gpc606_5 gpc784 (
      {stage0_20[68], stage0_20[69], stage0_20[70], stage0_20[71], stage0_20[72], stage0_20[73]},
      {stage0_22[15], stage0_22[16], stage0_22[17], stage0_22[18], stage0_22[19], stage0_22[20]},
      {stage1_24[8],stage1_23[49],stage1_22[49],stage1_21[81],stage1_20[152]}
   );
   gpc606_5 gpc785 (
      {stage0_20[74], stage0_20[75], stage0_20[76], stage0_20[77], stage0_20[78], stage0_20[79]},
      {stage0_22[21], stage0_22[22], stage0_22[23], stage0_22[24], stage0_22[25], stage0_22[26]},
      {stage1_24[9],stage1_23[50],stage1_22[50],stage1_21[82],stage1_20[153]}
   );
   gpc606_5 gpc786 (
      {stage0_20[80], stage0_20[81], stage0_20[82], stage0_20[83], stage0_20[84], stage0_20[85]},
      {stage0_22[27], stage0_22[28], stage0_22[29], stage0_22[30], stage0_22[31], stage0_22[32]},
      {stage1_24[10],stage1_23[51],stage1_22[51],stage1_21[83],stage1_20[154]}
   );
   gpc606_5 gpc787 (
      {stage0_20[86], stage0_20[87], stage0_20[88], stage0_20[89], stage0_20[90], stage0_20[91]},
      {stage0_22[33], stage0_22[34], stage0_22[35], stage0_22[36], stage0_22[37], stage0_22[38]},
      {stage1_24[11],stage1_23[52],stage1_22[52],stage1_21[84],stage1_20[155]}
   );
   gpc606_5 gpc788 (
      {stage0_20[92], stage0_20[93], stage0_20[94], stage0_20[95], stage0_20[96], stage0_20[97]},
      {stage0_22[39], stage0_22[40], stage0_22[41], stage0_22[42], stage0_22[43], stage0_22[44]},
      {stage1_24[12],stage1_23[53],stage1_22[53],stage1_21[85],stage1_20[156]}
   );
   gpc606_5 gpc789 (
      {stage0_20[98], stage0_20[99], stage0_20[100], stage0_20[101], stage0_20[102], stage0_20[103]},
      {stage0_22[45], stage0_22[46], stage0_22[47], stage0_22[48], stage0_22[49], stage0_22[50]},
      {stage1_24[13],stage1_23[54],stage1_22[54],stage1_21[86],stage1_20[157]}
   );
   gpc606_5 gpc790 (
      {stage0_20[104], stage0_20[105], stage0_20[106], stage0_20[107], stage0_20[108], stage0_20[109]},
      {stage0_22[51], stage0_22[52], stage0_22[53], stage0_22[54], stage0_22[55], stage0_22[56]},
      {stage1_24[14],stage1_23[55],stage1_22[55],stage1_21[87],stage1_20[158]}
   );
   gpc606_5 gpc791 (
      {stage0_20[110], stage0_20[111], stage0_20[112], stage0_20[113], stage0_20[114], stage0_20[115]},
      {stage0_22[57], stage0_22[58], stage0_22[59], stage0_22[60], stage0_22[61], stage0_22[62]},
      {stage1_24[15],stage1_23[56],stage1_22[56],stage1_21[88],stage1_20[159]}
   );
   gpc606_5 gpc792 (
      {stage0_20[116], stage0_20[117], stage0_20[118], stage0_20[119], stage0_20[120], stage0_20[121]},
      {stage0_22[63], stage0_22[64], stage0_22[65], stage0_22[66], stage0_22[67], stage0_22[68]},
      {stage1_24[16],stage1_23[57],stage1_22[57],stage1_21[89],stage1_20[160]}
   );
   gpc606_5 gpc793 (
      {stage0_20[122], stage0_20[123], stage0_20[124], stage0_20[125], stage0_20[126], stage0_20[127]},
      {stage0_22[69], stage0_22[70], stage0_22[71], stage0_22[72], stage0_22[73], stage0_22[74]},
      {stage1_24[17],stage1_23[58],stage1_22[58],stage1_21[90],stage1_20[161]}
   );
   gpc606_5 gpc794 (
      {stage0_20[128], stage0_20[129], stage0_20[130], stage0_20[131], stage0_20[132], stage0_20[133]},
      {stage0_22[75], stage0_22[76], stage0_22[77], stage0_22[78], stage0_22[79], stage0_22[80]},
      {stage1_24[18],stage1_23[59],stage1_22[59],stage1_21[91],stage1_20[162]}
   );
   gpc606_5 gpc795 (
      {stage0_20[134], stage0_20[135], stage0_20[136], stage0_20[137], stage0_20[138], stage0_20[139]},
      {stage0_22[81], stage0_22[82], stage0_22[83], stage0_22[84], stage0_22[85], stage0_22[86]},
      {stage1_24[19],stage1_23[60],stage1_22[60],stage1_21[92],stage1_20[163]}
   );
   gpc606_5 gpc796 (
      {stage0_20[140], stage0_20[141], stage0_20[142], stage0_20[143], stage0_20[144], stage0_20[145]},
      {stage0_22[87], stage0_22[88], stage0_22[89], stage0_22[90], stage0_22[91], stage0_22[92]},
      {stage1_24[20],stage1_23[61],stage1_22[61],stage1_21[93],stage1_20[164]}
   );
   gpc606_5 gpc797 (
      {stage0_20[146], stage0_20[147], stage0_20[148], stage0_20[149], stage0_20[150], stage0_20[151]},
      {stage0_22[93], stage0_22[94], stage0_22[95], stage0_22[96], stage0_22[97], stage0_22[98]},
      {stage1_24[21],stage1_23[62],stage1_22[62],stage1_21[94],stage1_20[165]}
   );
   gpc606_5 gpc798 (
      {stage0_20[152], stage0_20[153], stage0_20[154], stage0_20[155], stage0_20[156], stage0_20[157]},
      {stage0_22[99], stage0_22[100], stage0_22[101], stage0_22[102], stage0_22[103], stage0_22[104]},
      {stage1_24[22],stage1_23[63],stage1_22[63],stage1_21[95],stage1_20[166]}
   );
   gpc606_5 gpc799 (
      {stage0_20[158], stage0_20[159], stage0_20[160], stage0_20[161], stage0_20[162], stage0_20[163]},
      {stage0_22[105], stage0_22[106], stage0_22[107], stage0_22[108], stage0_22[109], stage0_22[110]},
      {stage1_24[23],stage1_23[64],stage1_22[64],stage1_21[96],stage1_20[167]}
   );
   gpc606_5 gpc800 (
      {stage0_20[164], stage0_20[165], stage0_20[166], stage0_20[167], stage0_20[168], stage0_20[169]},
      {stage0_22[111], stage0_22[112], stage0_22[113], stage0_22[114], stage0_22[115], stage0_22[116]},
      {stage1_24[24],stage1_23[65],stage1_22[65],stage1_21[97],stage1_20[168]}
   );
   gpc606_5 gpc801 (
      {stage0_20[170], stage0_20[171], stage0_20[172], stage0_20[173], stage0_20[174], stage0_20[175]},
      {stage0_22[117], stage0_22[118], stage0_22[119], stage0_22[120], stage0_22[121], stage0_22[122]},
      {stage1_24[25],stage1_23[66],stage1_22[66],stage1_21[98],stage1_20[169]}
   );
   gpc606_5 gpc802 (
      {stage0_20[176], stage0_20[177], stage0_20[178], stage0_20[179], stage0_20[180], stage0_20[181]},
      {stage0_22[123], stage0_22[124], stage0_22[125], stage0_22[126], stage0_22[127], stage0_22[128]},
      {stage1_24[26],stage1_23[67],stage1_22[67],stage1_21[99],stage1_20[170]}
   );
   gpc606_5 gpc803 (
      {stage0_20[182], stage0_20[183], stage0_20[184], stage0_20[185], stage0_20[186], stage0_20[187]},
      {stage0_22[129], stage0_22[130], stage0_22[131], stage0_22[132], stage0_22[133], stage0_22[134]},
      {stage1_24[27],stage1_23[68],stage1_22[68],stage1_21[100],stage1_20[171]}
   );
   gpc606_5 gpc804 (
      {stage0_20[188], stage0_20[189], stage0_20[190], stage0_20[191], stage0_20[192], stage0_20[193]},
      {stage0_22[135], stage0_22[136], stage0_22[137], stage0_22[138], stage0_22[139], stage0_22[140]},
      {stage1_24[28],stage1_23[69],stage1_22[69],stage1_21[101],stage1_20[172]}
   );
   gpc606_5 gpc805 (
      {stage0_20[194], stage0_20[195], stage0_20[196], stage0_20[197], stage0_20[198], stage0_20[199]},
      {stage0_22[141], stage0_22[142], stage0_22[143], stage0_22[144], stage0_22[145], stage0_22[146]},
      {stage1_24[29],stage1_23[70],stage1_22[70],stage1_21[102],stage1_20[173]}
   );
   gpc606_5 gpc806 (
      {stage0_20[200], stage0_20[201], stage0_20[202], stage0_20[203], stage0_20[204], stage0_20[205]},
      {stage0_22[147], stage0_22[148], stage0_22[149], stage0_22[150], stage0_22[151], stage0_22[152]},
      {stage1_24[30],stage1_23[71],stage1_22[71],stage1_21[103],stage1_20[174]}
   );
   gpc606_5 gpc807 (
      {stage0_20[206], stage0_20[207], stage0_20[208], stage0_20[209], stage0_20[210], stage0_20[211]},
      {stage0_22[153], stage0_22[154], stage0_22[155], stage0_22[156], stage0_22[157], stage0_22[158]},
      {stage1_24[31],stage1_23[72],stage1_22[72],stage1_21[104],stage1_20[175]}
   );
   gpc606_5 gpc808 (
      {stage0_20[212], stage0_20[213], stage0_20[214], stage0_20[215], stage0_20[216], stage0_20[217]},
      {stage0_22[159], stage0_22[160], stage0_22[161], stage0_22[162], stage0_22[163], stage0_22[164]},
      {stage1_24[32],stage1_23[73],stage1_22[73],stage1_21[105],stage1_20[176]}
   );
   gpc606_5 gpc809 (
      {stage0_20[218], stage0_20[219], stage0_20[220], stage0_20[221], stage0_20[222], stage0_20[223]},
      {stage0_22[165], stage0_22[166], stage0_22[167], stage0_22[168], stage0_22[169], stage0_22[170]},
      {stage1_24[33],stage1_23[74],stage1_22[74],stage1_21[106],stage1_20[177]}
   );
   gpc606_5 gpc810 (
      {stage0_20[224], stage0_20[225], stage0_20[226], stage0_20[227], stage0_20[228], stage0_20[229]},
      {stage0_22[171], stage0_22[172], stage0_22[173], stage0_22[174], stage0_22[175], stage0_22[176]},
      {stage1_24[34],stage1_23[75],stage1_22[75],stage1_21[107],stage1_20[178]}
   );
   gpc606_5 gpc811 (
      {stage0_20[230], stage0_20[231], stage0_20[232], stage0_20[233], stage0_20[234], stage0_20[235]},
      {stage0_22[177], stage0_22[178], stage0_22[179], stage0_22[180], stage0_22[181], stage0_22[182]},
      {stage1_24[35],stage1_23[76],stage1_22[76],stage1_21[108],stage1_20[179]}
   );
   gpc606_5 gpc812 (
      {stage0_20[236], stage0_20[237], stage0_20[238], stage0_20[239], stage0_20[240], stage0_20[241]},
      {stage0_22[183], stage0_22[184], stage0_22[185], stage0_22[186], stage0_22[187], stage0_22[188]},
      {stage1_24[36],stage1_23[77],stage1_22[77],stage1_21[109],stage1_20[180]}
   );
   gpc606_5 gpc813 (
      {stage0_20[242], stage0_20[243], stage0_20[244], stage0_20[245], stage0_20[246], stage0_20[247]},
      {stage0_22[189], stage0_22[190], stage0_22[191], stage0_22[192], stage0_22[193], stage0_22[194]},
      {stage1_24[37],stage1_23[78],stage1_22[78],stage1_21[110],stage1_20[181]}
   );
   gpc606_5 gpc814 (
      {stage0_20[248], stage0_20[249], stage0_20[250], stage0_20[251], stage0_20[252], stage0_20[253]},
      {stage0_22[195], stage0_22[196], stage0_22[197], stage0_22[198], stage0_22[199], stage0_22[200]},
      {stage1_24[38],stage1_23[79],stage1_22[79],stage1_21[111],stage1_20[182]}
   );
   gpc606_5 gpc815 (
      {stage0_20[254], stage0_20[255], stage0_20[256], stage0_20[257], stage0_20[258], stage0_20[259]},
      {stage0_22[201], stage0_22[202], stage0_22[203], stage0_22[204], stage0_22[205], stage0_22[206]},
      {stage1_24[39],stage1_23[80],stage1_22[80],stage1_21[112],stage1_20[183]}
   );
   gpc606_5 gpc816 (
      {stage0_20[260], stage0_20[261], stage0_20[262], stage0_20[263], stage0_20[264], stage0_20[265]},
      {stage0_22[207], stage0_22[208], stage0_22[209], stage0_22[210], stage0_22[211], stage0_22[212]},
      {stage1_24[40],stage1_23[81],stage1_22[81],stage1_21[113],stage1_20[184]}
   );
   gpc606_5 gpc817 (
      {stage0_20[266], stage0_20[267], stage0_20[268], stage0_20[269], stage0_20[270], stage0_20[271]},
      {stage0_22[213], stage0_22[214], stage0_22[215], stage0_22[216], stage0_22[217], stage0_22[218]},
      {stage1_24[41],stage1_23[82],stage1_22[82],stage1_21[114],stage1_20[185]}
   );
   gpc606_5 gpc818 (
      {stage0_20[272], stage0_20[273], stage0_20[274], stage0_20[275], stage0_20[276], stage0_20[277]},
      {stage0_22[219], stage0_22[220], stage0_22[221], stage0_22[222], stage0_22[223], stage0_22[224]},
      {stage1_24[42],stage1_23[83],stage1_22[83],stage1_21[115],stage1_20[186]}
   );
   gpc606_5 gpc819 (
      {stage0_20[278], stage0_20[279], stage0_20[280], stage0_20[281], stage0_20[282], stage0_20[283]},
      {stage0_22[225], stage0_22[226], stage0_22[227], stage0_22[228], stage0_22[229], stage0_22[230]},
      {stage1_24[43],stage1_23[84],stage1_22[84],stage1_21[116],stage1_20[187]}
   );
   gpc606_5 gpc820 (
      {stage0_20[284], stage0_20[285], stage0_20[286], stage0_20[287], stage0_20[288], stage0_20[289]},
      {stage0_22[231], stage0_22[232], stage0_22[233], stage0_22[234], stage0_22[235], stage0_22[236]},
      {stage1_24[44],stage1_23[85],stage1_22[85],stage1_21[117],stage1_20[188]}
   );
   gpc606_5 gpc821 (
      {stage0_20[290], stage0_20[291], stage0_20[292], stage0_20[293], stage0_20[294], stage0_20[295]},
      {stage0_22[237], stage0_22[238], stage0_22[239], stage0_22[240], stage0_22[241], stage0_22[242]},
      {stage1_24[45],stage1_23[86],stage1_22[86],stage1_21[118],stage1_20[189]}
   );
   gpc606_5 gpc822 (
      {stage0_20[296], stage0_20[297], stage0_20[298], stage0_20[299], stage0_20[300], stage0_20[301]},
      {stage0_22[243], stage0_22[244], stage0_22[245], stage0_22[246], stage0_22[247], stage0_22[248]},
      {stage1_24[46],stage1_23[87],stage1_22[87],stage1_21[119],stage1_20[190]}
   );
   gpc606_5 gpc823 (
      {stage0_20[302], stage0_20[303], stage0_20[304], stage0_20[305], stage0_20[306], stage0_20[307]},
      {stage0_22[249], stage0_22[250], stage0_22[251], stage0_22[252], stage0_22[253], stage0_22[254]},
      {stage1_24[47],stage1_23[88],stage1_22[88],stage1_21[120],stage1_20[191]}
   );
   gpc606_5 gpc824 (
      {stage0_20[308], stage0_20[309], stage0_20[310], stage0_20[311], stage0_20[312], stage0_20[313]},
      {stage0_22[255], stage0_22[256], stage0_22[257], stage0_22[258], stage0_22[259], stage0_22[260]},
      {stage1_24[48],stage1_23[89],stage1_22[89],stage1_21[121],stage1_20[192]}
   );
   gpc606_5 gpc825 (
      {stage0_20[314], stage0_20[315], stage0_20[316], stage0_20[317], stage0_20[318], stage0_20[319]},
      {stage0_22[261], stage0_22[262], stage0_22[263], stage0_22[264], stage0_22[265], stage0_22[266]},
      {stage1_24[49],stage1_23[90],stage1_22[90],stage1_21[122],stage1_20[193]}
   );
   gpc606_5 gpc826 (
      {stage0_20[320], stage0_20[321], stage0_20[322], stage0_20[323], stage0_20[324], stage0_20[325]},
      {stage0_22[267], stage0_22[268], stage0_22[269], stage0_22[270], stage0_22[271], stage0_22[272]},
      {stage1_24[50],stage1_23[91],stage1_22[91],stage1_21[123],stage1_20[194]}
   );
   gpc606_5 gpc827 (
      {stage0_20[326], stage0_20[327], stage0_20[328], stage0_20[329], stage0_20[330], stage0_20[331]},
      {stage0_22[273], stage0_22[274], stage0_22[275], stage0_22[276], stage0_22[277], stage0_22[278]},
      {stage1_24[51],stage1_23[92],stage1_22[92],stage1_21[124],stage1_20[195]}
   );
   gpc606_5 gpc828 (
      {stage0_20[332], stage0_20[333], stage0_20[334], stage0_20[335], stage0_20[336], stage0_20[337]},
      {stage0_22[279], stage0_22[280], stage0_22[281], stage0_22[282], stage0_22[283], stage0_22[284]},
      {stage1_24[52],stage1_23[93],stage1_22[93],stage1_21[125],stage1_20[196]}
   );
   gpc606_5 gpc829 (
      {stage0_20[338], stage0_20[339], stage0_20[340], stage0_20[341], stage0_20[342], stage0_20[343]},
      {stage0_22[285], stage0_22[286], stage0_22[287], stage0_22[288], stage0_22[289], stage0_22[290]},
      {stage1_24[53],stage1_23[94],stage1_22[94],stage1_21[126],stage1_20[197]}
   );
   gpc606_5 gpc830 (
      {stage0_20[344], stage0_20[345], stage0_20[346], stage0_20[347], stage0_20[348], stage0_20[349]},
      {stage0_22[291], stage0_22[292], stage0_22[293], stage0_22[294], stage0_22[295], stage0_22[296]},
      {stage1_24[54],stage1_23[95],stage1_22[95],stage1_21[127],stage1_20[198]}
   );
   gpc606_5 gpc831 (
      {stage0_20[350], stage0_20[351], stage0_20[352], stage0_20[353], stage0_20[354], stage0_20[355]},
      {stage0_22[297], stage0_22[298], stage0_22[299], stage0_22[300], stage0_22[301], stage0_22[302]},
      {stage1_24[55],stage1_23[96],stage1_22[96],stage1_21[128],stage1_20[199]}
   );
   gpc606_5 gpc832 (
      {stage0_20[356], stage0_20[357], stage0_20[358], stage0_20[359], stage0_20[360], stage0_20[361]},
      {stage0_22[303], stage0_22[304], stage0_22[305], stage0_22[306], stage0_22[307], stage0_22[308]},
      {stage1_24[56],stage1_23[97],stage1_22[97],stage1_21[129],stage1_20[200]}
   );
   gpc606_5 gpc833 (
      {stage0_20[362], stage0_20[363], stage0_20[364], stage0_20[365], stage0_20[366], stage0_20[367]},
      {stage0_22[309], stage0_22[310], stage0_22[311], stage0_22[312], stage0_22[313], stage0_22[314]},
      {stage1_24[57],stage1_23[98],stage1_22[98],stage1_21[130],stage1_20[201]}
   );
   gpc606_5 gpc834 (
      {stage0_20[368], stage0_20[369], stage0_20[370], stage0_20[371], stage0_20[372], stage0_20[373]},
      {stage0_22[315], stage0_22[316], stage0_22[317], stage0_22[318], stage0_22[319], stage0_22[320]},
      {stage1_24[58],stage1_23[99],stage1_22[99],stage1_21[131],stage1_20[202]}
   );
   gpc606_5 gpc835 (
      {stage0_20[374], stage0_20[375], stage0_20[376], stage0_20[377], stage0_20[378], stage0_20[379]},
      {stage0_22[321], stage0_22[322], stage0_22[323], stage0_22[324], stage0_22[325], stage0_22[326]},
      {stage1_24[59],stage1_23[100],stage1_22[100],stage1_21[132],stage1_20[203]}
   );
   gpc606_5 gpc836 (
      {stage0_20[380], stage0_20[381], stage0_20[382], stage0_20[383], stage0_20[384], stage0_20[385]},
      {stage0_22[327], stage0_22[328], stage0_22[329], stage0_22[330], stage0_22[331], stage0_22[332]},
      {stage1_24[60],stage1_23[101],stage1_22[101],stage1_21[133],stage1_20[204]}
   );
   gpc606_5 gpc837 (
      {stage0_20[386], stage0_20[387], stage0_20[388], stage0_20[389], stage0_20[390], stage0_20[391]},
      {stage0_22[333], stage0_22[334], stage0_22[335], stage0_22[336], stage0_22[337], stage0_22[338]},
      {stage1_24[61],stage1_23[102],stage1_22[102],stage1_21[134],stage1_20[205]}
   );
   gpc615_5 gpc838 (
      {stage0_20[392], stage0_20[393], stage0_20[394], stage0_20[395], stage0_20[396]},
      {stage0_21[286]},
      {stage0_22[339], stage0_22[340], stage0_22[341], stage0_22[342], stage0_22[343], stage0_22[344]},
      {stage1_24[62],stage1_23[103],stage1_22[103],stage1_21[135],stage1_20[206]}
   );
   gpc615_5 gpc839 (
      {stage0_20[397], stage0_20[398], stage0_20[399], stage0_20[400], stage0_20[401]},
      {stage0_21[287]},
      {stage0_22[345], stage0_22[346], stage0_22[347], stage0_22[348], stage0_22[349], stage0_22[350]},
      {stage1_24[63],stage1_23[104],stage1_22[104],stage1_21[136],stage1_20[207]}
   );
   gpc615_5 gpc840 (
      {stage0_20[402], stage0_20[403], stage0_20[404], stage0_20[405], stage0_20[406]},
      {stage0_21[288]},
      {stage0_22[351], stage0_22[352], stage0_22[353], stage0_22[354], stage0_22[355], stage0_22[356]},
      {stage1_24[64],stage1_23[105],stage1_22[105],stage1_21[137],stage1_20[208]}
   );
   gpc615_5 gpc841 (
      {stage0_20[407], stage0_20[408], stage0_20[409], stage0_20[410], stage0_20[411]},
      {stage0_21[289]},
      {stage0_22[357], stage0_22[358], stage0_22[359], stage0_22[360], stage0_22[361], stage0_22[362]},
      {stage1_24[65],stage1_23[106],stage1_22[106],stage1_21[138],stage1_20[209]}
   );
   gpc615_5 gpc842 (
      {stage0_20[412], stage0_20[413], stage0_20[414], stage0_20[415], stage0_20[416]},
      {stage0_21[290]},
      {stage0_22[363], stage0_22[364], stage0_22[365], stage0_22[366], stage0_22[367], stage0_22[368]},
      {stage1_24[66],stage1_23[107],stage1_22[107],stage1_21[139],stage1_20[210]}
   );
   gpc615_5 gpc843 (
      {stage0_20[417], stage0_20[418], stage0_20[419], stage0_20[420], stage0_20[421]},
      {stage0_21[291]},
      {stage0_22[369], stage0_22[370], stage0_22[371], stage0_22[372], stage0_22[373], stage0_22[374]},
      {stage1_24[67],stage1_23[108],stage1_22[108],stage1_21[140],stage1_20[211]}
   );
   gpc615_5 gpc844 (
      {stage0_20[422], stage0_20[423], stage0_20[424], stage0_20[425], stage0_20[426]},
      {stage0_21[292]},
      {stage0_22[375], stage0_22[376], stage0_22[377], stage0_22[378], stage0_22[379], stage0_22[380]},
      {stage1_24[68],stage1_23[109],stage1_22[109],stage1_21[141],stage1_20[212]}
   );
   gpc615_5 gpc845 (
      {stage0_20[427], stage0_20[428], stage0_20[429], stage0_20[430], stage0_20[431]},
      {stage0_21[293]},
      {stage0_22[381], stage0_22[382], stage0_22[383], stage0_22[384], stage0_22[385], stage0_22[386]},
      {stage1_24[69],stage1_23[110],stage1_22[110],stage1_21[142],stage1_20[213]}
   );
   gpc606_5 gpc846 (
      {stage0_21[294], stage0_21[295], stage0_21[296], stage0_21[297], stage0_21[298], stage0_21[299]},
      {stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11], stage0_23[12]},
      {stage1_25[0],stage1_24[70],stage1_23[111],stage1_22[111],stage1_21[143]}
   );
   gpc606_5 gpc847 (
      {stage0_21[300], stage0_21[301], stage0_21[302], stage0_21[303], stage0_21[304], stage0_21[305]},
      {stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17], stage0_23[18]},
      {stage1_25[1],stage1_24[71],stage1_23[112],stage1_22[112],stage1_21[144]}
   );
   gpc606_5 gpc848 (
      {stage0_21[306], stage0_21[307], stage0_21[308], stage0_21[309], stage0_21[310], stage0_21[311]},
      {stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23], stage0_23[24]},
      {stage1_25[2],stage1_24[72],stage1_23[113],stage1_22[113],stage1_21[145]}
   );
   gpc606_5 gpc849 (
      {stage0_21[312], stage0_21[313], stage0_21[314], stage0_21[315], stage0_21[316], stage0_21[317]},
      {stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29], stage0_23[30]},
      {stage1_25[3],stage1_24[73],stage1_23[114],stage1_22[114],stage1_21[146]}
   );
   gpc606_5 gpc850 (
      {stage0_21[318], stage0_21[319], stage0_21[320], stage0_21[321], stage0_21[322], stage0_21[323]},
      {stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34], stage0_23[35], stage0_23[36]},
      {stage1_25[4],stage1_24[74],stage1_23[115],stage1_22[115],stage1_21[147]}
   );
   gpc606_5 gpc851 (
      {stage0_21[324], stage0_21[325], stage0_21[326], stage0_21[327], stage0_21[328], stage0_21[329]},
      {stage0_23[37], stage0_23[38], stage0_23[39], stage0_23[40], stage0_23[41], stage0_23[42]},
      {stage1_25[5],stage1_24[75],stage1_23[116],stage1_22[116],stage1_21[148]}
   );
   gpc606_5 gpc852 (
      {stage0_21[330], stage0_21[331], stage0_21[332], stage0_21[333], stage0_21[334], stage0_21[335]},
      {stage0_23[43], stage0_23[44], stage0_23[45], stage0_23[46], stage0_23[47], stage0_23[48]},
      {stage1_25[6],stage1_24[76],stage1_23[117],stage1_22[117],stage1_21[149]}
   );
   gpc606_5 gpc853 (
      {stage0_21[336], stage0_21[337], stage0_21[338], stage0_21[339], stage0_21[340], stage0_21[341]},
      {stage0_23[49], stage0_23[50], stage0_23[51], stage0_23[52], stage0_23[53], stage0_23[54]},
      {stage1_25[7],stage1_24[77],stage1_23[118],stage1_22[118],stage1_21[150]}
   );
   gpc606_5 gpc854 (
      {stage0_21[342], stage0_21[343], stage0_21[344], stage0_21[345], stage0_21[346], stage0_21[347]},
      {stage0_23[55], stage0_23[56], stage0_23[57], stage0_23[58], stage0_23[59], stage0_23[60]},
      {stage1_25[8],stage1_24[78],stage1_23[119],stage1_22[119],stage1_21[151]}
   );
   gpc606_5 gpc855 (
      {stage0_21[348], stage0_21[349], stage0_21[350], stage0_21[351], stage0_21[352], stage0_21[353]},
      {stage0_23[61], stage0_23[62], stage0_23[63], stage0_23[64], stage0_23[65], stage0_23[66]},
      {stage1_25[9],stage1_24[79],stage1_23[120],stage1_22[120],stage1_21[152]}
   );
   gpc606_5 gpc856 (
      {stage0_21[354], stage0_21[355], stage0_21[356], stage0_21[357], stage0_21[358], stage0_21[359]},
      {stage0_23[67], stage0_23[68], stage0_23[69], stage0_23[70], stage0_23[71], stage0_23[72]},
      {stage1_25[10],stage1_24[80],stage1_23[121],stage1_22[121],stage1_21[153]}
   );
   gpc606_5 gpc857 (
      {stage0_21[360], stage0_21[361], stage0_21[362], stage0_21[363], stage0_21[364], stage0_21[365]},
      {stage0_23[73], stage0_23[74], stage0_23[75], stage0_23[76], stage0_23[77], stage0_23[78]},
      {stage1_25[11],stage1_24[81],stage1_23[122],stage1_22[122],stage1_21[154]}
   );
   gpc606_5 gpc858 (
      {stage0_21[366], stage0_21[367], stage0_21[368], stage0_21[369], stage0_21[370], stage0_21[371]},
      {stage0_23[79], stage0_23[80], stage0_23[81], stage0_23[82], stage0_23[83], stage0_23[84]},
      {stage1_25[12],stage1_24[82],stage1_23[123],stage1_22[123],stage1_21[155]}
   );
   gpc606_5 gpc859 (
      {stage0_21[372], stage0_21[373], stage0_21[374], stage0_21[375], stage0_21[376], stage0_21[377]},
      {stage0_23[85], stage0_23[86], stage0_23[87], stage0_23[88], stage0_23[89], stage0_23[90]},
      {stage1_25[13],stage1_24[83],stage1_23[124],stage1_22[124],stage1_21[156]}
   );
   gpc606_5 gpc860 (
      {stage0_21[378], stage0_21[379], stage0_21[380], stage0_21[381], stage0_21[382], stage0_21[383]},
      {stage0_23[91], stage0_23[92], stage0_23[93], stage0_23[94], stage0_23[95], stage0_23[96]},
      {stage1_25[14],stage1_24[84],stage1_23[125],stage1_22[125],stage1_21[157]}
   );
   gpc606_5 gpc861 (
      {stage0_21[384], stage0_21[385], stage0_21[386], stage0_21[387], stage0_21[388], stage0_21[389]},
      {stage0_23[97], stage0_23[98], stage0_23[99], stage0_23[100], stage0_23[101], stage0_23[102]},
      {stage1_25[15],stage1_24[85],stage1_23[126],stage1_22[126],stage1_21[158]}
   );
   gpc606_5 gpc862 (
      {stage0_21[390], stage0_21[391], stage0_21[392], stage0_21[393], stage0_21[394], stage0_21[395]},
      {stage0_23[103], stage0_23[104], stage0_23[105], stage0_23[106], stage0_23[107], stage0_23[108]},
      {stage1_25[16],stage1_24[86],stage1_23[127],stage1_22[127],stage1_21[159]}
   );
   gpc606_5 gpc863 (
      {stage0_21[396], stage0_21[397], stage0_21[398], stage0_21[399], stage0_21[400], stage0_21[401]},
      {stage0_23[109], stage0_23[110], stage0_23[111], stage0_23[112], stage0_23[113], stage0_23[114]},
      {stage1_25[17],stage1_24[87],stage1_23[128],stage1_22[128],stage1_21[160]}
   );
   gpc606_5 gpc864 (
      {stage0_21[402], stage0_21[403], stage0_21[404], stage0_21[405], stage0_21[406], stage0_21[407]},
      {stage0_23[115], stage0_23[116], stage0_23[117], stage0_23[118], stage0_23[119], stage0_23[120]},
      {stage1_25[18],stage1_24[88],stage1_23[129],stage1_22[129],stage1_21[161]}
   );
   gpc606_5 gpc865 (
      {stage0_21[408], stage0_21[409], stage0_21[410], stage0_21[411], stage0_21[412], stage0_21[413]},
      {stage0_23[121], stage0_23[122], stage0_23[123], stage0_23[124], stage0_23[125], stage0_23[126]},
      {stage1_25[19],stage1_24[89],stage1_23[130],stage1_22[130],stage1_21[162]}
   );
   gpc606_5 gpc866 (
      {stage0_21[414], stage0_21[415], stage0_21[416], stage0_21[417], stage0_21[418], stage0_21[419]},
      {stage0_23[127], stage0_23[128], stage0_23[129], stage0_23[130], stage0_23[131], stage0_23[132]},
      {stage1_25[20],stage1_24[90],stage1_23[131],stage1_22[131],stage1_21[163]}
   );
   gpc606_5 gpc867 (
      {stage0_21[420], stage0_21[421], stage0_21[422], stage0_21[423], stage0_21[424], stage0_21[425]},
      {stage0_23[133], stage0_23[134], stage0_23[135], stage0_23[136], stage0_23[137], stage0_23[138]},
      {stage1_25[21],stage1_24[91],stage1_23[132],stage1_22[132],stage1_21[164]}
   );
   gpc606_5 gpc868 (
      {stage0_21[426], stage0_21[427], stage0_21[428], stage0_21[429], stage0_21[430], stage0_21[431]},
      {stage0_23[139], stage0_23[140], stage0_23[141], stage0_23[142], stage0_23[143], stage0_23[144]},
      {stage1_25[22],stage1_24[92],stage1_23[133],stage1_22[133],stage1_21[165]}
   );
   gpc606_5 gpc869 (
      {stage0_21[432], stage0_21[433], stage0_21[434], stage0_21[435], stage0_21[436], stage0_21[437]},
      {stage0_23[145], stage0_23[146], stage0_23[147], stage0_23[148], stage0_23[149], stage0_23[150]},
      {stage1_25[23],stage1_24[93],stage1_23[134],stage1_22[134],stage1_21[166]}
   );
   gpc606_5 gpc870 (
      {stage0_21[438], stage0_21[439], stage0_21[440], stage0_21[441], stage0_21[442], stage0_21[443]},
      {stage0_23[151], stage0_23[152], stage0_23[153], stage0_23[154], stage0_23[155], stage0_23[156]},
      {stage1_25[24],stage1_24[94],stage1_23[135],stage1_22[135],stage1_21[167]}
   );
   gpc606_5 gpc871 (
      {stage0_21[444], stage0_21[445], stage0_21[446], stage0_21[447], stage0_21[448], stage0_21[449]},
      {stage0_23[157], stage0_23[158], stage0_23[159], stage0_23[160], stage0_23[161], stage0_23[162]},
      {stage1_25[25],stage1_24[95],stage1_23[136],stage1_22[136],stage1_21[168]}
   );
   gpc606_5 gpc872 (
      {stage0_21[450], stage0_21[451], stage0_21[452], stage0_21[453], stage0_21[454], stage0_21[455]},
      {stage0_23[163], stage0_23[164], stage0_23[165], stage0_23[166], stage0_23[167], stage0_23[168]},
      {stage1_25[26],stage1_24[96],stage1_23[137],stage1_22[137],stage1_21[169]}
   );
   gpc606_5 gpc873 (
      {stage0_21[456], stage0_21[457], stage0_21[458], stage0_21[459], stage0_21[460], stage0_21[461]},
      {stage0_23[169], stage0_23[170], stage0_23[171], stage0_23[172], stage0_23[173], stage0_23[174]},
      {stage1_25[27],stage1_24[97],stage1_23[138],stage1_22[138],stage1_21[170]}
   );
   gpc606_5 gpc874 (
      {stage0_21[462], stage0_21[463], stage0_21[464], stage0_21[465], stage0_21[466], stage0_21[467]},
      {stage0_23[175], stage0_23[176], stage0_23[177], stage0_23[178], stage0_23[179], stage0_23[180]},
      {stage1_25[28],stage1_24[98],stage1_23[139],stage1_22[139],stage1_21[171]}
   );
   gpc615_5 gpc875 (
      {stage0_22[387], stage0_22[388], stage0_22[389], stage0_22[390], stage0_22[391]},
      {stage0_23[181]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[29],stage1_24[99],stage1_23[140],stage1_22[140]}
   );
   gpc615_5 gpc876 (
      {stage0_22[392], stage0_22[393], stage0_22[394], stage0_22[395], stage0_22[396]},
      {stage0_23[182]},
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage1_26[1],stage1_25[30],stage1_24[100],stage1_23[141],stage1_22[141]}
   );
   gpc615_5 gpc877 (
      {stage0_22[397], stage0_22[398], stage0_22[399], stage0_22[400], stage0_22[401]},
      {stage0_23[183]},
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage1_26[2],stage1_25[31],stage1_24[101],stage1_23[142],stage1_22[142]}
   );
   gpc615_5 gpc878 (
      {stage0_22[402], stage0_22[403], stage0_22[404], stage0_22[405], stage0_22[406]},
      {stage0_23[184]},
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage1_26[3],stage1_25[32],stage1_24[102],stage1_23[143],stage1_22[143]}
   );
   gpc615_5 gpc879 (
      {stage0_22[407], stage0_22[408], stage0_22[409], stage0_22[410], stage0_22[411]},
      {stage0_23[185]},
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage1_26[4],stage1_25[33],stage1_24[103],stage1_23[144],stage1_22[144]}
   );
   gpc615_5 gpc880 (
      {stage0_22[412], stage0_22[413], stage0_22[414], stage0_22[415], stage0_22[416]},
      {stage0_23[186]},
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage1_26[5],stage1_25[34],stage1_24[104],stage1_23[145],stage1_22[145]}
   );
   gpc615_5 gpc881 (
      {stage0_22[417], stage0_22[418], stage0_22[419], stage0_22[420], stage0_22[421]},
      {stage0_23[187]},
      {stage0_24[36], stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41]},
      {stage1_26[6],stage1_25[35],stage1_24[105],stage1_23[146],stage1_22[146]}
   );
   gpc615_5 gpc882 (
      {stage0_22[422], stage0_22[423], stage0_22[424], stage0_22[425], stage0_22[426]},
      {stage0_23[188]},
      {stage0_24[42], stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47]},
      {stage1_26[7],stage1_25[36],stage1_24[106],stage1_23[147],stage1_22[147]}
   );
   gpc615_5 gpc883 (
      {stage0_22[427], stage0_22[428], stage0_22[429], stage0_22[430], stage0_22[431]},
      {stage0_23[189]},
      {stage0_24[48], stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53]},
      {stage1_26[8],stage1_25[37],stage1_24[107],stage1_23[148],stage1_22[148]}
   );
   gpc615_5 gpc884 (
      {stage0_22[432], stage0_22[433], stage0_22[434], stage0_22[435], stage0_22[436]},
      {stage0_23[190]},
      {stage0_24[54], stage0_24[55], stage0_24[56], stage0_24[57], stage0_24[58], stage0_24[59]},
      {stage1_26[9],stage1_25[38],stage1_24[108],stage1_23[149],stage1_22[149]}
   );
   gpc615_5 gpc885 (
      {stage0_22[437], stage0_22[438], stage0_22[439], stage0_22[440], stage0_22[441]},
      {stage0_23[191]},
      {stage0_24[60], stage0_24[61], stage0_24[62], stage0_24[63], stage0_24[64], stage0_24[65]},
      {stage1_26[10],stage1_25[39],stage1_24[109],stage1_23[150],stage1_22[150]}
   );
   gpc615_5 gpc886 (
      {stage0_22[442], stage0_22[443], stage0_22[444], stage0_22[445], stage0_22[446]},
      {stage0_23[192]},
      {stage0_24[66], stage0_24[67], stage0_24[68], stage0_24[69], stage0_24[70], stage0_24[71]},
      {stage1_26[11],stage1_25[40],stage1_24[110],stage1_23[151],stage1_22[151]}
   );
   gpc615_5 gpc887 (
      {stage0_22[447], stage0_22[448], stage0_22[449], stage0_22[450], stage0_22[451]},
      {stage0_23[193]},
      {stage0_24[72], stage0_24[73], stage0_24[74], stage0_24[75], stage0_24[76], stage0_24[77]},
      {stage1_26[12],stage1_25[41],stage1_24[111],stage1_23[152],stage1_22[152]}
   );
   gpc615_5 gpc888 (
      {stage0_22[452], stage0_22[453], stage0_22[454], stage0_22[455], stage0_22[456]},
      {stage0_23[194]},
      {stage0_24[78], stage0_24[79], stage0_24[80], stage0_24[81], stage0_24[82], stage0_24[83]},
      {stage1_26[13],stage1_25[42],stage1_24[112],stage1_23[153],stage1_22[153]}
   );
   gpc615_5 gpc889 (
      {stage0_22[457], stage0_22[458], stage0_22[459], stage0_22[460], stage0_22[461]},
      {stage0_23[195]},
      {stage0_24[84], stage0_24[85], stage0_24[86], stage0_24[87], stage0_24[88], stage0_24[89]},
      {stage1_26[14],stage1_25[43],stage1_24[113],stage1_23[154],stage1_22[154]}
   );
   gpc615_5 gpc890 (
      {stage0_22[462], stage0_22[463], stage0_22[464], stage0_22[465], stage0_22[466]},
      {stage0_23[196]},
      {stage0_24[90], stage0_24[91], stage0_24[92], stage0_24[93], stage0_24[94], stage0_24[95]},
      {stage1_26[15],stage1_25[44],stage1_24[114],stage1_23[155],stage1_22[155]}
   );
   gpc615_5 gpc891 (
      {stage0_22[467], stage0_22[468], stage0_22[469], stage0_22[470], stage0_22[471]},
      {stage0_23[197]},
      {stage0_24[96], stage0_24[97], stage0_24[98], stage0_24[99], stage0_24[100], stage0_24[101]},
      {stage1_26[16],stage1_25[45],stage1_24[115],stage1_23[156],stage1_22[156]}
   );
   gpc615_5 gpc892 (
      {stage0_23[198], stage0_23[199], stage0_23[200], stage0_23[201], stage0_23[202]},
      {stage0_24[102]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[17],stage1_25[46],stage1_24[116],stage1_23[157]}
   );
   gpc615_5 gpc893 (
      {stage0_23[203], stage0_23[204], stage0_23[205], stage0_23[206], stage0_23[207]},
      {stage0_24[103]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[18],stage1_25[47],stage1_24[117],stage1_23[158]}
   );
   gpc615_5 gpc894 (
      {stage0_23[208], stage0_23[209], stage0_23[210], stage0_23[211], stage0_23[212]},
      {stage0_24[104]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[19],stage1_25[48],stage1_24[118],stage1_23[159]}
   );
   gpc615_5 gpc895 (
      {stage0_23[213], stage0_23[214], stage0_23[215], stage0_23[216], stage0_23[217]},
      {stage0_24[105]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[20],stage1_25[49],stage1_24[119],stage1_23[160]}
   );
   gpc615_5 gpc896 (
      {stage0_23[218], stage0_23[219], stage0_23[220], stage0_23[221], stage0_23[222]},
      {stage0_24[106]},
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage1_27[4],stage1_26[21],stage1_25[50],stage1_24[120],stage1_23[161]}
   );
   gpc615_5 gpc897 (
      {stage0_23[223], stage0_23[224], stage0_23[225], stage0_23[226], stage0_23[227]},
      {stage0_24[107]},
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage1_27[5],stage1_26[22],stage1_25[51],stage1_24[121],stage1_23[162]}
   );
   gpc615_5 gpc898 (
      {stage0_23[228], stage0_23[229], stage0_23[230], stage0_23[231], stage0_23[232]},
      {stage0_24[108]},
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage1_27[6],stage1_26[23],stage1_25[52],stage1_24[122],stage1_23[163]}
   );
   gpc615_5 gpc899 (
      {stage0_23[233], stage0_23[234], stage0_23[235], stage0_23[236], stage0_23[237]},
      {stage0_24[109]},
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46], stage0_25[47]},
      {stage1_27[7],stage1_26[24],stage1_25[53],stage1_24[123],stage1_23[164]}
   );
   gpc615_5 gpc900 (
      {stage0_23[238], stage0_23[239], stage0_23[240], stage0_23[241], stage0_23[242]},
      {stage0_24[110]},
      {stage0_25[48], stage0_25[49], stage0_25[50], stage0_25[51], stage0_25[52], stage0_25[53]},
      {stage1_27[8],stage1_26[25],stage1_25[54],stage1_24[124],stage1_23[165]}
   );
   gpc615_5 gpc901 (
      {stage0_23[243], stage0_23[244], stage0_23[245], stage0_23[246], stage0_23[247]},
      {stage0_24[111]},
      {stage0_25[54], stage0_25[55], stage0_25[56], stage0_25[57], stage0_25[58], stage0_25[59]},
      {stage1_27[9],stage1_26[26],stage1_25[55],stage1_24[125],stage1_23[166]}
   );
   gpc615_5 gpc902 (
      {stage0_23[248], stage0_23[249], stage0_23[250], stage0_23[251], stage0_23[252]},
      {stage0_24[112]},
      {stage0_25[60], stage0_25[61], stage0_25[62], stage0_25[63], stage0_25[64], stage0_25[65]},
      {stage1_27[10],stage1_26[27],stage1_25[56],stage1_24[126],stage1_23[167]}
   );
   gpc615_5 gpc903 (
      {stage0_23[253], stage0_23[254], stage0_23[255], stage0_23[256], stage0_23[257]},
      {stage0_24[113]},
      {stage0_25[66], stage0_25[67], stage0_25[68], stage0_25[69], stage0_25[70], stage0_25[71]},
      {stage1_27[11],stage1_26[28],stage1_25[57],stage1_24[127],stage1_23[168]}
   );
   gpc615_5 gpc904 (
      {stage0_23[258], stage0_23[259], stage0_23[260], stage0_23[261], stage0_23[262]},
      {stage0_24[114]},
      {stage0_25[72], stage0_25[73], stage0_25[74], stage0_25[75], stage0_25[76], stage0_25[77]},
      {stage1_27[12],stage1_26[29],stage1_25[58],stage1_24[128],stage1_23[169]}
   );
   gpc615_5 gpc905 (
      {stage0_23[263], stage0_23[264], stage0_23[265], stage0_23[266], stage0_23[267]},
      {stage0_24[115]},
      {stage0_25[78], stage0_25[79], stage0_25[80], stage0_25[81], stage0_25[82], stage0_25[83]},
      {stage1_27[13],stage1_26[30],stage1_25[59],stage1_24[129],stage1_23[170]}
   );
   gpc615_5 gpc906 (
      {stage0_23[268], stage0_23[269], stage0_23[270], stage0_23[271], stage0_23[272]},
      {stage0_24[116]},
      {stage0_25[84], stage0_25[85], stage0_25[86], stage0_25[87], stage0_25[88], stage0_25[89]},
      {stage1_27[14],stage1_26[31],stage1_25[60],stage1_24[130],stage1_23[171]}
   );
   gpc615_5 gpc907 (
      {stage0_23[273], stage0_23[274], stage0_23[275], stage0_23[276], stage0_23[277]},
      {stage0_24[117]},
      {stage0_25[90], stage0_25[91], stage0_25[92], stage0_25[93], stage0_25[94], stage0_25[95]},
      {stage1_27[15],stage1_26[32],stage1_25[61],stage1_24[131],stage1_23[172]}
   );
   gpc615_5 gpc908 (
      {stage0_23[278], stage0_23[279], stage0_23[280], stage0_23[281], stage0_23[282]},
      {stage0_24[118]},
      {stage0_25[96], stage0_25[97], stage0_25[98], stage0_25[99], stage0_25[100], stage0_25[101]},
      {stage1_27[16],stage1_26[33],stage1_25[62],stage1_24[132],stage1_23[173]}
   );
   gpc615_5 gpc909 (
      {stage0_23[283], stage0_23[284], stage0_23[285], stage0_23[286], stage0_23[287]},
      {stage0_24[119]},
      {stage0_25[102], stage0_25[103], stage0_25[104], stage0_25[105], stage0_25[106], stage0_25[107]},
      {stage1_27[17],stage1_26[34],stage1_25[63],stage1_24[133],stage1_23[174]}
   );
   gpc615_5 gpc910 (
      {stage0_23[288], stage0_23[289], stage0_23[290], stage0_23[291], stage0_23[292]},
      {stage0_24[120]},
      {stage0_25[108], stage0_25[109], stage0_25[110], stage0_25[111], stage0_25[112], stage0_25[113]},
      {stage1_27[18],stage1_26[35],stage1_25[64],stage1_24[134],stage1_23[175]}
   );
   gpc615_5 gpc911 (
      {stage0_23[293], stage0_23[294], stage0_23[295], stage0_23[296], stage0_23[297]},
      {stage0_24[121]},
      {stage0_25[114], stage0_25[115], stage0_25[116], stage0_25[117], stage0_25[118], stage0_25[119]},
      {stage1_27[19],stage1_26[36],stage1_25[65],stage1_24[135],stage1_23[176]}
   );
   gpc615_5 gpc912 (
      {stage0_23[298], stage0_23[299], stage0_23[300], stage0_23[301], stage0_23[302]},
      {stage0_24[122]},
      {stage0_25[120], stage0_25[121], stage0_25[122], stage0_25[123], stage0_25[124], stage0_25[125]},
      {stage1_27[20],stage1_26[37],stage1_25[66],stage1_24[136],stage1_23[177]}
   );
   gpc615_5 gpc913 (
      {stage0_23[303], stage0_23[304], stage0_23[305], stage0_23[306], stage0_23[307]},
      {stage0_24[123]},
      {stage0_25[126], stage0_25[127], stage0_25[128], stage0_25[129], stage0_25[130], stage0_25[131]},
      {stage1_27[21],stage1_26[38],stage1_25[67],stage1_24[137],stage1_23[178]}
   );
   gpc615_5 gpc914 (
      {stage0_23[308], stage0_23[309], stage0_23[310], stage0_23[311], stage0_23[312]},
      {stage0_24[124]},
      {stage0_25[132], stage0_25[133], stage0_25[134], stage0_25[135], stage0_25[136], stage0_25[137]},
      {stage1_27[22],stage1_26[39],stage1_25[68],stage1_24[138],stage1_23[179]}
   );
   gpc615_5 gpc915 (
      {stage0_23[313], stage0_23[314], stage0_23[315], stage0_23[316], stage0_23[317]},
      {stage0_24[125]},
      {stage0_25[138], stage0_25[139], stage0_25[140], stage0_25[141], stage0_25[142], stage0_25[143]},
      {stage1_27[23],stage1_26[40],stage1_25[69],stage1_24[139],stage1_23[180]}
   );
   gpc615_5 gpc916 (
      {stage0_23[318], stage0_23[319], stage0_23[320], stage0_23[321], stage0_23[322]},
      {stage0_24[126]},
      {stage0_25[144], stage0_25[145], stage0_25[146], stage0_25[147], stage0_25[148], stage0_25[149]},
      {stage1_27[24],stage1_26[41],stage1_25[70],stage1_24[140],stage1_23[181]}
   );
   gpc615_5 gpc917 (
      {stage0_23[323], stage0_23[324], stage0_23[325], stage0_23[326], stage0_23[327]},
      {stage0_24[127]},
      {stage0_25[150], stage0_25[151], stage0_25[152], stage0_25[153], stage0_25[154], stage0_25[155]},
      {stage1_27[25],stage1_26[42],stage1_25[71],stage1_24[141],stage1_23[182]}
   );
   gpc615_5 gpc918 (
      {stage0_23[328], stage0_23[329], stage0_23[330], stage0_23[331], stage0_23[332]},
      {stage0_24[128]},
      {stage0_25[156], stage0_25[157], stage0_25[158], stage0_25[159], stage0_25[160], stage0_25[161]},
      {stage1_27[26],stage1_26[43],stage1_25[72],stage1_24[142],stage1_23[183]}
   );
   gpc615_5 gpc919 (
      {stage0_23[333], stage0_23[334], stage0_23[335], stage0_23[336], stage0_23[337]},
      {stage0_24[129]},
      {stage0_25[162], stage0_25[163], stage0_25[164], stage0_25[165], stage0_25[166], stage0_25[167]},
      {stage1_27[27],stage1_26[44],stage1_25[73],stage1_24[143],stage1_23[184]}
   );
   gpc615_5 gpc920 (
      {stage0_23[338], stage0_23[339], stage0_23[340], stage0_23[341], stage0_23[342]},
      {stage0_24[130]},
      {stage0_25[168], stage0_25[169], stage0_25[170], stage0_25[171], stage0_25[172], stage0_25[173]},
      {stage1_27[28],stage1_26[45],stage1_25[74],stage1_24[144],stage1_23[185]}
   );
   gpc615_5 gpc921 (
      {stage0_23[343], stage0_23[344], stage0_23[345], stage0_23[346], stage0_23[347]},
      {stage0_24[131]},
      {stage0_25[174], stage0_25[175], stage0_25[176], stage0_25[177], stage0_25[178], stage0_25[179]},
      {stage1_27[29],stage1_26[46],stage1_25[75],stage1_24[145],stage1_23[186]}
   );
   gpc615_5 gpc922 (
      {stage0_23[348], stage0_23[349], stage0_23[350], stage0_23[351], stage0_23[352]},
      {stage0_24[132]},
      {stage0_25[180], stage0_25[181], stage0_25[182], stage0_25[183], stage0_25[184], stage0_25[185]},
      {stage1_27[30],stage1_26[47],stage1_25[76],stage1_24[146],stage1_23[187]}
   );
   gpc615_5 gpc923 (
      {stage0_23[353], stage0_23[354], stage0_23[355], stage0_23[356], stage0_23[357]},
      {stage0_24[133]},
      {stage0_25[186], stage0_25[187], stage0_25[188], stage0_25[189], stage0_25[190], stage0_25[191]},
      {stage1_27[31],stage1_26[48],stage1_25[77],stage1_24[147],stage1_23[188]}
   );
   gpc615_5 gpc924 (
      {stage0_23[358], stage0_23[359], stage0_23[360], stage0_23[361], stage0_23[362]},
      {stage0_24[134]},
      {stage0_25[192], stage0_25[193], stage0_25[194], stage0_25[195], stage0_25[196], stage0_25[197]},
      {stage1_27[32],stage1_26[49],stage1_25[78],stage1_24[148],stage1_23[189]}
   );
   gpc615_5 gpc925 (
      {stage0_23[363], stage0_23[364], stage0_23[365], stage0_23[366], stage0_23[367]},
      {stage0_24[135]},
      {stage0_25[198], stage0_25[199], stage0_25[200], stage0_25[201], stage0_25[202], stage0_25[203]},
      {stage1_27[33],stage1_26[50],stage1_25[79],stage1_24[149],stage1_23[190]}
   );
   gpc615_5 gpc926 (
      {stage0_23[368], stage0_23[369], stage0_23[370], stage0_23[371], stage0_23[372]},
      {stage0_24[136]},
      {stage0_25[204], stage0_25[205], stage0_25[206], stage0_25[207], stage0_25[208], stage0_25[209]},
      {stage1_27[34],stage1_26[51],stage1_25[80],stage1_24[150],stage1_23[191]}
   );
   gpc615_5 gpc927 (
      {stage0_23[373], stage0_23[374], stage0_23[375], stage0_23[376], stage0_23[377]},
      {stage0_24[137]},
      {stage0_25[210], stage0_25[211], stage0_25[212], stage0_25[213], stage0_25[214], stage0_25[215]},
      {stage1_27[35],stage1_26[52],stage1_25[81],stage1_24[151],stage1_23[192]}
   );
   gpc615_5 gpc928 (
      {stage0_23[378], stage0_23[379], stage0_23[380], stage0_23[381], stage0_23[382]},
      {stage0_24[138]},
      {stage0_25[216], stage0_25[217], stage0_25[218], stage0_25[219], stage0_25[220], stage0_25[221]},
      {stage1_27[36],stage1_26[53],stage1_25[82],stage1_24[152],stage1_23[193]}
   );
   gpc615_5 gpc929 (
      {stage0_23[383], stage0_23[384], stage0_23[385], stage0_23[386], stage0_23[387]},
      {stage0_24[139]},
      {stage0_25[222], stage0_25[223], stage0_25[224], stage0_25[225], stage0_25[226], stage0_25[227]},
      {stage1_27[37],stage1_26[54],stage1_25[83],stage1_24[153],stage1_23[194]}
   );
   gpc615_5 gpc930 (
      {stage0_23[388], stage0_23[389], stage0_23[390], stage0_23[391], stage0_23[392]},
      {stage0_24[140]},
      {stage0_25[228], stage0_25[229], stage0_25[230], stage0_25[231], stage0_25[232], stage0_25[233]},
      {stage1_27[38],stage1_26[55],stage1_25[84],stage1_24[154],stage1_23[195]}
   );
   gpc623_5 gpc931 (
      {stage0_23[393], stage0_23[394], stage0_23[395]},
      {stage0_24[141], stage0_24[142]},
      {stage0_25[234], stage0_25[235], stage0_25[236], stage0_25[237], stage0_25[238], stage0_25[239]},
      {stage1_27[39],stage1_26[56],stage1_25[85],stage1_24[155],stage1_23[196]}
   );
   gpc606_5 gpc932 (
      {stage0_24[143], stage0_24[144], stage0_24[145], stage0_24[146], stage0_24[147], stage0_24[148]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[40],stage1_26[57],stage1_25[86],stage1_24[156]}
   );
   gpc606_5 gpc933 (
      {stage0_24[149], stage0_24[150], stage0_24[151], stage0_24[152], stage0_24[153], stage0_24[154]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[41],stage1_26[58],stage1_25[87],stage1_24[157]}
   );
   gpc606_5 gpc934 (
      {stage0_24[155], stage0_24[156], stage0_24[157], stage0_24[158], stage0_24[159], stage0_24[160]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[42],stage1_26[59],stage1_25[88],stage1_24[158]}
   );
   gpc606_5 gpc935 (
      {stage0_24[161], stage0_24[162], stage0_24[163], stage0_24[164], stage0_24[165], stage0_24[166]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[43],stage1_26[60],stage1_25[89],stage1_24[159]}
   );
   gpc606_5 gpc936 (
      {stage0_24[167], stage0_24[168], stage0_24[169], stage0_24[170], stage0_24[171], stage0_24[172]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[44],stage1_26[61],stage1_25[90],stage1_24[160]}
   );
   gpc606_5 gpc937 (
      {stage0_24[173], stage0_24[174], stage0_24[175], stage0_24[176], stage0_24[177], stage0_24[178]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[45],stage1_26[62],stage1_25[91],stage1_24[161]}
   );
   gpc606_5 gpc938 (
      {stage0_24[179], stage0_24[180], stage0_24[181], stage0_24[182], stage0_24[183], stage0_24[184]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[46],stage1_26[63],stage1_25[92],stage1_24[162]}
   );
   gpc606_5 gpc939 (
      {stage0_24[185], stage0_24[186], stage0_24[187], stage0_24[188], stage0_24[189], stage0_24[190]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[47],stage1_26[64],stage1_25[93],stage1_24[163]}
   );
   gpc606_5 gpc940 (
      {stage0_24[191], stage0_24[192], stage0_24[193], stage0_24[194], stage0_24[195], stage0_24[196]},
      {stage0_26[48], stage0_26[49], stage0_26[50], stage0_26[51], stage0_26[52], stage0_26[53]},
      {stage1_28[8],stage1_27[48],stage1_26[65],stage1_25[94],stage1_24[164]}
   );
   gpc606_5 gpc941 (
      {stage0_24[197], stage0_24[198], stage0_24[199], stage0_24[200], stage0_24[201], stage0_24[202]},
      {stage0_26[54], stage0_26[55], stage0_26[56], stage0_26[57], stage0_26[58], stage0_26[59]},
      {stage1_28[9],stage1_27[49],stage1_26[66],stage1_25[95],stage1_24[165]}
   );
   gpc606_5 gpc942 (
      {stage0_24[203], stage0_24[204], stage0_24[205], stage0_24[206], stage0_24[207], stage0_24[208]},
      {stage0_26[60], stage0_26[61], stage0_26[62], stage0_26[63], stage0_26[64], stage0_26[65]},
      {stage1_28[10],stage1_27[50],stage1_26[67],stage1_25[96],stage1_24[166]}
   );
   gpc606_5 gpc943 (
      {stage0_24[209], stage0_24[210], stage0_24[211], stage0_24[212], stage0_24[213], stage0_24[214]},
      {stage0_26[66], stage0_26[67], stage0_26[68], stage0_26[69], stage0_26[70], stage0_26[71]},
      {stage1_28[11],stage1_27[51],stage1_26[68],stage1_25[97],stage1_24[167]}
   );
   gpc606_5 gpc944 (
      {stage0_24[215], stage0_24[216], stage0_24[217], stage0_24[218], stage0_24[219], stage0_24[220]},
      {stage0_26[72], stage0_26[73], stage0_26[74], stage0_26[75], stage0_26[76], stage0_26[77]},
      {stage1_28[12],stage1_27[52],stage1_26[69],stage1_25[98],stage1_24[168]}
   );
   gpc606_5 gpc945 (
      {stage0_24[221], stage0_24[222], stage0_24[223], stage0_24[224], stage0_24[225], stage0_24[226]},
      {stage0_26[78], stage0_26[79], stage0_26[80], stage0_26[81], stage0_26[82], stage0_26[83]},
      {stage1_28[13],stage1_27[53],stage1_26[70],stage1_25[99],stage1_24[169]}
   );
   gpc606_5 gpc946 (
      {stage0_24[227], stage0_24[228], stage0_24[229], stage0_24[230], stage0_24[231], stage0_24[232]},
      {stage0_26[84], stage0_26[85], stage0_26[86], stage0_26[87], stage0_26[88], stage0_26[89]},
      {stage1_28[14],stage1_27[54],stage1_26[71],stage1_25[100],stage1_24[170]}
   );
   gpc606_5 gpc947 (
      {stage0_24[233], stage0_24[234], stage0_24[235], stage0_24[236], stage0_24[237], stage0_24[238]},
      {stage0_26[90], stage0_26[91], stage0_26[92], stage0_26[93], stage0_26[94], stage0_26[95]},
      {stage1_28[15],stage1_27[55],stage1_26[72],stage1_25[101],stage1_24[171]}
   );
   gpc606_5 gpc948 (
      {stage0_24[239], stage0_24[240], stage0_24[241], stage0_24[242], stage0_24[243], stage0_24[244]},
      {stage0_26[96], stage0_26[97], stage0_26[98], stage0_26[99], stage0_26[100], stage0_26[101]},
      {stage1_28[16],stage1_27[56],stage1_26[73],stage1_25[102],stage1_24[172]}
   );
   gpc606_5 gpc949 (
      {stage0_24[245], stage0_24[246], stage0_24[247], stage0_24[248], stage0_24[249], stage0_24[250]},
      {stage0_26[102], stage0_26[103], stage0_26[104], stage0_26[105], stage0_26[106], stage0_26[107]},
      {stage1_28[17],stage1_27[57],stage1_26[74],stage1_25[103],stage1_24[173]}
   );
   gpc606_5 gpc950 (
      {stage0_24[251], stage0_24[252], stage0_24[253], stage0_24[254], stage0_24[255], stage0_24[256]},
      {stage0_26[108], stage0_26[109], stage0_26[110], stage0_26[111], stage0_26[112], stage0_26[113]},
      {stage1_28[18],stage1_27[58],stage1_26[75],stage1_25[104],stage1_24[174]}
   );
   gpc606_5 gpc951 (
      {stage0_24[257], stage0_24[258], stage0_24[259], stage0_24[260], stage0_24[261], stage0_24[262]},
      {stage0_26[114], stage0_26[115], stage0_26[116], stage0_26[117], stage0_26[118], stage0_26[119]},
      {stage1_28[19],stage1_27[59],stage1_26[76],stage1_25[105],stage1_24[175]}
   );
   gpc606_5 gpc952 (
      {stage0_24[263], stage0_24[264], stage0_24[265], stage0_24[266], stage0_24[267], stage0_24[268]},
      {stage0_26[120], stage0_26[121], stage0_26[122], stage0_26[123], stage0_26[124], stage0_26[125]},
      {stage1_28[20],stage1_27[60],stage1_26[77],stage1_25[106],stage1_24[176]}
   );
   gpc606_5 gpc953 (
      {stage0_24[269], stage0_24[270], stage0_24[271], stage0_24[272], stage0_24[273], stage0_24[274]},
      {stage0_26[126], stage0_26[127], stage0_26[128], stage0_26[129], stage0_26[130], stage0_26[131]},
      {stage1_28[21],stage1_27[61],stage1_26[78],stage1_25[107],stage1_24[177]}
   );
   gpc606_5 gpc954 (
      {stage0_24[275], stage0_24[276], stage0_24[277], stage0_24[278], stage0_24[279], stage0_24[280]},
      {stage0_26[132], stage0_26[133], stage0_26[134], stage0_26[135], stage0_26[136], stage0_26[137]},
      {stage1_28[22],stage1_27[62],stage1_26[79],stage1_25[108],stage1_24[178]}
   );
   gpc606_5 gpc955 (
      {stage0_24[281], stage0_24[282], stage0_24[283], stage0_24[284], stage0_24[285], stage0_24[286]},
      {stage0_26[138], stage0_26[139], stage0_26[140], stage0_26[141], stage0_26[142], stage0_26[143]},
      {stage1_28[23],stage1_27[63],stage1_26[80],stage1_25[109],stage1_24[179]}
   );
   gpc606_5 gpc956 (
      {stage0_24[287], stage0_24[288], stage0_24[289], stage0_24[290], stage0_24[291], stage0_24[292]},
      {stage0_26[144], stage0_26[145], stage0_26[146], stage0_26[147], stage0_26[148], stage0_26[149]},
      {stage1_28[24],stage1_27[64],stage1_26[81],stage1_25[110],stage1_24[180]}
   );
   gpc606_5 gpc957 (
      {stage0_24[293], stage0_24[294], stage0_24[295], stage0_24[296], stage0_24[297], stage0_24[298]},
      {stage0_26[150], stage0_26[151], stage0_26[152], stage0_26[153], stage0_26[154], stage0_26[155]},
      {stage1_28[25],stage1_27[65],stage1_26[82],stage1_25[111],stage1_24[181]}
   );
   gpc606_5 gpc958 (
      {stage0_24[299], stage0_24[300], stage0_24[301], stage0_24[302], stage0_24[303], stage0_24[304]},
      {stage0_26[156], stage0_26[157], stage0_26[158], stage0_26[159], stage0_26[160], stage0_26[161]},
      {stage1_28[26],stage1_27[66],stage1_26[83],stage1_25[112],stage1_24[182]}
   );
   gpc606_5 gpc959 (
      {stage0_24[305], stage0_24[306], stage0_24[307], stage0_24[308], stage0_24[309], stage0_24[310]},
      {stage0_26[162], stage0_26[163], stage0_26[164], stage0_26[165], stage0_26[166], stage0_26[167]},
      {stage1_28[27],stage1_27[67],stage1_26[84],stage1_25[113],stage1_24[183]}
   );
   gpc606_5 gpc960 (
      {stage0_24[311], stage0_24[312], stage0_24[313], stage0_24[314], stage0_24[315], stage0_24[316]},
      {stage0_26[168], stage0_26[169], stage0_26[170], stage0_26[171], stage0_26[172], stage0_26[173]},
      {stage1_28[28],stage1_27[68],stage1_26[85],stage1_25[114],stage1_24[184]}
   );
   gpc606_5 gpc961 (
      {stage0_24[317], stage0_24[318], stage0_24[319], stage0_24[320], stage0_24[321], stage0_24[322]},
      {stage0_26[174], stage0_26[175], stage0_26[176], stage0_26[177], stage0_26[178], stage0_26[179]},
      {stage1_28[29],stage1_27[69],stage1_26[86],stage1_25[115],stage1_24[185]}
   );
   gpc606_5 gpc962 (
      {stage0_24[323], stage0_24[324], stage0_24[325], stage0_24[326], stage0_24[327], stage0_24[328]},
      {stage0_26[180], stage0_26[181], stage0_26[182], stage0_26[183], stage0_26[184], stage0_26[185]},
      {stage1_28[30],stage1_27[70],stage1_26[87],stage1_25[116],stage1_24[186]}
   );
   gpc606_5 gpc963 (
      {stage0_24[329], stage0_24[330], stage0_24[331], stage0_24[332], stage0_24[333], stage0_24[334]},
      {stage0_26[186], stage0_26[187], stage0_26[188], stage0_26[189], stage0_26[190], stage0_26[191]},
      {stage1_28[31],stage1_27[71],stage1_26[88],stage1_25[117],stage1_24[187]}
   );
   gpc606_5 gpc964 (
      {stage0_24[335], stage0_24[336], stage0_24[337], stage0_24[338], stage0_24[339], stage0_24[340]},
      {stage0_26[192], stage0_26[193], stage0_26[194], stage0_26[195], stage0_26[196], stage0_26[197]},
      {stage1_28[32],stage1_27[72],stage1_26[89],stage1_25[118],stage1_24[188]}
   );
   gpc606_5 gpc965 (
      {stage0_24[341], stage0_24[342], stage0_24[343], stage0_24[344], stage0_24[345], stage0_24[346]},
      {stage0_26[198], stage0_26[199], stage0_26[200], stage0_26[201], stage0_26[202], stage0_26[203]},
      {stage1_28[33],stage1_27[73],stage1_26[90],stage1_25[119],stage1_24[189]}
   );
   gpc606_5 gpc966 (
      {stage0_24[347], stage0_24[348], stage0_24[349], stage0_24[350], stage0_24[351], stage0_24[352]},
      {stage0_26[204], stage0_26[205], stage0_26[206], stage0_26[207], stage0_26[208], stage0_26[209]},
      {stage1_28[34],stage1_27[74],stage1_26[91],stage1_25[120],stage1_24[190]}
   );
   gpc606_5 gpc967 (
      {stage0_24[353], stage0_24[354], stage0_24[355], stage0_24[356], stage0_24[357], stage0_24[358]},
      {stage0_26[210], stage0_26[211], stage0_26[212], stage0_26[213], stage0_26[214], stage0_26[215]},
      {stage1_28[35],stage1_27[75],stage1_26[92],stage1_25[121],stage1_24[191]}
   );
   gpc606_5 gpc968 (
      {stage0_24[359], stage0_24[360], stage0_24[361], stage0_24[362], stage0_24[363], stage0_24[364]},
      {stage0_26[216], stage0_26[217], stage0_26[218], stage0_26[219], stage0_26[220], stage0_26[221]},
      {stage1_28[36],stage1_27[76],stage1_26[93],stage1_25[122],stage1_24[192]}
   );
   gpc606_5 gpc969 (
      {stage0_24[365], stage0_24[366], stage0_24[367], stage0_24[368], stage0_24[369], stage0_24[370]},
      {stage0_26[222], stage0_26[223], stage0_26[224], stage0_26[225], stage0_26[226], stage0_26[227]},
      {stage1_28[37],stage1_27[77],stage1_26[94],stage1_25[123],stage1_24[193]}
   );
   gpc606_5 gpc970 (
      {stage0_24[371], stage0_24[372], stage0_24[373], stage0_24[374], stage0_24[375], stage0_24[376]},
      {stage0_26[228], stage0_26[229], stage0_26[230], stage0_26[231], stage0_26[232], stage0_26[233]},
      {stage1_28[38],stage1_27[78],stage1_26[95],stage1_25[124],stage1_24[194]}
   );
   gpc606_5 gpc971 (
      {stage0_24[377], stage0_24[378], stage0_24[379], stage0_24[380], stage0_24[381], stage0_24[382]},
      {stage0_26[234], stage0_26[235], stage0_26[236], stage0_26[237], stage0_26[238], stage0_26[239]},
      {stage1_28[39],stage1_27[79],stage1_26[96],stage1_25[125],stage1_24[195]}
   );
   gpc606_5 gpc972 (
      {stage0_24[383], stage0_24[384], stage0_24[385], stage0_24[386], stage0_24[387], stage0_24[388]},
      {stage0_26[240], stage0_26[241], stage0_26[242], stage0_26[243], stage0_26[244], stage0_26[245]},
      {stage1_28[40],stage1_27[80],stage1_26[97],stage1_25[126],stage1_24[196]}
   );
   gpc606_5 gpc973 (
      {stage0_24[389], stage0_24[390], stage0_24[391], stage0_24[392], stage0_24[393], stage0_24[394]},
      {stage0_26[246], stage0_26[247], stage0_26[248], stage0_26[249], stage0_26[250], stage0_26[251]},
      {stage1_28[41],stage1_27[81],stage1_26[98],stage1_25[127],stage1_24[197]}
   );
   gpc606_5 gpc974 (
      {stage0_24[395], stage0_24[396], stage0_24[397], stage0_24[398], stage0_24[399], stage0_24[400]},
      {stage0_26[252], stage0_26[253], stage0_26[254], stage0_26[255], stage0_26[256], stage0_26[257]},
      {stage1_28[42],stage1_27[82],stage1_26[99],stage1_25[128],stage1_24[198]}
   );
   gpc606_5 gpc975 (
      {stage0_24[401], stage0_24[402], stage0_24[403], stage0_24[404], stage0_24[405], stage0_24[406]},
      {stage0_26[258], stage0_26[259], stage0_26[260], stage0_26[261], stage0_26[262], stage0_26[263]},
      {stage1_28[43],stage1_27[83],stage1_26[100],stage1_25[129],stage1_24[199]}
   );
   gpc606_5 gpc976 (
      {stage0_24[407], stage0_24[408], stage0_24[409], stage0_24[410], stage0_24[411], stage0_24[412]},
      {stage0_26[264], stage0_26[265], stage0_26[266], stage0_26[267], stage0_26[268], stage0_26[269]},
      {stage1_28[44],stage1_27[84],stage1_26[101],stage1_25[130],stage1_24[200]}
   );
   gpc606_5 gpc977 (
      {stage0_24[413], stage0_24[414], stage0_24[415], stage0_24[416], stage0_24[417], stage0_24[418]},
      {stage0_26[270], stage0_26[271], stage0_26[272], stage0_26[273], stage0_26[274], stage0_26[275]},
      {stage1_28[45],stage1_27[85],stage1_26[102],stage1_25[131],stage1_24[201]}
   );
   gpc606_5 gpc978 (
      {stage0_24[419], stage0_24[420], stage0_24[421], stage0_24[422], stage0_24[423], stage0_24[424]},
      {stage0_26[276], stage0_26[277], stage0_26[278], stage0_26[279], stage0_26[280], stage0_26[281]},
      {stage1_28[46],stage1_27[86],stage1_26[103],stage1_25[132],stage1_24[202]}
   );
   gpc606_5 gpc979 (
      {stage0_24[425], stage0_24[426], stage0_24[427], stage0_24[428], stage0_24[429], stage0_24[430]},
      {stage0_26[282], stage0_26[283], stage0_26[284], stage0_26[285], stage0_26[286], stage0_26[287]},
      {stage1_28[47],stage1_27[87],stage1_26[104],stage1_25[133],stage1_24[203]}
   );
   gpc606_5 gpc980 (
      {stage0_24[431], stage0_24[432], stage0_24[433], stage0_24[434], stage0_24[435], stage0_24[436]},
      {stage0_26[288], stage0_26[289], stage0_26[290], stage0_26[291], stage0_26[292], stage0_26[293]},
      {stage1_28[48],stage1_27[88],stage1_26[105],stage1_25[134],stage1_24[204]}
   );
   gpc606_5 gpc981 (
      {stage0_24[437], stage0_24[438], stage0_24[439], stage0_24[440], stage0_24[441], stage0_24[442]},
      {stage0_26[294], stage0_26[295], stage0_26[296], stage0_26[297], stage0_26[298], stage0_26[299]},
      {stage1_28[49],stage1_27[89],stage1_26[106],stage1_25[135],stage1_24[205]}
   );
   gpc606_5 gpc982 (
      {stage0_24[443], stage0_24[444], stage0_24[445], stage0_24[446], stage0_24[447], stage0_24[448]},
      {stage0_26[300], stage0_26[301], stage0_26[302], stage0_26[303], stage0_26[304], stage0_26[305]},
      {stage1_28[50],stage1_27[90],stage1_26[107],stage1_25[136],stage1_24[206]}
   );
   gpc606_5 gpc983 (
      {stage0_24[449], stage0_24[450], stage0_24[451], stage0_24[452], stage0_24[453], stage0_24[454]},
      {stage0_26[306], stage0_26[307], stage0_26[308], stage0_26[309], stage0_26[310], stage0_26[311]},
      {stage1_28[51],stage1_27[91],stage1_26[108],stage1_25[137],stage1_24[207]}
   );
   gpc606_5 gpc984 (
      {stage0_24[455], stage0_24[456], stage0_24[457], stage0_24[458], stage0_24[459], stage0_24[460]},
      {stage0_26[312], stage0_26[313], stage0_26[314], stage0_26[315], stage0_26[316], stage0_26[317]},
      {stage1_28[52],stage1_27[92],stage1_26[109],stage1_25[138],stage1_24[208]}
   );
   gpc606_5 gpc985 (
      {stage0_24[461], stage0_24[462], stage0_24[463], stage0_24[464], stage0_24[465], stage0_24[466]},
      {stage0_26[318], stage0_26[319], stage0_26[320], stage0_26[321], stage0_26[322], stage0_26[323]},
      {stage1_28[53],stage1_27[93],stage1_26[110],stage1_25[139],stage1_24[209]}
   );
   gpc606_5 gpc986 (
      {stage0_24[467], stage0_24[468], stage0_24[469], stage0_24[470], stage0_24[471], stage0_24[472]},
      {stage0_26[324], stage0_26[325], stage0_26[326], stage0_26[327], stage0_26[328], stage0_26[329]},
      {stage1_28[54],stage1_27[94],stage1_26[111],stage1_25[140],stage1_24[210]}
   );
   gpc606_5 gpc987 (
      {stage0_24[473], stage0_24[474], stage0_24[475], stage0_24[476], stage0_24[477], stage0_24[478]},
      {stage0_26[330], stage0_26[331], stage0_26[332], stage0_26[333], stage0_26[334], stage0_26[335]},
      {stage1_28[55],stage1_27[95],stage1_26[112],stage1_25[141],stage1_24[211]}
   );
   gpc606_5 gpc988 (
      {stage0_24[479], stage0_24[480], stage0_24[481], stage0_24[482], stage0_24[483], stage0_24[484]},
      {stage0_26[336], stage0_26[337], stage0_26[338], stage0_26[339], stage0_26[340], stage0_26[341]},
      {stage1_28[56],stage1_27[96],stage1_26[113],stage1_25[142],stage1_24[212]}
   );
   gpc606_5 gpc989 (
      {stage0_25[240], stage0_25[241], stage0_25[242], stage0_25[243], stage0_25[244], stage0_25[245]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[57],stage1_27[97],stage1_26[114],stage1_25[143]}
   );
   gpc606_5 gpc990 (
      {stage0_25[246], stage0_25[247], stage0_25[248], stage0_25[249], stage0_25[250], stage0_25[251]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[58],stage1_27[98],stage1_26[115],stage1_25[144]}
   );
   gpc606_5 gpc991 (
      {stage0_25[252], stage0_25[253], stage0_25[254], stage0_25[255], stage0_25[256], stage0_25[257]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[59],stage1_27[99],stage1_26[116],stage1_25[145]}
   );
   gpc606_5 gpc992 (
      {stage0_25[258], stage0_25[259], stage0_25[260], stage0_25[261], stage0_25[262], stage0_25[263]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[60],stage1_27[100],stage1_26[117],stage1_25[146]}
   );
   gpc606_5 gpc993 (
      {stage0_25[264], stage0_25[265], stage0_25[266], stage0_25[267], stage0_25[268], stage0_25[269]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[61],stage1_27[101],stage1_26[118],stage1_25[147]}
   );
   gpc606_5 gpc994 (
      {stage0_25[270], stage0_25[271], stage0_25[272], stage0_25[273], stage0_25[274], stage0_25[275]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[62],stage1_27[102],stage1_26[119],stage1_25[148]}
   );
   gpc606_5 gpc995 (
      {stage0_25[276], stage0_25[277], stage0_25[278], stage0_25[279], stage0_25[280], stage0_25[281]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[63],stage1_27[103],stage1_26[120],stage1_25[149]}
   );
   gpc606_5 gpc996 (
      {stage0_25[282], stage0_25[283], stage0_25[284], stage0_25[285], stage0_25[286], stage0_25[287]},
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage1_29[7],stage1_28[64],stage1_27[104],stage1_26[121],stage1_25[150]}
   );
   gpc606_5 gpc997 (
      {stage0_25[288], stage0_25[289], stage0_25[290], stage0_25[291], stage0_25[292], stage0_25[293]},
      {stage0_27[48], stage0_27[49], stage0_27[50], stage0_27[51], stage0_27[52], stage0_27[53]},
      {stage1_29[8],stage1_28[65],stage1_27[105],stage1_26[122],stage1_25[151]}
   );
   gpc606_5 gpc998 (
      {stage0_25[294], stage0_25[295], stage0_25[296], stage0_25[297], stage0_25[298], stage0_25[299]},
      {stage0_27[54], stage0_27[55], stage0_27[56], stage0_27[57], stage0_27[58], stage0_27[59]},
      {stage1_29[9],stage1_28[66],stage1_27[106],stage1_26[123],stage1_25[152]}
   );
   gpc606_5 gpc999 (
      {stage0_25[300], stage0_25[301], stage0_25[302], stage0_25[303], stage0_25[304], stage0_25[305]},
      {stage0_27[60], stage0_27[61], stage0_27[62], stage0_27[63], stage0_27[64], stage0_27[65]},
      {stage1_29[10],stage1_28[67],stage1_27[107],stage1_26[124],stage1_25[153]}
   );
   gpc606_5 gpc1000 (
      {stage0_25[306], stage0_25[307], stage0_25[308], stage0_25[309], stage0_25[310], stage0_25[311]},
      {stage0_27[66], stage0_27[67], stage0_27[68], stage0_27[69], stage0_27[70], stage0_27[71]},
      {stage1_29[11],stage1_28[68],stage1_27[108],stage1_26[125],stage1_25[154]}
   );
   gpc606_5 gpc1001 (
      {stage0_25[312], stage0_25[313], stage0_25[314], stage0_25[315], stage0_25[316], stage0_25[317]},
      {stage0_27[72], stage0_27[73], stage0_27[74], stage0_27[75], stage0_27[76], stage0_27[77]},
      {stage1_29[12],stage1_28[69],stage1_27[109],stage1_26[126],stage1_25[155]}
   );
   gpc606_5 gpc1002 (
      {stage0_25[318], stage0_25[319], stage0_25[320], stage0_25[321], stage0_25[322], stage0_25[323]},
      {stage0_27[78], stage0_27[79], stage0_27[80], stage0_27[81], stage0_27[82], stage0_27[83]},
      {stage1_29[13],stage1_28[70],stage1_27[110],stage1_26[127],stage1_25[156]}
   );
   gpc606_5 gpc1003 (
      {stage0_25[324], stage0_25[325], stage0_25[326], stage0_25[327], stage0_25[328], stage0_25[329]},
      {stage0_27[84], stage0_27[85], stage0_27[86], stage0_27[87], stage0_27[88], stage0_27[89]},
      {stage1_29[14],stage1_28[71],stage1_27[111],stage1_26[128],stage1_25[157]}
   );
   gpc606_5 gpc1004 (
      {stage0_25[330], stage0_25[331], stage0_25[332], stage0_25[333], stage0_25[334], stage0_25[335]},
      {stage0_27[90], stage0_27[91], stage0_27[92], stage0_27[93], stage0_27[94], stage0_27[95]},
      {stage1_29[15],stage1_28[72],stage1_27[112],stage1_26[129],stage1_25[158]}
   );
   gpc606_5 gpc1005 (
      {stage0_25[336], stage0_25[337], stage0_25[338], stage0_25[339], stage0_25[340], stage0_25[341]},
      {stage0_27[96], stage0_27[97], stage0_27[98], stage0_27[99], stage0_27[100], stage0_27[101]},
      {stage1_29[16],stage1_28[73],stage1_27[113],stage1_26[130],stage1_25[159]}
   );
   gpc606_5 gpc1006 (
      {stage0_25[342], stage0_25[343], stage0_25[344], stage0_25[345], stage0_25[346], stage0_25[347]},
      {stage0_27[102], stage0_27[103], stage0_27[104], stage0_27[105], stage0_27[106], stage0_27[107]},
      {stage1_29[17],stage1_28[74],stage1_27[114],stage1_26[131],stage1_25[160]}
   );
   gpc606_5 gpc1007 (
      {stage0_25[348], stage0_25[349], stage0_25[350], stage0_25[351], stage0_25[352], stage0_25[353]},
      {stage0_27[108], stage0_27[109], stage0_27[110], stage0_27[111], stage0_27[112], stage0_27[113]},
      {stage1_29[18],stage1_28[75],stage1_27[115],stage1_26[132],stage1_25[161]}
   );
   gpc606_5 gpc1008 (
      {stage0_25[354], stage0_25[355], stage0_25[356], stage0_25[357], stage0_25[358], stage0_25[359]},
      {stage0_27[114], stage0_27[115], stage0_27[116], stage0_27[117], stage0_27[118], stage0_27[119]},
      {stage1_29[19],stage1_28[76],stage1_27[116],stage1_26[133],stage1_25[162]}
   );
   gpc606_5 gpc1009 (
      {stage0_25[360], stage0_25[361], stage0_25[362], stage0_25[363], stage0_25[364], stage0_25[365]},
      {stage0_27[120], stage0_27[121], stage0_27[122], stage0_27[123], stage0_27[124], stage0_27[125]},
      {stage1_29[20],stage1_28[77],stage1_27[117],stage1_26[134],stage1_25[163]}
   );
   gpc606_5 gpc1010 (
      {stage0_25[366], stage0_25[367], stage0_25[368], stage0_25[369], stage0_25[370], stage0_25[371]},
      {stage0_27[126], stage0_27[127], stage0_27[128], stage0_27[129], stage0_27[130], stage0_27[131]},
      {stage1_29[21],stage1_28[78],stage1_27[118],stage1_26[135],stage1_25[164]}
   );
   gpc606_5 gpc1011 (
      {stage0_25[372], stage0_25[373], stage0_25[374], stage0_25[375], stage0_25[376], stage0_25[377]},
      {stage0_27[132], stage0_27[133], stage0_27[134], stage0_27[135], stage0_27[136], stage0_27[137]},
      {stage1_29[22],stage1_28[79],stage1_27[119],stage1_26[136],stage1_25[165]}
   );
   gpc606_5 gpc1012 (
      {stage0_25[378], stage0_25[379], stage0_25[380], stage0_25[381], stage0_25[382], stage0_25[383]},
      {stage0_27[138], stage0_27[139], stage0_27[140], stage0_27[141], stage0_27[142], stage0_27[143]},
      {stage1_29[23],stage1_28[80],stage1_27[120],stage1_26[137],stage1_25[166]}
   );
   gpc606_5 gpc1013 (
      {stage0_25[384], stage0_25[385], stage0_25[386], stage0_25[387], stage0_25[388], stage0_25[389]},
      {stage0_27[144], stage0_27[145], stage0_27[146], stage0_27[147], stage0_27[148], stage0_27[149]},
      {stage1_29[24],stage1_28[81],stage1_27[121],stage1_26[138],stage1_25[167]}
   );
   gpc606_5 gpc1014 (
      {stage0_25[390], stage0_25[391], stage0_25[392], stage0_25[393], stage0_25[394], stage0_25[395]},
      {stage0_27[150], stage0_27[151], stage0_27[152], stage0_27[153], stage0_27[154], stage0_27[155]},
      {stage1_29[25],stage1_28[82],stage1_27[122],stage1_26[139],stage1_25[168]}
   );
   gpc606_5 gpc1015 (
      {stage0_25[396], stage0_25[397], stage0_25[398], stage0_25[399], stage0_25[400], stage0_25[401]},
      {stage0_27[156], stage0_27[157], stage0_27[158], stage0_27[159], stage0_27[160], stage0_27[161]},
      {stage1_29[26],stage1_28[83],stage1_27[123],stage1_26[140],stage1_25[169]}
   );
   gpc606_5 gpc1016 (
      {stage0_25[402], stage0_25[403], stage0_25[404], stage0_25[405], stage0_25[406], stage0_25[407]},
      {stage0_27[162], stage0_27[163], stage0_27[164], stage0_27[165], stage0_27[166], stage0_27[167]},
      {stage1_29[27],stage1_28[84],stage1_27[124],stage1_26[141],stage1_25[170]}
   );
   gpc606_5 gpc1017 (
      {stage0_25[408], stage0_25[409], stage0_25[410], stage0_25[411], stage0_25[412], stage0_25[413]},
      {stage0_27[168], stage0_27[169], stage0_27[170], stage0_27[171], stage0_27[172], stage0_27[173]},
      {stage1_29[28],stage1_28[85],stage1_27[125],stage1_26[142],stage1_25[171]}
   );
   gpc606_5 gpc1018 (
      {stage0_25[414], stage0_25[415], stage0_25[416], stage0_25[417], stage0_25[418], stage0_25[419]},
      {stage0_27[174], stage0_27[175], stage0_27[176], stage0_27[177], stage0_27[178], stage0_27[179]},
      {stage1_29[29],stage1_28[86],stage1_27[126],stage1_26[143],stage1_25[172]}
   );
   gpc606_5 gpc1019 (
      {stage0_25[420], stage0_25[421], stage0_25[422], stage0_25[423], stage0_25[424], stage0_25[425]},
      {stage0_27[180], stage0_27[181], stage0_27[182], stage0_27[183], stage0_27[184], stage0_27[185]},
      {stage1_29[30],stage1_28[87],stage1_27[127],stage1_26[144],stage1_25[173]}
   );
   gpc606_5 gpc1020 (
      {stage0_25[426], stage0_25[427], stage0_25[428], stage0_25[429], stage0_25[430], stage0_25[431]},
      {stage0_27[186], stage0_27[187], stage0_27[188], stage0_27[189], stage0_27[190], stage0_27[191]},
      {stage1_29[31],stage1_28[88],stage1_27[128],stage1_26[145],stage1_25[174]}
   );
   gpc606_5 gpc1021 (
      {stage0_25[432], stage0_25[433], stage0_25[434], stage0_25[435], stage0_25[436], stage0_25[437]},
      {stage0_27[192], stage0_27[193], stage0_27[194], stage0_27[195], stage0_27[196], stage0_27[197]},
      {stage1_29[32],stage1_28[89],stage1_27[129],stage1_26[146],stage1_25[175]}
   );
   gpc606_5 gpc1022 (
      {stage0_25[438], stage0_25[439], stage0_25[440], stage0_25[441], stage0_25[442], stage0_25[443]},
      {stage0_27[198], stage0_27[199], stage0_27[200], stage0_27[201], stage0_27[202], stage0_27[203]},
      {stage1_29[33],stage1_28[90],stage1_27[130],stage1_26[147],stage1_25[176]}
   );
   gpc606_5 gpc1023 (
      {stage0_25[444], stage0_25[445], stage0_25[446], stage0_25[447], stage0_25[448], stage0_25[449]},
      {stage0_27[204], stage0_27[205], stage0_27[206], stage0_27[207], stage0_27[208], stage0_27[209]},
      {stage1_29[34],stage1_28[91],stage1_27[131],stage1_26[148],stage1_25[177]}
   );
   gpc606_5 gpc1024 (
      {stage0_25[450], stage0_25[451], stage0_25[452], stage0_25[453], stage0_25[454], stage0_25[455]},
      {stage0_27[210], stage0_27[211], stage0_27[212], stage0_27[213], stage0_27[214], stage0_27[215]},
      {stage1_29[35],stage1_28[92],stage1_27[132],stage1_26[149],stage1_25[178]}
   );
   gpc606_5 gpc1025 (
      {stage0_25[456], stage0_25[457], stage0_25[458], stage0_25[459], stage0_25[460], stage0_25[461]},
      {stage0_27[216], stage0_27[217], stage0_27[218], stage0_27[219], stage0_27[220], stage0_27[221]},
      {stage1_29[36],stage1_28[93],stage1_27[133],stage1_26[150],stage1_25[179]}
   );
   gpc606_5 gpc1026 (
      {stage0_25[462], stage0_25[463], stage0_25[464], stage0_25[465], stage0_25[466], stage0_25[467]},
      {stage0_27[222], stage0_27[223], stage0_27[224], stage0_27[225], stage0_27[226], stage0_27[227]},
      {stage1_29[37],stage1_28[94],stage1_27[134],stage1_26[151],stage1_25[180]}
   );
   gpc606_5 gpc1027 (
      {stage0_25[468], stage0_25[469], stage0_25[470], stage0_25[471], stage0_25[472], stage0_25[473]},
      {stage0_27[228], stage0_27[229], stage0_27[230], stage0_27[231], stage0_27[232], stage0_27[233]},
      {stage1_29[38],stage1_28[95],stage1_27[135],stage1_26[152],stage1_25[181]}
   );
   gpc606_5 gpc1028 (
      {stage0_25[474], stage0_25[475], stage0_25[476], stage0_25[477], stage0_25[478], stage0_25[479]},
      {stage0_27[234], stage0_27[235], stage0_27[236], stage0_27[237], stage0_27[238], stage0_27[239]},
      {stage1_29[39],stage1_28[96],stage1_27[136],stage1_26[153],stage1_25[182]}
   );
   gpc606_5 gpc1029 (
      {stage0_25[480], stage0_25[481], stage0_25[482], stage0_25[483], stage0_25[484], stage0_25[485]},
      {stage0_27[240], stage0_27[241], stage0_27[242], stage0_27[243], stage0_27[244], stage0_27[245]},
      {stage1_29[40],stage1_28[97],stage1_27[137],stage1_26[154],stage1_25[183]}
   );
   gpc615_5 gpc1030 (
      {stage0_26[342], stage0_26[343], stage0_26[344], stage0_26[345], stage0_26[346]},
      {stage0_27[246]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[41],stage1_28[98],stage1_27[138],stage1_26[155]}
   );
   gpc615_5 gpc1031 (
      {stage0_26[347], stage0_26[348], stage0_26[349], stage0_26[350], stage0_26[351]},
      {stage0_27[247]},
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage1_30[1],stage1_29[42],stage1_28[99],stage1_27[139],stage1_26[156]}
   );
   gpc615_5 gpc1032 (
      {stage0_26[352], stage0_26[353], stage0_26[354], stage0_26[355], stage0_26[356]},
      {stage0_27[248]},
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage1_30[2],stage1_29[43],stage1_28[100],stage1_27[140],stage1_26[157]}
   );
   gpc615_5 gpc1033 (
      {stage0_26[357], stage0_26[358], stage0_26[359], stage0_26[360], stage0_26[361]},
      {stage0_27[249]},
      {stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23]},
      {stage1_30[3],stage1_29[44],stage1_28[101],stage1_27[141],stage1_26[158]}
   );
   gpc615_5 gpc1034 (
      {stage0_26[362], stage0_26[363], stage0_26[364], stage0_26[365], stage0_26[366]},
      {stage0_27[250]},
      {stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29]},
      {stage1_30[4],stage1_29[45],stage1_28[102],stage1_27[142],stage1_26[159]}
   );
   gpc615_5 gpc1035 (
      {stage0_26[367], stage0_26[368], stage0_26[369], stage0_26[370], stage0_26[371]},
      {stage0_27[251]},
      {stage0_28[30], stage0_28[31], stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35]},
      {stage1_30[5],stage1_29[46],stage1_28[103],stage1_27[143],stage1_26[160]}
   );
   gpc615_5 gpc1036 (
      {stage0_26[372], stage0_26[373], stage0_26[374], stage0_26[375], stage0_26[376]},
      {stage0_27[252]},
      {stage0_28[36], stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41]},
      {stage1_30[6],stage1_29[47],stage1_28[104],stage1_27[144],stage1_26[161]}
   );
   gpc615_5 gpc1037 (
      {stage0_26[377], stage0_26[378], stage0_26[379], stage0_26[380], stage0_26[381]},
      {stage0_27[253]},
      {stage0_28[42], stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47]},
      {stage1_30[7],stage1_29[48],stage1_28[105],stage1_27[145],stage1_26[162]}
   );
   gpc615_5 gpc1038 (
      {stage0_26[382], stage0_26[383], stage0_26[384], stage0_26[385], stage0_26[386]},
      {stage0_27[254]},
      {stage0_28[48], stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53]},
      {stage1_30[8],stage1_29[49],stage1_28[106],stage1_27[146],stage1_26[163]}
   );
   gpc615_5 gpc1039 (
      {stage0_26[387], stage0_26[388], stage0_26[389], stage0_26[390], stage0_26[391]},
      {stage0_27[255]},
      {stage0_28[54], stage0_28[55], stage0_28[56], stage0_28[57], stage0_28[58], stage0_28[59]},
      {stage1_30[9],stage1_29[50],stage1_28[107],stage1_27[147],stage1_26[164]}
   );
   gpc615_5 gpc1040 (
      {stage0_26[392], stage0_26[393], stage0_26[394], stage0_26[395], stage0_26[396]},
      {stage0_27[256]},
      {stage0_28[60], stage0_28[61], stage0_28[62], stage0_28[63], stage0_28[64], stage0_28[65]},
      {stage1_30[10],stage1_29[51],stage1_28[108],stage1_27[148],stage1_26[165]}
   );
   gpc615_5 gpc1041 (
      {stage0_26[397], stage0_26[398], stage0_26[399], stage0_26[400], stage0_26[401]},
      {stage0_27[257]},
      {stage0_28[66], stage0_28[67], stage0_28[68], stage0_28[69], stage0_28[70], stage0_28[71]},
      {stage1_30[11],stage1_29[52],stage1_28[109],stage1_27[149],stage1_26[166]}
   );
   gpc615_5 gpc1042 (
      {stage0_27[258], stage0_27[259], stage0_27[260], stage0_27[261], stage0_27[262]},
      {stage0_28[72]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[12],stage1_29[53],stage1_28[110],stage1_27[150]}
   );
   gpc615_5 gpc1043 (
      {stage0_27[263], stage0_27[264], stage0_27[265], stage0_27[266], stage0_27[267]},
      {stage0_28[73]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[13],stage1_29[54],stage1_28[111],stage1_27[151]}
   );
   gpc615_5 gpc1044 (
      {stage0_27[268], stage0_27[269], stage0_27[270], stage0_27[271], stage0_27[272]},
      {stage0_28[74]},
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage1_31[2],stage1_30[14],stage1_29[55],stage1_28[112],stage1_27[152]}
   );
   gpc615_5 gpc1045 (
      {stage0_27[273], stage0_27[274], stage0_27[275], stage0_27[276], stage0_27[277]},
      {stage0_28[75]},
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage1_31[3],stage1_30[15],stage1_29[56],stage1_28[113],stage1_27[153]}
   );
   gpc615_5 gpc1046 (
      {stage0_27[278], stage0_27[279], stage0_27[280], stage0_27[281], stage0_27[282]},
      {stage0_28[76]},
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage1_31[4],stage1_30[16],stage1_29[57],stage1_28[114],stage1_27[154]}
   );
   gpc615_5 gpc1047 (
      {stage0_27[283], stage0_27[284], stage0_27[285], stage0_27[286], stage0_27[287]},
      {stage0_28[77]},
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage1_31[5],stage1_30[17],stage1_29[58],stage1_28[115],stage1_27[155]}
   );
   gpc615_5 gpc1048 (
      {stage0_27[288], stage0_27[289], stage0_27[290], stage0_27[291], stage0_27[292]},
      {stage0_28[78]},
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage1_31[6],stage1_30[18],stage1_29[59],stage1_28[116],stage1_27[156]}
   );
   gpc615_5 gpc1049 (
      {stage0_27[293], stage0_27[294], stage0_27[295], stage0_27[296], stage0_27[297]},
      {stage0_28[79]},
      {stage0_29[42], stage0_29[43], stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47]},
      {stage1_31[7],stage1_30[19],stage1_29[60],stage1_28[117],stage1_27[157]}
   );
   gpc615_5 gpc1050 (
      {stage0_27[298], stage0_27[299], stage0_27[300], stage0_27[301], stage0_27[302]},
      {stage0_28[80]},
      {stage0_29[48], stage0_29[49], stage0_29[50], stage0_29[51], stage0_29[52], stage0_29[53]},
      {stage1_31[8],stage1_30[20],stage1_29[61],stage1_28[118],stage1_27[158]}
   );
   gpc615_5 gpc1051 (
      {stage0_27[303], stage0_27[304], stage0_27[305], stage0_27[306], stage0_27[307]},
      {stage0_28[81]},
      {stage0_29[54], stage0_29[55], stage0_29[56], stage0_29[57], stage0_29[58], stage0_29[59]},
      {stage1_31[9],stage1_30[21],stage1_29[62],stage1_28[119],stage1_27[159]}
   );
   gpc615_5 gpc1052 (
      {stage0_27[308], stage0_27[309], stage0_27[310], stage0_27[311], stage0_27[312]},
      {stage0_28[82]},
      {stage0_29[60], stage0_29[61], stage0_29[62], stage0_29[63], stage0_29[64], stage0_29[65]},
      {stage1_31[10],stage1_30[22],stage1_29[63],stage1_28[120],stage1_27[160]}
   );
   gpc615_5 gpc1053 (
      {stage0_27[313], stage0_27[314], stage0_27[315], stage0_27[316], stage0_27[317]},
      {stage0_28[83]},
      {stage0_29[66], stage0_29[67], stage0_29[68], stage0_29[69], stage0_29[70], stage0_29[71]},
      {stage1_31[11],stage1_30[23],stage1_29[64],stage1_28[121],stage1_27[161]}
   );
   gpc615_5 gpc1054 (
      {stage0_27[318], stage0_27[319], stage0_27[320], stage0_27[321], stage0_27[322]},
      {stage0_28[84]},
      {stage0_29[72], stage0_29[73], stage0_29[74], stage0_29[75], stage0_29[76], stage0_29[77]},
      {stage1_31[12],stage1_30[24],stage1_29[65],stage1_28[122],stage1_27[162]}
   );
   gpc615_5 gpc1055 (
      {stage0_27[323], stage0_27[324], stage0_27[325], stage0_27[326], stage0_27[327]},
      {stage0_28[85]},
      {stage0_29[78], stage0_29[79], stage0_29[80], stage0_29[81], stage0_29[82], stage0_29[83]},
      {stage1_31[13],stage1_30[25],stage1_29[66],stage1_28[123],stage1_27[163]}
   );
   gpc615_5 gpc1056 (
      {stage0_27[328], stage0_27[329], stage0_27[330], stage0_27[331], stage0_27[332]},
      {stage0_28[86]},
      {stage0_29[84], stage0_29[85], stage0_29[86], stage0_29[87], stage0_29[88], stage0_29[89]},
      {stage1_31[14],stage1_30[26],stage1_29[67],stage1_28[124],stage1_27[164]}
   );
   gpc615_5 gpc1057 (
      {stage0_27[333], stage0_27[334], stage0_27[335], stage0_27[336], stage0_27[337]},
      {stage0_28[87]},
      {stage0_29[90], stage0_29[91], stage0_29[92], stage0_29[93], stage0_29[94], stage0_29[95]},
      {stage1_31[15],stage1_30[27],stage1_29[68],stage1_28[125],stage1_27[165]}
   );
   gpc615_5 gpc1058 (
      {stage0_27[338], stage0_27[339], stage0_27[340], stage0_27[341], stage0_27[342]},
      {stage0_28[88]},
      {stage0_29[96], stage0_29[97], stage0_29[98], stage0_29[99], stage0_29[100], stage0_29[101]},
      {stage1_31[16],stage1_30[28],stage1_29[69],stage1_28[126],stage1_27[166]}
   );
   gpc615_5 gpc1059 (
      {stage0_27[343], stage0_27[344], stage0_27[345], stage0_27[346], stage0_27[347]},
      {stage0_28[89]},
      {stage0_29[102], stage0_29[103], stage0_29[104], stage0_29[105], stage0_29[106], stage0_29[107]},
      {stage1_31[17],stage1_30[29],stage1_29[70],stage1_28[127],stage1_27[167]}
   );
   gpc615_5 gpc1060 (
      {stage0_27[348], stage0_27[349], stage0_27[350], stage0_27[351], stage0_27[352]},
      {stage0_28[90]},
      {stage0_29[108], stage0_29[109], stage0_29[110], stage0_29[111], stage0_29[112], stage0_29[113]},
      {stage1_31[18],stage1_30[30],stage1_29[71],stage1_28[128],stage1_27[168]}
   );
   gpc615_5 gpc1061 (
      {stage0_27[353], stage0_27[354], stage0_27[355], stage0_27[356], stage0_27[357]},
      {stage0_28[91]},
      {stage0_29[114], stage0_29[115], stage0_29[116], stage0_29[117], stage0_29[118], stage0_29[119]},
      {stage1_31[19],stage1_30[31],stage1_29[72],stage1_28[129],stage1_27[169]}
   );
   gpc615_5 gpc1062 (
      {stage0_27[358], stage0_27[359], stage0_27[360], stage0_27[361], stage0_27[362]},
      {stage0_28[92]},
      {stage0_29[120], stage0_29[121], stage0_29[122], stage0_29[123], stage0_29[124], stage0_29[125]},
      {stage1_31[20],stage1_30[32],stage1_29[73],stage1_28[130],stage1_27[170]}
   );
   gpc615_5 gpc1063 (
      {stage0_27[363], stage0_27[364], stage0_27[365], stage0_27[366], stage0_27[367]},
      {stage0_28[93]},
      {stage0_29[126], stage0_29[127], stage0_29[128], stage0_29[129], stage0_29[130], stage0_29[131]},
      {stage1_31[21],stage1_30[33],stage1_29[74],stage1_28[131],stage1_27[171]}
   );
   gpc615_5 gpc1064 (
      {stage0_27[368], stage0_27[369], stage0_27[370], stage0_27[371], stage0_27[372]},
      {stage0_28[94]},
      {stage0_29[132], stage0_29[133], stage0_29[134], stage0_29[135], stage0_29[136], stage0_29[137]},
      {stage1_31[22],stage1_30[34],stage1_29[75],stage1_28[132],stage1_27[172]}
   );
   gpc615_5 gpc1065 (
      {stage0_27[373], stage0_27[374], stage0_27[375], stage0_27[376], stage0_27[377]},
      {stage0_28[95]},
      {stage0_29[138], stage0_29[139], stage0_29[140], stage0_29[141], stage0_29[142], stage0_29[143]},
      {stage1_31[23],stage1_30[35],stage1_29[76],stage1_28[133],stage1_27[173]}
   );
   gpc615_5 gpc1066 (
      {stage0_27[378], stage0_27[379], stage0_27[380], stage0_27[381], stage0_27[382]},
      {stage0_28[96]},
      {stage0_29[144], stage0_29[145], stage0_29[146], stage0_29[147], stage0_29[148], stage0_29[149]},
      {stage1_31[24],stage1_30[36],stage1_29[77],stage1_28[134],stage1_27[174]}
   );
   gpc615_5 gpc1067 (
      {stage0_27[383], stage0_27[384], stage0_27[385], stage0_27[386], stage0_27[387]},
      {stage0_28[97]},
      {stage0_29[150], stage0_29[151], stage0_29[152], stage0_29[153], stage0_29[154], stage0_29[155]},
      {stage1_31[25],stage1_30[37],stage1_29[78],stage1_28[135],stage1_27[175]}
   );
   gpc615_5 gpc1068 (
      {stage0_27[388], stage0_27[389], stage0_27[390], stage0_27[391], stage0_27[392]},
      {stage0_28[98]},
      {stage0_29[156], stage0_29[157], stage0_29[158], stage0_29[159], stage0_29[160], stage0_29[161]},
      {stage1_31[26],stage1_30[38],stage1_29[79],stage1_28[136],stage1_27[176]}
   );
   gpc615_5 gpc1069 (
      {stage0_27[393], stage0_27[394], stage0_27[395], stage0_27[396], stage0_27[397]},
      {stage0_28[99]},
      {stage0_29[162], stage0_29[163], stage0_29[164], stage0_29[165], stage0_29[166], stage0_29[167]},
      {stage1_31[27],stage1_30[39],stage1_29[80],stage1_28[137],stage1_27[177]}
   );
   gpc615_5 gpc1070 (
      {stage0_27[398], stage0_27[399], stage0_27[400], stage0_27[401], stage0_27[402]},
      {stage0_28[100]},
      {stage0_29[168], stage0_29[169], stage0_29[170], stage0_29[171], stage0_29[172], stage0_29[173]},
      {stage1_31[28],stage1_30[40],stage1_29[81],stage1_28[138],stage1_27[178]}
   );
   gpc615_5 gpc1071 (
      {stage0_27[403], stage0_27[404], stage0_27[405], stage0_27[406], stage0_27[407]},
      {stage0_28[101]},
      {stage0_29[174], stage0_29[175], stage0_29[176], stage0_29[177], stage0_29[178], stage0_29[179]},
      {stage1_31[29],stage1_30[41],stage1_29[82],stage1_28[139],stage1_27[179]}
   );
   gpc615_5 gpc1072 (
      {stage0_27[408], stage0_27[409], stage0_27[410], stage0_27[411], stage0_27[412]},
      {stage0_28[102]},
      {stage0_29[180], stage0_29[181], stage0_29[182], stage0_29[183], stage0_29[184], stage0_29[185]},
      {stage1_31[30],stage1_30[42],stage1_29[83],stage1_28[140],stage1_27[180]}
   );
   gpc615_5 gpc1073 (
      {stage0_27[413], stage0_27[414], stage0_27[415], stage0_27[416], stage0_27[417]},
      {stage0_28[103]},
      {stage0_29[186], stage0_29[187], stage0_29[188], stage0_29[189], stage0_29[190], stage0_29[191]},
      {stage1_31[31],stage1_30[43],stage1_29[84],stage1_28[141],stage1_27[181]}
   );
   gpc615_5 gpc1074 (
      {stage0_27[418], stage0_27[419], stage0_27[420], stage0_27[421], stage0_27[422]},
      {stage0_28[104]},
      {stage0_29[192], stage0_29[193], stage0_29[194], stage0_29[195], stage0_29[196], stage0_29[197]},
      {stage1_31[32],stage1_30[44],stage1_29[85],stage1_28[142],stage1_27[182]}
   );
   gpc615_5 gpc1075 (
      {stage0_27[423], stage0_27[424], stage0_27[425], stage0_27[426], stage0_27[427]},
      {stage0_28[105]},
      {stage0_29[198], stage0_29[199], stage0_29[200], stage0_29[201], stage0_29[202], stage0_29[203]},
      {stage1_31[33],stage1_30[45],stage1_29[86],stage1_28[143],stage1_27[183]}
   );
   gpc615_5 gpc1076 (
      {stage0_27[428], stage0_27[429], stage0_27[430], stage0_27[431], stage0_27[432]},
      {stage0_28[106]},
      {stage0_29[204], stage0_29[205], stage0_29[206], stage0_29[207], stage0_29[208], stage0_29[209]},
      {stage1_31[34],stage1_30[46],stage1_29[87],stage1_28[144],stage1_27[184]}
   );
   gpc615_5 gpc1077 (
      {stage0_27[433], stage0_27[434], stage0_27[435], stage0_27[436], stage0_27[437]},
      {stage0_28[107]},
      {stage0_29[210], stage0_29[211], stage0_29[212], stage0_29[213], stage0_29[214], stage0_29[215]},
      {stage1_31[35],stage1_30[47],stage1_29[88],stage1_28[145],stage1_27[185]}
   );
   gpc615_5 gpc1078 (
      {stage0_27[438], stage0_27[439], stage0_27[440], stage0_27[441], stage0_27[442]},
      {stage0_28[108]},
      {stage0_29[216], stage0_29[217], stage0_29[218], stage0_29[219], stage0_29[220], stage0_29[221]},
      {stage1_31[36],stage1_30[48],stage1_29[89],stage1_28[146],stage1_27[186]}
   );
   gpc615_5 gpc1079 (
      {stage0_27[443], stage0_27[444], stage0_27[445], stage0_27[446], stage0_27[447]},
      {stage0_28[109]},
      {stage0_29[222], stage0_29[223], stage0_29[224], stage0_29[225], stage0_29[226], stage0_29[227]},
      {stage1_31[37],stage1_30[49],stage1_29[90],stage1_28[147],stage1_27[187]}
   );
   gpc615_5 gpc1080 (
      {stage0_27[448], stage0_27[449], stage0_27[450], stage0_27[451], stage0_27[452]},
      {stage0_28[110]},
      {stage0_29[228], stage0_29[229], stage0_29[230], stage0_29[231], stage0_29[232], stage0_29[233]},
      {stage1_31[38],stage1_30[50],stage1_29[91],stage1_28[148],stage1_27[188]}
   );
   gpc615_5 gpc1081 (
      {stage0_27[453], stage0_27[454], stage0_27[455], stage0_27[456], stage0_27[457]},
      {stage0_28[111]},
      {stage0_29[234], stage0_29[235], stage0_29[236], stage0_29[237], stage0_29[238], stage0_29[239]},
      {stage1_31[39],stage1_30[51],stage1_29[92],stage1_28[149],stage1_27[189]}
   );
   gpc615_5 gpc1082 (
      {stage0_27[458], stage0_27[459], stage0_27[460], stage0_27[461], stage0_27[462]},
      {stage0_28[112]},
      {stage0_29[240], stage0_29[241], stage0_29[242], stage0_29[243], stage0_29[244], stage0_29[245]},
      {stage1_31[40],stage1_30[52],stage1_29[93],stage1_28[150],stage1_27[190]}
   );
   gpc615_5 gpc1083 (
      {stage0_27[463], stage0_27[464], stage0_27[465], stage0_27[466], stage0_27[467]},
      {stage0_28[113]},
      {stage0_29[246], stage0_29[247], stage0_29[248], stage0_29[249], stage0_29[250], stage0_29[251]},
      {stage1_31[41],stage1_30[53],stage1_29[94],stage1_28[151],stage1_27[191]}
   );
   gpc615_5 gpc1084 (
      {stage0_27[468], stage0_27[469], stage0_27[470], stage0_27[471], stage0_27[472]},
      {stage0_28[114]},
      {stage0_29[252], stage0_29[253], stage0_29[254], stage0_29[255], stage0_29[256], stage0_29[257]},
      {stage1_31[42],stage1_30[54],stage1_29[95],stage1_28[152],stage1_27[192]}
   );
   gpc606_5 gpc1085 (
      {stage0_28[115], stage0_28[116], stage0_28[117], stage0_28[118], stage0_28[119], stage0_28[120]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[43],stage1_30[55],stage1_29[96],stage1_28[153]}
   );
   gpc606_5 gpc1086 (
      {stage0_28[121], stage0_28[122], stage0_28[123], stage0_28[124], stage0_28[125], stage0_28[126]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[44],stage1_30[56],stage1_29[97],stage1_28[154]}
   );
   gpc606_5 gpc1087 (
      {stage0_28[127], stage0_28[128], stage0_28[129], stage0_28[130], stage0_28[131], stage0_28[132]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[45],stage1_30[57],stage1_29[98],stage1_28[155]}
   );
   gpc606_5 gpc1088 (
      {stage0_28[133], stage0_28[134], stage0_28[135], stage0_28[136], stage0_28[137], stage0_28[138]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[46],stage1_30[58],stage1_29[99],stage1_28[156]}
   );
   gpc606_5 gpc1089 (
      {stage0_28[139], stage0_28[140], stage0_28[141], stage0_28[142], stage0_28[143], stage0_28[144]},
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage1_32[4],stage1_31[47],stage1_30[59],stage1_29[100],stage1_28[157]}
   );
   gpc606_5 gpc1090 (
      {stage0_28[145], stage0_28[146], stage0_28[147], stage0_28[148], stage0_28[149], stage0_28[150]},
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage1_32[5],stage1_31[48],stage1_30[60],stage1_29[101],stage1_28[158]}
   );
   gpc606_5 gpc1091 (
      {stage0_28[151], stage0_28[152], stage0_28[153], stage0_28[154], stage0_28[155], stage0_28[156]},
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage1_32[6],stage1_31[49],stage1_30[61],stage1_29[102],stage1_28[159]}
   );
   gpc606_5 gpc1092 (
      {stage0_28[157], stage0_28[158], stage0_28[159], stage0_28[160], stage0_28[161], stage0_28[162]},
      {stage0_30[42], stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47]},
      {stage1_32[7],stage1_31[50],stage1_30[62],stage1_29[103],stage1_28[160]}
   );
   gpc606_5 gpc1093 (
      {stage0_28[163], stage0_28[164], stage0_28[165], stage0_28[166], stage0_28[167], stage0_28[168]},
      {stage0_30[48], stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53]},
      {stage1_32[8],stage1_31[51],stage1_30[63],stage1_29[104],stage1_28[161]}
   );
   gpc606_5 gpc1094 (
      {stage0_28[169], stage0_28[170], stage0_28[171], stage0_28[172], stage0_28[173], stage0_28[174]},
      {stage0_30[54], stage0_30[55], stage0_30[56], stage0_30[57], stage0_30[58], stage0_30[59]},
      {stage1_32[9],stage1_31[52],stage1_30[64],stage1_29[105],stage1_28[162]}
   );
   gpc606_5 gpc1095 (
      {stage0_28[175], stage0_28[176], stage0_28[177], stage0_28[178], stage0_28[179], stage0_28[180]},
      {stage0_30[60], stage0_30[61], stage0_30[62], stage0_30[63], stage0_30[64], stage0_30[65]},
      {stage1_32[10],stage1_31[53],stage1_30[65],stage1_29[106],stage1_28[163]}
   );
   gpc606_5 gpc1096 (
      {stage0_28[181], stage0_28[182], stage0_28[183], stage0_28[184], stage0_28[185], stage0_28[186]},
      {stage0_30[66], stage0_30[67], stage0_30[68], stage0_30[69], stage0_30[70], stage0_30[71]},
      {stage1_32[11],stage1_31[54],stage1_30[66],stage1_29[107],stage1_28[164]}
   );
   gpc606_5 gpc1097 (
      {stage0_28[187], stage0_28[188], stage0_28[189], stage0_28[190], stage0_28[191], stage0_28[192]},
      {stage0_30[72], stage0_30[73], stage0_30[74], stage0_30[75], stage0_30[76], stage0_30[77]},
      {stage1_32[12],stage1_31[55],stage1_30[67],stage1_29[108],stage1_28[165]}
   );
   gpc606_5 gpc1098 (
      {stage0_28[193], stage0_28[194], stage0_28[195], stage0_28[196], stage0_28[197], stage0_28[198]},
      {stage0_30[78], stage0_30[79], stage0_30[80], stage0_30[81], stage0_30[82], stage0_30[83]},
      {stage1_32[13],stage1_31[56],stage1_30[68],stage1_29[109],stage1_28[166]}
   );
   gpc606_5 gpc1099 (
      {stage0_28[199], stage0_28[200], stage0_28[201], stage0_28[202], stage0_28[203], stage0_28[204]},
      {stage0_30[84], stage0_30[85], stage0_30[86], stage0_30[87], stage0_30[88], stage0_30[89]},
      {stage1_32[14],stage1_31[57],stage1_30[69],stage1_29[110],stage1_28[167]}
   );
   gpc606_5 gpc1100 (
      {stage0_28[205], stage0_28[206], stage0_28[207], stage0_28[208], stage0_28[209], stage0_28[210]},
      {stage0_30[90], stage0_30[91], stage0_30[92], stage0_30[93], stage0_30[94], stage0_30[95]},
      {stage1_32[15],stage1_31[58],stage1_30[70],stage1_29[111],stage1_28[168]}
   );
   gpc606_5 gpc1101 (
      {stage0_28[211], stage0_28[212], stage0_28[213], stage0_28[214], stage0_28[215], stage0_28[216]},
      {stage0_30[96], stage0_30[97], stage0_30[98], stage0_30[99], stage0_30[100], stage0_30[101]},
      {stage1_32[16],stage1_31[59],stage1_30[71],stage1_29[112],stage1_28[169]}
   );
   gpc606_5 gpc1102 (
      {stage0_28[217], stage0_28[218], stage0_28[219], stage0_28[220], stage0_28[221], stage0_28[222]},
      {stage0_30[102], stage0_30[103], stage0_30[104], stage0_30[105], stage0_30[106], stage0_30[107]},
      {stage1_32[17],stage1_31[60],stage1_30[72],stage1_29[113],stage1_28[170]}
   );
   gpc606_5 gpc1103 (
      {stage0_28[223], stage0_28[224], stage0_28[225], stage0_28[226], stage0_28[227], stage0_28[228]},
      {stage0_30[108], stage0_30[109], stage0_30[110], stage0_30[111], stage0_30[112], stage0_30[113]},
      {stage1_32[18],stage1_31[61],stage1_30[73],stage1_29[114],stage1_28[171]}
   );
   gpc606_5 gpc1104 (
      {stage0_28[229], stage0_28[230], stage0_28[231], stage0_28[232], stage0_28[233], stage0_28[234]},
      {stage0_30[114], stage0_30[115], stage0_30[116], stage0_30[117], stage0_30[118], stage0_30[119]},
      {stage1_32[19],stage1_31[62],stage1_30[74],stage1_29[115],stage1_28[172]}
   );
   gpc606_5 gpc1105 (
      {stage0_28[235], stage0_28[236], stage0_28[237], stage0_28[238], stage0_28[239], stage0_28[240]},
      {stage0_30[120], stage0_30[121], stage0_30[122], stage0_30[123], stage0_30[124], stage0_30[125]},
      {stage1_32[20],stage1_31[63],stage1_30[75],stage1_29[116],stage1_28[173]}
   );
   gpc606_5 gpc1106 (
      {stage0_28[241], stage0_28[242], stage0_28[243], stage0_28[244], stage0_28[245], stage0_28[246]},
      {stage0_30[126], stage0_30[127], stage0_30[128], stage0_30[129], stage0_30[130], stage0_30[131]},
      {stage1_32[21],stage1_31[64],stage1_30[76],stage1_29[117],stage1_28[174]}
   );
   gpc606_5 gpc1107 (
      {stage0_28[247], stage0_28[248], stage0_28[249], stage0_28[250], stage0_28[251], stage0_28[252]},
      {stage0_30[132], stage0_30[133], stage0_30[134], stage0_30[135], stage0_30[136], stage0_30[137]},
      {stage1_32[22],stage1_31[65],stage1_30[77],stage1_29[118],stage1_28[175]}
   );
   gpc606_5 gpc1108 (
      {stage0_28[253], stage0_28[254], stage0_28[255], stage0_28[256], stage0_28[257], stage0_28[258]},
      {stage0_30[138], stage0_30[139], stage0_30[140], stage0_30[141], stage0_30[142], stage0_30[143]},
      {stage1_32[23],stage1_31[66],stage1_30[78],stage1_29[119],stage1_28[176]}
   );
   gpc606_5 gpc1109 (
      {stage0_28[259], stage0_28[260], stage0_28[261], stage0_28[262], stage0_28[263], stage0_28[264]},
      {stage0_30[144], stage0_30[145], stage0_30[146], stage0_30[147], stage0_30[148], stage0_30[149]},
      {stage1_32[24],stage1_31[67],stage1_30[79],stage1_29[120],stage1_28[177]}
   );
   gpc606_5 gpc1110 (
      {stage0_28[265], stage0_28[266], stage0_28[267], stage0_28[268], stage0_28[269], stage0_28[270]},
      {stage0_30[150], stage0_30[151], stage0_30[152], stage0_30[153], stage0_30[154], stage0_30[155]},
      {stage1_32[25],stage1_31[68],stage1_30[80],stage1_29[121],stage1_28[178]}
   );
   gpc606_5 gpc1111 (
      {stage0_28[271], stage0_28[272], stage0_28[273], stage0_28[274], stage0_28[275], stage0_28[276]},
      {stage0_30[156], stage0_30[157], stage0_30[158], stage0_30[159], stage0_30[160], stage0_30[161]},
      {stage1_32[26],stage1_31[69],stage1_30[81],stage1_29[122],stage1_28[179]}
   );
   gpc606_5 gpc1112 (
      {stage0_28[277], stage0_28[278], stage0_28[279], stage0_28[280], stage0_28[281], stage0_28[282]},
      {stage0_30[162], stage0_30[163], stage0_30[164], stage0_30[165], stage0_30[166], stage0_30[167]},
      {stage1_32[27],stage1_31[70],stage1_30[82],stage1_29[123],stage1_28[180]}
   );
   gpc606_5 gpc1113 (
      {stage0_28[283], stage0_28[284], stage0_28[285], stage0_28[286], stage0_28[287], stage0_28[288]},
      {stage0_30[168], stage0_30[169], stage0_30[170], stage0_30[171], stage0_30[172], stage0_30[173]},
      {stage1_32[28],stage1_31[71],stage1_30[83],stage1_29[124],stage1_28[181]}
   );
   gpc606_5 gpc1114 (
      {stage0_28[289], stage0_28[290], stage0_28[291], stage0_28[292], stage0_28[293], stage0_28[294]},
      {stage0_30[174], stage0_30[175], stage0_30[176], stage0_30[177], stage0_30[178], stage0_30[179]},
      {stage1_32[29],stage1_31[72],stage1_30[84],stage1_29[125],stage1_28[182]}
   );
   gpc606_5 gpc1115 (
      {stage0_28[295], stage0_28[296], stage0_28[297], stage0_28[298], stage0_28[299], stage0_28[300]},
      {stage0_30[180], stage0_30[181], stage0_30[182], stage0_30[183], stage0_30[184], stage0_30[185]},
      {stage1_32[30],stage1_31[73],stage1_30[85],stage1_29[126],stage1_28[183]}
   );
   gpc606_5 gpc1116 (
      {stage0_28[301], stage0_28[302], stage0_28[303], stage0_28[304], stage0_28[305], stage0_28[306]},
      {stage0_30[186], stage0_30[187], stage0_30[188], stage0_30[189], stage0_30[190], stage0_30[191]},
      {stage1_32[31],stage1_31[74],stage1_30[86],stage1_29[127],stage1_28[184]}
   );
   gpc606_5 gpc1117 (
      {stage0_28[307], stage0_28[308], stage0_28[309], stage0_28[310], stage0_28[311], stage0_28[312]},
      {stage0_30[192], stage0_30[193], stage0_30[194], stage0_30[195], stage0_30[196], stage0_30[197]},
      {stage1_32[32],stage1_31[75],stage1_30[87],stage1_29[128],stage1_28[185]}
   );
   gpc606_5 gpc1118 (
      {stage0_28[313], stage0_28[314], stage0_28[315], stage0_28[316], stage0_28[317], stage0_28[318]},
      {stage0_30[198], stage0_30[199], stage0_30[200], stage0_30[201], stage0_30[202], stage0_30[203]},
      {stage1_32[33],stage1_31[76],stage1_30[88],stage1_29[129],stage1_28[186]}
   );
   gpc606_5 gpc1119 (
      {stage0_28[319], stage0_28[320], stage0_28[321], stage0_28[322], stage0_28[323], stage0_28[324]},
      {stage0_30[204], stage0_30[205], stage0_30[206], stage0_30[207], stage0_30[208], stage0_30[209]},
      {stage1_32[34],stage1_31[77],stage1_30[89],stage1_29[130],stage1_28[187]}
   );
   gpc606_5 gpc1120 (
      {stage0_28[325], stage0_28[326], stage0_28[327], stage0_28[328], stage0_28[329], stage0_28[330]},
      {stage0_30[210], stage0_30[211], stage0_30[212], stage0_30[213], stage0_30[214], stage0_30[215]},
      {stage1_32[35],stage1_31[78],stage1_30[90],stage1_29[131],stage1_28[188]}
   );
   gpc606_5 gpc1121 (
      {stage0_28[331], stage0_28[332], stage0_28[333], stage0_28[334], stage0_28[335], stage0_28[336]},
      {stage0_30[216], stage0_30[217], stage0_30[218], stage0_30[219], stage0_30[220], stage0_30[221]},
      {stage1_32[36],stage1_31[79],stage1_30[91],stage1_29[132],stage1_28[189]}
   );
   gpc606_5 gpc1122 (
      {stage0_28[337], stage0_28[338], stage0_28[339], stage0_28[340], stage0_28[341], stage0_28[342]},
      {stage0_30[222], stage0_30[223], stage0_30[224], stage0_30[225], stage0_30[226], stage0_30[227]},
      {stage1_32[37],stage1_31[80],stage1_30[92],stage1_29[133],stage1_28[190]}
   );
   gpc606_5 gpc1123 (
      {stage0_28[343], stage0_28[344], stage0_28[345], stage0_28[346], stage0_28[347], stage0_28[348]},
      {stage0_30[228], stage0_30[229], stage0_30[230], stage0_30[231], stage0_30[232], stage0_30[233]},
      {stage1_32[38],stage1_31[81],stage1_30[93],stage1_29[134],stage1_28[191]}
   );
   gpc606_5 gpc1124 (
      {stage0_28[349], stage0_28[350], stage0_28[351], stage0_28[352], stage0_28[353], stage0_28[354]},
      {stage0_30[234], stage0_30[235], stage0_30[236], stage0_30[237], stage0_30[238], stage0_30[239]},
      {stage1_32[39],stage1_31[82],stage1_30[94],stage1_29[135],stage1_28[192]}
   );
   gpc606_5 gpc1125 (
      {stage0_28[355], stage0_28[356], stage0_28[357], stage0_28[358], stage0_28[359], stage0_28[360]},
      {stage0_30[240], stage0_30[241], stage0_30[242], stage0_30[243], stage0_30[244], stage0_30[245]},
      {stage1_32[40],stage1_31[83],stage1_30[95],stage1_29[136],stage1_28[193]}
   );
   gpc606_5 gpc1126 (
      {stage0_28[361], stage0_28[362], stage0_28[363], stage0_28[364], stage0_28[365], stage0_28[366]},
      {stage0_30[246], stage0_30[247], stage0_30[248], stage0_30[249], stage0_30[250], stage0_30[251]},
      {stage1_32[41],stage1_31[84],stage1_30[96],stage1_29[137],stage1_28[194]}
   );
   gpc606_5 gpc1127 (
      {stage0_28[367], stage0_28[368], stage0_28[369], stage0_28[370], stage0_28[371], stage0_28[372]},
      {stage0_30[252], stage0_30[253], stage0_30[254], stage0_30[255], stage0_30[256], stage0_30[257]},
      {stage1_32[42],stage1_31[85],stage1_30[97],stage1_29[138],stage1_28[195]}
   );
   gpc606_5 gpc1128 (
      {stage0_28[373], stage0_28[374], stage0_28[375], stage0_28[376], stage0_28[377], stage0_28[378]},
      {stage0_30[258], stage0_30[259], stage0_30[260], stage0_30[261], stage0_30[262], stage0_30[263]},
      {stage1_32[43],stage1_31[86],stage1_30[98],stage1_29[139],stage1_28[196]}
   );
   gpc606_5 gpc1129 (
      {stage0_28[379], stage0_28[380], stage0_28[381], stage0_28[382], stage0_28[383], stage0_28[384]},
      {stage0_30[264], stage0_30[265], stage0_30[266], stage0_30[267], stage0_30[268], stage0_30[269]},
      {stage1_32[44],stage1_31[87],stage1_30[99],stage1_29[140],stage1_28[197]}
   );
   gpc606_5 gpc1130 (
      {stage0_28[385], stage0_28[386], stage0_28[387], stage0_28[388], stage0_28[389], stage0_28[390]},
      {stage0_30[270], stage0_30[271], stage0_30[272], stage0_30[273], stage0_30[274], stage0_30[275]},
      {stage1_32[45],stage1_31[88],stage1_30[100],stage1_29[141],stage1_28[198]}
   );
   gpc606_5 gpc1131 (
      {stage0_28[391], stage0_28[392], stage0_28[393], stage0_28[394], stage0_28[395], stage0_28[396]},
      {stage0_30[276], stage0_30[277], stage0_30[278], stage0_30[279], stage0_30[280], stage0_30[281]},
      {stage1_32[46],stage1_31[89],stage1_30[101],stage1_29[142],stage1_28[199]}
   );
   gpc606_5 gpc1132 (
      {stage0_28[397], stage0_28[398], stage0_28[399], stage0_28[400], stage0_28[401], stage0_28[402]},
      {stage0_30[282], stage0_30[283], stage0_30[284], stage0_30[285], stage0_30[286], stage0_30[287]},
      {stage1_32[47],stage1_31[90],stage1_30[102],stage1_29[143],stage1_28[200]}
   );
   gpc606_5 gpc1133 (
      {stage0_28[403], stage0_28[404], stage0_28[405], stage0_28[406], stage0_28[407], stage0_28[408]},
      {stage0_30[288], stage0_30[289], stage0_30[290], stage0_30[291], stage0_30[292], stage0_30[293]},
      {stage1_32[48],stage1_31[91],stage1_30[103],stage1_29[144],stage1_28[201]}
   );
   gpc606_5 gpc1134 (
      {stage0_28[409], stage0_28[410], stage0_28[411], stage0_28[412], stage0_28[413], stage0_28[414]},
      {stage0_30[294], stage0_30[295], stage0_30[296], stage0_30[297], stage0_30[298], stage0_30[299]},
      {stage1_32[49],stage1_31[92],stage1_30[104],stage1_29[145],stage1_28[202]}
   );
   gpc606_5 gpc1135 (
      {stage0_28[415], stage0_28[416], stage0_28[417], stage0_28[418], stage0_28[419], stage0_28[420]},
      {stage0_30[300], stage0_30[301], stage0_30[302], stage0_30[303], stage0_30[304], stage0_30[305]},
      {stage1_32[50],stage1_31[93],stage1_30[105],stage1_29[146],stage1_28[203]}
   );
   gpc606_5 gpc1136 (
      {stage0_28[421], stage0_28[422], stage0_28[423], stage0_28[424], stage0_28[425], stage0_28[426]},
      {stage0_30[306], stage0_30[307], stage0_30[308], stage0_30[309], stage0_30[310], stage0_30[311]},
      {stage1_32[51],stage1_31[94],stage1_30[106],stage1_29[147],stage1_28[204]}
   );
   gpc606_5 gpc1137 (
      {stage0_28[427], stage0_28[428], stage0_28[429], stage0_28[430], stage0_28[431], stage0_28[432]},
      {stage0_30[312], stage0_30[313], stage0_30[314], stage0_30[315], stage0_30[316], stage0_30[317]},
      {stage1_32[52],stage1_31[95],stage1_30[107],stage1_29[148],stage1_28[205]}
   );
   gpc606_5 gpc1138 (
      {stage0_28[433], stage0_28[434], stage0_28[435], stage0_28[436], stage0_28[437], stage0_28[438]},
      {stage0_30[318], stage0_30[319], stage0_30[320], stage0_30[321], stage0_30[322], stage0_30[323]},
      {stage1_32[53],stage1_31[96],stage1_30[108],stage1_29[149],stage1_28[206]}
   );
   gpc606_5 gpc1139 (
      {stage0_28[439], stage0_28[440], stage0_28[441], stage0_28[442], stage0_28[443], stage0_28[444]},
      {stage0_30[324], stage0_30[325], stage0_30[326], stage0_30[327], stage0_30[328], stage0_30[329]},
      {stage1_32[54],stage1_31[97],stage1_30[109],stage1_29[150],stage1_28[207]}
   );
   gpc606_5 gpc1140 (
      {stage0_28[445], stage0_28[446], stage0_28[447], stage0_28[448], stage0_28[449], stage0_28[450]},
      {stage0_30[330], stage0_30[331], stage0_30[332], stage0_30[333], stage0_30[334], stage0_30[335]},
      {stage1_32[55],stage1_31[98],stage1_30[110],stage1_29[151],stage1_28[208]}
   );
   gpc606_5 gpc1141 (
      {stage0_28[451], stage0_28[452], stage0_28[453], stage0_28[454], stage0_28[455], stage0_28[456]},
      {stage0_30[336], stage0_30[337], stage0_30[338], stage0_30[339], stage0_30[340], stage0_30[341]},
      {stage1_32[56],stage1_31[99],stage1_30[111],stage1_29[152],stage1_28[209]}
   );
   gpc606_5 gpc1142 (
      {stage0_28[457], stage0_28[458], stage0_28[459], stage0_28[460], stage0_28[461], stage0_28[462]},
      {stage0_30[342], stage0_30[343], stage0_30[344], stage0_30[345], stage0_30[346], stage0_30[347]},
      {stage1_32[57],stage1_31[100],stage1_30[112],stage1_29[153],stage1_28[210]}
   );
   gpc606_5 gpc1143 (
      {stage0_28[463], stage0_28[464], stage0_28[465], stage0_28[466], stage0_28[467], stage0_28[468]},
      {stage0_30[348], stage0_30[349], stage0_30[350], stage0_30[351], stage0_30[352], stage0_30[353]},
      {stage1_32[58],stage1_31[101],stage1_30[113],stage1_29[154],stage1_28[211]}
   );
   gpc606_5 gpc1144 (
      {stage0_28[469], stage0_28[470], stage0_28[471], stage0_28[472], stage0_28[473], stage0_28[474]},
      {stage0_30[354], stage0_30[355], stage0_30[356], stage0_30[357], stage0_30[358], stage0_30[359]},
      {stage1_32[59],stage1_31[102],stage1_30[114],stage1_29[155],stage1_28[212]}
   );
   gpc606_5 gpc1145 (
      {stage0_29[258], stage0_29[259], stage0_29[260], stage0_29[261], stage0_29[262], stage0_29[263]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[60],stage1_31[103],stage1_30[115],stage1_29[156]}
   );
   gpc606_5 gpc1146 (
      {stage0_29[264], stage0_29[265], stage0_29[266], stage0_29[267], stage0_29[268], stage0_29[269]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[61],stage1_31[104],stage1_30[116],stage1_29[157]}
   );
   gpc606_5 gpc1147 (
      {stage0_29[270], stage0_29[271], stage0_29[272], stage0_29[273], stage0_29[274], stage0_29[275]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[62],stage1_31[105],stage1_30[117],stage1_29[158]}
   );
   gpc606_5 gpc1148 (
      {stage0_29[276], stage0_29[277], stage0_29[278], stage0_29[279], stage0_29[280], stage0_29[281]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[63],stage1_31[106],stage1_30[118],stage1_29[159]}
   );
   gpc606_5 gpc1149 (
      {stage0_29[282], stage0_29[283], stage0_29[284], stage0_29[285], stage0_29[286], stage0_29[287]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[64],stage1_31[107],stage1_30[119],stage1_29[160]}
   );
   gpc606_5 gpc1150 (
      {stage0_29[288], stage0_29[289], stage0_29[290], stage0_29[291], stage0_29[292], stage0_29[293]},
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage1_33[5],stage1_32[65],stage1_31[108],stage1_30[120],stage1_29[161]}
   );
   gpc606_5 gpc1151 (
      {stage0_29[294], stage0_29[295], stage0_29[296], stage0_29[297], stage0_29[298], stage0_29[299]},
      {stage0_31[36], stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41]},
      {stage1_33[6],stage1_32[66],stage1_31[109],stage1_30[121],stage1_29[162]}
   );
   gpc606_5 gpc1152 (
      {stage0_29[300], stage0_29[301], stage0_29[302], stage0_29[303], stage0_29[304], stage0_29[305]},
      {stage0_31[42], stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47]},
      {stage1_33[7],stage1_32[67],stage1_31[110],stage1_30[122],stage1_29[163]}
   );
   gpc606_5 gpc1153 (
      {stage0_29[306], stage0_29[307], stage0_29[308], stage0_29[309], stage0_29[310], stage0_29[311]},
      {stage0_31[48], stage0_31[49], stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53]},
      {stage1_33[8],stage1_32[68],stage1_31[111],stage1_30[123],stage1_29[164]}
   );
   gpc606_5 gpc1154 (
      {stage0_29[312], stage0_29[313], stage0_29[314], stage0_29[315], stage0_29[316], stage0_29[317]},
      {stage0_31[54], stage0_31[55], stage0_31[56], stage0_31[57], stage0_31[58], stage0_31[59]},
      {stage1_33[9],stage1_32[69],stage1_31[112],stage1_30[124],stage1_29[165]}
   );
   gpc606_5 gpc1155 (
      {stage0_29[318], stage0_29[319], stage0_29[320], stage0_29[321], stage0_29[322], stage0_29[323]},
      {stage0_31[60], stage0_31[61], stage0_31[62], stage0_31[63], stage0_31[64], stage0_31[65]},
      {stage1_33[10],stage1_32[70],stage1_31[113],stage1_30[125],stage1_29[166]}
   );
   gpc606_5 gpc1156 (
      {stage0_29[324], stage0_29[325], stage0_29[326], stage0_29[327], stage0_29[328], stage0_29[329]},
      {stage0_31[66], stage0_31[67], stage0_31[68], stage0_31[69], stage0_31[70], stage0_31[71]},
      {stage1_33[11],stage1_32[71],stage1_31[114],stage1_30[126],stage1_29[167]}
   );
   gpc606_5 gpc1157 (
      {stage0_29[330], stage0_29[331], stage0_29[332], stage0_29[333], stage0_29[334], stage0_29[335]},
      {stage0_31[72], stage0_31[73], stage0_31[74], stage0_31[75], stage0_31[76], stage0_31[77]},
      {stage1_33[12],stage1_32[72],stage1_31[115],stage1_30[127],stage1_29[168]}
   );
   gpc606_5 gpc1158 (
      {stage0_29[336], stage0_29[337], stage0_29[338], stage0_29[339], stage0_29[340], stage0_29[341]},
      {stage0_31[78], stage0_31[79], stage0_31[80], stage0_31[81], stage0_31[82], stage0_31[83]},
      {stage1_33[13],stage1_32[73],stage1_31[116],stage1_30[128],stage1_29[169]}
   );
   gpc606_5 gpc1159 (
      {stage0_29[342], stage0_29[343], stage0_29[344], stage0_29[345], stage0_29[346], stage0_29[347]},
      {stage0_31[84], stage0_31[85], stage0_31[86], stage0_31[87], stage0_31[88], stage0_31[89]},
      {stage1_33[14],stage1_32[74],stage1_31[117],stage1_30[129],stage1_29[170]}
   );
   gpc606_5 gpc1160 (
      {stage0_29[348], stage0_29[349], stage0_29[350], stage0_29[351], stage0_29[352], stage0_29[353]},
      {stage0_31[90], stage0_31[91], stage0_31[92], stage0_31[93], stage0_31[94], stage0_31[95]},
      {stage1_33[15],stage1_32[75],stage1_31[118],stage1_30[130],stage1_29[171]}
   );
   gpc606_5 gpc1161 (
      {stage0_29[354], stage0_29[355], stage0_29[356], stage0_29[357], stage0_29[358], stage0_29[359]},
      {stage0_31[96], stage0_31[97], stage0_31[98], stage0_31[99], stage0_31[100], stage0_31[101]},
      {stage1_33[16],stage1_32[76],stage1_31[119],stage1_30[131],stage1_29[172]}
   );
   gpc606_5 gpc1162 (
      {stage0_29[360], stage0_29[361], stage0_29[362], stage0_29[363], stage0_29[364], stage0_29[365]},
      {stage0_31[102], stage0_31[103], stage0_31[104], stage0_31[105], stage0_31[106], stage0_31[107]},
      {stage1_33[17],stage1_32[77],stage1_31[120],stage1_30[132],stage1_29[173]}
   );
   gpc606_5 gpc1163 (
      {stage0_29[366], stage0_29[367], stage0_29[368], stage0_29[369], stage0_29[370], stage0_29[371]},
      {stage0_31[108], stage0_31[109], stage0_31[110], stage0_31[111], stage0_31[112], stage0_31[113]},
      {stage1_33[18],stage1_32[78],stage1_31[121],stage1_30[133],stage1_29[174]}
   );
   gpc606_5 gpc1164 (
      {stage0_29[372], stage0_29[373], stage0_29[374], stage0_29[375], stage0_29[376], stage0_29[377]},
      {stage0_31[114], stage0_31[115], stage0_31[116], stage0_31[117], stage0_31[118], stage0_31[119]},
      {stage1_33[19],stage1_32[79],stage1_31[122],stage1_30[134],stage1_29[175]}
   );
   gpc606_5 gpc1165 (
      {stage0_29[378], stage0_29[379], stage0_29[380], stage0_29[381], stage0_29[382], stage0_29[383]},
      {stage0_31[120], stage0_31[121], stage0_31[122], stage0_31[123], stage0_31[124], stage0_31[125]},
      {stage1_33[20],stage1_32[80],stage1_31[123],stage1_30[135],stage1_29[176]}
   );
   gpc606_5 gpc1166 (
      {stage0_29[384], stage0_29[385], stage0_29[386], stage0_29[387], stage0_29[388], stage0_29[389]},
      {stage0_31[126], stage0_31[127], stage0_31[128], stage0_31[129], stage0_31[130], stage0_31[131]},
      {stage1_33[21],stage1_32[81],stage1_31[124],stage1_30[136],stage1_29[177]}
   );
   gpc606_5 gpc1167 (
      {stage0_29[390], stage0_29[391], stage0_29[392], stage0_29[393], stage0_29[394], stage0_29[395]},
      {stage0_31[132], stage0_31[133], stage0_31[134], stage0_31[135], stage0_31[136], stage0_31[137]},
      {stage1_33[22],stage1_32[82],stage1_31[125],stage1_30[137],stage1_29[178]}
   );
   gpc606_5 gpc1168 (
      {stage0_29[396], stage0_29[397], stage0_29[398], stage0_29[399], stage0_29[400], stage0_29[401]},
      {stage0_31[138], stage0_31[139], stage0_31[140], stage0_31[141], stage0_31[142], stage0_31[143]},
      {stage1_33[23],stage1_32[83],stage1_31[126],stage1_30[138],stage1_29[179]}
   );
   gpc606_5 gpc1169 (
      {stage0_29[402], stage0_29[403], stage0_29[404], stage0_29[405], stage0_29[406], stage0_29[407]},
      {stage0_31[144], stage0_31[145], stage0_31[146], stage0_31[147], stage0_31[148], stage0_31[149]},
      {stage1_33[24],stage1_32[84],stage1_31[127],stage1_30[139],stage1_29[180]}
   );
   gpc606_5 gpc1170 (
      {stage0_29[408], stage0_29[409], stage0_29[410], stage0_29[411], stage0_29[412], stage0_29[413]},
      {stage0_31[150], stage0_31[151], stage0_31[152], stage0_31[153], stage0_31[154], stage0_31[155]},
      {stage1_33[25],stage1_32[85],stage1_31[128],stage1_30[140],stage1_29[181]}
   );
   gpc606_5 gpc1171 (
      {stage0_29[414], stage0_29[415], stage0_29[416], stage0_29[417], stage0_29[418], stage0_29[419]},
      {stage0_31[156], stage0_31[157], stage0_31[158], stage0_31[159], stage0_31[160], stage0_31[161]},
      {stage1_33[26],stage1_32[86],stage1_31[129],stage1_30[141],stage1_29[182]}
   );
   gpc606_5 gpc1172 (
      {stage0_29[420], stage0_29[421], stage0_29[422], stage0_29[423], stage0_29[424], stage0_29[425]},
      {stage0_31[162], stage0_31[163], stage0_31[164], stage0_31[165], stage0_31[166], stage0_31[167]},
      {stage1_33[27],stage1_32[87],stage1_31[130],stage1_30[142],stage1_29[183]}
   );
   gpc606_5 gpc1173 (
      {stage0_29[426], stage0_29[427], stage0_29[428], stage0_29[429], stage0_29[430], stage0_29[431]},
      {stage0_31[168], stage0_31[169], stage0_31[170], stage0_31[171], stage0_31[172], stage0_31[173]},
      {stage1_33[28],stage1_32[88],stage1_31[131],stage1_30[143],stage1_29[184]}
   );
   gpc606_5 gpc1174 (
      {stage0_29[432], stage0_29[433], stage0_29[434], stage0_29[435], stage0_29[436], stage0_29[437]},
      {stage0_31[174], stage0_31[175], stage0_31[176], stage0_31[177], stage0_31[178], stage0_31[179]},
      {stage1_33[29],stage1_32[89],stage1_31[132],stage1_30[144],stage1_29[185]}
   );
   gpc606_5 gpc1175 (
      {stage0_29[438], stage0_29[439], stage0_29[440], stage0_29[441], stage0_29[442], stage0_29[443]},
      {stage0_31[180], stage0_31[181], stage0_31[182], stage0_31[183], stage0_31[184], stage0_31[185]},
      {stage1_33[30],stage1_32[90],stage1_31[133],stage1_30[145],stage1_29[186]}
   );
   gpc615_5 gpc1176 (
      {stage0_30[360], stage0_30[361], stage0_30[362], stage0_30[363], stage0_30[364]},
      {stage0_31[186]},
      {stage0_32[0], stage0_32[1], stage0_32[2], stage0_32[3], stage0_32[4], stage0_32[5]},
      {stage1_34[0],stage1_33[31],stage1_32[91],stage1_31[134],stage1_30[146]}
   );
   gpc615_5 gpc1177 (
      {stage0_30[365], stage0_30[366], stage0_30[367], stage0_30[368], stage0_30[369]},
      {stage0_31[187]},
      {stage0_32[6], stage0_32[7], stage0_32[8], stage0_32[9], stage0_32[10], stage0_32[11]},
      {stage1_34[1],stage1_33[32],stage1_32[92],stage1_31[135],stage1_30[147]}
   );
   gpc615_5 gpc1178 (
      {stage0_30[370], stage0_30[371], stage0_30[372], stage0_30[373], stage0_30[374]},
      {stage0_31[188]},
      {stage0_32[12], stage0_32[13], stage0_32[14], stage0_32[15], stage0_32[16], stage0_32[17]},
      {stage1_34[2],stage1_33[33],stage1_32[93],stage1_31[136],stage1_30[148]}
   );
   gpc615_5 gpc1179 (
      {stage0_30[375], stage0_30[376], stage0_30[377], stage0_30[378], stage0_30[379]},
      {stage0_31[189]},
      {stage0_32[18], stage0_32[19], stage0_32[20], stage0_32[21], stage0_32[22], stage0_32[23]},
      {stage1_34[3],stage1_33[34],stage1_32[94],stage1_31[137],stage1_30[149]}
   );
   gpc615_5 gpc1180 (
      {stage0_30[380], stage0_30[381], stage0_30[382], stage0_30[383], stage0_30[384]},
      {stage0_31[190]},
      {stage0_32[24], stage0_32[25], stage0_32[26], stage0_32[27], stage0_32[28], stage0_32[29]},
      {stage1_34[4],stage1_33[35],stage1_32[95],stage1_31[138],stage1_30[150]}
   );
   gpc615_5 gpc1181 (
      {stage0_30[385], stage0_30[386], stage0_30[387], stage0_30[388], stage0_30[389]},
      {stage0_31[191]},
      {stage0_32[30], stage0_32[31], stage0_32[32], stage0_32[33], stage0_32[34], stage0_32[35]},
      {stage1_34[5],stage1_33[36],stage1_32[96],stage1_31[139],stage1_30[151]}
   );
   gpc615_5 gpc1182 (
      {stage0_30[390], stage0_30[391], stage0_30[392], stage0_30[393], stage0_30[394]},
      {stage0_31[192]},
      {stage0_32[36], stage0_32[37], stage0_32[38], stage0_32[39], stage0_32[40], stage0_32[41]},
      {stage1_34[6],stage1_33[37],stage1_32[97],stage1_31[140],stage1_30[152]}
   );
   gpc615_5 gpc1183 (
      {stage0_30[395], stage0_30[396], stage0_30[397], stage0_30[398], stage0_30[399]},
      {stage0_31[193]},
      {stage0_32[42], stage0_32[43], stage0_32[44], stage0_32[45], stage0_32[46], stage0_32[47]},
      {stage1_34[7],stage1_33[38],stage1_32[98],stage1_31[141],stage1_30[153]}
   );
   gpc615_5 gpc1184 (
      {stage0_30[400], stage0_30[401], stage0_30[402], stage0_30[403], stage0_30[404]},
      {stage0_31[194]},
      {stage0_32[48], stage0_32[49], stage0_32[50], stage0_32[51], stage0_32[52], stage0_32[53]},
      {stage1_34[8],stage1_33[39],stage1_32[99],stage1_31[142],stage1_30[154]}
   );
   gpc615_5 gpc1185 (
      {stage0_30[405], stage0_30[406], stage0_30[407], stage0_30[408], stage0_30[409]},
      {stage0_31[195]},
      {stage0_32[54], stage0_32[55], stage0_32[56], stage0_32[57], stage0_32[58], stage0_32[59]},
      {stage1_34[9],stage1_33[40],stage1_32[100],stage1_31[143],stage1_30[155]}
   );
   gpc615_5 gpc1186 (
      {stage0_30[410], stage0_30[411], stage0_30[412], stage0_30[413], stage0_30[414]},
      {stage0_31[196]},
      {stage0_32[60], stage0_32[61], stage0_32[62], stage0_32[63], stage0_32[64], stage0_32[65]},
      {stage1_34[10],stage1_33[41],stage1_32[101],stage1_31[144],stage1_30[156]}
   );
   gpc615_5 gpc1187 (
      {stage0_30[415], stage0_30[416], stage0_30[417], stage0_30[418], stage0_30[419]},
      {stage0_31[197]},
      {stage0_32[66], stage0_32[67], stage0_32[68], stage0_32[69], stage0_32[70], stage0_32[71]},
      {stage1_34[11],stage1_33[42],stage1_32[102],stage1_31[145],stage1_30[157]}
   );
   gpc615_5 gpc1188 (
      {stage0_30[420], stage0_30[421], stage0_30[422], stage0_30[423], stage0_30[424]},
      {stage0_31[198]},
      {stage0_32[72], stage0_32[73], stage0_32[74], stage0_32[75], stage0_32[76], stage0_32[77]},
      {stage1_34[12],stage1_33[43],stage1_32[103],stage1_31[146],stage1_30[158]}
   );
   gpc615_5 gpc1189 (
      {stage0_30[425], stage0_30[426], stage0_30[427], stage0_30[428], stage0_30[429]},
      {stage0_31[199]},
      {stage0_32[78], stage0_32[79], stage0_32[80], stage0_32[81], stage0_32[82], stage0_32[83]},
      {stage1_34[13],stage1_33[44],stage1_32[104],stage1_31[147],stage1_30[159]}
   );
   gpc615_5 gpc1190 (
      {stage0_30[430], stage0_30[431], stage0_30[432], stage0_30[433], stage0_30[434]},
      {stage0_31[200]},
      {stage0_32[84], stage0_32[85], stage0_32[86], stage0_32[87], stage0_32[88], stage0_32[89]},
      {stage1_34[14],stage1_33[45],stage1_32[105],stage1_31[148],stage1_30[160]}
   );
   gpc615_5 gpc1191 (
      {stage0_30[435], stage0_30[436], stage0_30[437], stage0_30[438], stage0_30[439]},
      {stage0_31[201]},
      {stage0_32[90], stage0_32[91], stage0_32[92], stage0_32[93], stage0_32[94], stage0_32[95]},
      {stage1_34[15],stage1_33[46],stage1_32[106],stage1_31[149],stage1_30[161]}
   );
   gpc615_5 gpc1192 (
      {stage0_30[440], stage0_30[441], stage0_30[442], stage0_30[443], stage0_30[444]},
      {stage0_31[202]},
      {stage0_32[96], stage0_32[97], stage0_32[98], stage0_32[99], stage0_32[100], stage0_32[101]},
      {stage1_34[16],stage1_33[47],stage1_32[107],stage1_31[150],stage1_30[162]}
   );
   gpc615_5 gpc1193 (
      {stage0_30[445], stage0_30[446], stage0_30[447], stage0_30[448], stage0_30[449]},
      {stage0_31[203]},
      {stage0_32[102], stage0_32[103], stage0_32[104], stage0_32[105], stage0_32[106], stage0_32[107]},
      {stage1_34[17],stage1_33[48],stage1_32[108],stage1_31[151],stage1_30[163]}
   );
   gpc615_5 gpc1194 (
      {stage0_30[450], stage0_30[451], stage0_30[452], stage0_30[453], stage0_30[454]},
      {stage0_31[204]},
      {stage0_32[108], stage0_32[109], stage0_32[110], stage0_32[111], stage0_32[112], stage0_32[113]},
      {stage1_34[18],stage1_33[49],stage1_32[109],stage1_31[152],stage1_30[164]}
   );
   gpc615_5 gpc1195 (
      {stage0_30[455], stage0_30[456], stage0_30[457], stage0_30[458], stage0_30[459]},
      {stage0_31[205]},
      {stage0_32[114], stage0_32[115], stage0_32[116], stage0_32[117], stage0_32[118], stage0_32[119]},
      {stage1_34[19],stage1_33[50],stage1_32[110],stage1_31[153],stage1_30[165]}
   );
   gpc615_5 gpc1196 (
      {stage0_31[206], stage0_31[207], stage0_31[208], stage0_31[209], stage0_31[210]},
      {stage0_32[120]},
      {stage0_33[0], stage0_33[1], stage0_33[2], stage0_33[3], stage0_33[4], stage0_33[5]},
      {stage1_35[0],stage1_34[20],stage1_33[51],stage1_32[111],stage1_31[154]}
   );
   gpc615_5 gpc1197 (
      {stage0_31[211], stage0_31[212], stage0_31[213], stage0_31[214], stage0_31[215]},
      {stage0_32[121]},
      {stage0_33[6], stage0_33[7], stage0_33[8], stage0_33[9], stage0_33[10], stage0_33[11]},
      {stage1_35[1],stage1_34[21],stage1_33[52],stage1_32[112],stage1_31[155]}
   );
   gpc615_5 gpc1198 (
      {stage0_31[216], stage0_31[217], stage0_31[218], stage0_31[219], stage0_31[220]},
      {stage0_32[122]},
      {stage0_33[12], stage0_33[13], stage0_33[14], stage0_33[15], stage0_33[16], stage0_33[17]},
      {stage1_35[2],stage1_34[22],stage1_33[53],stage1_32[113],stage1_31[156]}
   );
   gpc615_5 gpc1199 (
      {stage0_31[221], stage0_31[222], stage0_31[223], stage0_31[224], stage0_31[225]},
      {stage0_32[123]},
      {stage0_33[18], stage0_33[19], stage0_33[20], stage0_33[21], stage0_33[22], stage0_33[23]},
      {stage1_35[3],stage1_34[23],stage1_33[54],stage1_32[114],stage1_31[157]}
   );
   gpc615_5 gpc1200 (
      {stage0_31[226], stage0_31[227], stage0_31[228], stage0_31[229], stage0_31[230]},
      {stage0_32[124]},
      {stage0_33[24], stage0_33[25], stage0_33[26], stage0_33[27], stage0_33[28], stage0_33[29]},
      {stage1_35[4],stage1_34[24],stage1_33[55],stage1_32[115],stage1_31[158]}
   );
   gpc615_5 gpc1201 (
      {stage0_31[231], stage0_31[232], stage0_31[233], stage0_31[234], stage0_31[235]},
      {stage0_32[125]},
      {stage0_33[30], stage0_33[31], stage0_33[32], stage0_33[33], stage0_33[34], stage0_33[35]},
      {stage1_35[5],stage1_34[25],stage1_33[56],stage1_32[116],stage1_31[159]}
   );
   gpc615_5 gpc1202 (
      {stage0_31[236], stage0_31[237], stage0_31[238], stage0_31[239], stage0_31[240]},
      {stage0_32[126]},
      {stage0_33[36], stage0_33[37], stage0_33[38], stage0_33[39], stage0_33[40], stage0_33[41]},
      {stage1_35[6],stage1_34[26],stage1_33[57],stage1_32[117],stage1_31[160]}
   );
   gpc615_5 gpc1203 (
      {stage0_31[241], stage0_31[242], stage0_31[243], stage0_31[244], stage0_31[245]},
      {stage0_32[127]},
      {stage0_33[42], stage0_33[43], stage0_33[44], stage0_33[45], stage0_33[46], stage0_33[47]},
      {stage1_35[7],stage1_34[27],stage1_33[58],stage1_32[118],stage1_31[161]}
   );
   gpc615_5 gpc1204 (
      {stage0_31[246], stage0_31[247], stage0_31[248], stage0_31[249], stage0_31[250]},
      {stage0_32[128]},
      {stage0_33[48], stage0_33[49], stage0_33[50], stage0_33[51], stage0_33[52], stage0_33[53]},
      {stage1_35[8],stage1_34[28],stage1_33[59],stage1_32[119],stage1_31[162]}
   );
   gpc615_5 gpc1205 (
      {stage0_31[251], stage0_31[252], stage0_31[253], stage0_31[254], stage0_31[255]},
      {stage0_32[129]},
      {stage0_33[54], stage0_33[55], stage0_33[56], stage0_33[57], stage0_33[58], stage0_33[59]},
      {stage1_35[9],stage1_34[29],stage1_33[60],stage1_32[120],stage1_31[163]}
   );
   gpc615_5 gpc1206 (
      {stage0_31[256], stage0_31[257], stage0_31[258], stage0_31[259], stage0_31[260]},
      {stage0_32[130]},
      {stage0_33[60], stage0_33[61], stage0_33[62], stage0_33[63], stage0_33[64], stage0_33[65]},
      {stage1_35[10],stage1_34[30],stage1_33[61],stage1_32[121],stage1_31[164]}
   );
   gpc615_5 gpc1207 (
      {stage0_31[261], stage0_31[262], stage0_31[263], stage0_31[264], stage0_31[265]},
      {stage0_32[131]},
      {stage0_33[66], stage0_33[67], stage0_33[68], stage0_33[69], stage0_33[70], stage0_33[71]},
      {stage1_35[11],stage1_34[31],stage1_33[62],stage1_32[122],stage1_31[165]}
   );
   gpc615_5 gpc1208 (
      {stage0_31[266], stage0_31[267], stage0_31[268], stage0_31[269], stage0_31[270]},
      {stage0_32[132]},
      {stage0_33[72], stage0_33[73], stage0_33[74], stage0_33[75], stage0_33[76], stage0_33[77]},
      {stage1_35[12],stage1_34[32],stage1_33[63],stage1_32[123],stage1_31[166]}
   );
   gpc615_5 gpc1209 (
      {stage0_31[271], stage0_31[272], stage0_31[273], stage0_31[274], stage0_31[275]},
      {stage0_32[133]},
      {stage0_33[78], stage0_33[79], stage0_33[80], stage0_33[81], stage0_33[82], stage0_33[83]},
      {stage1_35[13],stage1_34[33],stage1_33[64],stage1_32[124],stage1_31[167]}
   );
   gpc615_5 gpc1210 (
      {stage0_31[276], stage0_31[277], stage0_31[278], stage0_31[279], stage0_31[280]},
      {stage0_32[134]},
      {stage0_33[84], stage0_33[85], stage0_33[86], stage0_33[87], stage0_33[88], stage0_33[89]},
      {stage1_35[14],stage1_34[34],stage1_33[65],stage1_32[125],stage1_31[168]}
   );
   gpc615_5 gpc1211 (
      {stage0_31[281], stage0_31[282], stage0_31[283], stage0_31[284], stage0_31[285]},
      {stage0_32[135]},
      {stage0_33[90], stage0_33[91], stage0_33[92], stage0_33[93], stage0_33[94], stage0_33[95]},
      {stage1_35[15],stage1_34[35],stage1_33[66],stage1_32[126],stage1_31[169]}
   );
   gpc615_5 gpc1212 (
      {stage0_31[286], stage0_31[287], stage0_31[288], stage0_31[289], stage0_31[290]},
      {stage0_32[136]},
      {stage0_33[96], stage0_33[97], stage0_33[98], stage0_33[99], stage0_33[100], stage0_33[101]},
      {stage1_35[16],stage1_34[36],stage1_33[67],stage1_32[127],stage1_31[170]}
   );
   gpc615_5 gpc1213 (
      {stage0_31[291], stage0_31[292], stage0_31[293], stage0_31[294], stage0_31[295]},
      {stage0_32[137]},
      {stage0_33[102], stage0_33[103], stage0_33[104], stage0_33[105], stage0_33[106], stage0_33[107]},
      {stage1_35[17],stage1_34[37],stage1_33[68],stage1_32[128],stage1_31[171]}
   );
   gpc615_5 gpc1214 (
      {stage0_31[296], stage0_31[297], stage0_31[298], stage0_31[299], stage0_31[300]},
      {stage0_32[138]},
      {stage0_33[108], stage0_33[109], stage0_33[110], stage0_33[111], stage0_33[112], stage0_33[113]},
      {stage1_35[18],stage1_34[38],stage1_33[69],stage1_32[129],stage1_31[172]}
   );
   gpc615_5 gpc1215 (
      {stage0_31[301], stage0_31[302], stage0_31[303], stage0_31[304], stage0_31[305]},
      {stage0_32[139]},
      {stage0_33[114], stage0_33[115], stage0_33[116], stage0_33[117], stage0_33[118], stage0_33[119]},
      {stage1_35[19],stage1_34[39],stage1_33[70],stage1_32[130],stage1_31[173]}
   );
   gpc615_5 gpc1216 (
      {stage0_31[306], stage0_31[307], stage0_31[308], stage0_31[309], stage0_31[310]},
      {stage0_32[140]},
      {stage0_33[120], stage0_33[121], stage0_33[122], stage0_33[123], stage0_33[124], stage0_33[125]},
      {stage1_35[20],stage1_34[40],stage1_33[71],stage1_32[131],stage1_31[174]}
   );
   gpc615_5 gpc1217 (
      {stage0_31[311], stage0_31[312], stage0_31[313], stage0_31[314], stage0_31[315]},
      {stage0_32[141]},
      {stage0_33[126], stage0_33[127], stage0_33[128], stage0_33[129], stage0_33[130], stage0_33[131]},
      {stage1_35[21],stage1_34[41],stage1_33[72],stage1_32[132],stage1_31[175]}
   );
   gpc615_5 gpc1218 (
      {stage0_31[316], stage0_31[317], stage0_31[318], stage0_31[319], stage0_31[320]},
      {stage0_32[142]},
      {stage0_33[132], stage0_33[133], stage0_33[134], stage0_33[135], stage0_33[136], stage0_33[137]},
      {stage1_35[22],stage1_34[42],stage1_33[73],stage1_32[133],stage1_31[176]}
   );
   gpc615_5 gpc1219 (
      {stage0_31[321], stage0_31[322], stage0_31[323], stage0_31[324], stage0_31[325]},
      {stage0_32[143]},
      {stage0_33[138], stage0_33[139], stage0_33[140], stage0_33[141], stage0_33[142], stage0_33[143]},
      {stage1_35[23],stage1_34[43],stage1_33[74],stage1_32[134],stage1_31[177]}
   );
   gpc615_5 gpc1220 (
      {stage0_31[326], stage0_31[327], stage0_31[328], stage0_31[329], stage0_31[330]},
      {stage0_32[144]},
      {stage0_33[144], stage0_33[145], stage0_33[146], stage0_33[147], stage0_33[148], stage0_33[149]},
      {stage1_35[24],stage1_34[44],stage1_33[75],stage1_32[135],stage1_31[178]}
   );
   gpc615_5 gpc1221 (
      {stage0_31[331], stage0_31[332], stage0_31[333], stage0_31[334], stage0_31[335]},
      {stage0_32[145]},
      {stage0_33[150], stage0_33[151], stage0_33[152], stage0_33[153], stage0_33[154], stage0_33[155]},
      {stage1_35[25],stage1_34[45],stage1_33[76],stage1_32[136],stage1_31[179]}
   );
   gpc615_5 gpc1222 (
      {stage0_31[336], stage0_31[337], stage0_31[338], stage0_31[339], stage0_31[340]},
      {stage0_32[146]},
      {stage0_33[156], stage0_33[157], stage0_33[158], stage0_33[159], stage0_33[160], stage0_33[161]},
      {stage1_35[26],stage1_34[46],stage1_33[77],stage1_32[137],stage1_31[180]}
   );
   gpc615_5 gpc1223 (
      {stage0_31[341], stage0_31[342], stage0_31[343], stage0_31[344], stage0_31[345]},
      {stage0_32[147]},
      {stage0_33[162], stage0_33[163], stage0_33[164], stage0_33[165], stage0_33[166], stage0_33[167]},
      {stage1_35[27],stage1_34[47],stage1_33[78],stage1_32[138],stage1_31[181]}
   );
   gpc615_5 gpc1224 (
      {stage0_31[346], stage0_31[347], stage0_31[348], stage0_31[349], stage0_31[350]},
      {stage0_32[148]},
      {stage0_33[168], stage0_33[169], stage0_33[170], stage0_33[171], stage0_33[172], stage0_33[173]},
      {stage1_35[28],stage1_34[48],stage1_33[79],stage1_32[139],stage1_31[182]}
   );
   gpc615_5 gpc1225 (
      {stage0_31[351], stage0_31[352], stage0_31[353], stage0_31[354], stage0_31[355]},
      {stage0_32[149]},
      {stage0_33[174], stage0_33[175], stage0_33[176], stage0_33[177], stage0_33[178], stage0_33[179]},
      {stage1_35[29],stage1_34[49],stage1_33[80],stage1_32[140],stage1_31[183]}
   );
   gpc615_5 gpc1226 (
      {stage0_31[356], stage0_31[357], stage0_31[358], stage0_31[359], stage0_31[360]},
      {stage0_32[150]},
      {stage0_33[180], stage0_33[181], stage0_33[182], stage0_33[183], stage0_33[184], stage0_33[185]},
      {stage1_35[30],stage1_34[50],stage1_33[81],stage1_32[141],stage1_31[184]}
   );
   gpc615_5 gpc1227 (
      {stage0_31[361], stage0_31[362], stage0_31[363], stage0_31[364], stage0_31[365]},
      {stage0_32[151]},
      {stage0_33[186], stage0_33[187], stage0_33[188], stage0_33[189], stage0_33[190], stage0_33[191]},
      {stage1_35[31],stage1_34[51],stage1_33[82],stage1_32[142],stage1_31[185]}
   );
   gpc615_5 gpc1228 (
      {stage0_31[366], stage0_31[367], stage0_31[368], stage0_31[369], stage0_31[370]},
      {stage0_32[152]},
      {stage0_33[192], stage0_33[193], stage0_33[194], stage0_33[195], stage0_33[196], stage0_33[197]},
      {stage1_35[32],stage1_34[52],stage1_33[83],stage1_32[143],stage1_31[186]}
   );
   gpc615_5 gpc1229 (
      {stage0_31[371], stage0_31[372], stage0_31[373], stage0_31[374], stage0_31[375]},
      {stage0_32[153]},
      {stage0_33[198], stage0_33[199], stage0_33[200], stage0_33[201], stage0_33[202], stage0_33[203]},
      {stage1_35[33],stage1_34[53],stage1_33[84],stage1_32[144],stage1_31[187]}
   );
   gpc615_5 gpc1230 (
      {stage0_31[376], stage0_31[377], stage0_31[378], stage0_31[379], stage0_31[380]},
      {stage0_32[154]},
      {stage0_33[204], stage0_33[205], stage0_33[206], stage0_33[207], stage0_33[208], stage0_33[209]},
      {stage1_35[34],stage1_34[54],stage1_33[85],stage1_32[145],stage1_31[188]}
   );
   gpc615_5 gpc1231 (
      {stage0_31[381], stage0_31[382], stage0_31[383], stage0_31[384], stage0_31[385]},
      {stage0_32[155]},
      {stage0_33[210], stage0_33[211], stage0_33[212], stage0_33[213], stage0_33[214], stage0_33[215]},
      {stage1_35[35],stage1_34[55],stage1_33[86],stage1_32[146],stage1_31[189]}
   );
   gpc615_5 gpc1232 (
      {stage0_31[386], stage0_31[387], stage0_31[388], stage0_31[389], stage0_31[390]},
      {stage0_32[156]},
      {stage0_33[216], stage0_33[217], stage0_33[218], stage0_33[219], stage0_33[220], stage0_33[221]},
      {stage1_35[36],stage1_34[56],stage1_33[87],stage1_32[147],stage1_31[190]}
   );
   gpc615_5 gpc1233 (
      {stage0_31[391], stage0_31[392], stage0_31[393], stage0_31[394], stage0_31[395]},
      {stage0_32[157]},
      {stage0_33[222], stage0_33[223], stage0_33[224], stage0_33[225], stage0_33[226], stage0_33[227]},
      {stage1_35[37],stage1_34[57],stage1_33[88],stage1_32[148],stage1_31[191]}
   );
   gpc615_5 gpc1234 (
      {stage0_31[396], stage0_31[397], stage0_31[398], stage0_31[399], stage0_31[400]},
      {stage0_32[158]},
      {stage0_33[228], stage0_33[229], stage0_33[230], stage0_33[231], stage0_33[232], stage0_33[233]},
      {stage1_35[38],stage1_34[58],stage1_33[89],stage1_32[149],stage1_31[192]}
   );
   gpc615_5 gpc1235 (
      {stage0_31[401], stage0_31[402], stage0_31[403], stage0_31[404], stage0_31[405]},
      {stage0_32[159]},
      {stage0_33[234], stage0_33[235], stage0_33[236], stage0_33[237], stage0_33[238], stage0_33[239]},
      {stage1_35[39],stage1_34[59],stage1_33[90],stage1_32[150],stage1_31[193]}
   );
   gpc615_5 gpc1236 (
      {stage0_31[406], stage0_31[407], stage0_31[408], stage0_31[409], stage0_31[410]},
      {stage0_32[160]},
      {stage0_33[240], stage0_33[241], stage0_33[242], stage0_33[243], stage0_33[244], stage0_33[245]},
      {stage1_35[40],stage1_34[60],stage1_33[91],stage1_32[151],stage1_31[194]}
   );
   gpc615_5 gpc1237 (
      {stage0_31[411], stage0_31[412], stage0_31[413], stage0_31[414], stage0_31[415]},
      {stage0_32[161]},
      {stage0_33[246], stage0_33[247], stage0_33[248], stage0_33[249], stage0_33[250], stage0_33[251]},
      {stage1_35[41],stage1_34[61],stage1_33[92],stage1_32[152],stage1_31[195]}
   );
   gpc615_5 gpc1238 (
      {stage0_31[416], stage0_31[417], stage0_31[418], stage0_31[419], stage0_31[420]},
      {stage0_32[162]},
      {stage0_33[252], stage0_33[253], stage0_33[254], stage0_33[255], stage0_33[256], stage0_33[257]},
      {stage1_35[42],stage1_34[62],stage1_33[93],stage1_32[153],stage1_31[196]}
   );
   gpc615_5 gpc1239 (
      {stage0_31[421], stage0_31[422], stage0_31[423], stage0_31[424], stage0_31[425]},
      {stage0_32[163]},
      {stage0_33[258], stage0_33[259], stage0_33[260], stage0_33[261], stage0_33[262], stage0_33[263]},
      {stage1_35[43],stage1_34[63],stage1_33[94],stage1_32[154],stage1_31[197]}
   );
   gpc615_5 gpc1240 (
      {stage0_31[426], stage0_31[427], stage0_31[428], stage0_31[429], stage0_31[430]},
      {stage0_32[164]},
      {stage0_33[264], stage0_33[265], stage0_33[266], stage0_33[267], stage0_33[268], stage0_33[269]},
      {stage1_35[44],stage1_34[64],stage1_33[95],stage1_32[155],stage1_31[198]}
   );
   gpc615_5 gpc1241 (
      {stage0_31[431], stage0_31[432], stage0_31[433], stage0_31[434], stage0_31[435]},
      {stage0_32[165]},
      {stage0_33[270], stage0_33[271], stage0_33[272], stage0_33[273], stage0_33[274], stage0_33[275]},
      {stage1_35[45],stage1_34[65],stage1_33[96],stage1_32[156],stage1_31[199]}
   );
   gpc615_5 gpc1242 (
      {stage0_31[436], stage0_31[437], stage0_31[438], stage0_31[439], stage0_31[440]},
      {stage0_32[166]},
      {stage0_33[276], stage0_33[277], stage0_33[278], stage0_33[279], stage0_33[280], stage0_33[281]},
      {stage1_35[46],stage1_34[66],stage1_33[97],stage1_32[157],stage1_31[200]}
   );
   gpc615_5 gpc1243 (
      {stage0_31[441], stage0_31[442], stage0_31[443], stage0_31[444], stage0_31[445]},
      {stage0_32[167]},
      {stage0_33[282], stage0_33[283], stage0_33[284], stage0_33[285], stage0_33[286], stage0_33[287]},
      {stage1_35[47],stage1_34[67],stage1_33[98],stage1_32[158],stage1_31[201]}
   );
   gpc615_5 gpc1244 (
      {stage0_31[446], stage0_31[447], stage0_31[448], stage0_31[449], stage0_31[450]},
      {stage0_32[168]},
      {stage0_33[288], stage0_33[289], stage0_33[290], stage0_33[291], stage0_33[292], stage0_33[293]},
      {stage1_35[48],stage1_34[68],stage1_33[99],stage1_32[159],stage1_31[202]}
   );
   gpc615_5 gpc1245 (
      {stage0_31[451], stage0_31[452], stage0_31[453], stage0_31[454], stage0_31[455]},
      {stage0_32[169]},
      {stage0_33[294], stage0_33[295], stage0_33[296], stage0_33[297], stage0_33[298], stage0_33[299]},
      {stage1_35[49],stage1_34[69],stage1_33[100],stage1_32[160],stage1_31[203]}
   );
   gpc615_5 gpc1246 (
      {stage0_31[456], stage0_31[457], stage0_31[458], stage0_31[459], stage0_31[460]},
      {stage0_32[170]},
      {stage0_33[300], stage0_33[301], stage0_33[302], stage0_33[303], stage0_33[304], stage0_33[305]},
      {stage1_35[50],stage1_34[70],stage1_33[101],stage1_32[161],stage1_31[204]}
   );
   gpc615_5 gpc1247 (
      {stage0_31[461], stage0_31[462], stage0_31[463], stage0_31[464], stage0_31[465]},
      {stage0_32[171]},
      {stage0_33[306], stage0_33[307], stage0_33[308], stage0_33[309], stage0_33[310], stage0_33[311]},
      {stage1_35[51],stage1_34[71],stage1_33[102],stage1_32[162],stage1_31[205]}
   );
   gpc615_5 gpc1248 (
      {stage0_31[466], stage0_31[467], stage0_31[468], stage0_31[469], stage0_31[470]},
      {stage0_32[172]},
      {stage0_33[312], stage0_33[313], stage0_33[314], stage0_33[315], stage0_33[316], stage0_33[317]},
      {stage1_35[52],stage1_34[72],stage1_33[103],stage1_32[163],stage1_31[206]}
   );
   gpc615_5 gpc1249 (
      {stage0_31[471], stage0_31[472], stage0_31[473], stage0_31[474], stage0_31[475]},
      {stage0_32[173]},
      {stage0_33[318], stage0_33[319], stage0_33[320], stage0_33[321], stage0_33[322], stage0_33[323]},
      {stage1_35[53],stage1_34[73],stage1_33[104],stage1_32[164],stage1_31[207]}
   );
   gpc606_5 gpc1250 (
      {stage0_32[174], stage0_32[175], stage0_32[176], stage0_32[177], stage0_32[178], stage0_32[179]},
      {stage0_34[0], stage0_34[1], stage0_34[2], stage0_34[3], stage0_34[4], stage0_34[5]},
      {stage1_36[0],stage1_35[54],stage1_34[74],stage1_33[105],stage1_32[165]}
   );
   gpc606_5 gpc1251 (
      {stage0_32[180], stage0_32[181], stage0_32[182], stage0_32[183], stage0_32[184], stage0_32[185]},
      {stage0_34[6], stage0_34[7], stage0_34[8], stage0_34[9], stage0_34[10], stage0_34[11]},
      {stage1_36[1],stage1_35[55],stage1_34[75],stage1_33[106],stage1_32[166]}
   );
   gpc606_5 gpc1252 (
      {stage0_32[186], stage0_32[187], stage0_32[188], stage0_32[189], stage0_32[190], stage0_32[191]},
      {stage0_34[12], stage0_34[13], stage0_34[14], stage0_34[15], stage0_34[16], stage0_34[17]},
      {stage1_36[2],stage1_35[56],stage1_34[76],stage1_33[107],stage1_32[167]}
   );
   gpc606_5 gpc1253 (
      {stage0_32[192], stage0_32[193], stage0_32[194], stage0_32[195], stage0_32[196], stage0_32[197]},
      {stage0_34[18], stage0_34[19], stage0_34[20], stage0_34[21], stage0_34[22], stage0_34[23]},
      {stage1_36[3],stage1_35[57],stage1_34[77],stage1_33[108],stage1_32[168]}
   );
   gpc606_5 gpc1254 (
      {stage0_32[198], stage0_32[199], stage0_32[200], stage0_32[201], stage0_32[202], stage0_32[203]},
      {stage0_34[24], stage0_34[25], stage0_34[26], stage0_34[27], stage0_34[28], stage0_34[29]},
      {stage1_36[4],stage1_35[58],stage1_34[78],stage1_33[109],stage1_32[169]}
   );
   gpc606_5 gpc1255 (
      {stage0_32[204], stage0_32[205], stage0_32[206], stage0_32[207], stage0_32[208], stage0_32[209]},
      {stage0_34[30], stage0_34[31], stage0_34[32], stage0_34[33], stage0_34[34], stage0_34[35]},
      {stage1_36[5],stage1_35[59],stage1_34[79],stage1_33[110],stage1_32[170]}
   );
   gpc606_5 gpc1256 (
      {stage0_32[210], stage0_32[211], stage0_32[212], stage0_32[213], stage0_32[214], stage0_32[215]},
      {stage0_34[36], stage0_34[37], stage0_34[38], stage0_34[39], stage0_34[40], stage0_34[41]},
      {stage1_36[6],stage1_35[60],stage1_34[80],stage1_33[111],stage1_32[171]}
   );
   gpc606_5 gpc1257 (
      {stage0_32[216], stage0_32[217], stage0_32[218], stage0_32[219], stage0_32[220], stage0_32[221]},
      {stage0_34[42], stage0_34[43], stage0_34[44], stage0_34[45], stage0_34[46], stage0_34[47]},
      {stage1_36[7],stage1_35[61],stage1_34[81],stage1_33[112],stage1_32[172]}
   );
   gpc606_5 gpc1258 (
      {stage0_32[222], stage0_32[223], stage0_32[224], stage0_32[225], stage0_32[226], stage0_32[227]},
      {stage0_34[48], stage0_34[49], stage0_34[50], stage0_34[51], stage0_34[52], stage0_34[53]},
      {stage1_36[8],stage1_35[62],stage1_34[82],stage1_33[113],stage1_32[173]}
   );
   gpc606_5 gpc1259 (
      {stage0_32[228], stage0_32[229], stage0_32[230], stage0_32[231], stage0_32[232], stage0_32[233]},
      {stage0_34[54], stage0_34[55], stage0_34[56], stage0_34[57], stage0_34[58], stage0_34[59]},
      {stage1_36[9],stage1_35[63],stage1_34[83],stage1_33[114],stage1_32[174]}
   );
   gpc606_5 gpc1260 (
      {stage0_32[234], stage0_32[235], stage0_32[236], stage0_32[237], stage0_32[238], stage0_32[239]},
      {stage0_34[60], stage0_34[61], stage0_34[62], stage0_34[63], stage0_34[64], stage0_34[65]},
      {stage1_36[10],stage1_35[64],stage1_34[84],stage1_33[115],stage1_32[175]}
   );
   gpc606_5 gpc1261 (
      {stage0_32[240], stage0_32[241], stage0_32[242], stage0_32[243], stage0_32[244], stage0_32[245]},
      {stage0_34[66], stage0_34[67], stage0_34[68], stage0_34[69], stage0_34[70], stage0_34[71]},
      {stage1_36[11],stage1_35[65],stage1_34[85],stage1_33[116],stage1_32[176]}
   );
   gpc606_5 gpc1262 (
      {stage0_32[246], stage0_32[247], stage0_32[248], stage0_32[249], stage0_32[250], stage0_32[251]},
      {stage0_34[72], stage0_34[73], stage0_34[74], stage0_34[75], stage0_34[76], stage0_34[77]},
      {stage1_36[12],stage1_35[66],stage1_34[86],stage1_33[117],stage1_32[177]}
   );
   gpc606_5 gpc1263 (
      {stage0_32[252], stage0_32[253], stage0_32[254], stage0_32[255], stage0_32[256], stage0_32[257]},
      {stage0_34[78], stage0_34[79], stage0_34[80], stage0_34[81], stage0_34[82], stage0_34[83]},
      {stage1_36[13],stage1_35[67],stage1_34[87],stage1_33[118],stage1_32[178]}
   );
   gpc606_5 gpc1264 (
      {stage0_32[258], stage0_32[259], stage0_32[260], stage0_32[261], stage0_32[262], stage0_32[263]},
      {stage0_34[84], stage0_34[85], stage0_34[86], stage0_34[87], stage0_34[88], stage0_34[89]},
      {stage1_36[14],stage1_35[68],stage1_34[88],stage1_33[119],stage1_32[179]}
   );
   gpc606_5 gpc1265 (
      {stage0_32[264], stage0_32[265], stage0_32[266], stage0_32[267], stage0_32[268], stage0_32[269]},
      {stage0_34[90], stage0_34[91], stage0_34[92], stage0_34[93], stage0_34[94], stage0_34[95]},
      {stage1_36[15],stage1_35[69],stage1_34[89],stage1_33[120],stage1_32[180]}
   );
   gpc606_5 gpc1266 (
      {stage0_32[270], stage0_32[271], stage0_32[272], stage0_32[273], stage0_32[274], stage0_32[275]},
      {stage0_34[96], stage0_34[97], stage0_34[98], stage0_34[99], stage0_34[100], stage0_34[101]},
      {stage1_36[16],stage1_35[70],stage1_34[90],stage1_33[121],stage1_32[181]}
   );
   gpc606_5 gpc1267 (
      {stage0_32[276], stage0_32[277], stage0_32[278], stage0_32[279], stage0_32[280], stage0_32[281]},
      {stage0_34[102], stage0_34[103], stage0_34[104], stage0_34[105], stage0_34[106], stage0_34[107]},
      {stage1_36[17],stage1_35[71],stage1_34[91],stage1_33[122],stage1_32[182]}
   );
   gpc606_5 gpc1268 (
      {stage0_32[282], stage0_32[283], stage0_32[284], stage0_32[285], stage0_32[286], stage0_32[287]},
      {stage0_34[108], stage0_34[109], stage0_34[110], stage0_34[111], stage0_34[112], stage0_34[113]},
      {stage1_36[18],stage1_35[72],stage1_34[92],stage1_33[123],stage1_32[183]}
   );
   gpc606_5 gpc1269 (
      {stage0_32[288], stage0_32[289], stage0_32[290], stage0_32[291], stage0_32[292], stage0_32[293]},
      {stage0_34[114], stage0_34[115], stage0_34[116], stage0_34[117], stage0_34[118], stage0_34[119]},
      {stage1_36[19],stage1_35[73],stage1_34[93],stage1_33[124],stage1_32[184]}
   );
   gpc606_5 gpc1270 (
      {stage0_32[294], stage0_32[295], stage0_32[296], stage0_32[297], stage0_32[298], stage0_32[299]},
      {stage0_34[120], stage0_34[121], stage0_34[122], stage0_34[123], stage0_34[124], stage0_34[125]},
      {stage1_36[20],stage1_35[74],stage1_34[94],stage1_33[125],stage1_32[185]}
   );
   gpc606_5 gpc1271 (
      {stage0_32[300], stage0_32[301], stage0_32[302], stage0_32[303], stage0_32[304], stage0_32[305]},
      {stage0_34[126], stage0_34[127], stage0_34[128], stage0_34[129], stage0_34[130], stage0_34[131]},
      {stage1_36[21],stage1_35[75],stage1_34[95],stage1_33[126],stage1_32[186]}
   );
   gpc606_5 gpc1272 (
      {stage0_32[306], stage0_32[307], stage0_32[308], stage0_32[309], stage0_32[310], stage0_32[311]},
      {stage0_34[132], stage0_34[133], stage0_34[134], stage0_34[135], stage0_34[136], stage0_34[137]},
      {stage1_36[22],stage1_35[76],stage1_34[96],stage1_33[127],stage1_32[187]}
   );
   gpc606_5 gpc1273 (
      {stage0_32[312], stage0_32[313], stage0_32[314], stage0_32[315], stage0_32[316], stage0_32[317]},
      {stage0_34[138], stage0_34[139], stage0_34[140], stage0_34[141], stage0_34[142], stage0_34[143]},
      {stage1_36[23],stage1_35[77],stage1_34[97],stage1_33[128],stage1_32[188]}
   );
   gpc606_5 gpc1274 (
      {stage0_32[318], stage0_32[319], stage0_32[320], stage0_32[321], stage0_32[322], stage0_32[323]},
      {stage0_34[144], stage0_34[145], stage0_34[146], stage0_34[147], stage0_34[148], stage0_34[149]},
      {stage1_36[24],stage1_35[78],stage1_34[98],stage1_33[129],stage1_32[189]}
   );
   gpc606_5 gpc1275 (
      {stage0_32[324], stage0_32[325], stage0_32[326], stage0_32[327], stage0_32[328], stage0_32[329]},
      {stage0_34[150], stage0_34[151], stage0_34[152], stage0_34[153], stage0_34[154], stage0_34[155]},
      {stage1_36[25],stage1_35[79],stage1_34[99],stage1_33[130],stage1_32[190]}
   );
   gpc606_5 gpc1276 (
      {stage0_32[330], stage0_32[331], stage0_32[332], stage0_32[333], stage0_32[334], stage0_32[335]},
      {stage0_34[156], stage0_34[157], stage0_34[158], stage0_34[159], stage0_34[160], stage0_34[161]},
      {stage1_36[26],stage1_35[80],stage1_34[100],stage1_33[131],stage1_32[191]}
   );
   gpc606_5 gpc1277 (
      {stage0_32[336], stage0_32[337], stage0_32[338], stage0_32[339], stage0_32[340], stage0_32[341]},
      {stage0_34[162], stage0_34[163], stage0_34[164], stage0_34[165], stage0_34[166], stage0_34[167]},
      {stage1_36[27],stage1_35[81],stage1_34[101],stage1_33[132],stage1_32[192]}
   );
   gpc606_5 gpc1278 (
      {stage0_32[342], stage0_32[343], stage0_32[344], stage0_32[345], stage0_32[346], stage0_32[347]},
      {stage0_34[168], stage0_34[169], stage0_34[170], stage0_34[171], stage0_34[172], stage0_34[173]},
      {stage1_36[28],stage1_35[82],stage1_34[102],stage1_33[133],stage1_32[193]}
   );
   gpc606_5 gpc1279 (
      {stage0_32[348], stage0_32[349], stage0_32[350], stage0_32[351], stage0_32[352], stage0_32[353]},
      {stage0_34[174], stage0_34[175], stage0_34[176], stage0_34[177], stage0_34[178], stage0_34[179]},
      {stage1_36[29],stage1_35[83],stage1_34[103],stage1_33[134],stage1_32[194]}
   );
   gpc606_5 gpc1280 (
      {stage0_32[354], stage0_32[355], stage0_32[356], stage0_32[357], stage0_32[358], stage0_32[359]},
      {stage0_34[180], stage0_34[181], stage0_34[182], stage0_34[183], stage0_34[184], stage0_34[185]},
      {stage1_36[30],stage1_35[84],stage1_34[104],stage1_33[135],stage1_32[195]}
   );
   gpc606_5 gpc1281 (
      {stage0_32[360], stage0_32[361], stage0_32[362], stage0_32[363], stage0_32[364], stage0_32[365]},
      {stage0_34[186], stage0_34[187], stage0_34[188], stage0_34[189], stage0_34[190], stage0_34[191]},
      {stage1_36[31],stage1_35[85],stage1_34[105],stage1_33[136],stage1_32[196]}
   );
   gpc606_5 gpc1282 (
      {stage0_32[366], stage0_32[367], stage0_32[368], stage0_32[369], stage0_32[370], stage0_32[371]},
      {stage0_34[192], stage0_34[193], stage0_34[194], stage0_34[195], stage0_34[196], stage0_34[197]},
      {stage1_36[32],stage1_35[86],stage1_34[106],stage1_33[137],stage1_32[197]}
   );
   gpc606_5 gpc1283 (
      {stage0_32[372], stage0_32[373], stage0_32[374], stage0_32[375], stage0_32[376], stage0_32[377]},
      {stage0_34[198], stage0_34[199], stage0_34[200], stage0_34[201], stage0_34[202], stage0_34[203]},
      {stage1_36[33],stage1_35[87],stage1_34[107],stage1_33[138],stage1_32[198]}
   );
   gpc606_5 gpc1284 (
      {stage0_32[378], stage0_32[379], stage0_32[380], stage0_32[381], stage0_32[382], stage0_32[383]},
      {stage0_34[204], stage0_34[205], stage0_34[206], stage0_34[207], stage0_34[208], stage0_34[209]},
      {stage1_36[34],stage1_35[88],stage1_34[108],stage1_33[139],stage1_32[199]}
   );
   gpc606_5 gpc1285 (
      {stage0_32[384], stage0_32[385], stage0_32[386], stage0_32[387], stage0_32[388], stage0_32[389]},
      {stage0_34[210], stage0_34[211], stage0_34[212], stage0_34[213], stage0_34[214], stage0_34[215]},
      {stage1_36[35],stage1_35[89],stage1_34[109],stage1_33[140],stage1_32[200]}
   );
   gpc606_5 gpc1286 (
      {stage0_32[390], stage0_32[391], stage0_32[392], stage0_32[393], stage0_32[394], stage0_32[395]},
      {stage0_34[216], stage0_34[217], stage0_34[218], stage0_34[219], stage0_34[220], stage0_34[221]},
      {stage1_36[36],stage1_35[90],stage1_34[110],stage1_33[141],stage1_32[201]}
   );
   gpc606_5 gpc1287 (
      {stage0_32[396], stage0_32[397], stage0_32[398], stage0_32[399], stage0_32[400], stage0_32[401]},
      {stage0_34[222], stage0_34[223], stage0_34[224], stage0_34[225], stage0_34[226], stage0_34[227]},
      {stage1_36[37],stage1_35[91],stage1_34[111],stage1_33[142],stage1_32[202]}
   );
   gpc606_5 gpc1288 (
      {stage0_32[402], stage0_32[403], stage0_32[404], stage0_32[405], stage0_32[406], stage0_32[407]},
      {stage0_34[228], stage0_34[229], stage0_34[230], stage0_34[231], stage0_34[232], stage0_34[233]},
      {stage1_36[38],stage1_35[92],stage1_34[112],stage1_33[143],stage1_32[203]}
   );
   gpc606_5 gpc1289 (
      {stage0_32[408], stage0_32[409], stage0_32[410], stage0_32[411], stage0_32[412], stage0_32[413]},
      {stage0_34[234], stage0_34[235], stage0_34[236], stage0_34[237], stage0_34[238], stage0_34[239]},
      {stage1_36[39],stage1_35[93],stage1_34[113],stage1_33[144],stage1_32[204]}
   );
   gpc606_5 gpc1290 (
      {stage0_32[414], stage0_32[415], stage0_32[416], stage0_32[417], stage0_32[418], stage0_32[419]},
      {stage0_34[240], stage0_34[241], stage0_34[242], stage0_34[243], stage0_34[244], stage0_34[245]},
      {stage1_36[40],stage1_35[94],stage1_34[114],stage1_33[145],stage1_32[205]}
   );
   gpc606_5 gpc1291 (
      {stage0_32[420], stage0_32[421], stage0_32[422], stage0_32[423], stage0_32[424], stage0_32[425]},
      {stage0_34[246], stage0_34[247], stage0_34[248], stage0_34[249], stage0_34[250], stage0_34[251]},
      {stage1_36[41],stage1_35[95],stage1_34[115],stage1_33[146],stage1_32[206]}
   );
   gpc606_5 gpc1292 (
      {stage0_32[426], stage0_32[427], stage0_32[428], stage0_32[429], stage0_32[430], stage0_32[431]},
      {stage0_34[252], stage0_34[253], stage0_34[254], stage0_34[255], stage0_34[256], stage0_34[257]},
      {stage1_36[42],stage1_35[96],stage1_34[116],stage1_33[147],stage1_32[207]}
   );
   gpc606_5 gpc1293 (
      {stage0_32[432], stage0_32[433], stage0_32[434], stage0_32[435], stage0_32[436], stage0_32[437]},
      {stage0_34[258], stage0_34[259], stage0_34[260], stage0_34[261], stage0_34[262], stage0_34[263]},
      {stage1_36[43],stage1_35[97],stage1_34[117],stage1_33[148],stage1_32[208]}
   );
   gpc606_5 gpc1294 (
      {stage0_32[438], stage0_32[439], stage0_32[440], stage0_32[441], stage0_32[442], stage0_32[443]},
      {stage0_34[264], stage0_34[265], stage0_34[266], stage0_34[267], stage0_34[268], stage0_34[269]},
      {stage1_36[44],stage1_35[98],stage1_34[118],stage1_33[149],stage1_32[209]}
   );
   gpc606_5 gpc1295 (
      {stage0_32[444], stage0_32[445], stage0_32[446], stage0_32[447], stage0_32[448], stage0_32[449]},
      {stage0_34[270], stage0_34[271], stage0_34[272], stage0_34[273], stage0_34[274], stage0_34[275]},
      {stage1_36[45],stage1_35[99],stage1_34[119],stage1_33[150],stage1_32[210]}
   );
   gpc606_5 gpc1296 (
      {stage0_32[450], stage0_32[451], stage0_32[452], stage0_32[453], stage0_32[454], stage0_32[455]},
      {stage0_34[276], stage0_34[277], stage0_34[278], stage0_34[279], stage0_34[280], stage0_34[281]},
      {stage1_36[46],stage1_35[100],stage1_34[120],stage1_33[151],stage1_32[211]}
   );
   gpc606_5 gpc1297 (
      {stage0_32[456], stage0_32[457], stage0_32[458], stage0_32[459], stage0_32[460], stage0_32[461]},
      {stage0_34[282], stage0_34[283], stage0_34[284], stage0_34[285], stage0_34[286], stage0_34[287]},
      {stage1_36[47],stage1_35[101],stage1_34[121],stage1_33[152],stage1_32[212]}
   );
   gpc606_5 gpc1298 (
      {stage0_32[462], stage0_32[463], stage0_32[464], stage0_32[465], stage0_32[466], stage0_32[467]},
      {stage0_34[288], stage0_34[289], stage0_34[290], stage0_34[291], stage0_34[292], stage0_34[293]},
      {stage1_36[48],stage1_35[102],stage1_34[122],stage1_33[153],stage1_32[213]}
   );
   gpc606_5 gpc1299 (
      {stage0_32[468], stage0_32[469], stage0_32[470], stage0_32[471], stage0_32[472], stage0_32[473]},
      {stage0_34[294], stage0_34[295], stage0_34[296], stage0_34[297], stage0_34[298], stage0_34[299]},
      {stage1_36[49],stage1_35[103],stage1_34[123],stage1_33[154],stage1_32[214]}
   );
   gpc606_5 gpc1300 (
      {stage0_32[474], stage0_32[475], stage0_32[476], stage0_32[477], stage0_32[478], stage0_32[479]},
      {stage0_34[300], stage0_34[301], stage0_34[302], stage0_34[303], stage0_34[304], stage0_34[305]},
      {stage1_36[50],stage1_35[104],stage1_34[124],stage1_33[155],stage1_32[215]}
   );
   gpc606_5 gpc1301 (
      {stage0_32[480], stage0_32[481], stage0_32[482], stage0_32[483], stage0_32[484], stage0_32[485]},
      {stage0_34[306], stage0_34[307], stage0_34[308], stage0_34[309], stage0_34[310], stage0_34[311]},
      {stage1_36[51],stage1_35[105],stage1_34[125],stage1_33[156],stage1_32[216]}
   );
   gpc606_5 gpc1302 (
      {stage0_33[324], stage0_33[325], stage0_33[326], stage0_33[327], stage0_33[328], stage0_33[329]},
      {stage0_35[0], stage0_35[1], stage0_35[2], stage0_35[3], stage0_35[4], stage0_35[5]},
      {stage1_37[0],stage1_36[52],stage1_35[106],stage1_34[126],stage1_33[157]}
   );
   gpc606_5 gpc1303 (
      {stage0_33[330], stage0_33[331], stage0_33[332], stage0_33[333], stage0_33[334], stage0_33[335]},
      {stage0_35[6], stage0_35[7], stage0_35[8], stage0_35[9], stage0_35[10], stage0_35[11]},
      {stage1_37[1],stage1_36[53],stage1_35[107],stage1_34[127],stage1_33[158]}
   );
   gpc606_5 gpc1304 (
      {stage0_33[336], stage0_33[337], stage0_33[338], stage0_33[339], stage0_33[340], stage0_33[341]},
      {stage0_35[12], stage0_35[13], stage0_35[14], stage0_35[15], stage0_35[16], stage0_35[17]},
      {stage1_37[2],stage1_36[54],stage1_35[108],stage1_34[128],stage1_33[159]}
   );
   gpc606_5 gpc1305 (
      {stage0_33[342], stage0_33[343], stage0_33[344], stage0_33[345], stage0_33[346], stage0_33[347]},
      {stage0_35[18], stage0_35[19], stage0_35[20], stage0_35[21], stage0_35[22], stage0_35[23]},
      {stage1_37[3],stage1_36[55],stage1_35[109],stage1_34[129],stage1_33[160]}
   );
   gpc606_5 gpc1306 (
      {stage0_33[348], stage0_33[349], stage0_33[350], stage0_33[351], stage0_33[352], stage0_33[353]},
      {stage0_35[24], stage0_35[25], stage0_35[26], stage0_35[27], stage0_35[28], stage0_35[29]},
      {stage1_37[4],stage1_36[56],stage1_35[110],stage1_34[130],stage1_33[161]}
   );
   gpc606_5 gpc1307 (
      {stage0_33[354], stage0_33[355], stage0_33[356], stage0_33[357], stage0_33[358], stage0_33[359]},
      {stage0_35[30], stage0_35[31], stage0_35[32], stage0_35[33], stage0_35[34], stage0_35[35]},
      {stage1_37[5],stage1_36[57],stage1_35[111],stage1_34[131],stage1_33[162]}
   );
   gpc606_5 gpc1308 (
      {stage0_33[360], stage0_33[361], stage0_33[362], stage0_33[363], stage0_33[364], stage0_33[365]},
      {stage0_35[36], stage0_35[37], stage0_35[38], stage0_35[39], stage0_35[40], stage0_35[41]},
      {stage1_37[6],stage1_36[58],stage1_35[112],stage1_34[132],stage1_33[163]}
   );
   gpc606_5 gpc1309 (
      {stage0_33[366], stage0_33[367], stage0_33[368], stage0_33[369], stage0_33[370], stage0_33[371]},
      {stage0_35[42], stage0_35[43], stage0_35[44], stage0_35[45], stage0_35[46], stage0_35[47]},
      {stage1_37[7],stage1_36[59],stage1_35[113],stage1_34[133],stage1_33[164]}
   );
   gpc606_5 gpc1310 (
      {stage0_33[372], stage0_33[373], stage0_33[374], stage0_33[375], stage0_33[376], stage0_33[377]},
      {stage0_35[48], stage0_35[49], stage0_35[50], stage0_35[51], stage0_35[52], stage0_35[53]},
      {stage1_37[8],stage1_36[60],stage1_35[114],stage1_34[134],stage1_33[165]}
   );
   gpc606_5 gpc1311 (
      {stage0_33[378], stage0_33[379], stage0_33[380], stage0_33[381], stage0_33[382], stage0_33[383]},
      {stage0_35[54], stage0_35[55], stage0_35[56], stage0_35[57], stage0_35[58], stage0_35[59]},
      {stage1_37[9],stage1_36[61],stage1_35[115],stage1_34[135],stage1_33[166]}
   );
   gpc606_5 gpc1312 (
      {stage0_33[384], stage0_33[385], stage0_33[386], stage0_33[387], stage0_33[388], stage0_33[389]},
      {stage0_35[60], stage0_35[61], stage0_35[62], stage0_35[63], stage0_35[64], stage0_35[65]},
      {stage1_37[10],stage1_36[62],stage1_35[116],stage1_34[136],stage1_33[167]}
   );
   gpc606_5 gpc1313 (
      {stage0_33[390], stage0_33[391], stage0_33[392], stage0_33[393], stage0_33[394], stage0_33[395]},
      {stage0_35[66], stage0_35[67], stage0_35[68], stage0_35[69], stage0_35[70], stage0_35[71]},
      {stage1_37[11],stage1_36[63],stage1_35[117],stage1_34[137],stage1_33[168]}
   );
   gpc1163_5 gpc1314 (
      {stage0_34[312], stage0_34[313], stage0_34[314]},
      {stage0_35[72], stage0_35[73], stage0_35[74], stage0_35[75], stage0_35[76], stage0_35[77]},
      {stage0_36[0]},
      {stage0_37[0]},
      {stage1_38[0],stage1_37[12],stage1_36[64],stage1_35[118],stage1_34[138]}
   );
   gpc1163_5 gpc1315 (
      {stage0_34[315], stage0_34[316], stage0_34[317]},
      {stage0_35[78], stage0_35[79], stage0_35[80], stage0_35[81], stage0_35[82], stage0_35[83]},
      {stage0_36[1]},
      {stage0_37[1]},
      {stage1_38[1],stage1_37[13],stage1_36[65],stage1_35[119],stage1_34[139]}
   );
   gpc1163_5 gpc1316 (
      {stage0_34[318], stage0_34[319], stage0_34[320]},
      {stage0_35[84], stage0_35[85], stage0_35[86], stage0_35[87], stage0_35[88], stage0_35[89]},
      {stage0_36[2]},
      {stage0_37[2]},
      {stage1_38[2],stage1_37[14],stage1_36[66],stage1_35[120],stage1_34[140]}
   );
   gpc1163_5 gpc1317 (
      {stage0_34[321], stage0_34[322], stage0_34[323]},
      {stage0_35[90], stage0_35[91], stage0_35[92], stage0_35[93], stage0_35[94], stage0_35[95]},
      {stage0_36[3]},
      {stage0_37[3]},
      {stage1_38[3],stage1_37[15],stage1_36[67],stage1_35[121],stage1_34[141]}
   );
   gpc1163_5 gpc1318 (
      {stage0_34[324], stage0_34[325], stage0_34[326]},
      {stage0_35[96], stage0_35[97], stage0_35[98], stage0_35[99], stage0_35[100], stage0_35[101]},
      {stage0_36[4]},
      {stage0_37[4]},
      {stage1_38[4],stage1_37[16],stage1_36[68],stage1_35[122],stage1_34[142]}
   );
   gpc1163_5 gpc1319 (
      {stage0_34[327], stage0_34[328], stage0_34[329]},
      {stage0_35[102], stage0_35[103], stage0_35[104], stage0_35[105], stage0_35[106], stage0_35[107]},
      {stage0_36[5]},
      {stage0_37[5]},
      {stage1_38[5],stage1_37[17],stage1_36[69],stage1_35[123],stage1_34[143]}
   );
   gpc1163_5 gpc1320 (
      {stage0_34[330], stage0_34[331], stage0_34[332]},
      {stage0_35[108], stage0_35[109], stage0_35[110], stage0_35[111], stage0_35[112], stage0_35[113]},
      {stage0_36[6]},
      {stage0_37[6]},
      {stage1_38[6],stage1_37[18],stage1_36[70],stage1_35[124],stage1_34[144]}
   );
   gpc1163_5 gpc1321 (
      {stage0_34[333], stage0_34[334], stage0_34[335]},
      {stage0_35[114], stage0_35[115], stage0_35[116], stage0_35[117], stage0_35[118], stage0_35[119]},
      {stage0_36[7]},
      {stage0_37[7]},
      {stage1_38[7],stage1_37[19],stage1_36[71],stage1_35[125],stage1_34[145]}
   );
   gpc1163_5 gpc1322 (
      {stage0_34[336], stage0_34[337], stage0_34[338]},
      {stage0_35[120], stage0_35[121], stage0_35[122], stage0_35[123], stage0_35[124], stage0_35[125]},
      {stage0_36[8]},
      {stage0_37[8]},
      {stage1_38[8],stage1_37[20],stage1_36[72],stage1_35[126],stage1_34[146]}
   );
   gpc1163_5 gpc1323 (
      {stage0_34[339], stage0_34[340], stage0_34[341]},
      {stage0_35[126], stage0_35[127], stage0_35[128], stage0_35[129], stage0_35[130], stage0_35[131]},
      {stage0_36[9]},
      {stage0_37[9]},
      {stage1_38[9],stage1_37[21],stage1_36[73],stage1_35[127],stage1_34[147]}
   );
   gpc1163_5 gpc1324 (
      {stage0_34[342], stage0_34[343], stage0_34[344]},
      {stage0_35[132], stage0_35[133], stage0_35[134], stage0_35[135], stage0_35[136], stage0_35[137]},
      {stage0_36[10]},
      {stage0_37[10]},
      {stage1_38[10],stage1_37[22],stage1_36[74],stage1_35[128],stage1_34[148]}
   );
   gpc1163_5 gpc1325 (
      {stage0_34[345], stage0_34[346], stage0_34[347]},
      {stage0_35[138], stage0_35[139], stage0_35[140], stage0_35[141], stage0_35[142], stage0_35[143]},
      {stage0_36[11]},
      {stage0_37[11]},
      {stage1_38[11],stage1_37[23],stage1_36[75],stage1_35[129],stage1_34[149]}
   );
   gpc1163_5 gpc1326 (
      {stage0_34[348], stage0_34[349], stage0_34[350]},
      {stage0_35[144], stage0_35[145], stage0_35[146], stage0_35[147], stage0_35[148], stage0_35[149]},
      {stage0_36[12]},
      {stage0_37[12]},
      {stage1_38[12],stage1_37[24],stage1_36[76],stage1_35[130],stage1_34[150]}
   );
   gpc1163_5 gpc1327 (
      {stage0_34[351], stage0_34[352], stage0_34[353]},
      {stage0_35[150], stage0_35[151], stage0_35[152], stage0_35[153], stage0_35[154], stage0_35[155]},
      {stage0_36[13]},
      {stage0_37[13]},
      {stage1_38[13],stage1_37[25],stage1_36[77],stage1_35[131],stage1_34[151]}
   );
   gpc1163_5 gpc1328 (
      {stage0_34[354], stage0_34[355], stage0_34[356]},
      {stage0_35[156], stage0_35[157], stage0_35[158], stage0_35[159], stage0_35[160], stage0_35[161]},
      {stage0_36[14]},
      {stage0_37[14]},
      {stage1_38[14],stage1_37[26],stage1_36[78],stage1_35[132],stage1_34[152]}
   );
   gpc1163_5 gpc1329 (
      {stage0_34[357], stage0_34[358], stage0_34[359]},
      {stage0_35[162], stage0_35[163], stage0_35[164], stage0_35[165], stage0_35[166], stage0_35[167]},
      {stage0_36[15]},
      {stage0_37[15]},
      {stage1_38[15],stage1_37[27],stage1_36[79],stage1_35[133],stage1_34[153]}
   );
   gpc1163_5 gpc1330 (
      {stage0_34[360], stage0_34[361], stage0_34[362]},
      {stage0_35[168], stage0_35[169], stage0_35[170], stage0_35[171], stage0_35[172], stage0_35[173]},
      {stage0_36[16]},
      {stage0_37[16]},
      {stage1_38[16],stage1_37[28],stage1_36[80],stage1_35[134],stage1_34[154]}
   );
   gpc1163_5 gpc1331 (
      {stage0_34[363], stage0_34[364], stage0_34[365]},
      {stage0_35[174], stage0_35[175], stage0_35[176], stage0_35[177], stage0_35[178], stage0_35[179]},
      {stage0_36[17]},
      {stage0_37[17]},
      {stage1_38[17],stage1_37[29],stage1_36[81],stage1_35[135],stage1_34[155]}
   );
   gpc1163_5 gpc1332 (
      {stage0_34[366], stage0_34[367], stage0_34[368]},
      {stage0_35[180], stage0_35[181], stage0_35[182], stage0_35[183], stage0_35[184], stage0_35[185]},
      {stage0_36[18]},
      {stage0_37[18]},
      {stage1_38[18],stage1_37[30],stage1_36[82],stage1_35[136],stage1_34[156]}
   );
   gpc1163_5 gpc1333 (
      {stage0_34[369], stage0_34[370], stage0_34[371]},
      {stage0_35[186], stage0_35[187], stage0_35[188], stage0_35[189], stage0_35[190], stage0_35[191]},
      {stage0_36[19]},
      {stage0_37[19]},
      {stage1_38[19],stage1_37[31],stage1_36[83],stage1_35[137],stage1_34[157]}
   );
   gpc1163_5 gpc1334 (
      {stage0_34[372], stage0_34[373], stage0_34[374]},
      {stage0_35[192], stage0_35[193], stage0_35[194], stage0_35[195], stage0_35[196], stage0_35[197]},
      {stage0_36[20]},
      {stage0_37[20]},
      {stage1_38[20],stage1_37[32],stage1_36[84],stage1_35[138],stage1_34[158]}
   );
   gpc1163_5 gpc1335 (
      {stage0_34[375], stage0_34[376], stage0_34[377]},
      {stage0_35[198], stage0_35[199], stage0_35[200], stage0_35[201], stage0_35[202], stage0_35[203]},
      {stage0_36[21]},
      {stage0_37[21]},
      {stage1_38[21],stage1_37[33],stage1_36[85],stage1_35[139],stage1_34[159]}
   );
   gpc1163_5 gpc1336 (
      {stage0_34[378], stage0_34[379], stage0_34[380]},
      {stage0_35[204], stage0_35[205], stage0_35[206], stage0_35[207], stage0_35[208], stage0_35[209]},
      {stage0_36[22]},
      {stage0_37[22]},
      {stage1_38[22],stage1_37[34],stage1_36[86],stage1_35[140],stage1_34[160]}
   );
   gpc1163_5 gpc1337 (
      {stage0_34[381], stage0_34[382], stage0_34[383]},
      {stage0_35[210], stage0_35[211], stage0_35[212], stage0_35[213], stage0_35[214], stage0_35[215]},
      {stage0_36[23]},
      {stage0_37[23]},
      {stage1_38[23],stage1_37[35],stage1_36[87],stage1_35[141],stage1_34[161]}
   );
   gpc1163_5 gpc1338 (
      {stage0_34[384], stage0_34[385], stage0_34[386]},
      {stage0_35[216], stage0_35[217], stage0_35[218], stage0_35[219], stage0_35[220], stage0_35[221]},
      {stage0_36[24]},
      {stage0_37[24]},
      {stage1_38[24],stage1_37[36],stage1_36[88],stage1_35[142],stage1_34[162]}
   );
   gpc1163_5 gpc1339 (
      {stage0_34[387], stage0_34[388], stage0_34[389]},
      {stage0_35[222], stage0_35[223], stage0_35[224], stage0_35[225], stage0_35[226], stage0_35[227]},
      {stage0_36[25]},
      {stage0_37[25]},
      {stage1_38[25],stage1_37[37],stage1_36[89],stage1_35[143],stage1_34[163]}
   );
   gpc1163_5 gpc1340 (
      {stage0_34[390], stage0_34[391], stage0_34[392]},
      {stage0_35[228], stage0_35[229], stage0_35[230], stage0_35[231], stage0_35[232], stage0_35[233]},
      {stage0_36[26]},
      {stage0_37[26]},
      {stage1_38[26],stage1_37[38],stage1_36[90],stage1_35[144],stage1_34[164]}
   );
   gpc1163_5 gpc1341 (
      {stage0_34[393], stage0_34[394], stage0_34[395]},
      {stage0_35[234], stage0_35[235], stage0_35[236], stage0_35[237], stage0_35[238], stage0_35[239]},
      {stage0_36[27]},
      {stage0_37[27]},
      {stage1_38[27],stage1_37[39],stage1_36[91],stage1_35[145],stage1_34[165]}
   );
   gpc1163_5 gpc1342 (
      {stage0_34[396], stage0_34[397], stage0_34[398]},
      {stage0_35[240], stage0_35[241], stage0_35[242], stage0_35[243], stage0_35[244], stage0_35[245]},
      {stage0_36[28]},
      {stage0_37[28]},
      {stage1_38[28],stage1_37[40],stage1_36[92],stage1_35[146],stage1_34[166]}
   );
   gpc1163_5 gpc1343 (
      {stage0_34[399], stage0_34[400], stage0_34[401]},
      {stage0_35[246], stage0_35[247], stage0_35[248], stage0_35[249], stage0_35[250], stage0_35[251]},
      {stage0_36[29]},
      {stage0_37[29]},
      {stage1_38[29],stage1_37[41],stage1_36[93],stage1_35[147],stage1_34[167]}
   );
   gpc1163_5 gpc1344 (
      {stage0_34[402], stage0_34[403], stage0_34[404]},
      {stage0_35[252], stage0_35[253], stage0_35[254], stage0_35[255], stage0_35[256], stage0_35[257]},
      {stage0_36[30]},
      {stage0_37[30]},
      {stage1_38[30],stage1_37[42],stage1_36[94],stage1_35[148],stage1_34[168]}
   );
   gpc1163_5 gpc1345 (
      {stage0_34[405], stage0_34[406], stage0_34[407]},
      {stage0_35[258], stage0_35[259], stage0_35[260], stage0_35[261], stage0_35[262], stage0_35[263]},
      {stage0_36[31]},
      {stage0_37[31]},
      {stage1_38[31],stage1_37[43],stage1_36[95],stage1_35[149],stage1_34[169]}
   );
   gpc1163_5 gpc1346 (
      {stage0_34[408], stage0_34[409], stage0_34[410]},
      {stage0_35[264], stage0_35[265], stage0_35[266], stage0_35[267], stage0_35[268], stage0_35[269]},
      {stage0_36[32]},
      {stage0_37[32]},
      {stage1_38[32],stage1_37[44],stage1_36[96],stage1_35[150],stage1_34[170]}
   );
   gpc1163_5 gpc1347 (
      {stage0_34[411], stage0_34[412], stage0_34[413]},
      {stage0_35[270], stage0_35[271], stage0_35[272], stage0_35[273], stage0_35[274], stage0_35[275]},
      {stage0_36[33]},
      {stage0_37[33]},
      {stage1_38[33],stage1_37[45],stage1_36[97],stage1_35[151],stage1_34[171]}
   );
   gpc1163_5 gpc1348 (
      {stage0_34[414], stage0_34[415], stage0_34[416]},
      {stage0_35[276], stage0_35[277], stage0_35[278], stage0_35[279], stage0_35[280], stage0_35[281]},
      {stage0_36[34]},
      {stage0_37[34]},
      {stage1_38[34],stage1_37[46],stage1_36[98],stage1_35[152],stage1_34[172]}
   );
   gpc1163_5 gpc1349 (
      {stage0_34[417], stage0_34[418], stage0_34[419]},
      {stage0_35[282], stage0_35[283], stage0_35[284], stage0_35[285], stage0_35[286], stage0_35[287]},
      {stage0_36[35]},
      {stage0_37[35]},
      {stage1_38[35],stage1_37[47],stage1_36[99],stage1_35[153],stage1_34[173]}
   );
   gpc1163_5 gpc1350 (
      {stage0_34[420], stage0_34[421], stage0_34[422]},
      {stage0_35[288], stage0_35[289], stage0_35[290], stage0_35[291], stage0_35[292], stage0_35[293]},
      {stage0_36[36]},
      {stage0_37[36]},
      {stage1_38[36],stage1_37[48],stage1_36[100],stage1_35[154],stage1_34[174]}
   );
   gpc1163_5 gpc1351 (
      {stage0_34[423], stage0_34[424], stage0_34[425]},
      {stage0_35[294], stage0_35[295], stage0_35[296], stage0_35[297], stage0_35[298], stage0_35[299]},
      {stage0_36[37]},
      {stage0_37[37]},
      {stage1_38[37],stage1_37[49],stage1_36[101],stage1_35[155],stage1_34[175]}
   );
   gpc1163_5 gpc1352 (
      {stage0_34[426], stage0_34[427], stage0_34[428]},
      {stage0_35[300], stage0_35[301], stage0_35[302], stage0_35[303], stage0_35[304], stage0_35[305]},
      {stage0_36[38]},
      {stage0_37[38]},
      {stage1_38[38],stage1_37[50],stage1_36[102],stage1_35[156],stage1_34[176]}
   );
   gpc1163_5 gpc1353 (
      {stage0_34[429], stage0_34[430], stage0_34[431]},
      {stage0_35[306], stage0_35[307], stage0_35[308], stage0_35[309], stage0_35[310], stage0_35[311]},
      {stage0_36[39]},
      {stage0_37[39]},
      {stage1_38[39],stage1_37[51],stage1_36[103],stage1_35[157],stage1_34[177]}
   );
   gpc1163_5 gpc1354 (
      {stage0_34[432], stage0_34[433], stage0_34[434]},
      {stage0_35[312], stage0_35[313], stage0_35[314], stage0_35[315], stage0_35[316], stage0_35[317]},
      {stage0_36[40]},
      {stage0_37[40]},
      {stage1_38[40],stage1_37[52],stage1_36[104],stage1_35[158],stage1_34[178]}
   );
   gpc1163_5 gpc1355 (
      {stage0_34[435], stage0_34[436], stage0_34[437]},
      {stage0_35[318], stage0_35[319], stage0_35[320], stage0_35[321], stage0_35[322], stage0_35[323]},
      {stage0_36[41]},
      {stage0_37[41]},
      {stage1_38[41],stage1_37[53],stage1_36[105],stage1_35[159],stage1_34[179]}
   );
   gpc1163_5 gpc1356 (
      {stage0_34[438], stage0_34[439], stage0_34[440]},
      {stage0_35[324], stage0_35[325], stage0_35[326], stage0_35[327], stage0_35[328], stage0_35[329]},
      {stage0_36[42]},
      {stage0_37[42]},
      {stage1_38[42],stage1_37[54],stage1_36[106],stage1_35[160],stage1_34[180]}
   );
   gpc615_5 gpc1357 (
      {stage0_34[441], stage0_34[442], stage0_34[443], stage0_34[444], stage0_34[445]},
      {stage0_35[330]},
      {stage0_36[43], stage0_36[44], stage0_36[45], stage0_36[46], stage0_36[47], stage0_36[48]},
      {stage1_38[43],stage1_37[55],stage1_36[107],stage1_35[161],stage1_34[181]}
   );
   gpc615_5 gpc1358 (
      {stage0_34[446], stage0_34[447], stage0_34[448], stage0_34[449], stage0_34[450]},
      {stage0_35[331]},
      {stage0_36[49], stage0_36[50], stage0_36[51], stage0_36[52], stage0_36[53], stage0_36[54]},
      {stage1_38[44],stage1_37[56],stage1_36[108],stage1_35[162],stage1_34[182]}
   );
   gpc615_5 gpc1359 (
      {stage0_34[451], stage0_34[452], stage0_34[453], stage0_34[454], stage0_34[455]},
      {stage0_35[332]},
      {stage0_36[55], stage0_36[56], stage0_36[57], stage0_36[58], stage0_36[59], stage0_36[60]},
      {stage1_38[45],stage1_37[57],stage1_36[109],stage1_35[163],stage1_34[183]}
   );
   gpc615_5 gpc1360 (
      {stage0_34[456], stage0_34[457], stage0_34[458], stage0_34[459], stage0_34[460]},
      {stage0_35[333]},
      {stage0_36[61], stage0_36[62], stage0_36[63], stage0_36[64], stage0_36[65], stage0_36[66]},
      {stage1_38[46],stage1_37[58],stage1_36[110],stage1_35[164],stage1_34[184]}
   );
   gpc615_5 gpc1361 (
      {stage0_34[461], stage0_34[462], stage0_34[463], stage0_34[464], stage0_34[465]},
      {stage0_35[334]},
      {stage0_36[67], stage0_36[68], stage0_36[69], stage0_36[70], stage0_36[71], stage0_36[72]},
      {stage1_38[47],stage1_37[59],stage1_36[111],stage1_35[165],stage1_34[185]}
   );
   gpc615_5 gpc1362 (
      {stage0_34[466], stage0_34[467], stage0_34[468], stage0_34[469], stage0_34[470]},
      {stage0_35[335]},
      {stage0_36[73], stage0_36[74], stage0_36[75], stage0_36[76], stage0_36[77], stage0_36[78]},
      {stage1_38[48],stage1_37[60],stage1_36[112],stage1_35[166],stage1_34[186]}
   );
   gpc615_5 gpc1363 (
      {stage0_34[471], stage0_34[472], stage0_34[473], stage0_34[474], stage0_34[475]},
      {stage0_35[336]},
      {stage0_36[79], stage0_36[80], stage0_36[81], stage0_36[82], stage0_36[83], stage0_36[84]},
      {stage1_38[49],stage1_37[61],stage1_36[113],stage1_35[167],stage1_34[187]}
   );
   gpc615_5 gpc1364 (
      {stage0_34[476], stage0_34[477], stage0_34[478], stage0_34[479], stage0_34[480]},
      {stage0_35[337]},
      {stage0_36[85], stage0_36[86], stage0_36[87], stage0_36[88], stage0_36[89], stage0_36[90]},
      {stage1_38[50],stage1_37[62],stage1_36[114],stage1_35[168],stage1_34[188]}
   );
   gpc615_5 gpc1365 (
      {stage0_34[481], stage0_34[482], stage0_34[483], stage0_34[484], stage0_34[485]},
      {stage0_35[338]},
      {stage0_36[91], stage0_36[92], stage0_36[93], stage0_36[94], stage0_36[95], stage0_36[96]},
      {stage1_38[51],stage1_37[63],stage1_36[115],stage1_35[169],stage1_34[189]}
   );
   gpc615_5 gpc1366 (
      {stage0_35[339], stage0_35[340], stage0_35[341], stage0_35[342], stage0_35[343]},
      {stage0_36[97]},
      {stage0_37[43], stage0_37[44], stage0_37[45], stage0_37[46], stage0_37[47], stage0_37[48]},
      {stage1_39[0],stage1_38[52],stage1_37[64],stage1_36[116],stage1_35[170]}
   );
   gpc615_5 gpc1367 (
      {stage0_35[344], stage0_35[345], stage0_35[346], stage0_35[347], stage0_35[348]},
      {stage0_36[98]},
      {stage0_37[49], stage0_37[50], stage0_37[51], stage0_37[52], stage0_37[53], stage0_37[54]},
      {stage1_39[1],stage1_38[53],stage1_37[65],stage1_36[117],stage1_35[171]}
   );
   gpc615_5 gpc1368 (
      {stage0_35[349], stage0_35[350], stage0_35[351], stage0_35[352], stage0_35[353]},
      {stage0_36[99]},
      {stage0_37[55], stage0_37[56], stage0_37[57], stage0_37[58], stage0_37[59], stage0_37[60]},
      {stage1_39[2],stage1_38[54],stage1_37[66],stage1_36[118],stage1_35[172]}
   );
   gpc615_5 gpc1369 (
      {stage0_35[354], stage0_35[355], stage0_35[356], stage0_35[357], stage0_35[358]},
      {stage0_36[100]},
      {stage0_37[61], stage0_37[62], stage0_37[63], stage0_37[64], stage0_37[65], stage0_37[66]},
      {stage1_39[3],stage1_38[55],stage1_37[67],stage1_36[119],stage1_35[173]}
   );
   gpc615_5 gpc1370 (
      {stage0_35[359], stage0_35[360], stage0_35[361], stage0_35[362], stage0_35[363]},
      {stage0_36[101]},
      {stage0_37[67], stage0_37[68], stage0_37[69], stage0_37[70], stage0_37[71], stage0_37[72]},
      {stage1_39[4],stage1_38[56],stage1_37[68],stage1_36[120],stage1_35[174]}
   );
   gpc615_5 gpc1371 (
      {stage0_35[364], stage0_35[365], stage0_35[366], stage0_35[367], stage0_35[368]},
      {stage0_36[102]},
      {stage0_37[73], stage0_37[74], stage0_37[75], stage0_37[76], stage0_37[77], stage0_37[78]},
      {stage1_39[5],stage1_38[57],stage1_37[69],stage1_36[121],stage1_35[175]}
   );
   gpc615_5 gpc1372 (
      {stage0_35[369], stage0_35[370], stage0_35[371], stage0_35[372], stage0_35[373]},
      {stage0_36[103]},
      {stage0_37[79], stage0_37[80], stage0_37[81], stage0_37[82], stage0_37[83], stage0_37[84]},
      {stage1_39[6],stage1_38[58],stage1_37[70],stage1_36[122],stage1_35[176]}
   );
   gpc615_5 gpc1373 (
      {stage0_35[374], stage0_35[375], stage0_35[376], stage0_35[377], stage0_35[378]},
      {stage0_36[104]},
      {stage0_37[85], stage0_37[86], stage0_37[87], stage0_37[88], stage0_37[89], stage0_37[90]},
      {stage1_39[7],stage1_38[59],stage1_37[71],stage1_36[123],stage1_35[177]}
   );
   gpc615_5 gpc1374 (
      {stage0_35[379], stage0_35[380], stage0_35[381], stage0_35[382], stage0_35[383]},
      {stage0_36[105]},
      {stage0_37[91], stage0_37[92], stage0_37[93], stage0_37[94], stage0_37[95], stage0_37[96]},
      {stage1_39[8],stage1_38[60],stage1_37[72],stage1_36[124],stage1_35[178]}
   );
   gpc615_5 gpc1375 (
      {stage0_35[384], stage0_35[385], stage0_35[386], stage0_35[387], stage0_35[388]},
      {stage0_36[106]},
      {stage0_37[97], stage0_37[98], stage0_37[99], stage0_37[100], stage0_37[101], stage0_37[102]},
      {stage1_39[9],stage1_38[61],stage1_37[73],stage1_36[125],stage1_35[179]}
   );
   gpc615_5 gpc1376 (
      {stage0_35[389], stage0_35[390], stage0_35[391], stage0_35[392], stage0_35[393]},
      {stage0_36[107]},
      {stage0_37[103], stage0_37[104], stage0_37[105], stage0_37[106], stage0_37[107], stage0_37[108]},
      {stage1_39[10],stage1_38[62],stage1_37[74],stage1_36[126],stage1_35[180]}
   );
   gpc615_5 gpc1377 (
      {stage0_35[394], stage0_35[395], stage0_35[396], stage0_35[397], stage0_35[398]},
      {stage0_36[108]},
      {stage0_37[109], stage0_37[110], stage0_37[111], stage0_37[112], stage0_37[113], stage0_37[114]},
      {stage1_39[11],stage1_38[63],stage1_37[75],stage1_36[127],stage1_35[181]}
   );
   gpc615_5 gpc1378 (
      {stage0_35[399], stage0_35[400], stage0_35[401], stage0_35[402], stage0_35[403]},
      {stage0_36[109]},
      {stage0_37[115], stage0_37[116], stage0_37[117], stage0_37[118], stage0_37[119], stage0_37[120]},
      {stage1_39[12],stage1_38[64],stage1_37[76],stage1_36[128],stage1_35[182]}
   );
   gpc615_5 gpc1379 (
      {stage0_35[404], stage0_35[405], stage0_35[406], stage0_35[407], stage0_35[408]},
      {stage0_36[110]},
      {stage0_37[121], stage0_37[122], stage0_37[123], stage0_37[124], stage0_37[125], stage0_37[126]},
      {stage1_39[13],stage1_38[65],stage1_37[77],stage1_36[129],stage1_35[183]}
   );
   gpc615_5 gpc1380 (
      {stage0_35[409], stage0_35[410], stage0_35[411], stage0_35[412], stage0_35[413]},
      {stage0_36[111]},
      {stage0_37[127], stage0_37[128], stage0_37[129], stage0_37[130], stage0_37[131], stage0_37[132]},
      {stage1_39[14],stage1_38[66],stage1_37[78],stage1_36[130],stage1_35[184]}
   );
   gpc615_5 gpc1381 (
      {stage0_35[414], stage0_35[415], stage0_35[416], stage0_35[417], stage0_35[418]},
      {stage0_36[112]},
      {stage0_37[133], stage0_37[134], stage0_37[135], stage0_37[136], stage0_37[137], stage0_37[138]},
      {stage1_39[15],stage1_38[67],stage1_37[79],stage1_36[131],stage1_35[185]}
   );
   gpc615_5 gpc1382 (
      {stage0_35[419], stage0_35[420], stage0_35[421], stage0_35[422], stage0_35[423]},
      {stage0_36[113]},
      {stage0_37[139], stage0_37[140], stage0_37[141], stage0_37[142], stage0_37[143], stage0_37[144]},
      {stage1_39[16],stage1_38[68],stage1_37[80],stage1_36[132],stage1_35[186]}
   );
   gpc615_5 gpc1383 (
      {stage0_35[424], stage0_35[425], stage0_35[426], stage0_35[427], stage0_35[428]},
      {stage0_36[114]},
      {stage0_37[145], stage0_37[146], stage0_37[147], stage0_37[148], stage0_37[149], stage0_37[150]},
      {stage1_39[17],stage1_38[69],stage1_37[81],stage1_36[133],stage1_35[187]}
   );
   gpc615_5 gpc1384 (
      {stage0_35[429], stage0_35[430], stage0_35[431], stage0_35[432], stage0_35[433]},
      {stage0_36[115]},
      {stage0_37[151], stage0_37[152], stage0_37[153], stage0_37[154], stage0_37[155], stage0_37[156]},
      {stage1_39[18],stage1_38[70],stage1_37[82],stage1_36[134],stage1_35[188]}
   );
   gpc615_5 gpc1385 (
      {stage0_35[434], stage0_35[435], stage0_35[436], stage0_35[437], stage0_35[438]},
      {stage0_36[116]},
      {stage0_37[157], stage0_37[158], stage0_37[159], stage0_37[160], stage0_37[161], stage0_37[162]},
      {stage1_39[19],stage1_38[71],stage1_37[83],stage1_36[135],stage1_35[189]}
   );
   gpc615_5 gpc1386 (
      {stage0_35[439], stage0_35[440], stage0_35[441], stage0_35[442], stage0_35[443]},
      {stage0_36[117]},
      {stage0_37[163], stage0_37[164], stage0_37[165], stage0_37[166], stage0_37[167], stage0_37[168]},
      {stage1_39[20],stage1_38[72],stage1_37[84],stage1_36[136],stage1_35[190]}
   );
   gpc615_5 gpc1387 (
      {stage0_35[444], stage0_35[445], stage0_35[446], stage0_35[447], stage0_35[448]},
      {stage0_36[118]},
      {stage0_37[169], stage0_37[170], stage0_37[171], stage0_37[172], stage0_37[173], stage0_37[174]},
      {stage1_39[21],stage1_38[73],stage1_37[85],stage1_36[137],stage1_35[191]}
   );
   gpc615_5 gpc1388 (
      {stage0_35[449], stage0_35[450], stage0_35[451], stage0_35[452], stage0_35[453]},
      {stage0_36[119]},
      {stage0_37[175], stage0_37[176], stage0_37[177], stage0_37[178], stage0_37[179], stage0_37[180]},
      {stage1_39[22],stage1_38[74],stage1_37[86],stage1_36[138],stage1_35[192]}
   );
   gpc615_5 gpc1389 (
      {stage0_35[454], stage0_35[455], stage0_35[456], stage0_35[457], stage0_35[458]},
      {stage0_36[120]},
      {stage0_37[181], stage0_37[182], stage0_37[183], stage0_37[184], stage0_37[185], stage0_37[186]},
      {stage1_39[23],stage1_38[75],stage1_37[87],stage1_36[139],stage1_35[193]}
   );
   gpc615_5 gpc1390 (
      {stage0_35[459], stage0_35[460], stage0_35[461], stage0_35[462], stage0_35[463]},
      {stage0_36[121]},
      {stage0_37[187], stage0_37[188], stage0_37[189], stage0_37[190], stage0_37[191], stage0_37[192]},
      {stage1_39[24],stage1_38[76],stage1_37[88],stage1_36[140],stage1_35[194]}
   );
   gpc606_5 gpc1391 (
      {stage0_36[122], stage0_36[123], stage0_36[124], stage0_36[125], stage0_36[126], stage0_36[127]},
      {stage0_38[0], stage0_38[1], stage0_38[2], stage0_38[3], stage0_38[4], stage0_38[5]},
      {stage1_40[0],stage1_39[25],stage1_38[77],stage1_37[89],stage1_36[141]}
   );
   gpc606_5 gpc1392 (
      {stage0_36[128], stage0_36[129], stage0_36[130], stage0_36[131], stage0_36[132], stage0_36[133]},
      {stage0_38[6], stage0_38[7], stage0_38[8], stage0_38[9], stage0_38[10], stage0_38[11]},
      {stage1_40[1],stage1_39[26],stage1_38[78],stage1_37[90],stage1_36[142]}
   );
   gpc606_5 gpc1393 (
      {stage0_36[134], stage0_36[135], stage0_36[136], stage0_36[137], stage0_36[138], stage0_36[139]},
      {stage0_38[12], stage0_38[13], stage0_38[14], stage0_38[15], stage0_38[16], stage0_38[17]},
      {stage1_40[2],stage1_39[27],stage1_38[79],stage1_37[91],stage1_36[143]}
   );
   gpc606_5 gpc1394 (
      {stage0_36[140], stage0_36[141], stage0_36[142], stage0_36[143], stage0_36[144], stage0_36[145]},
      {stage0_38[18], stage0_38[19], stage0_38[20], stage0_38[21], stage0_38[22], stage0_38[23]},
      {stage1_40[3],stage1_39[28],stage1_38[80],stage1_37[92],stage1_36[144]}
   );
   gpc606_5 gpc1395 (
      {stage0_36[146], stage0_36[147], stage0_36[148], stage0_36[149], stage0_36[150], stage0_36[151]},
      {stage0_38[24], stage0_38[25], stage0_38[26], stage0_38[27], stage0_38[28], stage0_38[29]},
      {stage1_40[4],stage1_39[29],stage1_38[81],stage1_37[93],stage1_36[145]}
   );
   gpc606_5 gpc1396 (
      {stage0_36[152], stage0_36[153], stage0_36[154], stage0_36[155], stage0_36[156], stage0_36[157]},
      {stage0_38[30], stage0_38[31], stage0_38[32], stage0_38[33], stage0_38[34], stage0_38[35]},
      {stage1_40[5],stage1_39[30],stage1_38[82],stage1_37[94],stage1_36[146]}
   );
   gpc606_5 gpc1397 (
      {stage0_36[158], stage0_36[159], stage0_36[160], stage0_36[161], stage0_36[162], stage0_36[163]},
      {stage0_38[36], stage0_38[37], stage0_38[38], stage0_38[39], stage0_38[40], stage0_38[41]},
      {stage1_40[6],stage1_39[31],stage1_38[83],stage1_37[95],stage1_36[147]}
   );
   gpc606_5 gpc1398 (
      {stage0_36[164], stage0_36[165], stage0_36[166], stage0_36[167], stage0_36[168], stage0_36[169]},
      {stage0_38[42], stage0_38[43], stage0_38[44], stage0_38[45], stage0_38[46], stage0_38[47]},
      {stage1_40[7],stage1_39[32],stage1_38[84],stage1_37[96],stage1_36[148]}
   );
   gpc606_5 gpc1399 (
      {stage0_36[170], stage0_36[171], stage0_36[172], stage0_36[173], stage0_36[174], stage0_36[175]},
      {stage0_38[48], stage0_38[49], stage0_38[50], stage0_38[51], stage0_38[52], stage0_38[53]},
      {stage1_40[8],stage1_39[33],stage1_38[85],stage1_37[97],stage1_36[149]}
   );
   gpc606_5 gpc1400 (
      {stage0_36[176], stage0_36[177], stage0_36[178], stage0_36[179], stage0_36[180], stage0_36[181]},
      {stage0_38[54], stage0_38[55], stage0_38[56], stage0_38[57], stage0_38[58], stage0_38[59]},
      {stage1_40[9],stage1_39[34],stage1_38[86],stage1_37[98],stage1_36[150]}
   );
   gpc606_5 gpc1401 (
      {stage0_36[182], stage0_36[183], stage0_36[184], stage0_36[185], stage0_36[186], stage0_36[187]},
      {stage0_38[60], stage0_38[61], stage0_38[62], stage0_38[63], stage0_38[64], stage0_38[65]},
      {stage1_40[10],stage1_39[35],stage1_38[87],stage1_37[99],stage1_36[151]}
   );
   gpc606_5 gpc1402 (
      {stage0_36[188], stage0_36[189], stage0_36[190], stage0_36[191], stage0_36[192], stage0_36[193]},
      {stage0_38[66], stage0_38[67], stage0_38[68], stage0_38[69], stage0_38[70], stage0_38[71]},
      {stage1_40[11],stage1_39[36],stage1_38[88],stage1_37[100],stage1_36[152]}
   );
   gpc606_5 gpc1403 (
      {stage0_36[194], stage0_36[195], stage0_36[196], stage0_36[197], stage0_36[198], stage0_36[199]},
      {stage0_38[72], stage0_38[73], stage0_38[74], stage0_38[75], stage0_38[76], stage0_38[77]},
      {stage1_40[12],stage1_39[37],stage1_38[89],stage1_37[101],stage1_36[153]}
   );
   gpc606_5 gpc1404 (
      {stage0_36[200], stage0_36[201], stage0_36[202], stage0_36[203], stage0_36[204], stage0_36[205]},
      {stage0_38[78], stage0_38[79], stage0_38[80], stage0_38[81], stage0_38[82], stage0_38[83]},
      {stage1_40[13],stage1_39[38],stage1_38[90],stage1_37[102],stage1_36[154]}
   );
   gpc606_5 gpc1405 (
      {stage0_36[206], stage0_36[207], stage0_36[208], stage0_36[209], stage0_36[210], stage0_36[211]},
      {stage0_38[84], stage0_38[85], stage0_38[86], stage0_38[87], stage0_38[88], stage0_38[89]},
      {stage1_40[14],stage1_39[39],stage1_38[91],stage1_37[103],stage1_36[155]}
   );
   gpc606_5 gpc1406 (
      {stage0_36[212], stage0_36[213], stage0_36[214], stage0_36[215], stage0_36[216], stage0_36[217]},
      {stage0_38[90], stage0_38[91], stage0_38[92], stage0_38[93], stage0_38[94], stage0_38[95]},
      {stage1_40[15],stage1_39[40],stage1_38[92],stage1_37[104],stage1_36[156]}
   );
   gpc606_5 gpc1407 (
      {stage0_36[218], stage0_36[219], stage0_36[220], stage0_36[221], stage0_36[222], stage0_36[223]},
      {stage0_38[96], stage0_38[97], stage0_38[98], stage0_38[99], stage0_38[100], stage0_38[101]},
      {stage1_40[16],stage1_39[41],stage1_38[93],stage1_37[105],stage1_36[157]}
   );
   gpc606_5 gpc1408 (
      {stage0_36[224], stage0_36[225], stage0_36[226], stage0_36[227], stage0_36[228], stage0_36[229]},
      {stage0_38[102], stage0_38[103], stage0_38[104], stage0_38[105], stage0_38[106], stage0_38[107]},
      {stage1_40[17],stage1_39[42],stage1_38[94],stage1_37[106],stage1_36[158]}
   );
   gpc606_5 gpc1409 (
      {stage0_36[230], stage0_36[231], stage0_36[232], stage0_36[233], stage0_36[234], stage0_36[235]},
      {stage0_38[108], stage0_38[109], stage0_38[110], stage0_38[111], stage0_38[112], stage0_38[113]},
      {stage1_40[18],stage1_39[43],stage1_38[95],stage1_37[107],stage1_36[159]}
   );
   gpc606_5 gpc1410 (
      {stage0_36[236], stage0_36[237], stage0_36[238], stage0_36[239], stage0_36[240], stage0_36[241]},
      {stage0_38[114], stage0_38[115], stage0_38[116], stage0_38[117], stage0_38[118], stage0_38[119]},
      {stage1_40[19],stage1_39[44],stage1_38[96],stage1_37[108],stage1_36[160]}
   );
   gpc606_5 gpc1411 (
      {stage0_36[242], stage0_36[243], stage0_36[244], stage0_36[245], stage0_36[246], stage0_36[247]},
      {stage0_38[120], stage0_38[121], stage0_38[122], stage0_38[123], stage0_38[124], stage0_38[125]},
      {stage1_40[20],stage1_39[45],stage1_38[97],stage1_37[109],stage1_36[161]}
   );
   gpc606_5 gpc1412 (
      {stage0_36[248], stage0_36[249], stage0_36[250], stage0_36[251], stage0_36[252], stage0_36[253]},
      {stage0_38[126], stage0_38[127], stage0_38[128], stage0_38[129], stage0_38[130], stage0_38[131]},
      {stage1_40[21],stage1_39[46],stage1_38[98],stage1_37[110],stage1_36[162]}
   );
   gpc606_5 gpc1413 (
      {stage0_36[254], stage0_36[255], stage0_36[256], stage0_36[257], stage0_36[258], stage0_36[259]},
      {stage0_38[132], stage0_38[133], stage0_38[134], stage0_38[135], stage0_38[136], stage0_38[137]},
      {stage1_40[22],stage1_39[47],stage1_38[99],stage1_37[111],stage1_36[163]}
   );
   gpc606_5 gpc1414 (
      {stage0_36[260], stage0_36[261], stage0_36[262], stage0_36[263], stage0_36[264], stage0_36[265]},
      {stage0_38[138], stage0_38[139], stage0_38[140], stage0_38[141], stage0_38[142], stage0_38[143]},
      {stage1_40[23],stage1_39[48],stage1_38[100],stage1_37[112],stage1_36[164]}
   );
   gpc606_5 gpc1415 (
      {stage0_36[266], stage0_36[267], stage0_36[268], stage0_36[269], stage0_36[270], stage0_36[271]},
      {stage0_38[144], stage0_38[145], stage0_38[146], stage0_38[147], stage0_38[148], stage0_38[149]},
      {stage1_40[24],stage1_39[49],stage1_38[101],stage1_37[113],stage1_36[165]}
   );
   gpc606_5 gpc1416 (
      {stage0_36[272], stage0_36[273], stage0_36[274], stage0_36[275], stage0_36[276], stage0_36[277]},
      {stage0_38[150], stage0_38[151], stage0_38[152], stage0_38[153], stage0_38[154], stage0_38[155]},
      {stage1_40[25],stage1_39[50],stage1_38[102],stage1_37[114],stage1_36[166]}
   );
   gpc606_5 gpc1417 (
      {stage0_36[278], stage0_36[279], stage0_36[280], stage0_36[281], stage0_36[282], stage0_36[283]},
      {stage0_38[156], stage0_38[157], stage0_38[158], stage0_38[159], stage0_38[160], stage0_38[161]},
      {stage1_40[26],stage1_39[51],stage1_38[103],stage1_37[115],stage1_36[167]}
   );
   gpc606_5 gpc1418 (
      {stage0_36[284], stage0_36[285], stage0_36[286], stage0_36[287], stage0_36[288], stage0_36[289]},
      {stage0_38[162], stage0_38[163], stage0_38[164], stage0_38[165], stage0_38[166], stage0_38[167]},
      {stage1_40[27],stage1_39[52],stage1_38[104],stage1_37[116],stage1_36[168]}
   );
   gpc606_5 gpc1419 (
      {stage0_36[290], stage0_36[291], stage0_36[292], stage0_36[293], stage0_36[294], stage0_36[295]},
      {stage0_38[168], stage0_38[169], stage0_38[170], stage0_38[171], stage0_38[172], stage0_38[173]},
      {stage1_40[28],stage1_39[53],stage1_38[105],stage1_37[117],stage1_36[169]}
   );
   gpc606_5 gpc1420 (
      {stage0_36[296], stage0_36[297], stage0_36[298], stage0_36[299], stage0_36[300], stage0_36[301]},
      {stage0_38[174], stage0_38[175], stage0_38[176], stage0_38[177], stage0_38[178], stage0_38[179]},
      {stage1_40[29],stage1_39[54],stage1_38[106],stage1_37[118],stage1_36[170]}
   );
   gpc606_5 gpc1421 (
      {stage0_36[302], stage0_36[303], stage0_36[304], stage0_36[305], stage0_36[306], stage0_36[307]},
      {stage0_38[180], stage0_38[181], stage0_38[182], stage0_38[183], stage0_38[184], stage0_38[185]},
      {stage1_40[30],stage1_39[55],stage1_38[107],stage1_37[119],stage1_36[171]}
   );
   gpc606_5 gpc1422 (
      {stage0_36[308], stage0_36[309], stage0_36[310], stage0_36[311], stage0_36[312], stage0_36[313]},
      {stage0_38[186], stage0_38[187], stage0_38[188], stage0_38[189], stage0_38[190], stage0_38[191]},
      {stage1_40[31],stage1_39[56],stage1_38[108],stage1_37[120],stage1_36[172]}
   );
   gpc606_5 gpc1423 (
      {stage0_36[314], stage0_36[315], stage0_36[316], stage0_36[317], stage0_36[318], stage0_36[319]},
      {stage0_38[192], stage0_38[193], stage0_38[194], stage0_38[195], stage0_38[196], stage0_38[197]},
      {stage1_40[32],stage1_39[57],stage1_38[109],stage1_37[121],stage1_36[173]}
   );
   gpc606_5 gpc1424 (
      {stage0_36[320], stage0_36[321], stage0_36[322], stage0_36[323], stage0_36[324], stage0_36[325]},
      {stage0_38[198], stage0_38[199], stage0_38[200], stage0_38[201], stage0_38[202], stage0_38[203]},
      {stage1_40[33],stage1_39[58],stage1_38[110],stage1_37[122],stage1_36[174]}
   );
   gpc606_5 gpc1425 (
      {stage0_36[326], stage0_36[327], stage0_36[328], stage0_36[329], stage0_36[330], stage0_36[331]},
      {stage0_38[204], stage0_38[205], stage0_38[206], stage0_38[207], stage0_38[208], stage0_38[209]},
      {stage1_40[34],stage1_39[59],stage1_38[111],stage1_37[123],stage1_36[175]}
   );
   gpc606_5 gpc1426 (
      {stage0_36[332], stage0_36[333], stage0_36[334], stage0_36[335], stage0_36[336], stage0_36[337]},
      {stage0_38[210], stage0_38[211], stage0_38[212], stage0_38[213], stage0_38[214], stage0_38[215]},
      {stage1_40[35],stage1_39[60],stage1_38[112],stage1_37[124],stage1_36[176]}
   );
   gpc606_5 gpc1427 (
      {stage0_36[338], stage0_36[339], stage0_36[340], stage0_36[341], stage0_36[342], stage0_36[343]},
      {stage0_38[216], stage0_38[217], stage0_38[218], stage0_38[219], stage0_38[220], stage0_38[221]},
      {stage1_40[36],stage1_39[61],stage1_38[113],stage1_37[125],stage1_36[177]}
   );
   gpc606_5 gpc1428 (
      {stage0_36[344], stage0_36[345], stage0_36[346], stage0_36[347], stage0_36[348], stage0_36[349]},
      {stage0_38[222], stage0_38[223], stage0_38[224], stage0_38[225], stage0_38[226], stage0_38[227]},
      {stage1_40[37],stage1_39[62],stage1_38[114],stage1_37[126],stage1_36[178]}
   );
   gpc606_5 gpc1429 (
      {stage0_36[350], stage0_36[351], stage0_36[352], stage0_36[353], stage0_36[354], stage0_36[355]},
      {stage0_38[228], stage0_38[229], stage0_38[230], stage0_38[231], stage0_38[232], stage0_38[233]},
      {stage1_40[38],stage1_39[63],stage1_38[115],stage1_37[127],stage1_36[179]}
   );
   gpc606_5 gpc1430 (
      {stage0_36[356], stage0_36[357], stage0_36[358], stage0_36[359], stage0_36[360], stage0_36[361]},
      {stage0_38[234], stage0_38[235], stage0_38[236], stage0_38[237], stage0_38[238], stage0_38[239]},
      {stage1_40[39],stage1_39[64],stage1_38[116],stage1_37[128],stage1_36[180]}
   );
   gpc606_5 gpc1431 (
      {stage0_36[362], stage0_36[363], stage0_36[364], stage0_36[365], stage0_36[366], stage0_36[367]},
      {stage0_38[240], stage0_38[241], stage0_38[242], stage0_38[243], stage0_38[244], stage0_38[245]},
      {stage1_40[40],stage1_39[65],stage1_38[117],stage1_37[129],stage1_36[181]}
   );
   gpc606_5 gpc1432 (
      {stage0_36[368], stage0_36[369], stage0_36[370], stage0_36[371], stage0_36[372], stage0_36[373]},
      {stage0_38[246], stage0_38[247], stage0_38[248], stage0_38[249], stage0_38[250], stage0_38[251]},
      {stage1_40[41],stage1_39[66],stage1_38[118],stage1_37[130],stage1_36[182]}
   );
   gpc606_5 gpc1433 (
      {stage0_36[374], stage0_36[375], stage0_36[376], stage0_36[377], stage0_36[378], stage0_36[379]},
      {stage0_38[252], stage0_38[253], stage0_38[254], stage0_38[255], stage0_38[256], stage0_38[257]},
      {stage1_40[42],stage1_39[67],stage1_38[119],stage1_37[131],stage1_36[183]}
   );
   gpc606_5 gpc1434 (
      {stage0_36[380], stage0_36[381], stage0_36[382], stage0_36[383], stage0_36[384], stage0_36[385]},
      {stage0_38[258], stage0_38[259], stage0_38[260], stage0_38[261], stage0_38[262], stage0_38[263]},
      {stage1_40[43],stage1_39[68],stage1_38[120],stage1_37[132],stage1_36[184]}
   );
   gpc606_5 gpc1435 (
      {stage0_36[386], stage0_36[387], stage0_36[388], stage0_36[389], stage0_36[390], stage0_36[391]},
      {stage0_38[264], stage0_38[265], stage0_38[266], stage0_38[267], stage0_38[268], stage0_38[269]},
      {stage1_40[44],stage1_39[69],stage1_38[121],stage1_37[133],stage1_36[185]}
   );
   gpc606_5 gpc1436 (
      {stage0_36[392], stage0_36[393], stage0_36[394], stage0_36[395], stage0_36[396], stage0_36[397]},
      {stage0_38[270], stage0_38[271], stage0_38[272], stage0_38[273], stage0_38[274], stage0_38[275]},
      {stage1_40[45],stage1_39[70],stage1_38[122],stage1_37[134],stage1_36[186]}
   );
   gpc606_5 gpc1437 (
      {stage0_36[398], stage0_36[399], stage0_36[400], stage0_36[401], stage0_36[402], stage0_36[403]},
      {stage0_38[276], stage0_38[277], stage0_38[278], stage0_38[279], stage0_38[280], stage0_38[281]},
      {stage1_40[46],stage1_39[71],stage1_38[123],stage1_37[135],stage1_36[187]}
   );
   gpc606_5 gpc1438 (
      {stage0_36[404], stage0_36[405], stage0_36[406], stage0_36[407], stage0_36[408], stage0_36[409]},
      {stage0_38[282], stage0_38[283], stage0_38[284], stage0_38[285], stage0_38[286], stage0_38[287]},
      {stage1_40[47],stage1_39[72],stage1_38[124],stage1_37[136],stage1_36[188]}
   );
   gpc606_5 gpc1439 (
      {stage0_36[410], stage0_36[411], stage0_36[412], stage0_36[413], stage0_36[414], stage0_36[415]},
      {stage0_38[288], stage0_38[289], stage0_38[290], stage0_38[291], stage0_38[292], stage0_38[293]},
      {stage1_40[48],stage1_39[73],stage1_38[125],stage1_37[137],stage1_36[189]}
   );
   gpc606_5 gpc1440 (
      {stage0_36[416], stage0_36[417], stage0_36[418], stage0_36[419], stage0_36[420], stage0_36[421]},
      {stage0_38[294], stage0_38[295], stage0_38[296], stage0_38[297], stage0_38[298], stage0_38[299]},
      {stage1_40[49],stage1_39[74],stage1_38[126],stage1_37[138],stage1_36[190]}
   );
   gpc606_5 gpc1441 (
      {stage0_36[422], stage0_36[423], stage0_36[424], stage0_36[425], stage0_36[426], stage0_36[427]},
      {stage0_38[300], stage0_38[301], stage0_38[302], stage0_38[303], stage0_38[304], stage0_38[305]},
      {stage1_40[50],stage1_39[75],stage1_38[127],stage1_37[139],stage1_36[191]}
   );
   gpc606_5 gpc1442 (
      {stage0_36[428], stage0_36[429], stage0_36[430], stage0_36[431], stage0_36[432], stage0_36[433]},
      {stage0_38[306], stage0_38[307], stage0_38[308], stage0_38[309], stage0_38[310], stage0_38[311]},
      {stage1_40[51],stage1_39[76],stage1_38[128],stage1_37[140],stage1_36[192]}
   );
   gpc606_5 gpc1443 (
      {stage0_36[434], stage0_36[435], stage0_36[436], stage0_36[437], stage0_36[438], stage0_36[439]},
      {stage0_38[312], stage0_38[313], stage0_38[314], stage0_38[315], stage0_38[316], stage0_38[317]},
      {stage1_40[52],stage1_39[77],stage1_38[129],stage1_37[141],stage1_36[193]}
   );
   gpc606_5 gpc1444 (
      {stage0_36[440], stage0_36[441], stage0_36[442], stage0_36[443], stage0_36[444], stage0_36[445]},
      {stage0_38[318], stage0_38[319], stage0_38[320], stage0_38[321], stage0_38[322], stage0_38[323]},
      {stage1_40[53],stage1_39[78],stage1_38[130],stage1_37[142],stage1_36[194]}
   );
   gpc606_5 gpc1445 (
      {stage0_36[446], stage0_36[447], stage0_36[448], stage0_36[449], stage0_36[450], stage0_36[451]},
      {stage0_38[324], stage0_38[325], stage0_38[326], stage0_38[327], stage0_38[328], stage0_38[329]},
      {stage1_40[54],stage1_39[79],stage1_38[131],stage1_37[143],stage1_36[195]}
   );
   gpc606_5 gpc1446 (
      {stage0_36[452], stage0_36[453], stage0_36[454], stage0_36[455], stage0_36[456], stage0_36[457]},
      {stage0_38[330], stage0_38[331], stage0_38[332], stage0_38[333], stage0_38[334], stage0_38[335]},
      {stage1_40[55],stage1_39[80],stage1_38[132],stage1_37[144],stage1_36[196]}
   );
   gpc606_5 gpc1447 (
      {stage0_36[458], stage0_36[459], stage0_36[460], stage0_36[461], stage0_36[462], stage0_36[463]},
      {stage0_38[336], stage0_38[337], stage0_38[338], stage0_38[339], stage0_38[340], stage0_38[341]},
      {stage1_40[56],stage1_39[81],stage1_38[133],stage1_37[145],stage1_36[197]}
   );
   gpc606_5 gpc1448 (
      {stage0_36[464], stage0_36[465], stage0_36[466], stage0_36[467], stage0_36[468], stage0_36[469]},
      {stage0_38[342], stage0_38[343], stage0_38[344], stage0_38[345], stage0_38[346], stage0_38[347]},
      {stage1_40[57],stage1_39[82],stage1_38[134],stage1_37[146],stage1_36[198]}
   );
   gpc606_5 gpc1449 (
      {stage0_36[470], stage0_36[471], stage0_36[472], stage0_36[473], stage0_36[474], stage0_36[475]},
      {stage0_38[348], stage0_38[349], stage0_38[350], stage0_38[351], stage0_38[352], stage0_38[353]},
      {stage1_40[58],stage1_39[83],stage1_38[135],stage1_37[147],stage1_36[199]}
   );
   gpc606_5 gpc1450 (
      {stage0_36[476], stage0_36[477], stage0_36[478], stage0_36[479], stage0_36[480], stage0_36[481]},
      {stage0_38[354], stage0_38[355], stage0_38[356], stage0_38[357], stage0_38[358], stage0_38[359]},
      {stage1_40[59],stage1_39[84],stage1_38[136],stage1_37[148],stage1_36[200]}
   );
   gpc606_5 gpc1451 (
      {stage0_36[482], stage0_36[483], stage0_36[484], stage0_36[485], 1'b0, 1'b0},
      {stage0_38[360], stage0_38[361], stage0_38[362], stage0_38[363], stage0_38[364], stage0_38[365]},
      {stage1_40[60],stage1_39[85],stage1_38[137],stage1_37[149],stage1_36[201]}
   );
   gpc606_5 gpc1452 (
      {stage0_37[193], stage0_37[194], stage0_37[195], stage0_37[196], stage0_37[197], stage0_37[198]},
      {stage0_39[0], stage0_39[1], stage0_39[2], stage0_39[3], stage0_39[4], stage0_39[5]},
      {stage1_41[0],stage1_40[61],stage1_39[86],stage1_38[138],stage1_37[150]}
   );
   gpc606_5 gpc1453 (
      {stage0_37[199], stage0_37[200], stage0_37[201], stage0_37[202], stage0_37[203], stage0_37[204]},
      {stage0_39[6], stage0_39[7], stage0_39[8], stage0_39[9], stage0_39[10], stage0_39[11]},
      {stage1_41[1],stage1_40[62],stage1_39[87],stage1_38[139],stage1_37[151]}
   );
   gpc606_5 gpc1454 (
      {stage0_37[205], stage0_37[206], stage0_37[207], stage0_37[208], stage0_37[209], stage0_37[210]},
      {stage0_39[12], stage0_39[13], stage0_39[14], stage0_39[15], stage0_39[16], stage0_39[17]},
      {stage1_41[2],stage1_40[63],stage1_39[88],stage1_38[140],stage1_37[152]}
   );
   gpc606_5 gpc1455 (
      {stage0_37[211], stage0_37[212], stage0_37[213], stage0_37[214], stage0_37[215], stage0_37[216]},
      {stage0_39[18], stage0_39[19], stage0_39[20], stage0_39[21], stage0_39[22], stage0_39[23]},
      {stage1_41[3],stage1_40[64],stage1_39[89],stage1_38[141],stage1_37[153]}
   );
   gpc606_5 gpc1456 (
      {stage0_37[217], stage0_37[218], stage0_37[219], stage0_37[220], stage0_37[221], stage0_37[222]},
      {stage0_39[24], stage0_39[25], stage0_39[26], stage0_39[27], stage0_39[28], stage0_39[29]},
      {stage1_41[4],stage1_40[65],stage1_39[90],stage1_38[142],stage1_37[154]}
   );
   gpc606_5 gpc1457 (
      {stage0_37[223], stage0_37[224], stage0_37[225], stage0_37[226], stage0_37[227], stage0_37[228]},
      {stage0_39[30], stage0_39[31], stage0_39[32], stage0_39[33], stage0_39[34], stage0_39[35]},
      {stage1_41[5],stage1_40[66],stage1_39[91],stage1_38[143],stage1_37[155]}
   );
   gpc606_5 gpc1458 (
      {stage0_37[229], stage0_37[230], stage0_37[231], stage0_37[232], stage0_37[233], stage0_37[234]},
      {stage0_39[36], stage0_39[37], stage0_39[38], stage0_39[39], stage0_39[40], stage0_39[41]},
      {stage1_41[6],stage1_40[67],stage1_39[92],stage1_38[144],stage1_37[156]}
   );
   gpc606_5 gpc1459 (
      {stage0_37[235], stage0_37[236], stage0_37[237], stage0_37[238], stage0_37[239], stage0_37[240]},
      {stage0_39[42], stage0_39[43], stage0_39[44], stage0_39[45], stage0_39[46], stage0_39[47]},
      {stage1_41[7],stage1_40[68],stage1_39[93],stage1_38[145],stage1_37[157]}
   );
   gpc606_5 gpc1460 (
      {stage0_37[241], stage0_37[242], stage0_37[243], stage0_37[244], stage0_37[245], stage0_37[246]},
      {stage0_39[48], stage0_39[49], stage0_39[50], stage0_39[51], stage0_39[52], stage0_39[53]},
      {stage1_41[8],stage1_40[69],stage1_39[94],stage1_38[146],stage1_37[158]}
   );
   gpc606_5 gpc1461 (
      {stage0_37[247], stage0_37[248], stage0_37[249], stage0_37[250], stage0_37[251], stage0_37[252]},
      {stage0_39[54], stage0_39[55], stage0_39[56], stage0_39[57], stage0_39[58], stage0_39[59]},
      {stage1_41[9],stage1_40[70],stage1_39[95],stage1_38[147],stage1_37[159]}
   );
   gpc606_5 gpc1462 (
      {stage0_37[253], stage0_37[254], stage0_37[255], stage0_37[256], stage0_37[257], stage0_37[258]},
      {stage0_39[60], stage0_39[61], stage0_39[62], stage0_39[63], stage0_39[64], stage0_39[65]},
      {stage1_41[10],stage1_40[71],stage1_39[96],stage1_38[148],stage1_37[160]}
   );
   gpc606_5 gpc1463 (
      {stage0_37[259], stage0_37[260], stage0_37[261], stage0_37[262], stage0_37[263], stage0_37[264]},
      {stage0_39[66], stage0_39[67], stage0_39[68], stage0_39[69], stage0_39[70], stage0_39[71]},
      {stage1_41[11],stage1_40[72],stage1_39[97],stage1_38[149],stage1_37[161]}
   );
   gpc606_5 gpc1464 (
      {stage0_37[265], stage0_37[266], stage0_37[267], stage0_37[268], stage0_37[269], stage0_37[270]},
      {stage0_39[72], stage0_39[73], stage0_39[74], stage0_39[75], stage0_39[76], stage0_39[77]},
      {stage1_41[12],stage1_40[73],stage1_39[98],stage1_38[150],stage1_37[162]}
   );
   gpc606_5 gpc1465 (
      {stage0_37[271], stage0_37[272], stage0_37[273], stage0_37[274], stage0_37[275], stage0_37[276]},
      {stage0_39[78], stage0_39[79], stage0_39[80], stage0_39[81], stage0_39[82], stage0_39[83]},
      {stage1_41[13],stage1_40[74],stage1_39[99],stage1_38[151],stage1_37[163]}
   );
   gpc606_5 gpc1466 (
      {stage0_37[277], stage0_37[278], stage0_37[279], stage0_37[280], stage0_37[281], stage0_37[282]},
      {stage0_39[84], stage0_39[85], stage0_39[86], stage0_39[87], stage0_39[88], stage0_39[89]},
      {stage1_41[14],stage1_40[75],stage1_39[100],stage1_38[152],stage1_37[164]}
   );
   gpc606_5 gpc1467 (
      {stage0_37[283], stage0_37[284], stage0_37[285], stage0_37[286], stage0_37[287], stage0_37[288]},
      {stage0_39[90], stage0_39[91], stage0_39[92], stage0_39[93], stage0_39[94], stage0_39[95]},
      {stage1_41[15],stage1_40[76],stage1_39[101],stage1_38[153],stage1_37[165]}
   );
   gpc606_5 gpc1468 (
      {stage0_37[289], stage0_37[290], stage0_37[291], stage0_37[292], stage0_37[293], stage0_37[294]},
      {stage0_39[96], stage0_39[97], stage0_39[98], stage0_39[99], stage0_39[100], stage0_39[101]},
      {stage1_41[16],stage1_40[77],stage1_39[102],stage1_38[154],stage1_37[166]}
   );
   gpc606_5 gpc1469 (
      {stage0_37[295], stage0_37[296], stage0_37[297], stage0_37[298], stage0_37[299], stage0_37[300]},
      {stage0_39[102], stage0_39[103], stage0_39[104], stage0_39[105], stage0_39[106], stage0_39[107]},
      {stage1_41[17],stage1_40[78],stage1_39[103],stage1_38[155],stage1_37[167]}
   );
   gpc606_5 gpc1470 (
      {stage0_37[301], stage0_37[302], stage0_37[303], stage0_37[304], stage0_37[305], stage0_37[306]},
      {stage0_39[108], stage0_39[109], stage0_39[110], stage0_39[111], stage0_39[112], stage0_39[113]},
      {stage1_41[18],stage1_40[79],stage1_39[104],stage1_38[156],stage1_37[168]}
   );
   gpc606_5 gpc1471 (
      {stage0_37[307], stage0_37[308], stage0_37[309], stage0_37[310], stage0_37[311], stage0_37[312]},
      {stage0_39[114], stage0_39[115], stage0_39[116], stage0_39[117], stage0_39[118], stage0_39[119]},
      {stage1_41[19],stage1_40[80],stage1_39[105],stage1_38[157],stage1_37[169]}
   );
   gpc606_5 gpc1472 (
      {stage0_37[313], stage0_37[314], stage0_37[315], stage0_37[316], stage0_37[317], stage0_37[318]},
      {stage0_39[120], stage0_39[121], stage0_39[122], stage0_39[123], stage0_39[124], stage0_39[125]},
      {stage1_41[20],stage1_40[81],stage1_39[106],stage1_38[158],stage1_37[170]}
   );
   gpc606_5 gpc1473 (
      {stage0_37[319], stage0_37[320], stage0_37[321], stage0_37[322], stage0_37[323], stage0_37[324]},
      {stage0_39[126], stage0_39[127], stage0_39[128], stage0_39[129], stage0_39[130], stage0_39[131]},
      {stage1_41[21],stage1_40[82],stage1_39[107],stage1_38[159],stage1_37[171]}
   );
   gpc606_5 gpc1474 (
      {stage0_37[325], stage0_37[326], stage0_37[327], stage0_37[328], stage0_37[329], stage0_37[330]},
      {stage0_39[132], stage0_39[133], stage0_39[134], stage0_39[135], stage0_39[136], stage0_39[137]},
      {stage1_41[22],stage1_40[83],stage1_39[108],stage1_38[160],stage1_37[172]}
   );
   gpc606_5 gpc1475 (
      {stage0_37[331], stage0_37[332], stage0_37[333], stage0_37[334], stage0_37[335], stage0_37[336]},
      {stage0_39[138], stage0_39[139], stage0_39[140], stage0_39[141], stage0_39[142], stage0_39[143]},
      {stage1_41[23],stage1_40[84],stage1_39[109],stage1_38[161],stage1_37[173]}
   );
   gpc606_5 gpc1476 (
      {stage0_37[337], stage0_37[338], stage0_37[339], stage0_37[340], stage0_37[341], stage0_37[342]},
      {stage0_39[144], stage0_39[145], stage0_39[146], stage0_39[147], stage0_39[148], stage0_39[149]},
      {stage1_41[24],stage1_40[85],stage1_39[110],stage1_38[162],stage1_37[174]}
   );
   gpc606_5 gpc1477 (
      {stage0_37[343], stage0_37[344], stage0_37[345], stage0_37[346], stage0_37[347], stage0_37[348]},
      {stage0_39[150], stage0_39[151], stage0_39[152], stage0_39[153], stage0_39[154], stage0_39[155]},
      {stage1_41[25],stage1_40[86],stage1_39[111],stage1_38[163],stage1_37[175]}
   );
   gpc606_5 gpc1478 (
      {stage0_37[349], stage0_37[350], stage0_37[351], stage0_37[352], stage0_37[353], stage0_37[354]},
      {stage0_39[156], stage0_39[157], stage0_39[158], stage0_39[159], stage0_39[160], stage0_39[161]},
      {stage1_41[26],stage1_40[87],stage1_39[112],stage1_38[164],stage1_37[176]}
   );
   gpc615_5 gpc1479 (
      {stage0_38[366], stage0_38[367], stage0_38[368], stage0_38[369], stage0_38[370]},
      {stage0_39[162]},
      {stage0_40[0], stage0_40[1], stage0_40[2], stage0_40[3], stage0_40[4], stage0_40[5]},
      {stage1_42[0],stage1_41[27],stage1_40[88],stage1_39[113],stage1_38[165]}
   );
   gpc615_5 gpc1480 (
      {stage0_38[371], stage0_38[372], stage0_38[373], stage0_38[374], stage0_38[375]},
      {stage0_39[163]},
      {stage0_40[6], stage0_40[7], stage0_40[8], stage0_40[9], stage0_40[10], stage0_40[11]},
      {stage1_42[1],stage1_41[28],stage1_40[89],stage1_39[114],stage1_38[166]}
   );
   gpc615_5 gpc1481 (
      {stage0_38[376], stage0_38[377], stage0_38[378], stage0_38[379], stage0_38[380]},
      {stage0_39[164]},
      {stage0_40[12], stage0_40[13], stage0_40[14], stage0_40[15], stage0_40[16], stage0_40[17]},
      {stage1_42[2],stage1_41[29],stage1_40[90],stage1_39[115],stage1_38[167]}
   );
   gpc615_5 gpc1482 (
      {stage0_38[381], stage0_38[382], stage0_38[383], stage0_38[384], stage0_38[385]},
      {stage0_39[165]},
      {stage0_40[18], stage0_40[19], stage0_40[20], stage0_40[21], stage0_40[22], stage0_40[23]},
      {stage1_42[3],stage1_41[30],stage1_40[91],stage1_39[116],stage1_38[168]}
   );
   gpc615_5 gpc1483 (
      {stage0_38[386], stage0_38[387], stage0_38[388], stage0_38[389], stage0_38[390]},
      {stage0_39[166]},
      {stage0_40[24], stage0_40[25], stage0_40[26], stage0_40[27], stage0_40[28], stage0_40[29]},
      {stage1_42[4],stage1_41[31],stage1_40[92],stage1_39[117],stage1_38[169]}
   );
   gpc615_5 gpc1484 (
      {stage0_39[167], stage0_39[168], stage0_39[169], stage0_39[170], stage0_39[171]},
      {stage0_40[30]},
      {stage0_41[0], stage0_41[1], stage0_41[2], stage0_41[3], stage0_41[4], stage0_41[5]},
      {stage1_43[0],stage1_42[5],stage1_41[32],stage1_40[93],stage1_39[118]}
   );
   gpc615_5 gpc1485 (
      {stage0_39[172], stage0_39[173], stage0_39[174], stage0_39[175], stage0_39[176]},
      {stage0_40[31]},
      {stage0_41[6], stage0_41[7], stage0_41[8], stage0_41[9], stage0_41[10], stage0_41[11]},
      {stage1_43[1],stage1_42[6],stage1_41[33],stage1_40[94],stage1_39[119]}
   );
   gpc615_5 gpc1486 (
      {stage0_39[177], stage0_39[178], stage0_39[179], stage0_39[180], stage0_39[181]},
      {stage0_40[32]},
      {stage0_41[12], stage0_41[13], stage0_41[14], stage0_41[15], stage0_41[16], stage0_41[17]},
      {stage1_43[2],stage1_42[7],stage1_41[34],stage1_40[95],stage1_39[120]}
   );
   gpc615_5 gpc1487 (
      {stage0_39[182], stage0_39[183], stage0_39[184], stage0_39[185], stage0_39[186]},
      {stage0_40[33]},
      {stage0_41[18], stage0_41[19], stage0_41[20], stage0_41[21], stage0_41[22], stage0_41[23]},
      {stage1_43[3],stage1_42[8],stage1_41[35],stage1_40[96],stage1_39[121]}
   );
   gpc615_5 gpc1488 (
      {stage0_39[187], stage0_39[188], stage0_39[189], stage0_39[190], stage0_39[191]},
      {stage0_40[34]},
      {stage0_41[24], stage0_41[25], stage0_41[26], stage0_41[27], stage0_41[28], stage0_41[29]},
      {stage1_43[4],stage1_42[9],stage1_41[36],stage1_40[97],stage1_39[122]}
   );
   gpc615_5 gpc1489 (
      {stage0_39[192], stage0_39[193], stage0_39[194], stage0_39[195], stage0_39[196]},
      {stage0_40[35]},
      {stage0_41[30], stage0_41[31], stage0_41[32], stage0_41[33], stage0_41[34], stage0_41[35]},
      {stage1_43[5],stage1_42[10],stage1_41[37],stage1_40[98],stage1_39[123]}
   );
   gpc615_5 gpc1490 (
      {stage0_39[197], stage0_39[198], stage0_39[199], stage0_39[200], stage0_39[201]},
      {stage0_40[36]},
      {stage0_41[36], stage0_41[37], stage0_41[38], stage0_41[39], stage0_41[40], stage0_41[41]},
      {stage1_43[6],stage1_42[11],stage1_41[38],stage1_40[99],stage1_39[124]}
   );
   gpc615_5 gpc1491 (
      {stage0_39[202], stage0_39[203], stage0_39[204], stage0_39[205], stage0_39[206]},
      {stage0_40[37]},
      {stage0_41[42], stage0_41[43], stage0_41[44], stage0_41[45], stage0_41[46], stage0_41[47]},
      {stage1_43[7],stage1_42[12],stage1_41[39],stage1_40[100],stage1_39[125]}
   );
   gpc615_5 gpc1492 (
      {stage0_39[207], stage0_39[208], stage0_39[209], stage0_39[210], stage0_39[211]},
      {stage0_40[38]},
      {stage0_41[48], stage0_41[49], stage0_41[50], stage0_41[51], stage0_41[52], stage0_41[53]},
      {stage1_43[8],stage1_42[13],stage1_41[40],stage1_40[101],stage1_39[126]}
   );
   gpc615_5 gpc1493 (
      {stage0_39[212], stage0_39[213], stage0_39[214], stage0_39[215], stage0_39[216]},
      {stage0_40[39]},
      {stage0_41[54], stage0_41[55], stage0_41[56], stage0_41[57], stage0_41[58], stage0_41[59]},
      {stage1_43[9],stage1_42[14],stage1_41[41],stage1_40[102],stage1_39[127]}
   );
   gpc615_5 gpc1494 (
      {stage0_39[217], stage0_39[218], stage0_39[219], stage0_39[220], stage0_39[221]},
      {stage0_40[40]},
      {stage0_41[60], stage0_41[61], stage0_41[62], stage0_41[63], stage0_41[64], stage0_41[65]},
      {stage1_43[10],stage1_42[15],stage1_41[42],stage1_40[103],stage1_39[128]}
   );
   gpc615_5 gpc1495 (
      {stage0_39[222], stage0_39[223], stage0_39[224], stage0_39[225], stage0_39[226]},
      {stage0_40[41]},
      {stage0_41[66], stage0_41[67], stage0_41[68], stage0_41[69], stage0_41[70], stage0_41[71]},
      {stage1_43[11],stage1_42[16],stage1_41[43],stage1_40[104],stage1_39[129]}
   );
   gpc615_5 gpc1496 (
      {stage0_39[227], stage0_39[228], stage0_39[229], stage0_39[230], stage0_39[231]},
      {stage0_40[42]},
      {stage0_41[72], stage0_41[73], stage0_41[74], stage0_41[75], stage0_41[76], stage0_41[77]},
      {stage1_43[12],stage1_42[17],stage1_41[44],stage1_40[105],stage1_39[130]}
   );
   gpc615_5 gpc1497 (
      {stage0_39[232], stage0_39[233], stage0_39[234], stage0_39[235], stage0_39[236]},
      {stage0_40[43]},
      {stage0_41[78], stage0_41[79], stage0_41[80], stage0_41[81], stage0_41[82], stage0_41[83]},
      {stage1_43[13],stage1_42[18],stage1_41[45],stage1_40[106],stage1_39[131]}
   );
   gpc615_5 gpc1498 (
      {stage0_39[237], stage0_39[238], stage0_39[239], stage0_39[240], stage0_39[241]},
      {stage0_40[44]},
      {stage0_41[84], stage0_41[85], stage0_41[86], stage0_41[87], stage0_41[88], stage0_41[89]},
      {stage1_43[14],stage1_42[19],stage1_41[46],stage1_40[107],stage1_39[132]}
   );
   gpc615_5 gpc1499 (
      {stage0_39[242], stage0_39[243], stage0_39[244], stage0_39[245], stage0_39[246]},
      {stage0_40[45]},
      {stage0_41[90], stage0_41[91], stage0_41[92], stage0_41[93], stage0_41[94], stage0_41[95]},
      {stage1_43[15],stage1_42[20],stage1_41[47],stage1_40[108],stage1_39[133]}
   );
   gpc615_5 gpc1500 (
      {stage0_39[247], stage0_39[248], stage0_39[249], stage0_39[250], stage0_39[251]},
      {stage0_40[46]},
      {stage0_41[96], stage0_41[97], stage0_41[98], stage0_41[99], stage0_41[100], stage0_41[101]},
      {stage1_43[16],stage1_42[21],stage1_41[48],stage1_40[109],stage1_39[134]}
   );
   gpc615_5 gpc1501 (
      {stage0_39[252], stage0_39[253], stage0_39[254], stage0_39[255], stage0_39[256]},
      {stage0_40[47]},
      {stage0_41[102], stage0_41[103], stage0_41[104], stage0_41[105], stage0_41[106], stage0_41[107]},
      {stage1_43[17],stage1_42[22],stage1_41[49],stage1_40[110],stage1_39[135]}
   );
   gpc615_5 gpc1502 (
      {stage0_39[257], stage0_39[258], stage0_39[259], stage0_39[260], stage0_39[261]},
      {stage0_40[48]},
      {stage0_41[108], stage0_41[109], stage0_41[110], stage0_41[111], stage0_41[112], stage0_41[113]},
      {stage1_43[18],stage1_42[23],stage1_41[50],stage1_40[111],stage1_39[136]}
   );
   gpc615_5 gpc1503 (
      {stage0_39[262], stage0_39[263], stage0_39[264], stage0_39[265], stage0_39[266]},
      {stage0_40[49]},
      {stage0_41[114], stage0_41[115], stage0_41[116], stage0_41[117], stage0_41[118], stage0_41[119]},
      {stage1_43[19],stage1_42[24],stage1_41[51],stage1_40[112],stage1_39[137]}
   );
   gpc615_5 gpc1504 (
      {stage0_39[267], stage0_39[268], stage0_39[269], stage0_39[270], stage0_39[271]},
      {stage0_40[50]},
      {stage0_41[120], stage0_41[121], stage0_41[122], stage0_41[123], stage0_41[124], stage0_41[125]},
      {stage1_43[20],stage1_42[25],stage1_41[52],stage1_40[113],stage1_39[138]}
   );
   gpc615_5 gpc1505 (
      {stage0_39[272], stage0_39[273], stage0_39[274], stage0_39[275], stage0_39[276]},
      {stage0_40[51]},
      {stage0_41[126], stage0_41[127], stage0_41[128], stage0_41[129], stage0_41[130], stage0_41[131]},
      {stage1_43[21],stage1_42[26],stage1_41[53],stage1_40[114],stage1_39[139]}
   );
   gpc615_5 gpc1506 (
      {stage0_39[277], stage0_39[278], stage0_39[279], stage0_39[280], stage0_39[281]},
      {stage0_40[52]},
      {stage0_41[132], stage0_41[133], stage0_41[134], stage0_41[135], stage0_41[136], stage0_41[137]},
      {stage1_43[22],stage1_42[27],stage1_41[54],stage1_40[115],stage1_39[140]}
   );
   gpc615_5 gpc1507 (
      {stage0_39[282], stage0_39[283], stage0_39[284], stage0_39[285], stage0_39[286]},
      {stage0_40[53]},
      {stage0_41[138], stage0_41[139], stage0_41[140], stage0_41[141], stage0_41[142], stage0_41[143]},
      {stage1_43[23],stage1_42[28],stage1_41[55],stage1_40[116],stage1_39[141]}
   );
   gpc615_5 gpc1508 (
      {stage0_39[287], stage0_39[288], stage0_39[289], stage0_39[290], stage0_39[291]},
      {stage0_40[54]},
      {stage0_41[144], stage0_41[145], stage0_41[146], stage0_41[147], stage0_41[148], stage0_41[149]},
      {stage1_43[24],stage1_42[29],stage1_41[56],stage1_40[117],stage1_39[142]}
   );
   gpc615_5 gpc1509 (
      {stage0_39[292], stage0_39[293], stage0_39[294], stage0_39[295], stage0_39[296]},
      {stage0_40[55]},
      {stage0_41[150], stage0_41[151], stage0_41[152], stage0_41[153], stage0_41[154], stage0_41[155]},
      {stage1_43[25],stage1_42[30],stage1_41[57],stage1_40[118],stage1_39[143]}
   );
   gpc615_5 gpc1510 (
      {stage0_39[297], stage0_39[298], stage0_39[299], stage0_39[300], stage0_39[301]},
      {stage0_40[56]},
      {stage0_41[156], stage0_41[157], stage0_41[158], stage0_41[159], stage0_41[160], stage0_41[161]},
      {stage1_43[26],stage1_42[31],stage1_41[58],stage1_40[119],stage1_39[144]}
   );
   gpc615_5 gpc1511 (
      {stage0_39[302], stage0_39[303], stage0_39[304], stage0_39[305], stage0_39[306]},
      {stage0_40[57]},
      {stage0_41[162], stage0_41[163], stage0_41[164], stage0_41[165], stage0_41[166], stage0_41[167]},
      {stage1_43[27],stage1_42[32],stage1_41[59],stage1_40[120],stage1_39[145]}
   );
   gpc615_5 gpc1512 (
      {stage0_39[307], stage0_39[308], stage0_39[309], stage0_39[310], stage0_39[311]},
      {stage0_40[58]},
      {stage0_41[168], stage0_41[169], stage0_41[170], stage0_41[171], stage0_41[172], stage0_41[173]},
      {stage1_43[28],stage1_42[33],stage1_41[60],stage1_40[121],stage1_39[146]}
   );
   gpc615_5 gpc1513 (
      {stage0_39[312], stage0_39[313], stage0_39[314], stage0_39[315], stage0_39[316]},
      {stage0_40[59]},
      {stage0_41[174], stage0_41[175], stage0_41[176], stage0_41[177], stage0_41[178], stage0_41[179]},
      {stage1_43[29],stage1_42[34],stage1_41[61],stage1_40[122],stage1_39[147]}
   );
   gpc615_5 gpc1514 (
      {stage0_39[317], stage0_39[318], stage0_39[319], stage0_39[320], stage0_39[321]},
      {stage0_40[60]},
      {stage0_41[180], stage0_41[181], stage0_41[182], stage0_41[183], stage0_41[184], stage0_41[185]},
      {stage1_43[30],stage1_42[35],stage1_41[62],stage1_40[123],stage1_39[148]}
   );
   gpc615_5 gpc1515 (
      {stage0_39[322], stage0_39[323], stage0_39[324], stage0_39[325], stage0_39[326]},
      {stage0_40[61]},
      {stage0_41[186], stage0_41[187], stage0_41[188], stage0_41[189], stage0_41[190], stage0_41[191]},
      {stage1_43[31],stage1_42[36],stage1_41[63],stage1_40[124],stage1_39[149]}
   );
   gpc615_5 gpc1516 (
      {stage0_39[327], stage0_39[328], stage0_39[329], stage0_39[330], stage0_39[331]},
      {stage0_40[62]},
      {stage0_41[192], stage0_41[193], stage0_41[194], stage0_41[195], stage0_41[196], stage0_41[197]},
      {stage1_43[32],stage1_42[37],stage1_41[64],stage1_40[125],stage1_39[150]}
   );
   gpc615_5 gpc1517 (
      {stage0_39[332], stage0_39[333], stage0_39[334], stage0_39[335], stage0_39[336]},
      {stage0_40[63]},
      {stage0_41[198], stage0_41[199], stage0_41[200], stage0_41[201], stage0_41[202], stage0_41[203]},
      {stage1_43[33],stage1_42[38],stage1_41[65],stage1_40[126],stage1_39[151]}
   );
   gpc615_5 gpc1518 (
      {stage0_39[337], stage0_39[338], stage0_39[339], stage0_39[340], stage0_39[341]},
      {stage0_40[64]},
      {stage0_41[204], stage0_41[205], stage0_41[206], stage0_41[207], stage0_41[208], stage0_41[209]},
      {stage1_43[34],stage1_42[39],stage1_41[66],stage1_40[127],stage1_39[152]}
   );
   gpc615_5 gpc1519 (
      {stage0_39[342], stage0_39[343], stage0_39[344], stage0_39[345], stage0_39[346]},
      {stage0_40[65]},
      {stage0_41[210], stage0_41[211], stage0_41[212], stage0_41[213], stage0_41[214], stage0_41[215]},
      {stage1_43[35],stage1_42[40],stage1_41[67],stage1_40[128],stage1_39[153]}
   );
   gpc615_5 gpc1520 (
      {stage0_39[347], stage0_39[348], stage0_39[349], stage0_39[350], stage0_39[351]},
      {stage0_40[66]},
      {stage0_41[216], stage0_41[217], stage0_41[218], stage0_41[219], stage0_41[220], stage0_41[221]},
      {stage1_43[36],stage1_42[41],stage1_41[68],stage1_40[129],stage1_39[154]}
   );
   gpc615_5 gpc1521 (
      {stage0_39[352], stage0_39[353], stage0_39[354], stage0_39[355], stage0_39[356]},
      {stage0_40[67]},
      {stage0_41[222], stage0_41[223], stage0_41[224], stage0_41[225], stage0_41[226], stage0_41[227]},
      {stage1_43[37],stage1_42[42],stage1_41[69],stage1_40[130],stage1_39[155]}
   );
   gpc615_5 gpc1522 (
      {stage0_39[357], stage0_39[358], stage0_39[359], stage0_39[360], stage0_39[361]},
      {stage0_40[68]},
      {stage0_41[228], stage0_41[229], stage0_41[230], stage0_41[231], stage0_41[232], stage0_41[233]},
      {stage1_43[38],stage1_42[43],stage1_41[70],stage1_40[131],stage1_39[156]}
   );
   gpc615_5 gpc1523 (
      {stage0_39[362], stage0_39[363], stage0_39[364], stage0_39[365], stage0_39[366]},
      {stage0_40[69]},
      {stage0_41[234], stage0_41[235], stage0_41[236], stage0_41[237], stage0_41[238], stage0_41[239]},
      {stage1_43[39],stage1_42[44],stage1_41[71],stage1_40[132],stage1_39[157]}
   );
   gpc615_5 gpc1524 (
      {stage0_39[367], stage0_39[368], stage0_39[369], stage0_39[370], stage0_39[371]},
      {stage0_40[70]},
      {stage0_41[240], stage0_41[241], stage0_41[242], stage0_41[243], stage0_41[244], stage0_41[245]},
      {stage1_43[40],stage1_42[45],stage1_41[72],stage1_40[133],stage1_39[158]}
   );
   gpc615_5 gpc1525 (
      {stage0_39[372], stage0_39[373], stage0_39[374], stage0_39[375], stage0_39[376]},
      {stage0_40[71]},
      {stage0_41[246], stage0_41[247], stage0_41[248], stage0_41[249], stage0_41[250], stage0_41[251]},
      {stage1_43[41],stage1_42[46],stage1_41[73],stage1_40[134],stage1_39[159]}
   );
   gpc615_5 gpc1526 (
      {stage0_39[377], stage0_39[378], stage0_39[379], stage0_39[380], stage0_39[381]},
      {stage0_40[72]},
      {stage0_41[252], stage0_41[253], stage0_41[254], stage0_41[255], stage0_41[256], stage0_41[257]},
      {stage1_43[42],stage1_42[47],stage1_41[74],stage1_40[135],stage1_39[160]}
   );
   gpc615_5 gpc1527 (
      {stage0_39[382], stage0_39[383], stage0_39[384], stage0_39[385], stage0_39[386]},
      {stage0_40[73]},
      {stage0_41[258], stage0_41[259], stage0_41[260], stage0_41[261], stage0_41[262], stage0_41[263]},
      {stage1_43[43],stage1_42[48],stage1_41[75],stage1_40[136],stage1_39[161]}
   );
   gpc615_5 gpc1528 (
      {stage0_39[387], stage0_39[388], stage0_39[389], stage0_39[390], stage0_39[391]},
      {stage0_40[74]},
      {stage0_41[264], stage0_41[265], stage0_41[266], stage0_41[267], stage0_41[268], stage0_41[269]},
      {stage1_43[44],stage1_42[49],stage1_41[76],stage1_40[137],stage1_39[162]}
   );
   gpc615_5 gpc1529 (
      {stage0_39[392], stage0_39[393], stage0_39[394], stage0_39[395], stage0_39[396]},
      {stage0_40[75]},
      {stage0_41[270], stage0_41[271], stage0_41[272], stage0_41[273], stage0_41[274], stage0_41[275]},
      {stage1_43[45],stage1_42[50],stage1_41[77],stage1_40[138],stage1_39[163]}
   );
   gpc615_5 gpc1530 (
      {stage0_39[397], stage0_39[398], stage0_39[399], stage0_39[400], stage0_39[401]},
      {stage0_40[76]},
      {stage0_41[276], stage0_41[277], stage0_41[278], stage0_41[279], stage0_41[280], stage0_41[281]},
      {stage1_43[46],stage1_42[51],stage1_41[78],stage1_40[139],stage1_39[164]}
   );
   gpc615_5 gpc1531 (
      {stage0_39[402], stage0_39[403], stage0_39[404], stage0_39[405], stage0_39[406]},
      {stage0_40[77]},
      {stage0_41[282], stage0_41[283], stage0_41[284], stage0_41[285], stage0_41[286], stage0_41[287]},
      {stage1_43[47],stage1_42[52],stage1_41[79],stage1_40[140],stage1_39[165]}
   );
   gpc615_5 gpc1532 (
      {stage0_39[407], stage0_39[408], stage0_39[409], stage0_39[410], stage0_39[411]},
      {stage0_40[78]},
      {stage0_41[288], stage0_41[289], stage0_41[290], stage0_41[291], stage0_41[292], stage0_41[293]},
      {stage1_43[48],stage1_42[53],stage1_41[80],stage1_40[141],stage1_39[166]}
   );
   gpc615_5 gpc1533 (
      {stage0_39[412], stage0_39[413], stage0_39[414], stage0_39[415], stage0_39[416]},
      {stage0_40[79]},
      {stage0_41[294], stage0_41[295], stage0_41[296], stage0_41[297], stage0_41[298], stage0_41[299]},
      {stage1_43[49],stage1_42[54],stage1_41[81],stage1_40[142],stage1_39[167]}
   );
   gpc615_5 gpc1534 (
      {stage0_39[417], stage0_39[418], stage0_39[419], stage0_39[420], stage0_39[421]},
      {stage0_40[80]},
      {stage0_41[300], stage0_41[301], stage0_41[302], stage0_41[303], stage0_41[304], stage0_41[305]},
      {stage1_43[50],stage1_42[55],stage1_41[82],stage1_40[143],stage1_39[168]}
   );
   gpc615_5 gpc1535 (
      {stage0_39[422], stage0_39[423], stage0_39[424], stage0_39[425], stage0_39[426]},
      {stage0_40[81]},
      {stage0_41[306], stage0_41[307], stage0_41[308], stage0_41[309], stage0_41[310], stage0_41[311]},
      {stage1_43[51],stage1_42[56],stage1_41[83],stage1_40[144],stage1_39[169]}
   );
   gpc615_5 gpc1536 (
      {stage0_39[427], stage0_39[428], stage0_39[429], stage0_39[430], stage0_39[431]},
      {stage0_40[82]},
      {stage0_41[312], stage0_41[313], stage0_41[314], stage0_41[315], stage0_41[316], stage0_41[317]},
      {stage1_43[52],stage1_42[57],stage1_41[84],stage1_40[145],stage1_39[170]}
   );
   gpc615_5 gpc1537 (
      {stage0_39[432], stage0_39[433], stage0_39[434], stage0_39[435], stage0_39[436]},
      {stage0_40[83]},
      {stage0_41[318], stage0_41[319], stage0_41[320], stage0_41[321], stage0_41[322], stage0_41[323]},
      {stage1_43[53],stage1_42[58],stage1_41[85],stage1_40[146],stage1_39[171]}
   );
   gpc615_5 gpc1538 (
      {stage0_39[437], stage0_39[438], stage0_39[439], stage0_39[440], stage0_39[441]},
      {stage0_40[84]},
      {stage0_41[324], stage0_41[325], stage0_41[326], stage0_41[327], stage0_41[328], stage0_41[329]},
      {stage1_43[54],stage1_42[59],stage1_41[86],stage1_40[147],stage1_39[172]}
   );
   gpc615_5 gpc1539 (
      {stage0_39[442], stage0_39[443], stage0_39[444], stage0_39[445], stage0_39[446]},
      {stage0_40[85]},
      {stage0_41[330], stage0_41[331], stage0_41[332], stage0_41[333], stage0_41[334], stage0_41[335]},
      {stage1_43[55],stage1_42[60],stage1_41[87],stage1_40[148],stage1_39[173]}
   );
   gpc606_5 gpc1540 (
      {stage0_40[86], stage0_40[87], stage0_40[88], stage0_40[89], stage0_40[90], stage0_40[91]},
      {stage0_42[0], stage0_42[1], stage0_42[2], stage0_42[3], stage0_42[4], stage0_42[5]},
      {stage1_44[0],stage1_43[56],stage1_42[61],stage1_41[88],stage1_40[149]}
   );
   gpc606_5 gpc1541 (
      {stage0_40[92], stage0_40[93], stage0_40[94], stage0_40[95], stage0_40[96], stage0_40[97]},
      {stage0_42[6], stage0_42[7], stage0_42[8], stage0_42[9], stage0_42[10], stage0_42[11]},
      {stage1_44[1],stage1_43[57],stage1_42[62],stage1_41[89],stage1_40[150]}
   );
   gpc606_5 gpc1542 (
      {stage0_40[98], stage0_40[99], stage0_40[100], stage0_40[101], stage0_40[102], stage0_40[103]},
      {stage0_42[12], stage0_42[13], stage0_42[14], stage0_42[15], stage0_42[16], stage0_42[17]},
      {stage1_44[2],stage1_43[58],stage1_42[63],stage1_41[90],stage1_40[151]}
   );
   gpc606_5 gpc1543 (
      {stage0_40[104], stage0_40[105], stage0_40[106], stage0_40[107], stage0_40[108], stage0_40[109]},
      {stage0_42[18], stage0_42[19], stage0_42[20], stage0_42[21], stage0_42[22], stage0_42[23]},
      {stage1_44[3],stage1_43[59],stage1_42[64],stage1_41[91],stage1_40[152]}
   );
   gpc606_5 gpc1544 (
      {stage0_40[110], stage0_40[111], stage0_40[112], stage0_40[113], stage0_40[114], stage0_40[115]},
      {stage0_42[24], stage0_42[25], stage0_42[26], stage0_42[27], stage0_42[28], stage0_42[29]},
      {stage1_44[4],stage1_43[60],stage1_42[65],stage1_41[92],stage1_40[153]}
   );
   gpc606_5 gpc1545 (
      {stage0_40[116], stage0_40[117], stage0_40[118], stage0_40[119], stage0_40[120], stage0_40[121]},
      {stage0_42[30], stage0_42[31], stage0_42[32], stage0_42[33], stage0_42[34], stage0_42[35]},
      {stage1_44[5],stage1_43[61],stage1_42[66],stage1_41[93],stage1_40[154]}
   );
   gpc606_5 gpc1546 (
      {stage0_40[122], stage0_40[123], stage0_40[124], stage0_40[125], stage0_40[126], stage0_40[127]},
      {stage0_42[36], stage0_42[37], stage0_42[38], stage0_42[39], stage0_42[40], stage0_42[41]},
      {stage1_44[6],stage1_43[62],stage1_42[67],stage1_41[94],stage1_40[155]}
   );
   gpc606_5 gpc1547 (
      {stage0_40[128], stage0_40[129], stage0_40[130], stage0_40[131], stage0_40[132], stage0_40[133]},
      {stage0_42[42], stage0_42[43], stage0_42[44], stage0_42[45], stage0_42[46], stage0_42[47]},
      {stage1_44[7],stage1_43[63],stage1_42[68],stage1_41[95],stage1_40[156]}
   );
   gpc606_5 gpc1548 (
      {stage0_40[134], stage0_40[135], stage0_40[136], stage0_40[137], stage0_40[138], stage0_40[139]},
      {stage0_42[48], stage0_42[49], stage0_42[50], stage0_42[51], stage0_42[52], stage0_42[53]},
      {stage1_44[8],stage1_43[64],stage1_42[69],stage1_41[96],stage1_40[157]}
   );
   gpc606_5 gpc1549 (
      {stage0_40[140], stage0_40[141], stage0_40[142], stage0_40[143], stage0_40[144], stage0_40[145]},
      {stage0_42[54], stage0_42[55], stage0_42[56], stage0_42[57], stage0_42[58], stage0_42[59]},
      {stage1_44[9],stage1_43[65],stage1_42[70],stage1_41[97],stage1_40[158]}
   );
   gpc606_5 gpc1550 (
      {stage0_40[146], stage0_40[147], stage0_40[148], stage0_40[149], stage0_40[150], stage0_40[151]},
      {stage0_42[60], stage0_42[61], stage0_42[62], stage0_42[63], stage0_42[64], stage0_42[65]},
      {stage1_44[10],stage1_43[66],stage1_42[71],stage1_41[98],stage1_40[159]}
   );
   gpc606_5 gpc1551 (
      {stage0_40[152], stage0_40[153], stage0_40[154], stage0_40[155], stage0_40[156], stage0_40[157]},
      {stage0_42[66], stage0_42[67], stage0_42[68], stage0_42[69], stage0_42[70], stage0_42[71]},
      {stage1_44[11],stage1_43[67],stage1_42[72],stage1_41[99],stage1_40[160]}
   );
   gpc606_5 gpc1552 (
      {stage0_40[158], stage0_40[159], stage0_40[160], stage0_40[161], stage0_40[162], stage0_40[163]},
      {stage0_42[72], stage0_42[73], stage0_42[74], stage0_42[75], stage0_42[76], stage0_42[77]},
      {stage1_44[12],stage1_43[68],stage1_42[73],stage1_41[100],stage1_40[161]}
   );
   gpc606_5 gpc1553 (
      {stage0_40[164], stage0_40[165], stage0_40[166], stage0_40[167], stage0_40[168], stage0_40[169]},
      {stage0_42[78], stage0_42[79], stage0_42[80], stage0_42[81], stage0_42[82], stage0_42[83]},
      {stage1_44[13],stage1_43[69],stage1_42[74],stage1_41[101],stage1_40[162]}
   );
   gpc606_5 gpc1554 (
      {stage0_40[170], stage0_40[171], stage0_40[172], stage0_40[173], stage0_40[174], stage0_40[175]},
      {stage0_42[84], stage0_42[85], stage0_42[86], stage0_42[87], stage0_42[88], stage0_42[89]},
      {stage1_44[14],stage1_43[70],stage1_42[75],stage1_41[102],stage1_40[163]}
   );
   gpc606_5 gpc1555 (
      {stage0_40[176], stage0_40[177], stage0_40[178], stage0_40[179], stage0_40[180], stage0_40[181]},
      {stage0_42[90], stage0_42[91], stage0_42[92], stage0_42[93], stage0_42[94], stage0_42[95]},
      {stage1_44[15],stage1_43[71],stage1_42[76],stage1_41[103],stage1_40[164]}
   );
   gpc606_5 gpc1556 (
      {stage0_40[182], stage0_40[183], stage0_40[184], stage0_40[185], stage0_40[186], stage0_40[187]},
      {stage0_42[96], stage0_42[97], stage0_42[98], stage0_42[99], stage0_42[100], stage0_42[101]},
      {stage1_44[16],stage1_43[72],stage1_42[77],stage1_41[104],stage1_40[165]}
   );
   gpc606_5 gpc1557 (
      {stage0_40[188], stage0_40[189], stage0_40[190], stage0_40[191], stage0_40[192], stage0_40[193]},
      {stage0_42[102], stage0_42[103], stage0_42[104], stage0_42[105], stage0_42[106], stage0_42[107]},
      {stage1_44[17],stage1_43[73],stage1_42[78],stage1_41[105],stage1_40[166]}
   );
   gpc606_5 gpc1558 (
      {stage0_40[194], stage0_40[195], stage0_40[196], stage0_40[197], stage0_40[198], stage0_40[199]},
      {stage0_42[108], stage0_42[109], stage0_42[110], stage0_42[111], stage0_42[112], stage0_42[113]},
      {stage1_44[18],stage1_43[74],stage1_42[79],stage1_41[106],stage1_40[167]}
   );
   gpc606_5 gpc1559 (
      {stage0_40[200], stage0_40[201], stage0_40[202], stage0_40[203], stage0_40[204], stage0_40[205]},
      {stage0_42[114], stage0_42[115], stage0_42[116], stage0_42[117], stage0_42[118], stage0_42[119]},
      {stage1_44[19],stage1_43[75],stage1_42[80],stage1_41[107],stage1_40[168]}
   );
   gpc606_5 gpc1560 (
      {stage0_40[206], stage0_40[207], stage0_40[208], stage0_40[209], stage0_40[210], stage0_40[211]},
      {stage0_42[120], stage0_42[121], stage0_42[122], stage0_42[123], stage0_42[124], stage0_42[125]},
      {stage1_44[20],stage1_43[76],stage1_42[81],stage1_41[108],stage1_40[169]}
   );
   gpc606_5 gpc1561 (
      {stage0_40[212], stage0_40[213], stage0_40[214], stage0_40[215], stage0_40[216], stage0_40[217]},
      {stage0_42[126], stage0_42[127], stage0_42[128], stage0_42[129], stage0_42[130], stage0_42[131]},
      {stage1_44[21],stage1_43[77],stage1_42[82],stage1_41[109],stage1_40[170]}
   );
   gpc606_5 gpc1562 (
      {stage0_40[218], stage0_40[219], stage0_40[220], stage0_40[221], stage0_40[222], stage0_40[223]},
      {stage0_42[132], stage0_42[133], stage0_42[134], stage0_42[135], stage0_42[136], stage0_42[137]},
      {stage1_44[22],stage1_43[78],stage1_42[83],stage1_41[110],stage1_40[171]}
   );
   gpc606_5 gpc1563 (
      {stage0_40[224], stage0_40[225], stage0_40[226], stage0_40[227], stage0_40[228], stage0_40[229]},
      {stage0_42[138], stage0_42[139], stage0_42[140], stage0_42[141], stage0_42[142], stage0_42[143]},
      {stage1_44[23],stage1_43[79],stage1_42[84],stage1_41[111],stage1_40[172]}
   );
   gpc606_5 gpc1564 (
      {stage0_40[230], stage0_40[231], stage0_40[232], stage0_40[233], stage0_40[234], stage0_40[235]},
      {stage0_42[144], stage0_42[145], stage0_42[146], stage0_42[147], stage0_42[148], stage0_42[149]},
      {stage1_44[24],stage1_43[80],stage1_42[85],stage1_41[112],stage1_40[173]}
   );
   gpc606_5 gpc1565 (
      {stage0_40[236], stage0_40[237], stage0_40[238], stage0_40[239], stage0_40[240], stage0_40[241]},
      {stage0_42[150], stage0_42[151], stage0_42[152], stage0_42[153], stage0_42[154], stage0_42[155]},
      {stage1_44[25],stage1_43[81],stage1_42[86],stage1_41[113],stage1_40[174]}
   );
   gpc606_5 gpc1566 (
      {stage0_40[242], stage0_40[243], stage0_40[244], stage0_40[245], stage0_40[246], stage0_40[247]},
      {stage0_42[156], stage0_42[157], stage0_42[158], stage0_42[159], stage0_42[160], stage0_42[161]},
      {stage1_44[26],stage1_43[82],stage1_42[87],stage1_41[114],stage1_40[175]}
   );
   gpc606_5 gpc1567 (
      {stage0_40[248], stage0_40[249], stage0_40[250], stage0_40[251], stage0_40[252], stage0_40[253]},
      {stage0_42[162], stage0_42[163], stage0_42[164], stage0_42[165], stage0_42[166], stage0_42[167]},
      {stage1_44[27],stage1_43[83],stage1_42[88],stage1_41[115],stage1_40[176]}
   );
   gpc606_5 gpc1568 (
      {stage0_40[254], stage0_40[255], stage0_40[256], stage0_40[257], stage0_40[258], stage0_40[259]},
      {stage0_42[168], stage0_42[169], stage0_42[170], stage0_42[171], stage0_42[172], stage0_42[173]},
      {stage1_44[28],stage1_43[84],stage1_42[89],stage1_41[116],stage1_40[177]}
   );
   gpc606_5 gpc1569 (
      {stage0_40[260], stage0_40[261], stage0_40[262], stage0_40[263], stage0_40[264], stage0_40[265]},
      {stage0_42[174], stage0_42[175], stage0_42[176], stage0_42[177], stage0_42[178], stage0_42[179]},
      {stage1_44[29],stage1_43[85],stage1_42[90],stage1_41[117],stage1_40[178]}
   );
   gpc606_5 gpc1570 (
      {stage0_40[266], stage0_40[267], stage0_40[268], stage0_40[269], stage0_40[270], stage0_40[271]},
      {stage0_42[180], stage0_42[181], stage0_42[182], stage0_42[183], stage0_42[184], stage0_42[185]},
      {stage1_44[30],stage1_43[86],stage1_42[91],stage1_41[118],stage1_40[179]}
   );
   gpc606_5 gpc1571 (
      {stage0_40[272], stage0_40[273], stage0_40[274], stage0_40[275], stage0_40[276], stage0_40[277]},
      {stage0_42[186], stage0_42[187], stage0_42[188], stage0_42[189], stage0_42[190], stage0_42[191]},
      {stage1_44[31],stage1_43[87],stage1_42[92],stage1_41[119],stage1_40[180]}
   );
   gpc606_5 gpc1572 (
      {stage0_40[278], stage0_40[279], stage0_40[280], stage0_40[281], stage0_40[282], stage0_40[283]},
      {stage0_42[192], stage0_42[193], stage0_42[194], stage0_42[195], stage0_42[196], stage0_42[197]},
      {stage1_44[32],stage1_43[88],stage1_42[93],stage1_41[120],stage1_40[181]}
   );
   gpc606_5 gpc1573 (
      {stage0_40[284], stage0_40[285], stage0_40[286], stage0_40[287], stage0_40[288], stage0_40[289]},
      {stage0_42[198], stage0_42[199], stage0_42[200], stage0_42[201], stage0_42[202], stage0_42[203]},
      {stage1_44[33],stage1_43[89],stage1_42[94],stage1_41[121],stage1_40[182]}
   );
   gpc606_5 gpc1574 (
      {stage0_40[290], stage0_40[291], stage0_40[292], stage0_40[293], stage0_40[294], stage0_40[295]},
      {stage0_42[204], stage0_42[205], stage0_42[206], stage0_42[207], stage0_42[208], stage0_42[209]},
      {stage1_44[34],stage1_43[90],stage1_42[95],stage1_41[122],stage1_40[183]}
   );
   gpc606_5 gpc1575 (
      {stage0_40[296], stage0_40[297], stage0_40[298], stage0_40[299], stage0_40[300], stage0_40[301]},
      {stage0_42[210], stage0_42[211], stage0_42[212], stage0_42[213], stage0_42[214], stage0_42[215]},
      {stage1_44[35],stage1_43[91],stage1_42[96],stage1_41[123],stage1_40[184]}
   );
   gpc606_5 gpc1576 (
      {stage0_40[302], stage0_40[303], stage0_40[304], stage0_40[305], stage0_40[306], stage0_40[307]},
      {stage0_42[216], stage0_42[217], stage0_42[218], stage0_42[219], stage0_42[220], stage0_42[221]},
      {stage1_44[36],stage1_43[92],stage1_42[97],stage1_41[124],stage1_40[185]}
   );
   gpc606_5 gpc1577 (
      {stage0_40[308], stage0_40[309], stage0_40[310], stage0_40[311], stage0_40[312], stage0_40[313]},
      {stage0_42[222], stage0_42[223], stage0_42[224], stage0_42[225], stage0_42[226], stage0_42[227]},
      {stage1_44[37],stage1_43[93],stage1_42[98],stage1_41[125],stage1_40[186]}
   );
   gpc606_5 gpc1578 (
      {stage0_40[314], stage0_40[315], stage0_40[316], stage0_40[317], stage0_40[318], stage0_40[319]},
      {stage0_42[228], stage0_42[229], stage0_42[230], stage0_42[231], stage0_42[232], stage0_42[233]},
      {stage1_44[38],stage1_43[94],stage1_42[99],stage1_41[126],stage1_40[187]}
   );
   gpc606_5 gpc1579 (
      {stage0_40[320], stage0_40[321], stage0_40[322], stage0_40[323], stage0_40[324], stage0_40[325]},
      {stage0_42[234], stage0_42[235], stage0_42[236], stage0_42[237], stage0_42[238], stage0_42[239]},
      {stage1_44[39],stage1_43[95],stage1_42[100],stage1_41[127],stage1_40[188]}
   );
   gpc606_5 gpc1580 (
      {stage0_40[326], stage0_40[327], stage0_40[328], stage0_40[329], stage0_40[330], stage0_40[331]},
      {stage0_42[240], stage0_42[241], stage0_42[242], stage0_42[243], stage0_42[244], stage0_42[245]},
      {stage1_44[40],stage1_43[96],stage1_42[101],stage1_41[128],stage1_40[189]}
   );
   gpc606_5 gpc1581 (
      {stage0_40[332], stage0_40[333], stage0_40[334], stage0_40[335], stage0_40[336], stage0_40[337]},
      {stage0_42[246], stage0_42[247], stage0_42[248], stage0_42[249], stage0_42[250], stage0_42[251]},
      {stage1_44[41],stage1_43[97],stage1_42[102],stage1_41[129],stage1_40[190]}
   );
   gpc606_5 gpc1582 (
      {stage0_40[338], stage0_40[339], stage0_40[340], stage0_40[341], stage0_40[342], stage0_40[343]},
      {stage0_42[252], stage0_42[253], stage0_42[254], stage0_42[255], stage0_42[256], stage0_42[257]},
      {stage1_44[42],stage1_43[98],stage1_42[103],stage1_41[130],stage1_40[191]}
   );
   gpc606_5 gpc1583 (
      {stage0_40[344], stage0_40[345], stage0_40[346], stage0_40[347], stage0_40[348], stage0_40[349]},
      {stage0_42[258], stage0_42[259], stage0_42[260], stage0_42[261], stage0_42[262], stage0_42[263]},
      {stage1_44[43],stage1_43[99],stage1_42[104],stage1_41[131],stage1_40[192]}
   );
   gpc606_5 gpc1584 (
      {stage0_40[350], stage0_40[351], stage0_40[352], stage0_40[353], stage0_40[354], stage0_40[355]},
      {stage0_42[264], stage0_42[265], stage0_42[266], stage0_42[267], stage0_42[268], stage0_42[269]},
      {stage1_44[44],stage1_43[100],stage1_42[105],stage1_41[132],stage1_40[193]}
   );
   gpc606_5 gpc1585 (
      {stage0_40[356], stage0_40[357], stage0_40[358], stage0_40[359], stage0_40[360], stage0_40[361]},
      {stage0_42[270], stage0_42[271], stage0_42[272], stage0_42[273], stage0_42[274], stage0_42[275]},
      {stage1_44[45],stage1_43[101],stage1_42[106],stage1_41[133],stage1_40[194]}
   );
   gpc606_5 gpc1586 (
      {stage0_40[362], stage0_40[363], stage0_40[364], stage0_40[365], stage0_40[366], stage0_40[367]},
      {stage0_42[276], stage0_42[277], stage0_42[278], stage0_42[279], stage0_42[280], stage0_42[281]},
      {stage1_44[46],stage1_43[102],stage1_42[107],stage1_41[134],stage1_40[195]}
   );
   gpc606_5 gpc1587 (
      {stage0_40[368], stage0_40[369], stage0_40[370], stage0_40[371], stage0_40[372], stage0_40[373]},
      {stage0_42[282], stage0_42[283], stage0_42[284], stage0_42[285], stage0_42[286], stage0_42[287]},
      {stage1_44[47],stage1_43[103],stage1_42[108],stage1_41[135],stage1_40[196]}
   );
   gpc606_5 gpc1588 (
      {stage0_40[374], stage0_40[375], stage0_40[376], stage0_40[377], stage0_40[378], stage0_40[379]},
      {stage0_42[288], stage0_42[289], stage0_42[290], stage0_42[291], stage0_42[292], stage0_42[293]},
      {stage1_44[48],stage1_43[104],stage1_42[109],stage1_41[136],stage1_40[197]}
   );
   gpc606_5 gpc1589 (
      {stage0_41[336], stage0_41[337], stage0_41[338], stage0_41[339], stage0_41[340], stage0_41[341]},
      {stage0_43[0], stage0_43[1], stage0_43[2], stage0_43[3], stage0_43[4], stage0_43[5]},
      {stage1_45[0],stage1_44[49],stage1_43[105],stage1_42[110],stage1_41[137]}
   );
   gpc606_5 gpc1590 (
      {stage0_41[342], stage0_41[343], stage0_41[344], stage0_41[345], stage0_41[346], stage0_41[347]},
      {stage0_43[6], stage0_43[7], stage0_43[8], stage0_43[9], stage0_43[10], stage0_43[11]},
      {stage1_45[1],stage1_44[50],stage1_43[106],stage1_42[111],stage1_41[138]}
   );
   gpc606_5 gpc1591 (
      {stage0_41[348], stage0_41[349], stage0_41[350], stage0_41[351], stage0_41[352], stage0_41[353]},
      {stage0_43[12], stage0_43[13], stage0_43[14], stage0_43[15], stage0_43[16], stage0_43[17]},
      {stage1_45[2],stage1_44[51],stage1_43[107],stage1_42[112],stage1_41[139]}
   );
   gpc606_5 gpc1592 (
      {stage0_41[354], stage0_41[355], stage0_41[356], stage0_41[357], stage0_41[358], stage0_41[359]},
      {stage0_43[18], stage0_43[19], stage0_43[20], stage0_43[21], stage0_43[22], stage0_43[23]},
      {stage1_45[3],stage1_44[52],stage1_43[108],stage1_42[113],stage1_41[140]}
   );
   gpc606_5 gpc1593 (
      {stage0_41[360], stage0_41[361], stage0_41[362], stage0_41[363], stage0_41[364], stage0_41[365]},
      {stage0_43[24], stage0_43[25], stage0_43[26], stage0_43[27], stage0_43[28], stage0_43[29]},
      {stage1_45[4],stage1_44[53],stage1_43[109],stage1_42[114],stage1_41[141]}
   );
   gpc606_5 gpc1594 (
      {stage0_41[366], stage0_41[367], stage0_41[368], stage0_41[369], stage0_41[370], stage0_41[371]},
      {stage0_43[30], stage0_43[31], stage0_43[32], stage0_43[33], stage0_43[34], stage0_43[35]},
      {stage1_45[5],stage1_44[54],stage1_43[110],stage1_42[115],stage1_41[142]}
   );
   gpc606_5 gpc1595 (
      {stage0_41[372], stage0_41[373], stage0_41[374], stage0_41[375], stage0_41[376], stage0_41[377]},
      {stage0_43[36], stage0_43[37], stage0_43[38], stage0_43[39], stage0_43[40], stage0_43[41]},
      {stage1_45[6],stage1_44[55],stage1_43[111],stage1_42[116],stage1_41[143]}
   );
   gpc606_5 gpc1596 (
      {stage0_41[378], stage0_41[379], stage0_41[380], stage0_41[381], stage0_41[382], stage0_41[383]},
      {stage0_43[42], stage0_43[43], stage0_43[44], stage0_43[45], stage0_43[46], stage0_43[47]},
      {stage1_45[7],stage1_44[56],stage1_43[112],stage1_42[117],stage1_41[144]}
   );
   gpc606_5 gpc1597 (
      {stage0_41[384], stage0_41[385], stage0_41[386], stage0_41[387], stage0_41[388], stage0_41[389]},
      {stage0_43[48], stage0_43[49], stage0_43[50], stage0_43[51], stage0_43[52], stage0_43[53]},
      {stage1_45[8],stage1_44[57],stage1_43[113],stage1_42[118],stage1_41[145]}
   );
   gpc606_5 gpc1598 (
      {stage0_41[390], stage0_41[391], stage0_41[392], stage0_41[393], stage0_41[394], stage0_41[395]},
      {stage0_43[54], stage0_43[55], stage0_43[56], stage0_43[57], stage0_43[58], stage0_43[59]},
      {stage1_45[9],stage1_44[58],stage1_43[114],stage1_42[119],stage1_41[146]}
   );
   gpc606_5 gpc1599 (
      {stage0_41[396], stage0_41[397], stage0_41[398], stage0_41[399], stage0_41[400], stage0_41[401]},
      {stage0_43[60], stage0_43[61], stage0_43[62], stage0_43[63], stage0_43[64], stage0_43[65]},
      {stage1_45[10],stage1_44[59],stage1_43[115],stage1_42[120],stage1_41[147]}
   );
   gpc606_5 gpc1600 (
      {stage0_41[402], stage0_41[403], stage0_41[404], stage0_41[405], stage0_41[406], stage0_41[407]},
      {stage0_43[66], stage0_43[67], stage0_43[68], stage0_43[69], stage0_43[70], stage0_43[71]},
      {stage1_45[11],stage1_44[60],stage1_43[116],stage1_42[121],stage1_41[148]}
   );
   gpc606_5 gpc1601 (
      {stage0_41[408], stage0_41[409], stage0_41[410], stage0_41[411], stage0_41[412], stage0_41[413]},
      {stage0_43[72], stage0_43[73], stage0_43[74], stage0_43[75], stage0_43[76], stage0_43[77]},
      {stage1_45[12],stage1_44[61],stage1_43[117],stage1_42[122],stage1_41[149]}
   );
   gpc606_5 gpc1602 (
      {stage0_41[414], stage0_41[415], stage0_41[416], stage0_41[417], stage0_41[418], stage0_41[419]},
      {stage0_43[78], stage0_43[79], stage0_43[80], stage0_43[81], stage0_43[82], stage0_43[83]},
      {stage1_45[13],stage1_44[62],stage1_43[118],stage1_42[123],stage1_41[150]}
   );
   gpc606_5 gpc1603 (
      {stage0_41[420], stage0_41[421], stage0_41[422], stage0_41[423], stage0_41[424], stage0_41[425]},
      {stage0_43[84], stage0_43[85], stage0_43[86], stage0_43[87], stage0_43[88], stage0_43[89]},
      {stage1_45[14],stage1_44[63],stage1_43[119],stage1_42[124],stage1_41[151]}
   );
   gpc606_5 gpc1604 (
      {stage0_41[426], stage0_41[427], stage0_41[428], stage0_41[429], stage0_41[430], stage0_41[431]},
      {stage0_43[90], stage0_43[91], stage0_43[92], stage0_43[93], stage0_43[94], stage0_43[95]},
      {stage1_45[15],stage1_44[64],stage1_43[120],stage1_42[125],stage1_41[152]}
   );
   gpc615_5 gpc1605 (
      {stage0_41[432], stage0_41[433], stage0_41[434], stage0_41[435], stage0_41[436]},
      {stage0_42[294]},
      {stage0_43[96], stage0_43[97], stage0_43[98], stage0_43[99], stage0_43[100], stage0_43[101]},
      {stage1_45[16],stage1_44[65],stage1_43[121],stage1_42[126],stage1_41[153]}
   );
   gpc615_5 gpc1606 (
      {stage0_41[437], stage0_41[438], stage0_41[439], stage0_41[440], stage0_41[441]},
      {stage0_42[295]},
      {stage0_43[102], stage0_43[103], stage0_43[104], stage0_43[105], stage0_43[106], stage0_43[107]},
      {stage1_45[17],stage1_44[66],stage1_43[122],stage1_42[127],stage1_41[154]}
   );
   gpc615_5 gpc1607 (
      {stage0_41[442], stage0_41[443], stage0_41[444], stage0_41[445], stage0_41[446]},
      {stage0_42[296]},
      {stage0_43[108], stage0_43[109], stage0_43[110], stage0_43[111], stage0_43[112], stage0_43[113]},
      {stage1_45[18],stage1_44[67],stage1_43[123],stage1_42[128],stage1_41[155]}
   );
   gpc615_5 gpc1608 (
      {stage0_41[447], stage0_41[448], stage0_41[449], stage0_41[450], stage0_41[451]},
      {stage0_42[297]},
      {stage0_43[114], stage0_43[115], stage0_43[116], stage0_43[117], stage0_43[118], stage0_43[119]},
      {stage1_45[19],stage1_44[68],stage1_43[124],stage1_42[129],stage1_41[156]}
   );
   gpc615_5 gpc1609 (
      {stage0_41[452], stage0_41[453], stage0_41[454], stage0_41[455], stage0_41[456]},
      {stage0_42[298]},
      {stage0_43[120], stage0_43[121], stage0_43[122], stage0_43[123], stage0_43[124], stage0_43[125]},
      {stage1_45[20],stage1_44[69],stage1_43[125],stage1_42[130],stage1_41[157]}
   );
   gpc615_5 gpc1610 (
      {stage0_41[457], stage0_41[458], stage0_41[459], stage0_41[460], stage0_41[461]},
      {stage0_42[299]},
      {stage0_43[126], stage0_43[127], stage0_43[128], stage0_43[129], stage0_43[130], stage0_43[131]},
      {stage1_45[21],stage1_44[70],stage1_43[126],stage1_42[131],stage1_41[158]}
   );
   gpc615_5 gpc1611 (
      {stage0_41[462], stage0_41[463], stage0_41[464], stage0_41[465], stage0_41[466]},
      {stage0_42[300]},
      {stage0_43[132], stage0_43[133], stage0_43[134], stage0_43[135], stage0_43[136], stage0_43[137]},
      {stage1_45[22],stage1_44[71],stage1_43[127],stage1_42[132],stage1_41[159]}
   );
   gpc615_5 gpc1612 (
      {stage0_41[467], stage0_41[468], stage0_41[469], stage0_41[470], stage0_41[471]},
      {stage0_42[301]},
      {stage0_43[138], stage0_43[139], stage0_43[140], stage0_43[141], stage0_43[142], stage0_43[143]},
      {stage1_45[23],stage1_44[72],stage1_43[128],stage1_42[133],stage1_41[160]}
   );
   gpc615_5 gpc1613 (
      {stage0_41[472], stage0_41[473], stage0_41[474], stage0_41[475], stage0_41[476]},
      {stage0_42[302]},
      {stage0_43[144], stage0_43[145], stage0_43[146], stage0_43[147], stage0_43[148], stage0_43[149]},
      {stage1_45[24],stage1_44[73],stage1_43[129],stage1_42[134],stage1_41[161]}
   );
   gpc615_5 gpc1614 (
      {stage0_42[303], stage0_42[304], stage0_42[305], stage0_42[306], stage0_42[307]},
      {stage0_43[150]},
      {stage0_44[0], stage0_44[1], stage0_44[2], stage0_44[3], stage0_44[4], stage0_44[5]},
      {stage1_46[0],stage1_45[25],stage1_44[74],stage1_43[130],stage1_42[135]}
   );
   gpc615_5 gpc1615 (
      {stage0_42[308], stage0_42[309], stage0_42[310], stage0_42[311], stage0_42[312]},
      {stage0_43[151]},
      {stage0_44[6], stage0_44[7], stage0_44[8], stage0_44[9], stage0_44[10], stage0_44[11]},
      {stage1_46[1],stage1_45[26],stage1_44[75],stage1_43[131],stage1_42[136]}
   );
   gpc615_5 gpc1616 (
      {stage0_42[313], stage0_42[314], stage0_42[315], stage0_42[316], stage0_42[317]},
      {stage0_43[152]},
      {stage0_44[12], stage0_44[13], stage0_44[14], stage0_44[15], stage0_44[16], stage0_44[17]},
      {stage1_46[2],stage1_45[27],stage1_44[76],stage1_43[132],stage1_42[137]}
   );
   gpc615_5 gpc1617 (
      {stage0_42[318], stage0_42[319], stage0_42[320], stage0_42[321], stage0_42[322]},
      {stage0_43[153]},
      {stage0_44[18], stage0_44[19], stage0_44[20], stage0_44[21], stage0_44[22], stage0_44[23]},
      {stage1_46[3],stage1_45[28],stage1_44[77],stage1_43[133],stage1_42[138]}
   );
   gpc615_5 gpc1618 (
      {stage0_42[323], stage0_42[324], stage0_42[325], stage0_42[326], stage0_42[327]},
      {stage0_43[154]},
      {stage0_44[24], stage0_44[25], stage0_44[26], stage0_44[27], stage0_44[28], stage0_44[29]},
      {stage1_46[4],stage1_45[29],stage1_44[78],stage1_43[134],stage1_42[139]}
   );
   gpc615_5 gpc1619 (
      {stage0_42[328], stage0_42[329], stage0_42[330], stage0_42[331], stage0_42[332]},
      {stage0_43[155]},
      {stage0_44[30], stage0_44[31], stage0_44[32], stage0_44[33], stage0_44[34], stage0_44[35]},
      {stage1_46[5],stage1_45[30],stage1_44[79],stage1_43[135],stage1_42[140]}
   );
   gpc615_5 gpc1620 (
      {stage0_42[333], stage0_42[334], stage0_42[335], stage0_42[336], stage0_42[337]},
      {stage0_43[156]},
      {stage0_44[36], stage0_44[37], stage0_44[38], stage0_44[39], stage0_44[40], stage0_44[41]},
      {stage1_46[6],stage1_45[31],stage1_44[80],stage1_43[136],stage1_42[141]}
   );
   gpc615_5 gpc1621 (
      {stage0_42[338], stage0_42[339], stage0_42[340], stage0_42[341], stage0_42[342]},
      {stage0_43[157]},
      {stage0_44[42], stage0_44[43], stage0_44[44], stage0_44[45], stage0_44[46], stage0_44[47]},
      {stage1_46[7],stage1_45[32],stage1_44[81],stage1_43[137],stage1_42[142]}
   );
   gpc615_5 gpc1622 (
      {stage0_42[343], stage0_42[344], stage0_42[345], stage0_42[346], stage0_42[347]},
      {stage0_43[158]},
      {stage0_44[48], stage0_44[49], stage0_44[50], stage0_44[51], stage0_44[52], stage0_44[53]},
      {stage1_46[8],stage1_45[33],stage1_44[82],stage1_43[138],stage1_42[143]}
   );
   gpc615_5 gpc1623 (
      {stage0_42[348], stage0_42[349], stage0_42[350], stage0_42[351], stage0_42[352]},
      {stage0_43[159]},
      {stage0_44[54], stage0_44[55], stage0_44[56], stage0_44[57], stage0_44[58], stage0_44[59]},
      {stage1_46[9],stage1_45[34],stage1_44[83],stage1_43[139],stage1_42[144]}
   );
   gpc615_5 gpc1624 (
      {stage0_42[353], stage0_42[354], stage0_42[355], stage0_42[356], stage0_42[357]},
      {stage0_43[160]},
      {stage0_44[60], stage0_44[61], stage0_44[62], stage0_44[63], stage0_44[64], stage0_44[65]},
      {stage1_46[10],stage1_45[35],stage1_44[84],stage1_43[140],stage1_42[145]}
   );
   gpc615_5 gpc1625 (
      {stage0_42[358], stage0_42[359], stage0_42[360], stage0_42[361], stage0_42[362]},
      {stage0_43[161]},
      {stage0_44[66], stage0_44[67], stage0_44[68], stage0_44[69], stage0_44[70], stage0_44[71]},
      {stage1_46[11],stage1_45[36],stage1_44[85],stage1_43[141],stage1_42[146]}
   );
   gpc615_5 gpc1626 (
      {stage0_42[363], stage0_42[364], stage0_42[365], stage0_42[366], stage0_42[367]},
      {stage0_43[162]},
      {stage0_44[72], stage0_44[73], stage0_44[74], stage0_44[75], stage0_44[76], stage0_44[77]},
      {stage1_46[12],stage1_45[37],stage1_44[86],stage1_43[142],stage1_42[147]}
   );
   gpc615_5 gpc1627 (
      {stage0_42[368], stage0_42[369], stage0_42[370], stage0_42[371], stage0_42[372]},
      {stage0_43[163]},
      {stage0_44[78], stage0_44[79], stage0_44[80], stage0_44[81], stage0_44[82], stage0_44[83]},
      {stage1_46[13],stage1_45[38],stage1_44[87],stage1_43[143],stage1_42[148]}
   );
   gpc615_5 gpc1628 (
      {stage0_42[373], stage0_42[374], stage0_42[375], stage0_42[376], stage0_42[377]},
      {stage0_43[164]},
      {stage0_44[84], stage0_44[85], stage0_44[86], stage0_44[87], stage0_44[88], stage0_44[89]},
      {stage1_46[14],stage1_45[39],stage1_44[88],stage1_43[144],stage1_42[149]}
   );
   gpc615_5 gpc1629 (
      {stage0_42[378], stage0_42[379], stage0_42[380], stage0_42[381], stage0_42[382]},
      {stage0_43[165]},
      {stage0_44[90], stage0_44[91], stage0_44[92], stage0_44[93], stage0_44[94], stage0_44[95]},
      {stage1_46[15],stage1_45[40],stage1_44[89],stage1_43[145],stage1_42[150]}
   );
   gpc615_5 gpc1630 (
      {stage0_42[383], stage0_42[384], stage0_42[385], stage0_42[386], stage0_42[387]},
      {stage0_43[166]},
      {stage0_44[96], stage0_44[97], stage0_44[98], stage0_44[99], stage0_44[100], stage0_44[101]},
      {stage1_46[16],stage1_45[41],stage1_44[90],stage1_43[146],stage1_42[151]}
   );
   gpc615_5 gpc1631 (
      {stage0_42[388], stage0_42[389], stage0_42[390], stage0_42[391], stage0_42[392]},
      {stage0_43[167]},
      {stage0_44[102], stage0_44[103], stage0_44[104], stage0_44[105], stage0_44[106], stage0_44[107]},
      {stage1_46[17],stage1_45[42],stage1_44[91],stage1_43[147],stage1_42[152]}
   );
   gpc615_5 gpc1632 (
      {stage0_42[393], stage0_42[394], stage0_42[395], stage0_42[396], stage0_42[397]},
      {stage0_43[168]},
      {stage0_44[108], stage0_44[109], stage0_44[110], stage0_44[111], stage0_44[112], stage0_44[113]},
      {stage1_46[18],stage1_45[43],stage1_44[92],stage1_43[148],stage1_42[153]}
   );
   gpc615_5 gpc1633 (
      {stage0_42[398], stage0_42[399], stage0_42[400], stage0_42[401], stage0_42[402]},
      {stage0_43[169]},
      {stage0_44[114], stage0_44[115], stage0_44[116], stage0_44[117], stage0_44[118], stage0_44[119]},
      {stage1_46[19],stage1_45[44],stage1_44[93],stage1_43[149],stage1_42[154]}
   );
   gpc615_5 gpc1634 (
      {stage0_42[403], stage0_42[404], stage0_42[405], stage0_42[406], stage0_42[407]},
      {stage0_43[170]},
      {stage0_44[120], stage0_44[121], stage0_44[122], stage0_44[123], stage0_44[124], stage0_44[125]},
      {stage1_46[20],stage1_45[45],stage1_44[94],stage1_43[150],stage1_42[155]}
   );
   gpc615_5 gpc1635 (
      {stage0_42[408], stage0_42[409], stage0_42[410], stage0_42[411], stage0_42[412]},
      {stage0_43[171]},
      {stage0_44[126], stage0_44[127], stage0_44[128], stage0_44[129], stage0_44[130], stage0_44[131]},
      {stage1_46[21],stage1_45[46],stage1_44[95],stage1_43[151],stage1_42[156]}
   );
   gpc615_5 gpc1636 (
      {stage0_42[413], stage0_42[414], stage0_42[415], stage0_42[416], stage0_42[417]},
      {stage0_43[172]},
      {stage0_44[132], stage0_44[133], stage0_44[134], stage0_44[135], stage0_44[136], stage0_44[137]},
      {stage1_46[22],stage1_45[47],stage1_44[96],stage1_43[152],stage1_42[157]}
   );
   gpc615_5 gpc1637 (
      {stage0_42[418], stage0_42[419], stage0_42[420], stage0_42[421], stage0_42[422]},
      {stage0_43[173]},
      {stage0_44[138], stage0_44[139], stage0_44[140], stage0_44[141], stage0_44[142], stage0_44[143]},
      {stage1_46[23],stage1_45[48],stage1_44[97],stage1_43[153],stage1_42[158]}
   );
   gpc615_5 gpc1638 (
      {stage0_42[423], stage0_42[424], stage0_42[425], stage0_42[426], stage0_42[427]},
      {stage0_43[174]},
      {stage0_44[144], stage0_44[145], stage0_44[146], stage0_44[147], stage0_44[148], stage0_44[149]},
      {stage1_46[24],stage1_45[49],stage1_44[98],stage1_43[154],stage1_42[159]}
   );
   gpc615_5 gpc1639 (
      {stage0_42[428], stage0_42[429], stage0_42[430], stage0_42[431], stage0_42[432]},
      {stage0_43[175]},
      {stage0_44[150], stage0_44[151], stage0_44[152], stage0_44[153], stage0_44[154], stage0_44[155]},
      {stage1_46[25],stage1_45[50],stage1_44[99],stage1_43[155],stage1_42[160]}
   );
   gpc615_5 gpc1640 (
      {stage0_42[433], stage0_42[434], stage0_42[435], stage0_42[436], stage0_42[437]},
      {stage0_43[176]},
      {stage0_44[156], stage0_44[157], stage0_44[158], stage0_44[159], stage0_44[160], stage0_44[161]},
      {stage1_46[26],stage1_45[51],stage1_44[100],stage1_43[156],stage1_42[161]}
   );
   gpc615_5 gpc1641 (
      {stage0_42[438], stage0_42[439], stage0_42[440], stage0_42[441], stage0_42[442]},
      {stage0_43[177]},
      {stage0_44[162], stage0_44[163], stage0_44[164], stage0_44[165], stage0_44[166], stage0_44[167]},
      {stage1_46[27],stage1_45[52],stage1_44[101],stage1_43[157],stage1_42[162]}
   );
   gpc615_5 gpc1642 (
      {stage0_42[443], stage0_42[444], stage0_42[445], stage0_42[446], stage0_42[447]},
      {stage0_43[178]},
      {stage0_44[168], stage0_44[169], stage0_44[170], stage0_44[171], stage0_44[172], stage0_44[173]},
      {stage1_46[28],stage1_45[53],stage1_44[102],stage1_43[158],stage1_42[163]}
   );
   gpc615_5 gpc1643 (
      {stage0_42[448], stage0_42[449], stage0_42[450], stage0_42[451], stage0_42[452]},
      {stage0_43[179]},
      {stage0_44[174], stage0_44[175], stage0_44[176], stage0_44[177], stage0_44[178], stage0_44[179]},
      {stage1_46[29],stage1_45[54],stage1_44[103],stage1_43[159],stage1_42[164]}
   );
   gpc615_5 gpc1644 (
      {stage0_42[453], stage0_42[454], stage0_42[455], stage0_42[456], stage0_42[457]},
      {stage0_43[180]},
      {stage0_44[180], stage0_44[181], stage0_44[182], stage0_44[183], stage0_44[184], stage0_44[185]},
      {stage1_46[30],stage1_45[55],stage1_44[104],stage1_43[160],stage1_42[165]}
   );
   gpc615_5 gpc1645 (
      {stage0_42[458], stage0_42[459], stage0_42[460], stage0_42[461], stage0_42[462]},
      {stage0_43[181]},
      {stage0_44[186], stage0_44[187], stage0_44[188], stage0_44[189], stage0_44[190], stage0_44[191]},
      {stage1_46[31],stage1_45[56],stage1_44[105],stage1_43[161],stage1_42[166]}
   );
   gpc615_5 gpc1646 (
      {stage0_42[463], stage0_42[464], stage0_42[465], stage0_42[466], stage0_42[467]},
      {stage0_43[182]},
      {stage0_44[192], stage0_44[193], stage0_44[194], stage0_44[195], stage0_44[196], stage0_44[197]},
      {stage1_46[32],stage1_45[57],stage1_44[106],stage1_43[162],stage1_42[167]}
   );
   gpc615_5 gpc1647 (
      {stage0_42[468], stage0_42[469], stage0_42[470], stage0_42[471], stage0_42[472]},
      {stage0_43[183]},
      {stage0_44[198], stage0_44[199], stage0_44[200], stage0_44[201], stage0_44[202], stage0_44[203]},
      {stage1_46[33],stage1_45[58],stage1_44[107],stage1_43[163],stage1_42[168]}
   );
   gpc615_5 gpc1648 (
      {stage0_42[473], stage0_42[474], stage0_42[475], stage0_42[476], stage0_42[477]},
      {stage0_43[184]},
      {stage0_44[204], stage0_44[205], stage0_44[206], stage0_44[207], stage0_44[208], stage0_44[209]},
      {stage1_46[34],stage1_45[59],stage1_44[108],stage1_43[164],stage1_42[169]}
   );
   gpc615_5 gpc1649 (
      {stage0_42[478], stage0_42[479], stage0_42[480], stage0_42[481], stage0_42[482]},
      {stage0_43[185]},
      {stage0_44[210], stage0_44[211], stage0_44[212], stage0_44[213], stage0_44[214], stage0_44[215]},
      {stage1_46[35],stage1_45[60],stage1_44[109],stage1_43[165],stage1_42[170]}
   );
   gpc615_5 gpc1650 (
      {stage0_43[186], stage0_43[187], stage0_43[188], stage0_43[189], stage0_43[190]},
      {stage0_44[216]},
      {stage0_45[0], stage0_45[1], stage0_45[2], stage0_45[3], stage0_45[4], stage0_45[5]},
      {stage1_47[0],stage1_46[36],stage1_45[61],stage1_44[110],stage1_43[166]}
   );
   gpc615_5 gpc1651 (
      {stage0_43[191], stage0_43[192], stage0_43[193], stage0_43[194], stage0_43[195]},
      {stage0_44[217]},
      {stage0_45[6], stage0_45[7], stage0_45[8], stage0_45[9], stage0_45[10], stage0_45[11]},
      {stage1_47[1],stage1_46[37],stage1_45[62],stage1_44[111],stage1_43[167]}
   );
   gpc615_5 gpc1652 (
      {stage0_43[196], stage0_43[197], stage0_43[198], stage0_43[199], stage0_43[200]},
      {stage0_44[218]},
      {stage0_45[12], stage0_45[13], stage0_45[14], stage0_45[15], stage0_45[16], stage0_45[17]},
      {stage1_47[2],stage1_46[38],stage1_45[63],stage1_44[112],stage1_43[168]}
   );
   gpc615_5 gpc1653 (
      {stage0_43[201], stage0_43[202], stage0_43[203], stage0_43[204], stage0_43[205]},
      {stage0_44[219]},
      {stage0_45[18], stage0_45[19], stage0_45[20], stage0_45[21], stage0_45[22], stage0_45[23]},
      {stage1_47[3],stage1_46[39],stage1_45[64],stage1_44[113],stage1_43[169]}
   );
   gpc615_5 gpc1654 (
      {stage0_43[206], stage0_43[207], stage0_43[208], stage0_43[209], stage0_43[210]},
      {stage0_44[220]},
      {stage0_45[24], stage0_45[25], stage0_45[26], stage0_45[27], stage0_45[28], stage0_45[29]},
      {stage1_47[4],stage1_46[40],stage1_45[65],stage1_44[114],stage1_43[170]}
   );
   gpc615_5 gpc1655 (
      {stage0_43[211], stage0_43[212], stage0_43[213], stage0_43[214], stage0_43[215]},
      {stage0_44[221]},
      {stage0_45[30], stage0_45[31], stage0_45[32], stage0_45[33], stage0_45[34], stage0_45[35]},
      {stage1_47[5],stage1_46[41],stage1_45[66],stage1_44[115],stage1_43[171]}
   );
   gpc615_5 gpc1656 (
      {stage0_43[216], stage0_43[217], stage0_43[218], stage0_43[219], stage0_43[220]},
      {stage0_44[222]},
      {stage0_45[36], stage0_45[37], stage0_45[38], stage0_45[39], stage0_45[40], stage0_45[41]},
      {stage1_47[6],stage1_46[42],stage1_45[67],stage1_44[116],stage1_43[172]}
   );
   gpc615_5 gpc1657 (
      {stage0_43[221], stage0_43[222], stage0_43[223], stage0_43[224], stage0_43[225]},
      {stage0_44[223]},
      {stage0_45[42], stage0_45[43], stage0_45[44], stage0_45[45], stage0_45[46], stage0_45[47]},
      {stage1_47[7],stage1_46[43],stage1_45[68],stage1_44[117],stage1_43[173]}
   );
   gpc615_5 gpc1658 (
      {stage0_43[226], stage0_43[227], stage0_43[228], stage0_43[229], stage0_43[230]},
      {stage0_44[224]},
      {stage0_45[48], stage0_45[49], stage0_45[50], stage0_45[51], stage0_45[52], stage0_45[53]},
      {stage1_47[8],stage1_46[44],stage1_45[69],stage1_44[118],stage1_43[174]}
   );
   gpc615_5 gpc1659 (
      {stage0_43[231], stage0_43[232], stage0_43[233], stage0_43[234], stage0_43[235]},
      {stage0_44[225]},
      {stage0_45[54], stage0_45[55], stage0_45[56], stage0_45[57], stage0_45[58], stage0_45[59]},
      {stage1_47[9],stage1_46[45],stage1_45[70],stage1_44[119],stage1_43[175]}
   );
   gpc615_5 gpc1660 (
      {stage0_43[236], stage0_43[237], stage0_43[238], stage0_43[239], stage0_43[240]},
      {stage0_44[226]},
      {stage0_45[60], stage0_45[61], stage0_45[62], stage0_45[63], stage0_45[64], stage0_45[65]},
      {stage1_47[10],stage1_46[46],stage1_45[71],stage1_44[120],stage1_43[176]}
   );
   gpc615_5 gpc1661 (
      {stage0_43[241], stage0_43[242], stage0_43[243], stage0_43[244], stage0_43[245]},
      {stage0_44[227]},
      {stage0_45[66], stage0_45[67], stage0_45[68], stage0_45[69], stage0_45[70], stage0_45[71]},
      {stage1_47[11],stage1_46[47],stage1_45[72],stage1_44[121],stage1_43[177]}
   );
   gpc615_5 gpc1662 (
      {stage0_43[246], stage0_43[247], stage0_43[248], stage0_43[249], stage0_43[250]},
      {stage0_44[228]},
      {stage0_45[72], stage0_45[73], stage0_45[74], stage0_45[75], stage0_45[76], stage0_45[77]},
      {stage1_47[12],stage1_46[48],stage1_45[73],stage1_44[122],stage1_43[178]}
   );
   gpc615_5 gpc1663 (
      {stage0_43[251], stage0_43[252], stage0_43[253], stage0_43[254], stage0_43[255]},
      {stage0_44[229]},
      {stage0_45[78], stage0_45[79], stage0_45[80], stage0_45[81], stage0_45[82], stage0_45[83]},
      {stage1_47[13],stage1_46[49],stage1_45[74],stage1_44[123],stage1_43[179]}
   );
   gpc615_5 gpc1664 (
      {stage0_43[256], stage0_43[257], stage0_43[258], stage0_43[259], stage0_43[260]},
      {stage0_44[230]},
      {stage0_45[84], stage0_45[85], stage0_45[86], stage0_45[87], stage0_45[88], stage0_45[89]},
      {stage1_47[14],stage1_46[50],stage1_45[75],stage1_44[124],stage1_43[180]}
   );
   gpc615_5 gpc1665 (
      {stage0_43[261], stage0_43[262], stage0_43[263], stage0_43[264], stage0_43[265]},
      {stage0_44[231]},
      {stage0_45[90], stage0_45[91], stage0_45[92], stage0_45[93], stage0_45[94], stage0_45[95]},
      {stage1_47[15],stage1_46[51],stage1_45[76],stage1_44[125],stage1_43[181]}
   );
   gpc615_5 gpc1666 (
      {stage0_43[266], stage0_43[267], stage0_43[268], stage0_43[269], stage0_43[270]},
      {stage0_44[232]},
      {stage0_45[96], stage0_45[97], stage0_45[98], stage0_45[99], stage0_45[100], stage0_45[101]},
      {stage1_47[16],stage1_46[52],stage1_45[77],stage1_44[126],stage1_43[182]}
   );
   gpc615_5 gpc1667 (
      {stage0_43[271], stage0_43[272], stage0_43[273], stage0_43[274], stage0_43[275]},
      {stage0_44[233]},
      {stage0_45[102], stage0_45[103], stage0_45[104], stage0_45[105], stage0_45[106], stage0_45[107]},
      {stage1_47[17],stage1_46[53],stage1_45[78],stage1_44[127],stage1_43[183]}
   );
   gpc615_5 gpc1668 (
      {stage0_43[276], stage0_43[277], stage0_43[278], stage0_43[279], stage0_43[280]},
      {stage0_44[234]},
      {stage0_45[108], stage0_45[109], stage0_45[110], stage0_45[111], stage0_45[112], stage0_45[113]},
      {stage1_47[18],stage1_46[54],stage1_45[79],stage1_44[128],stage1_43[184]}
   );
   gpc615_5 gpc1669 (
      {stage0_43[281], stage0_43[282], stage0_43[283], stage0_43[284], stage0_43[285]},
      {stage0_44[235]},
      {stage0_45[114], stage0_45[115], stage0_45[116], stage0_45[117], stage0_45[118], stage0_45[119]},
      {stage1_47[19],stage1_46[55],stage1_45[80],stage1_44[129],stage1_43[185]}
   );
   gpc615_5 gpc1670 (
      {stage0_43[286], stage0_43[287], stage0_43[288], stage0_43[289], stage0_43[290]},
      {stage0_44[236]},
      {stage0_45[120], stage0_45[121], stage0_45[122], stage0_45[123], stage0_45[124], stage0_45[125]},
      {stage1_47[20],stage1_46[56],stage1_45[81],stage1_44[130],stage1_43[186]}
   );
   gpc615_5 gpc1671 (
      {stage0_43[291], stage0_43[292], stage0_43[293], stage0_43[294], stage0_43[295]},
      {stage0_44[237]},
      {stage0_45[126], stage0_45[127], stage0_45[128], stage0_45[129], stage0_45[130], stage0_45[131]},
      {stage1_47[21],stage1_46[57],stage1_45[82],stage1_44[131],stage1_43[187]}
   );
   gpc615_5 gpc1672 (
      {stage0_43[296], stage0_43[297], stage0_43[298], stage0_43[299], stage0_43[300]},
      {stage0_44[238]},
      {stage0_45[132], stage0_45[133], stage0_45[134], stage0_45[135], stage0_45[136], stage0_45[137]},
      {stage1_47[22],stage1_46[58],stage1_45[83],stage1_44[132],stage1_43[188]}
   );
   gpc615_5 gpc1673 (
      {stage0_43[301], stage0_43[302], stage0_43[303], stage0_43[304], stage0_43[305]},
      {stage0_44[239]},
      {stage0_45[138], stage0_45[139], stage0_45[140], stage0_45[141], stage0_45[142], stage0_45[143]},
      {stage1_47[23],stage1_46[59],stage1_45[84],stage1_44[133],stage1_43[189]}
   );
   gpc615_5 gpc1674 (
      {stage0_43[306], stage0_43[307], stage0_43[308], stage0_43[309], stage0_43[310]},
      {stage0_44[240]},
      {stage0_45[144], stage0_45[145], stage0_45[146], stage0_45[147], stage0_45[148], stage0_45[149]},
      {stage1_47[24],stage1_46[60],stage1_45[85],stage1_44[134],stage1_43[190]}
   );
   gpc615_5 gpc1675 (
      {stage0_43[311], stage0_43[312], stage0_43[313], stage0_43[314], stage0_43[315]},
      {stage0_44[241]},
      {stage0_45[150], stage0_45[151], stage0_45[152], stage0_45[153], stage0_45[154], stage0_45[155]},
      {stage1_47[25],stage1_46[61],stage1_45[86],stage1_44[135],stage1_43[191]}
   );
   gpc615_5 gpc1676 (
      {stage0_43[316], stage0_43[317], stage0_43[318], stage0_43[319], stage0_43[320]},
      {stage0_44[242]},
      {stage0_45[156], stage0_45[157], stage0_45[158], stage0_45[159], stage0_45[160], stage0_45[161]},
      {stage1_47[26],stage1_46[62],stage1_45[87],stage1_44[136],stage1_43[192]}
   );
   gpc615_5 gpc1677 (
      {stage0_43[321], stage0_43[322], stage0_43[323], stage0_43[324], stage0_43[325]},
      {stage0_44[243]},
      {stage0_45[162], stage0_45[163], stage0_45[164], stage0_45[165], stage0_45[166], stage0_45[167]},
      {stage1_47[27],stage1_46[63],stage1_45[88],stage1_44[137],stage1_43[193]}
   );
   gpc615_5 gpc1678 (
      {stage0_43[326], stage0_43[327], stage0_43[328], stage0_43[329], stage0_43[330]},
      {stage0_44[244]},
      {stage0_45[168], stage0_45[169], stage0_45[170], stage0_45[171], stage0_45[172], stage0_45[173]},
      {stage1_47[28],stage1_46[64],stage1_45[89],stage1_44[138],stage1_43[194]}
   );
   gpc615_5 gpc1679 (
      {stage0_43[331], stage0_43[332], stage0_43[333], stage0_43[334], stage0_43[335]},
      {stage0_44[245]},
      {stage0_45[174], stage0_45[175], stage0_45[176], stage0_45[177], stage0_45[178], stage0_45[179]},
      {stage1_47[29],stage1_46[65],stage1_45[90],stage1_44[139],stage1_43[195]}
   );
   gpc615_5 gpc1680 (
      {stage0_43[336], stage0_43[337], stage0_43[338], stage0_43[339], stage0_43[340]},
      {stage0_44[246]},
      {stage0_45[180], stage0_45[181], stage0_45[182], stage0_45[183], stage0_45[184], stage0_45[185]},
      {stage1_47[30],stage1_46[66],stage1_45[91],stage1_44[140],stage1_43[196]}
   );
   gpc615_5 gpc1681 (
      {stage0_43[341], stage0_43[342], stage0_43[343], stage0_43[344], stage0_43[345]},
      {stage0_44[247]},
      {stage0_45[186], stage0_45[187], stage0_45[188], stage0_45[189], stage0_45[190], stage0_45[191]},
      {stage1_47[31],stage1_46[67],stage1_45[92],stage1_44[141],stage1_43[197]}
   );
   gpc615_5 gpc1682 (
      {stage0_43[346], stage0_43[347], stage0_43[348], stage0_43[349], stage0_43[350]},
      {stage0_44[248]},
      {stage0_45[192], stage0_45[193], stage0_45[194], stage0_45[195], stage0_45[196], stage0_45[197]},
      {stage1_47[32],stage1_46[68],stage1_45[93],stage1_44[142],stage1_43[198]}
   );
   gpc615_5 gpc1683 (
      {stage0_43[351], stage0_43[352], stage0_43[353], stage0_43[354], stage0_43[355]},
      {stage0_44[249]},
      {stage0_45[198], stage0_45[199], stage0_45[200], stage0_45[201], stage0_45[202], stage0_45[203]},
      {stage1_47[33],stage1_46[69],stage1_45[94],stage1_44[143],stage1_43[199]}
   );
   gpc615_5 gpc1684 (
      {stage0_43[356], stage0_43[357], stage0_43[358], stage0_43[359], stage0_43[360]},
      {stage0_44[250]},
      {stage0_45[204], stage0_45[205], stage0_45[206], stage0_45[207], stage0_45[208], stage0_45[209]},
      {stage1_47[34],stage1_46[70],stage1_45[95],stage1_44[144],stage1_43[200]}
   );
   gpc615_5 gpc1685 (
      {stage0_43[361], stage0_43[362], stage0_43[363], stage0_43[364], stage0_43[365]},
      {stage0_44[251]},
      {stage0_45[210], stage0_45[211], stage0_45[212], stage0_45[213], stage0_45[214], stage0_45[215]},
      {stage1_47[35],stage1_46[71],stage1_45[96],stage1_44[145],stage1_43[201]}
   );
   gpc615_5 gpc1686 (
      {stage0_43[366], stage0_43[367], stage0_43[368], stage0_43[369], stage0_43[370]},
      {stage0_44[252]},
      {stage0_45[216], stage0_45[217], stage0_45[218], stage0_45[219], stage0_45[220], stage0_45[221]},
      {stage1_47[36],stage1_46[72],stage1_45[97],stage1_44[146],stage1_43[202]}
   );
   gpc615_5 gpc1687 (
      {stage0_43[371], stage0_43[372], stage0_43[373], stage0_43[374], stage0_43[375]},
      {stage0_44[253]},
      {stage0_45[222], stage0_45[223], stage0_45[224], stage0_45[225], stage0_45[226], stage0_45[227]},
      {stage1_47[37],stage1_46[73],stage1_45[98],stage1_44[147],stage1_43[203]}
   );
   gpc615_5 gpc1688 (
      {stage0_43[376], stage0_43[377], stage0_43[378], stage0_43[379], stage0_43[380]},
      {stage0_44[254]},
      {stage0_45[228], stage0_45[229], stage0_45[230], stage0_45[231], stage0_45[232], stage0_45[233]},
      {stage1_47[38],stage1_46[74],stage1_45[99],stage1_44[148],stage1_43[204]}
   );
   gpc615_5 gpc1689 (
      {stage0_43[381], stage0_43[382], stage0_43[383], stage0_43[384], stage0_43[385]},
      {stage0_44[255]},
      {stage0_45[234], stage0_45[235], stage0_45[236], stage0_45[237], stage0_45[238], stage0_45[239]},
      {stage1_47[39],stage1_46[75],stage1_45[100],stage1_44[149],stage1_43[205]}
   );
   gpc615_5 gpc1690 (
      {stage0_43[386], stage0_43[387], stage0_43[388], stage0_43[389], stage0_43[390]},
      {stage0_44[256]},
      {stage0_45[240], stage0_45[241], stage0_45[242], stage0_45[243], stage0_45[244], stage0_45[245]},
      {stage1_47[40],stage1_46[76],stage1_45[101],stage1_44[150],stage1_43[206]}
   );
   gpc615_5 gpc1691 (
      {stage0_43[391], stage0_43[392], stage0_43[393], stage0_43[394], stage0_43[395]},
      {stage0_44[257]},
      {stage0_45[246], stage0_45[247], stage0_45[248], stage0_45[249], stage0_45[250], stage0_45[251]},
      {stage1_47[41],stage1_46[77],stage1_45[102],stage1_44[151],stage1_43[207]}
   );
   gpc615_5 gpc1692 (
      {stage0_43[396], stage0_43[397], stage0_43[398], stage0_43[399], stage0_43[400]},
      {stage0_44[258]},
      {stage0_45[252], stage0_45[253], stage0_45[254], stage0_45[255], stage0_45[256], stage0_45[257]},
      {stage1_47[42],stage1_46[78],stage1_45[103],stage1_44[152],stage1_43[208]}
   );
   gpc615_5 gpc1693 (
      {stage0_43[401], stage0_43[402], stage0_43[403], stage0_43[404], stage0_43[405]},
      {stage0_44[259]},
      {stage0_45[258], stage0_45[259], stage0_45[260], stage0_45[261], stage0_45[262], stage0_45[263]},
      {stage1_47[43],stage1_46[79],stage1_45[104],stage1_44[153],stage1_43[209]}
   );
   gpc615_5 gpc1694 (
      {stage0_43[406], stage0_43[407], stage0_43[408], stage0_43[409], stage0_43[410]},
      {stage0_44[260]},
      {stage0_45[264], stage0_45[265], stage0_45[266], stage0_45[267], stage0_45[268], stage0_45[269]},
      {stage1_47[44],stage1_46[80],stage1_45[105],stage1_44[154],stage1_43[210]}
   );
   gpc615_5 gpc1695 (
      {stage0_43[411], stage0_43[412], stage0_43[413], stage0_43[414], stage0_43[415]},
      {stage0_44[261]},
      {stage0_45[270], stage0_45[271], stage0_45[272], stage0_45[273], stage0_45[274], stage0_45[275]},
      {stage1_47[45],stage1_46[81],stage1_45[106],stage1_44[155],stage1_43[211]}
   );
   gpc615_5 gpc1696 (
      {stage0_43[416], stage0_43[417], stage0_43[418], stage0_43[419], stage0_43[420]},
      {stage0_44[262]},
      {stage0_45[276], stage0_45[277], stage0_45[278], stage0_45[279], stage0_45[280], stage0_45[281]},
      {stage1_47[46],stage1_46[82],stage1_45[107],stage1_44[156],stage1_43[212]}
   );
   gpc615_5 gpc1697 (
      {stage0_43[421], stage0_43[422], stage0_43[423], stage0_43[424], stage0_43[425]},
      {stage0_44[263]},
      {stage0_45[282], stage0_45[283], stage0_45[284], stage0_45[285], stage0_45[286], stage0_45[287]},
      {stage1_47[47],stage1_46[83],stage1_45[108],stage1_44[157],stage1_43[213]}
   );
   gpc615_5 gpc1698 (
      {stage0_43[426], stage0_43[427], stage0_43[428], stage0_43[429], stage0_43[430]},
      {stage0_44[264]},
      {stage0_45[288], stage0_45[289], stage0_45[290], stage0_45[291], stage0_45[292], stage0_45[293]},
      {stage1_47[48],stage1_46[84],stage1_45[109],stage1_44[158],stage1_43[214]}
   );
   gpc615_5 gpc1699 (
      {stage0_43[431], stage0_43[432], stage0_43[433], stage0_43[434], stage0_43[435]},
      {stage0_44[265]},
      {stage0_45[294], stage0_45[295], stage0_45[296], stage0_45[297], stage0_45[298], stage0_45[299]},
      {stage1_47[49],stage1_46[85],stage1_45[110],stage1_44[159],stage1_43[215]}
   );
   gpc615_5 gpc1700 (
      {stage0_43[436], stage0_43[437], stage0_43[438], stage0_43[439], stage0_43[440]},
      {stage0_44[266]},
      {stage0_45[300], stage0_45[301], stage0_45[302], stage0_45[303], stage0_45[304], stage0_45[305]},
      {stage1_47[50],stage1_46[86],stage1_45[111],stage1_44[160],stage1_43[216]}
   );
   gpc615_5 gpc1701 (
      {stage0_43[441], stage0_43[442], stage0_43[443], stage0_43[444], stage0_43[445]},
      {stage0_44[267]},
      {stage0_45[306], stage0_45[307], stage0_45[308], stage0_45[309], stage0_45[310], stage0_45[311]},
      {stage1_47[51],stage1_46[87],stage1_45[112],stage1_44[161],stage1_43[217]}
   );
   gpc615_5 gpc1702 (
      {stage0_43[446], stage0_43[447], stage0_43[448], stage0_43[449], stage0_43[450]},
      {stage0_44[268]},
      {stage0_45[312], stage0_45[313], stage0_45[314], stage0_45[315], stage0_45[316], stage0_45[317]},
      {stage1_47[52],stage1_46[88],stage1_45[113],stage1_44[162],stage1_43[218]}
   );
   gpc615_5 gpc1703 (
      {stage0_44[269], stage0_44[270], stage0_44[271], stage0_44[272], stage0_44[273]},
      {stage0_45[318]},
      {stage0_46[0], stage0_46[1], stage0_46[2], stage0_46[3], stage0_46[4], stage0_46[5]},
      {stage1_48[0],stage1_47[53],stage1_46[89],stage1_45[114],stage1_44[163]}
   );
   gpc615_5 gpc1704 (
      {stage0_44[274], stage0_44[275], stage0_44[276], stage0_44[277], stage0_44[278]},
      {stage0_45[319]},
      {stage0_46[6], stage0_46[7], stage0_46[8], stage0_46[9], stage0_46[10], stage0_46[11]},
      {stage1_48[1],stage1_47[54],stage1_46[90],stage1_45[115],stage1_44[164]}
   );
   gpc615_5 gpc1705 (
      {stage0_44[279], stage0_44[280], stage0_44[281], stage0_44[282], stage0_44[283]},
      {stage0_45[320]},
      {stage0_46[12], stage0_46[13], stage0_46[14], stage0_46[15], stage0_46[16], stage0_46[17]},
      {stage1_48[2],stage1_47[55],stage1_46[91],stage1_45[116],stage1_44[165]}
   );
   gpc615_5 gpc1706 (
      {stage0_44[284], stage0_44[285], stage0_44[286], stage0_44[287], stage0_44[288]},
      {stage0_45[321]},
      {stage0_46[18], stage0_46[19], stage0_46[20], stage0_46[21], stage0_46[22], stage0_46[23]},
      {stage1_48[3],stage1_47[56],stage1_46[92],stage1_45[117],stage1_44[166]}
   );
   gpc615_5 gpc1707 (
      {stage0_44[289], stage0_44[290], stage0_44[291], stage0_44[292], stage0_44[293]},
      {stage0_45[322]},
      {stage0_46[24], stage0_46[25], stage0_46[26], stage0_46[27], stage0_46[28], stage0_46[29]},
      {stage1_48[4],stage1_47[57],stage1_46[93],stage1_45[118],stage1_44[167]}
   );
   gpc615_5 gpc1708 (
      {stage0_44[294], stage0_44[295], stage0_44[296], stage0_44[297], stage0_44[298]},
      {stage0_45[323]},
      {stage0_46[30], stage0_46[31], stage0_46[32], stage0_46[33], stage0_46[34], stage0_46[35]},
      {stage1_48[5],stage1_47[58],stage1_46[94],stage1_45[119],stage1_44[168]}
   );
   gpc615_5 gpc1709 (
      {stage0_44[299], stage0_44[300], stage0_44[301], stage0_44[302], stage0_44[303]},
      {stage0_45[324]},
      {stage0_46[36], stage0_46[37], stage0_46[38], stage0_46[39], stage0_46[40], stage0_46[41]},
      {stage1_48[6],stage1_47[59],stage1_46[95],stage1_45[120],stage1_44[169]}
   );
   gpc615_5 gpc1710 (
      {stage0_44[304], stage0_44[305], stage0_44[306], stage0_44[307], stage0_44[308]},
      {stage0_45[325]},
      {stage0_46[42], stage0_46[43], stage0_46[44], stage0_46[45], stage0_46[46], stage0_46[47]},
      {stage1_48[7],stage1_47[60],stage1_46[96],stage1_45[121],stage1_44[170]}
   );
   gpc615_5 gpc1711 (
      {stage0_44[309], stage0_44[310], stage0_44[311], stage0_44[312], stage0_44[313]},
      {stage0_45[326]},
      {stage0_46[48], stage0_46[49], stage0_46[50], stage0_46[51], stage0_46[52], stage0_46[53]},
      {stage1_48[8],stage1_47[61],stage1_46[97],stage1_45[122],stage1_44[171]}
   );
   gpc615_5 gpc1712 (
      {stage0_44[314], stage0_44[315], stage0_44[316], stage0_44[317], stage0_44[318]},
      {stage0_45[327]},
      {stage0_46[54], stage0_46[55], stage0_46[56], stage0_46[57], stage0_46[58], stage0_46[59]},
      {stage1_48[9],stage1_47[62],stage1_46[98],stage1_45[123],stage1_44[172]}
   );
   gpc615_5 gpc1713 (
      {stage0_44[319], stage0_44[320], stage0_44[321], stage0_44[322], stage0_44[323]},
      {stage0_45[328]},
      {stage0_46[60], stage0_46[61], stage0_46[62], stage0_46[63], stage0_46[64], stage0_46[65]},
      {stage1_48[10],stage1_47[63],stage1_46[99],stage1_45[124],stage1_44[173]}
   );
   gpc615_5 gpc1714 (
      {stage0_44[324], stage0_44[325], stage0_44[326], stage0_44[327], stage0_44[328]},
      {stage0_45[329]},
      {stage0_46[66], stage0_46[67], stage0_46[68], stage0_46[69], stage0_46[70], stage0_46[71]},
      {stage1_48[11],stage1_47[64],stage1_46[100],stage1_45[125],stage1_44[174]}
   );
   gpc615_5 gpc1715 (
      {stage0_44[329], stage0_44[330], stage0_44[331], stage0_44[332], stage0_44[333]},
      {stage0_45[330]},
      {stage0_46[72], stage0_46[73], stage0_46[74], stage0_46[75], stage0_46[76], stage0_46[77]},
      {stage1_48[12],stage1_47[65],stage1_46[101],stage1_45[126],stage1_44[175]}
   );
   gpc615_5 gpc1716 (
      {stage0_44[334], stage0_44[335], stage0_44[336], stage0_44[337], stage0_44[338]},
      {stage0_45[331]},
      {stage0_46[78], stage0_46[79], stage0_46[80], stage0_46[81], stage0_46[82], stage0_46[83]},
      {stage1_48[13],stage1_47[66],stage1_46[102],stage1_45[127],stage1_44[176]}
   );
   gpc615_5 gpc1717 (
      {stage0_44[339], stage0_44[340], stage0_44[341], stage0_44[342], stage0_44[343]},
      {stage0_45[332]},
      {stage0_46[84], stage0_46[85], stage0_46[86], stage0_46[87], stage0_46[88], stage0_46[89]},
      {stage1_48[14],stage1_47[67],stage1_46[103],stage1_45[128],stage1_44[177]}
   );
   gpc615_5 gpc1718 (
      {stage0_44[344], stage0_44[345], stage0_44[346], stage0_44[347], stage0_44[348]},
      {stage0_45[333]},
      {stage0_46[90], stage0_46[91], stage0_46[92], stage0_46[93], stage0_46[94], stage0_46[95]},
      {stage1_48[15],stage1_47[68],stage1_46[104],stage1_45[129],stage1_44[178]}
   );
   gpc615_5 gpc1719 (
      {stage0_44[349], stage0_44[350], stage0_44[351], stage0_44[352], stage0_44[353]},
      {stage0_45[334]},
      {stage0_46[96], stage0_46[97], stage0_46[98], stage0_46[99], stage0_46[100], stage0_46[101]},
      {stage1_48[16],stage1_47[69],stage1_46[105],stage1_45[130],stage1_44[179]}
   );
   gpc615_5 gpc1720 (
      {stage0_44[354], stage0_44[355], stage0_44[356], stage0_44[357], stage0_44[358]},
      {stage0_45[335]},
      {stage0_46[102], stage0_46[103], stage0_46[104], stage0_46[105], stage0_46[106], stage0_46[107]},
      {stage1_48[17],stage1_47[70],stage1_46[106],stage1_45[131],stage1_44[180]}
   );
   gpc615_5 gpc1721 (
      {stage0_44[359], stage0_44[360], stage0_44[361], stage0_44[362], stage0_44[363]},
      {stage0_45[336]},
      {stage0_46[108], stage0_46[109], stage0_46[110], stage0_46[111], stage0_46[112], stage0_46[113]},
      {stage1_48[18],stage1_47[71],stage1_46[107],stage1_45[132],stage1_44[181]}
   );
   gpc615_5 gpc1722 (
      {stage0_44[364], stage0_44[365], stage0_44[366], stage0_44[367], stage0_44[368]},
      {stage0_45[337]},
      {stage0_46[114], stage0_46[115], stage0_46[116], stage0_46[117], stage0_46[118], stage0_46[119]},
      {stage1_48[19],stage1_47[72],stage1_46[108],stage1_45[133],stage1_44[182]}
   );
   gpc615_5 gpc1723 (
      {stage0_44[369], stage0_44[370], stage0_44[371], stage0_44[372], stage0_44[373]},
      {stage0_45[338]},
      {stage0_46[120], stage0_46[121], stage0_46[122], stage0_46[123], stage0_46[124], stage0_46[125]},
      {stage1_48[20],stage1_47[73],stage1_46[109],stage1_45[134],stage1_44[183]}
   );
   gpc615_5 gpc1724 (
      {stage0_44[374], stage0_44[375], stage0_44[376], stage0_44[377], stage0_44[378]},
      {stage0_45[339]},
      {stage0_46[126], stage0_46[127], stage0_46[128], stage0_46[129], stage0_46[130], stage0_46[131]},
      {stage1_48[21],stage1_47[74],stage1_46[110],stage1_45[135],stage1_44[184]}
   );
   gpc615_5 gpc1725 (
      {stage0_44[379], stage0_44[380], stage0_44[381], stage0_44[382], stage0_44[383]},
      {stage0_45[340]},
      {stage0_46[132], stage0_46[133], stage0_46[134], stage0_46[135], stage0_46[136], stage0_46[137]},
      {stage1_48[22],stage1_47[75],stage1_46[111],stage1_45[136],stage1_44[185]}
   );
   gpc615_5 gpc1726 (
      {stage0_44[384], stage0_44[385], stage0_44[386], stage0_44[387], stage0_44[388]},
      {stage0_45[341]},
      {stage0_46[138], stage0_46[139], stage0_46[140], stage0_46[141], stage0_46[142], stage0_46[143]},
      {stage1_48[23],stage1_47[76],stage1_46[112],stage1_45[137],stage1_44[186]}
   );
   gpc615_5 gpc1727 (
      {stage0_44[389], stage0_44[390], stage0_44[391], stage0_44[392], stage0_44[393]},
      {stage0_45[342]},
      {stage0_46[144], stage0_46[145], stage0_46[146], stage0_46[147], stage0_46[148], stage0_46[149]},
      {stage1_48[24],stage1_47[77],stage1_46[113],stage1_45[138],stage1_44[187]}
   );
   gpc615_5 gpc1728 (
      {stage0_44[394], stage0_44[395], stage0_44[396], stage0_44[397], stage0_44[398]},
      {stage0_45[343]},
      {stage0_46[150], stage0_46[151], stage0_46[152], stage0_46[153], stage0_46[154], stage0_46[155]},
      {stage1_48[25],stage1_47[78],stage1_46[114],stage1_45[139],stage1_44[188]}
   );
   gpc615_5 gpc1729 (
      {stage0_44[399], stage0_44[400], stage0_44[401], stage0_44[402], stage0_44[403]},
      {stage0_45[344]},
      {stage0_46[156], stage0_46[157], stage0_46[158], stage0_46[159], stage0_46[160], stage0_46[161]},
      {stage1_48[26],stage1_47[79],stage1_46[115],stage1_45[140],stage1_44[189]}
   );
   gpc615_5 gpc1730 (
      {stage0_44[404], stage0_44[405], stage0_44[406], stage0_44[407], stage0_44[408]},
      {stage0_45[345]},
      {stage0_46[162], stage0_46[163], stage0_46[164], stage0_46[165], stage0_46[166], stage0_46[167]},
      {stage1_48[27],stage1_47[80],stage1_46[116],stage1_45[141],stage1_44[190]}
   );
   gpc615_5 gpc1731 (
      {stage0_44[409], stage0_44[410], stage0_44[411], stage0_44[412], stage0_44[413]},
      {stage0_45[346]},
      {stage0_46[168], stage0_46[169], stage0_46[170], stage0_46[171], stage0_46[172], stage0_46[173]},
      {stage1_48[28],stage1_47[81],stage1_46[117],stage1_45[142],stage1_44[191]}
   );
   gpc615_5 gpc1732 (
      {stage0_44[414], stage0_44[415], stage0_44[416], stage0_44[417], stage0_44[418]},
      {stage0_45[347]},
      {stage0_46[174], stage0_46[175], stage0_46[176], stage0_46[177], stage0_46[178], stage0_46[179]},
      {stage1_48[29],stage1_47[82],stage1_46[118],stage1_45[143],stage1_44[192]}
   );
   gpc615_5 gpc1733 (
      {stage0_44[419], stage0_44[420], stage0_44[421], stage0_44[422], stage0_44[423]},
      {stage0_45[348]},
      {stage0_46[180], stage0_46[181], stage0_46[182], stage0_46[183], stage0_46[184], stage0_46[185]},
      {stage1_48[30],stage1_47[83],stage1_46[119],stage1_45[144],stage1_44[193]}
   );
   gpc606_5 gpc1734 (
      {stage0_45[349], stage0_45[350], stage0_45[351], stage0_45[352], stage0_45[353], stage0_45[354]},
      {stage0_47[0], stage0_47[1], stage0_47[2], stage0_47[3], stage0_47[4], stage0_47[5]},
      {stage1_49[0],stage1_48[31],stage1_47[84],stage1_46[120],stage1_45[145]}
   );
   gpc606_5 gpc1735 (
      {stage0_45[355], stage0_45[356], stage0_45[357], stage0_45[358], stage0_45[359], stage0_45[360]},
      {stage0_47[6], stage0_47[7], stage0_47[8], stage0_47[9], stage0_47[10], stage0_47[11]},
      {stage1_49[1],stage1_48[32],stage1_47[85],stage1_46[121],stage1_45[146]}
   );
   gpc606_5 gpc1736 (
      {stage0_45[361], stage0_45[362], stage0_45[363], stage0_45[364], stage0_45[365], stage0_45[366]},
      {stage0_47[12], stage0_47[13], stage0_47[14], stage0_47[15], stage0_47[16], stage0_47[17]},
      {stage1_49[2],stage1_48[33],stage1_47[86],stage1_46[122],stage1_45[147]}
   );
   gpc606_5 gpc1737 (
      {stage0_45[367], stage0_45[368], stage0_45[369], stage0_45[370], stage0_45[371], stage0_45[372]},
      {stage0_47[18], stage0_47[19], stage0_47[20], stage0_47[21], stage0_47[22], stage0_47[23]},
      {stage1_49[3],stage1_48[34],stage1_47[87],stage1_46[123],stage1_45[148]}
   );
   gpc606_5 gpc1738 (
      {stage0_45[373], stage0_45[374], stage0_45[375], stage0_45[376], stage0_45[377], stage0_45[378]},
      {stage0_47[24], stage0_47[25], stage0_47[26], stage0_47[27], stage0_47[28], stage0_47[29]},
      {stage1_49[4],stage1_48[35],stage1_47[88],stage1_46[124],stage1_45[149]}
   );
   gpc606_5 gpc1739 (
      {stage0_45[379], stage0_45[380], stage0_45[381], stage0_45[382], stage0_45[383], stage0_45[384]},
      {stage0_47[30], stage0_47[31], stage0_47[32], stage0_47[33], stage0_47[34], stage0_47[35]},
      {stage1_49[5],stage1_48[36],stage1_47[89],stage1_46[125],stage1_45[150]}
   );
   gpc606_5 gpc1740 (
      {stage0_45[385], stage0_45[386], stage0_45[387], stage0_45[388], stage0_45[389], stage0_45[390]},
      {stage0_47[36], stage0_47[37], stage0_47[38], stage0_47[39], stage0_47[40], stage0_47[41]},
      {stage1_49[6],stage1_48[37],stage1_47[90],stage1_46[126],stage1_45[151]}
   );
   gpc606_5 gpc1741 (
      {stage0_45[391], stage0_45[392], stage0_45[393], stage0_45[394], stage0_45[395], stage0_45[396]},
      {stage0_47[42], stage0_47[43], stage0_47[44], stage0_47[45], stage0_47[46], stage0_47[47]},
      {stage1_49[7],stage1_48[38],stage1_47[91],stage1_46[127],stage1_45[152]}
   );
   gpc606_5 gpc1742 (
      {stage0_45[397], stage0_45[398], stage0_45[399], stage0_45[400], stage0_45[401], stage0_45[402]},
      {stage0_47[48], stage0_47[49], stage0_47[50], stage0_47[51], stage0_47[52], stage0_47[53]},
      {stage1_49[8],stage1_48[39],stage1_47[92],stage1_46[128],stage1_45[153]}
   );
   gpc606_5 gpc1743 (
      {stage0_45[403], stage0_45[404], stage0_45[405], stage0_45[406], stage0_45[407], stage0_45[408]},
      {stage0_47[54], stage0_47[55], stage0_47[56], stage0_47[57], stage0_47[58], stage0_47[59]},
      {stage1_49[9],stage1_48[40],stage1_47[93],stage1_46[129],stage1_45[154]}
   );
   gpc606_5 gpc1744 (
      {stage0_45[409], stage0_45[410], stage0_45[411], stage0_45[412], stage0_45[413], stage0_45[414]},
      {stage0_47[60], stage0_47[61], stage0_47[62], stage0_47[63], stage0_47[64], stage0_47[65]},
      {stage1_49[10],stage1_48[41],stage1_47[94],stage1_46[130],stage1_45[155]}
   );
   gpc606_5 gpc1745 (
      {stage0_45[415], stage0_45[416], stage0_45[417], stage0_45[418], stage0_45[419], stage0_45[420]},
      {stage0_47[66], stage0_47[67], stage0_47[68], stage0_47[69], stage0_47[70], stage0_47[71]},
      {stage1_49[11],stage1_48[42],stage1_47[95],stage1_46[131],stage1_45[156]}
   );
   gpc606_5 gpc1746 (
      {stage0_45[421], stage0_45[422], stage0_45[423], stage0_45[424], stage0_45[425], stage0_45[426]},
      {stage0_47[72], stage0_47[73], stage0_47[74], stage0_47[75], stage0_47[76], stage0_47[77]},
      {stage1_49[12],stage1_48[43],stage1_47[96],stage1_46[132],stage1_45[157]}
   );
   gpc606_5 gpc1747 (
      {stage0_45[427], stage0_45[428], stage0_45[429], stage0_45[430], stage0_45[431], stage0_45[432]},
      {stage0_47[78], stage0_47[79], stage0_47[80], stage0_47[81], stage0_47[82], stage0_47[83]},
      {stage1_49[13],stage1_48[44],stage1_47[97],stage1_46[133],stage1_45[158]}
   );
   gpc135_4 gpc1748 (
      {stage0_46[186], stage0_46[187], stage0_46[188], stage0_46[189], stage0_46[190]},
      {stage0_47[84], stage0_47[85], stage0_47[86]},
      {stage0_48[0]},
      {stage1_49[14],stage1_48[45],stage1_47[98],stage1_46[134]}
   );
   gpc135_4 gpc1749 (
      {stage0_46[191], stage0_46[192], stage0_46[193], stage0_46[194], stage0_46[195]},
      {stage0_47[87], stage0_47[88], stage0_47[89]},
      {stage0_48[1]},
      {stage1_49[15],stage1_48[46],stage1_47[99],stage1_46[135]}
   );
   gpc135_4 gpc1750 (
      {stage0_46[196], stage0_46[197], stage0_46[198], stage0_46[199], stage0_46[200]},
      {stage0_47[90], stage0_47[91], stage0_47[92]},
      {stage0_48[2]},
      {stage1_49[16],stage1_48[47],stage1_47[100],stage1_46[136]}
   );
   gpc135_4 gpc1751 (
      {stage0_46[201], stage0_46[202], stage0_46[203], stage0_46[204], stage0_46[205]},
      {stage0_47[93], stage0_47[94], stage0_47[95]},
      {stage0_48[3]},
      {stage1_49[17],stage1_48[48],stage1_47[101],stage1_46[137]}
   );
   gpc135_4 gpc1752 (
      {stage0_46[206], stage0_46[207], stage0_46[208], stage0_46[209], stage0_46[210]},
      {stage0_47[96], stage0_47[97], stage0_47[98]},
      {stage0_48[4]},
      {stage1_49[18],stage1_48[49],stage1_47[102],stage1_46[138]}
   );
   gpc135_4 gpc1753 (
      {stage0_46[211], stage0_46[212], stage0_46[213], stage0_46[214], stage0_46[215]},
      {stage0_47[99], stage0_47[100], stage0_47[101]},
      {stage0_48[5]},
      {stage1_49[19],stage1_48[50],stage1_47[103],stage1_46[139]}
   );
   gpc135_4 gpc1754 (
      {stage0_46[216], stage0_46[217], stage0_46[218], stage0_46[219], stage0_46[220]},
      {stage0_47[102], stage0_47[103], stage0_47[104]},
      {stage0_48[6]},
      {stage1_49[20],stage1_48[51],stage1_47[104],stage1_46[140]}
   );
   gpc135_4 gpc1755 (
      {stage0_46[221], stage0_46[222], stage0_46[223], stage0_46[224], stage0_46[225]},
      {stage0_47[105], stage0_47[106], stage0_47[107]},
      {stage0_48[7]},
      {stage1_49[21],stage1_48[52],stage1_47[105],stage1_46[141]}
   );
   gpc135_4 gpc1756 (
      {stage0_46[226], stage0_46[227], stage0_46[228], stage0_46[229], stage0_46[230]},
      {stage0_47[108], stage0_47[109], stage0_47[110]},
      {stage0_48[8]},
      {stage1_49[22],stage1_48[53],stage1_47[106],stage1_46[142]}
   );
   gpc135_4 gpc1757 (
      {stage0_46[231], stage0_46[232], stage0_46[233], stage0_46[234], stage0_46[235]},
      {stage0_47[111], stage0_47[112], stage0_47[113]},
      {stage0_48[9]},
      {stage1_49[23],stage1_48[54],stage1_47[107],stage1_46[143]}
   );
   gpc615_5 gpc1758 (
      {stage0_46[236], stage0_46[237], stage0_46[238], stage0_46[239], stage0_46[240]},
      {stage0_47[114]},
      {stage0_48[10], stage0_48[11], stage0_48[12], stage0_48[13], stage0_48[14], stage0_48[15]},
      {stage1_50[0],stage1_49[24],stage1_48[55],stage1_47[108],stage1_46[144]}
   );
   gpc615_5 gpc1759 (
      {stage0_46[241], stage0_46[242], stage0_46[243], stage0_46[244], stage0_46[245]},
      {stage0_47[115]},
      {stage0_48[16], stage0_48[17], stage0_48[18], stage0_48[19], stage0_48[20], stage0_48[21]},
      {stage1_50[1],stage1_49[25],stage1_48[56],stage1_47[109],stage1_46[145]}
   );
   gpc615_5 gpc1760 (
      {stage0_46[246], stage0_46[247], stage0_46[248], stage0_46[249], stage0_46[250]},
      {stage0_47[116]},
      {stage0_48[22], stage0_48[23], stage0_48[24], stage0_48[25], stage0_48[26], stage0_48[27]},
      {stage1_50[2],stage1_49[26],stage1_48[57],stage1_47[110],stage1_46[146]}
   );
   gpc615_5 gpc1761 (
      {stage0_46[251], stage0_46[252], stage0_46[253], stage0_46[254], stage0_46[255]},
      {stage0_47[117]},
      {stage0_48[28], stage0_48[29], stage0_48[30], stage0_48[31], stage0_48[32], stage0_48[33]},
      {stage1_50[3],stage1_49[27],stage1_48[58],stage1_47[111],stage1_46[147]}
   );
   gpc615_5 gpc1762 (
      {stage0_46[256], stage0_46[257], stage0_46[258], stage0_46[259], stage0_46[260]},
      {stage0_47[118]},
      {stage0_48[34], stage0_48[35], stage0_48[36], stage0_48[37], stage0_48[38], stage0_48[39]},
      {stage1_50[4],stage1_49[28],stage1_48[59],stage1_47[112],stage1_46[148]}
   );
   gpc615_5 gpc1763 (
      {stage0_46[261], stage0_46[262], stage0_46[263], stage0_46[264], stage0_46[265]},
      {stage0_47[119]},
      {stage0_48[40], stage0_48[41], stage0_48[42], stage0_48[43], stage0_48[44], stage0_48[45]},
      {stage1_50[5],stage1_49[29],stage1_48[60],stage1_47[113],stage1_46[149]}
   );
   gpc615_5 gpc1764 (
      {stage0_46[266], stage0_46[267], stage0_46[268], stage0_46[269], stage0_46[270]},
      {stage0_47[120]},
      {stage0_48[46], stage0_48[47], stage0_48[48], stage0_48[49], stage0_48[50], stage0_48[51]},
      {stage1_50[6],stage1_49[30],stage1_48[61],stage1_47[114],stage1_46[150]}
   );
   gpc615_5 gpc1765 (
      {stage0_46[271], stage0_46[272], stage0_46[273], stage0_46[274], stage0_46[275]},
      {stage0_47[121]},
      {stage0_48[52], stage0_48[53], stage0_48[54], stage0_48[55], stage0_48[56], stage0_48[57]},
      {stage1_50[7],stage1_49[31],stage1_48[62],stage1_47[115],stage1_46[151]}
   );
   gpc615_5 gpc1766 (
      {stage0_46[276], stage0_46[277], stage0_46[278], stage0_46[279], stage0_46[280]},
      {stage0_47[122]},
      {stage0_48[58], stage0_48[59], stage0_48[60], stage0_48[61], stage0_48[62], stage0_48[63]},
      {stage1_50[8],stage1_49[32],stage1_48[63],stage1_47[116],stage1_46[152]}
   );
   gpc615_5 gpc1767 (
      {stage0_46[281], stage0_46[282], stage0_46[283], stage0_46[284], stage0_46[285]},
      {stage0_47[123]},
      {stage0_48[64], stage0_48[65], stage0_48[66], stage0_48[67], stage0_48[68], stage0_48[69]},
      {stage1_50[9],stage1_49[33],stage1_48[64],stage1_47[117],stage1_46[153]}
   );
   gpc615_5 gpc1768 (
      {stage0_46[286], stage0_46[287], stage0_46[288], stage0_46[289], stage0_46[290]},
      {stage0_47[124]},
      {stage0_48[70], stage0_48[71], stage0_48[72], stage0_48[73], stage0_48[74], stage0_48[75]},
      {stage1_50[10],stage1_49[34],stage1_48[65],stage1_47[118],stage1_46[154]}
   );
   gpc615_5 gpc1769 (
      {stage0_46[291], stage0_46[292], stage0_46[293], stage0_46[294], stage0_46[295]},
      {stage0_47[125]},
      {stage0_48[76], stage0_48[77], stage0_48[78], stage0_48[79], stage0_48[80], stage0_48[81]},
      {stage1_50[11],stage1_49[35],stage1_48[66],stage1_47[119],stage1_46[155]}
   );
   gpc615_5 gpc1770 (
      {stage0_46[296], stage0_46[297], stage0_46[298], stage0_46[299], stage0_46[300]},
      {stage0_47[126]},
      {stage0_48[82], stage0_48[83], stage0_48[84], stage0_48[85], stage0_48[86], stage0_48[87]},
      {stage1_50[12],stage1_49[36],stage1_48[67],stage1_47[120],stage1_46[156]}
   );
   gpc615_5 gpc1771 (
      {stage0_46[301], stage0_46[302], stage0_46[303], stage0_46[304], stage0_46[305]},
      {stage0_47[127]},
      {stage0_48[88], stage0_48[89], stage0_48[90], stage0_48[91], stage0_48[92], stage0_48[93]},
      {stage1_50[13],stage1_49[37],stage1_48[68],stage1_47[121],stage1_46[157]}
   );
   gpc615_5 gpc1772 (
      {stage0_46[306], stage0_46[307], stage0_46[308], stage0_46[309], stage0_46[310]},
      {stage0_47[128]},
      {stage0_48[94], stage0_48[95], stage0_48[96], stage0_48[97], stage0_48[98], stage0_48[99]},
      {stage1_50[14],stage1_49[38],stage1_48[69],stage1_47[122],stage1_46[158]}
   );
   gpc615_5 gpc1773 (
      {stage0_46[311], stage0_46[312], stage0_46[313], stage0_46[314], stage0_46[315]},
      {stage0_47[129]},
      {stage0_48[100], stage0_48[101], stage0_48[102], stage0_48[103], stage0_48[104], stage0_48[105]},
      {stage1_50[15],stage1_49[39],stage1_48[70],stage1_47[123],stage1_46[159]}
   );
   gpc615_5 gpc1774 (
      {stage0_46[316], stage0_46[317], stage0_46[318], stage0_46[319], stage0_46[320]},
      {stage0_47[130]},
      {stage0_48[106], stage0_48[107], stage0_48[108], stage0_48[109], stage0_48[110], stage0_48[111]},
      {stage1_50[16],stage1_49[40],stage1_48[71],stage1_47[124],stage1_46[160]}
   );
   gpc615_5 gpc1775 (
      {stage0_46[321], stage0_46[322], stage0_46[323], stage0_46[324], stage0_46[325]},
      {stage0_47[131]},
      {stage0_48[112], stage0_48[113], stage0_48[114], stage0_48[115], stage0_48[116], stage0_48[117]},
      {stage1_50[17],stage1_49[41],stage1_48[72],stage1_47[125],stage1_46[161]}
   );
   gpc615_5 gpc1776 (
      {stage0_46[326], stage0_46[327], stage0_46[328], stage0_46[329], stage0_46[330]},
      {stage0_47[132]},
      {stage0_48[118], stage0_48[119], stage0_48[120], stage0_48[121], stage0_48[122], stage0_48[123]},
      {stage1_50[18],stage1_49[42],stage1_48[73],stage1_47[126],stage1_46[162]}
   );
   gpc615_5 gpc1777 (
      {stage0_46[331], stage0_46[332], stage0_46[333], stage0_46[334], stage0_46[335]},
      {stage0_47[133]},
      {stage0_48[124], stage0_48[125], stage0_48[126], stage0_48[127], stage0_48[128], stage0_48[129]},
      {stage1_50[19],stage1_49[43],stage1_48[74],stage1_47[127],stage1_46[163]}
   );
   gpc615_5 gpc1778 (
      {stage0_46[336], stage0_46[337], stage0_46[338], stage0_46[339], stage0_46[340]},
      {stage0_47[134]},
      {stage0_48[130], stage0_48[131], stage0_48[132], stage0_48[133], stage0_48[134], stage0_48[135]},
      {stage1_50[20],stage1_49[44],stage1_48[75],stage1_47[128],stage1_46[164]}
   );
   gpc615_5 gpc1779 (
      {stage0_46[341], stage0_46[342], stage0_46[343], stage0_46[344], stage0_46[345]},
      {stage0_47[135]},
      {stage0_48[136], stage0_48[137], stage0_48[138], stage0_48[139], stage0_48[140], stage0_48[141]},
      {stage1_50[21],stage1_49[45],stage1_48[76],stage1_47[129],stage1_46[165]}
   );
   gpc615_5 gpc1780 (
      {stage0_46[346], stage0_46[347], stage0_46[348], stage0_46[349], stage0_46[350]},
      {stage0_47[136]},
      {stage0_48[142], stage0_48[143], stage0_48[144], stage0_48[145], stage0_48[146], stage0_48[147]},
      {stage1_50[22],stage1_49[46],stage1_48[77],stage1_47[130],stage1_46[166]}
   );
   gpc615_5 gpc1781 (
      {stage0_46[351], stage0_46[352], stage0_46[353], stage0_46[354], stage0_46[355]},
      {stage0_47[137]},
      {stage0_48[148], stage0_48[149], stage0_48[150], stage0_48[151], stage0_48[152], stage0_48[153]},
      {stage1_50[23],stage1_49[47],stage1_48[78],stage1_47[131],stage1_46[167]}
   );
   gpc615_5 gpc1782 (
      {stage0_47[138], stage0_47[139], stage0_47[140], stage0_47[141], stage0_47[142]},
      {stage0_48[154]},
      {stage0_49[0], stage0_49[1], stage0_49[2], stage0_49[3], stage0_49[4], stage0_49[5]},
      {stage1_51[0],stage1_50[24],stage1_49[48],stage1_48[79],stage1_47[132]}
   );
   gpc615_5 gpc1783 (
      {stage0_47[143], stage0_47[144], stage0_47[145], stage0_47[146], stage0_47[147]},
      {stage0_48[155]},
      {stage0_49[6], stage0_49[7], stage0_49[8], stage0_49[9], stage0_49[10], stage0_49[11]},
      {stage1_51[1],stage1_50[25],stage1_49[49],stage1_48[80],stage1_47[133]}
   );
   gpc615_5 gpc1784 (
      {stage0_47[148], stage0_47[149], stage0_47[150], stage0_47[151], stage0_47[152]},
      {stage0_48[156]},
      {stage0_49[12], stage0_49[13], stage0_49[14], stage0_49[15], stage0_49[16], stage0_49[17]},
      {stage1_51[2],stage1_50[26],stage1_49[50],stage1_48[81],stage1_47[134]}
   );
   gpc615_5 gpc1785 (
      {stage0_47[153], stage0_47[154], stage0_47[155], stage0_47[156], stage0_47[157]},
      {stage0_48[157]},
      {stage0_49[18], stage0_49[19], stage0_49[20], stage0_49[21], stage0_49[22], stage0_49[23]},
      {stage1_51[3],stage1_50[27],stage1_49[51],stage1_48[82],stage1_47[135]}
   );
   gpc615_5 gpc1786 (
      {stage0_47[158], stage0_47[159], stage0_47[160], stage0_47[161], stage0_47[162]},
      {stage0_48[158]},
      {stage0_49[24], stage0_49[25], stage0_49[26], stage0_49[27], stage0_49[28], stage0_49[29]},
      {stage1_51[4],stage1_50[28],stage1_49[52],stage1_48[83],stage1_47[136]}
   );
   gpc615_5 gpc1787 (
      {stage0_47[163], stage0_47[164], stage0_47[165], stage0_47[166], stage0_47[167]},
      {stage0_48[159]},
      {stage0_49[30], stage0_49[31], stage0_49[32], stage0_49[33], stage0_49[34], stage0_49[35]},
      {stage1_51[5],stage1_50[29],stage1_49[53],stage1_48[84],stage1_47[137]}
   );
   gpc615_5 gpc1788 (
      {stage0_47[168], stage0_47[169], stage0_47[170], stage0_47[171], stage0_47[172]},
      {stage0_48[160]},
      {stage0_49[36], stage0_49[37], stage0_49[38], stage0_49[39], stage0_49[40], stage0_49[41]},
      {stage1_51[6],stage1_50[30],stage1_49[54],stage1_48[85],stage1_47[138]}
   );
   gpc615_5 gpc1789 (
      {stage0_47[173], stage0_47[174], stage0_47[175], stage0_47[176], stage0_47[177]},
      {stage0_48[161]},
      {stage0_49[42], stage0_49[43], stage0_49[44], stage0_49[45], stage0_49[46], stage0_49[47]},
      {stage1_51[7],stage1_50[31],stage1_49[55],stage1_48[86],stage1_47[139]}
   );
   gpc615_5 gpc1790 (
      {stage0_47[178], stage0_47[179], stage0_47[180], stage0_47[181], stage0_47[182]},
      {stage0_48[162]},
      {stage0_49[48], stage0_49[49], stage0_49[50], stage0_49[51], stage0_49[52], stage0_49[53]},
      {stage1_51[8],stage1_50[32],stage1_49[56],stage1_48[87],stage1_47[140]}
   );
   gpc615_5 gpc1791 (
      {stage0_47[183], stage0_47[184], stage0_47[185], stage0_47[186], stage0_47[187]},
      {stage0_48[163]},
      {stage0_49[54], stage0_49[55], stage0_49[56], stage0_49[57], stage0_49[58], stage0_49[59]},
      {stage1_51[9],stage1_50[33],stage1_49[57],stage1_48[88],stage1_47[141]}
   );
   gpc615_5 gpc1792 (
      {stage0_47[188], stage0_47[189], stage0_47[190], stage0_47[191], stage0_47[192]},
      {stage0_48[164]},
      {stage0_49[60], stage0_49[61], stage0_49[62], stage0_49[63], stage0_49[64], stage0_49[65]},
      {stage1_51[10],stage1_50[34],stage1_49[58],stage1_48[89],stage1_47[142]}
   );
   gpc615_5 gpc1793 (
      {stage0_47[193], stage0_47[194], stage0_47[195], stage0_47[196], stage0_47[197]},
      {stage0_48[165]},
      {stage0_49[66], stage0_49[67], stage0_49[68], stage0_49[69], stage0_49[70], stage0_49[71]},
      {stage1_51[11],stage1_50[35],stage1_49[59],stage1_48[90],stage1_47[143]}
   );
   gpc615_5 gpc1794 (
      {stage0_47[198], stage0_47[199], stage0_47[200], stage0_47[201], stage0_47[202]},
      {stage0_48[166]},
      {stage0_49[72], stage0_49[73], stage0_49[74], stage0_49[75], stage0_49[76], stage0_49[77]},
      {stage1_51[12],stage1_50[36],stage1_49[60],stage1_48[91],stage1_47[144]}
   );
   gpc615_5 gpc1795 (
      {stage0_47[203], stage0_47[204], stage0_47[205], stage0_47[206], stage0_47[207]},
      {stage0_48[167]},
      {stage0_49[78], stage0_49[79], stage0_49[80], stage0_49[81], stage0_49[82], stage0_49[83]},
      {stage1_51[13],stage1_50[37],stage1_49[61],stage1_48[92],stage1_47[145]}
   );
   gpc615_5 gpc1796 (
      {stage0_47[208], stage0_47[209], stage0_47[210], stage0_47[211], stage0_47[212]},
      {stage0_48[168]},
      {stage0_49[84], stage0_49[85], stage0_49[86], stage0_49[87], stage0_49[88], stage0_49[89]},
      {stage1_51[14],stage1_50[38],stage1_49[62],stage1_48[93],stage1_47[146]}
   );
   gpc615_5 gpc1797 (
      {stage0_47[213], stage0_47[214], stage0_47[215], stage0_47[216], stage0_47[217]},
      {stage0_48[169]},
      {stage0_49[90], stage0_49[91], stage0_49[92], stage0_49[93], stage0_49[94], stage0_49[95]},
      {stage1_51[15],stage1_50[39],stage1_49[63],stage1_48[94],stage1_47[147]}
   );
   gpc615_5 gpc1798 (
      {stage0_47[218], stage0_47[219], stage0_47[220], stage0_47[221], stage0_47[222]},
      {stage0_48[170]},
      {stage0_49[96], stage0_49[97], stage0_49[98], stage0_49[99], stage0_49[100], stage0_49[101]},
      {stage1_51[16],stage1_50[40],stage1_49[64],stage1_48[95],stage1_47[148]}
   );
   gpc615_5 gpc1799 (
      {stage0_47[223], stage0_47[224], stage0_47[225], stage0_47[226], stage0_47[227]},
      {stage0_48[171]},
      {stage0_49[102], stage0_49[103], stage0_49[104], stage0_49[105], stage0_49[106], stage0_49[107]},
      {stage1_51[17],stage1_50[41],stage1_49[65],stage1_48[96],stage1_47[149]}
   );
   gpc615_5 gpc1800 (
      {stage0_47[228], stage0_47[229], stage0_47[230], stage0_47[231], stage0_47[232]},
      {stage0_48[172]},
      {stage0_49[108], stage0_49[109], stage0_49[110], stage0_49[111], stage0_49[112], stage0_49[113]},
      {stage1_51[18],stage1_50[42],stage1_49[66],stage1_48[97],stage1_47[150]}
   );
   gpc615_5 gpc1801 (
      {stage0_47[233], stage0_47[234], stage0_47[235], stage0_47[236], stage0_47[237]},
      {stage0_48[173]},
      {stage0_49[114], stage0_49[115], stage0_49[116], stage0_49[117], stage0_49[118], stage0_49[119]},
      {stage1_51[19],stage1_50[43],stage1_49[67],stage1_48[98],stage1_47[151]}
   );
   gpc615_5 gpc1802 (
      {stage0_47[238], stage0_47[239], stage0_47[240], stage0_47[241], stage0_47[242]},
      {stage0_48[174]},
      {stage0_49[120], stage0_49[121], stage0_49[122], stage0_49[123], stage0_49[124], stage0_49[125]},
      {stage1_51[20],stage1_50[44],stage1_49[68],stage1_48[99],stage1_47[152]}
   );
   gpc615_5 gpc1803 (
      {stage0_47[243], stage0_47[244], stage0_47[245], stage0_47[246], stage0_47[247]},
      {stage0_48[175]},
      {stage0_49[126], stage0_49[127], stage0_49[128], stage0_49[129], stage0_49[130], stage0_49[131]},
      {stage1_51[21],stage1_50[45],stage1_49[69],stage1_48[100],stage1_47[153]}
   );
   gpc615_5 gpc1804 (
      {stage0_47[248], stage0_47[249], stage0_47[250], stage0_47[251], stage0_47[252]},
      {stage0_48[176]},
      {stage0_49[132], stage0_49[133], stage0_49[134], stage0_49[135], stage0_49[136], stage0_49[137]},
      {stage1_51[22],stage1_50[46],stage1_49[70],stage1_48[101],stage1_47[154]}
   );
   gpc615_5 gpc1805 (
      {stage0_47[253], stage0_47[254], stage0_47[255], stage0_47[256], stage0_47[257]},
      {stage0_48[177]},
      {stage0_49[138], stage0_49[139], stage0_49[140], stage0_49[141], stage0_49[142], stage0_49[143]},
      {stage1_51[23],stage1_50[47],stage1_49[71],stage1_48[102],stage1_47[155]}
   );
   gpc615_5 gpc1806 (
      {stage0_47[258], stage0_47[259], stage0_47[260], stage0_47[261], stage0_47[262]},
      {stage0_48[178]},
      {stage0_49[144], stage0_49[145], stage0_49[146], stage0_49[147], stage0_49[148], stage0_49[149]},
      {stage1_51[24],stage1_50[48],stage1_49[72],stage1_48[103],stage1_47[156]}
   );
   gpc615_5 gpc1807 (
      {stage0_47[263], stage0_47[264], stage0_47[265], stage0_47[266], stage0_47[267]},
      {stage0_48[179]},
      {stage0_49[150], stage0_49[151], stage0_49[152], stage0_49[153], stage0_49[154], stage0_49[155]},
      {stage1_51[25],stage1_50[49],stage1_49[73],stage1_48[104],stage1_47[157]}
   );
   gpc615_5 gpc1808 (
      {stage0_47[268], stage0_47[269], stage0_47[270], stage0_47[271], stage0_47[272]},
      {stage0_48[180]},
      {stage0_49[156], stage0_49[157], stage0_49[158], stage0_49[159], stage0_49[160], stage0_49[161]},
      {stage1_51[26],stage1_50[50],stage1_49[74],stage1_48[105],stage1_47[158]}
   );
   gpc615_5 gpc1809 (
      {stage0_47[273], stage0_47[274], stage0_47[275], stage0_47[276], stage0_47[277]},
      {stage0_48[181]},
      {stage0_49[162], stage0_49[163], stage0_49[164], stage0_49[165], stage0_49[166], stage0_49[167]},
      {stage1_51[27],stage1_50[51],stage1_49[75],stage1_48[106],stage1_47[159]}
   );
   gpc615_5 gpc1810 (
      {stage0_47[278], stage0_47[279], stage0_47[280], stage0_47[281], stage0_47[282]},
      {stage0_48[182]},
      {stage0_49[168], stage0_49[169], stage0_49[170], stage0_49[171], stage0_49[172], stage0_49[173]},
      {stage1_51[28],stage1_50[52],stage1_49[76],stage1_48[107],stage1_47[160]}
   );
   gpc615_5 gpc1811 (
      {stage0_47[283], stage0_47[284], stage0_47[285], stage0_47[286], stage0_47[287]},
      {stage0_48[183]},
      {stage0_49[174], stage0_49[175], stage0_49[176], stage0_49[177], stage0_49[178], stage0_49[179]},
      {stage1_51[29],stage1_50[53],stage1_49[77],stage1_48[108],stage1_47[161]}
   );
   gpc615_5 gpc1812 (
      {stage0_47[288], stage0_47[289], stage0_47[290], stage0_47[291], stage0_47[292]},
      {stage0_48[184]},
      {stage0_49[180], stage0_49[181], stage0_49[182], stage0_49[183], stage0_49[184], stage0_49[185]},
      {stage1_51[30],stage1_50[54],stage1_49[78],stage1_48[109],stage1_47[162]}
   );
   gpc615_5 gpc1813 (
      {stage0_47[293], stage0_47[294], stage0_47[295], stage0_47[296], stage0_47[297]},
      {stage0_48[185]},
      {stage0_49[186], stage0_49[187], stage0_49[188], stage0_49[189], stage0_49[190], stage0_49[191]},
      {stage1_51[31],stage1_50[55],stage1_49[79],stage1_48[110],stage1_47[163]}
   );
   gpc615_5 gpc1814 (
      {stage0_47[298], stage0_47[299], stage0_47[300], stage0_47[301], stage0_47[302]},
      {stage0_48[186]},
      {stage0_49[192], stage0_49[193], stage0_49[194], stage0_49[195], stage0_49[196], stage0_49[197]},
      {stage1_51[32],stage1_50[56],stage1_49[80],stage1_48[111],stage1_47[164]}
   );
   gpc615_5 gpc1815 (
      {stage0_47[303], stage0_47[304], stage0_47[305], stage0_47[306], stage0_47[307]},
      {stage0_48[187]},
      {stage0_49[198], stage0_49[199], stage0_49[200], stage0_49[201], stage0_49[202], stage0_49[203]},
      {stage1_51[33],stage1_50[57],stage1_49[81],stage1_48[112],stage1_47[165]}
   );
   gpc615_5 gpc1816 (
      {stage0_47[308], stage0_47[309], stage0_47[310], stage0_47[311], stage0_47[312]},
      {stage0_48[188]},
      {stage0_49[204], stage0_49[205], stage0_49[206], stage0_49[207], stage0_49[208], stage0_49[209]},
      {stage1_51[34],stage1_50[58],stage1_49[82],stage1_48[113],stage1_47[166]}
   );
   gpc615_5 gpc1817 (
      {stage0_47[313], stage0_47[314], stage0_47[315], stage0_47[316], stage0_47[317]},
      {stage0_48[189]},
      {stage0_49[210], stage0_49[211], stage0_49[212], stage0_49[213], stage0_49[214], stage0_49[215]},
      {stage1_51[35],stage1_50[59],stage1_49[83],stage1_48[114],stage1_47[167]}
   );
   gpc615_5 gpc1818 (
      {stage0_47[318], stage0_47[319], stage0_47[320], stage0_47[321], stage0_47[322]},
      {stage0_48[190]},
      {stage0_49[216], stage0_49[217], stage0_49[218], stage0_49[219], stage0_49[220], stage0_49[221]},
      {stage1_51[36],stage1_50[60],stage1_49[84],stage1_48[115],stage1_47[168]}
   );
   gpc615_5 gpc1819 (
      {stage0_47[323], stage0_47[324], stage0_47[325], stage0_47[326], stage0_47[327]},
      {stage0_48[191]},
      {stage0_49[222], stage0_49[223], stage0_49[224], stage0_49[225], stage0_49[226], stage0_49[227]},
      {stage1_51[37],stage1_50[61],stage1_49[85],stage1_48[116],stage1_47[169]}
   );
   gpc615_5 gpc1820 (
      {stage0_47[328], stage0_47[329], stage0_47[330], stage0_47[331], stage0_47[332]},
      {stage0_48[192]},
      {stage0_49[228], stage0_49[229], stage0_49[230], stage0_49[231], stage0_49[232], stage0_49[233]},
      {stage1_51[38],stage1_50[62],stage1_49[86],stage1_48[117],stage1_47[170]}
   );
   gpc615_5 gpc1821 (
      {stage0_47[333], stage0_47[334], stage0_47[335], stage0_47[336], stage0_47[337]},
      {stage0_48[193]},
      {stage0_49[234], stage0_49[235], stage0_49[236], stage0_49[237], stage0_49[238], stage0_49[239]},
      {stage1_51[39],stage1_50[63],stage1_49[87],stage1_48[118],stage1_47[171]}
   );
   gpc615_5 gpc1822 (
      {stage0_47[338], stage0_47[339], stage0_47[340], stage0_47[341], stage0_47[342]},
      {stage0_48[194]},
      {stage0_49[240], stage0_49[241], stage0_49[242], stage0_49[243], stage0_49[244], stage0_49[245]},
      {stage1_51[40],stage1_50[64],stage1_49[88],stage1_48[119],stage1_47[172]}
   );
   gpc615_5 gpc1823 (
      {stage0_47[343], stage0_47[344], stage0_47[345], stage0_47[346], stage0_47[347]},
      {stage0_48[195]},
      {stage0_49[246], stage0_49[247], stage0_49[248], stage0_49[249], stage0_49[250], stage0_49[251]},
      {stage1_51[41],stage1_50[65],stage1_49[89],stage1_48[120],stage1_47[173]}
   );
   gpc615_5 gpc1824 (
      {stage0_47[348], stage0_47[349], stage0_47[350], stage0_47[351], stage0_47[352]},
      {stage0_48[196]},
      {stage0_49[252], stage0_49[253], stage0_49[254], stage0_49[255], stage0_49[256], stage0_49[257]},
      {stage1_51[42],stage1_50[66],stage1_49[90],stage1_48[121],stage1_47[174]}
   );
   gpc615_5 gpc1825 (
      {stage0_47[353], stage0_47[354], stage0_47[355], stage0_47[356], stage0_47[357]},
      {stage0_48[197]},
      {stage0_49[258], stage0_49[259], stage0_49[260], stage0_49[261], stage0_49[262], stage0_49[263]},
      {stage1_51[43],stage1_50[67],stage1_49[91],stage1_48[122],stage1_47[175]}
   );
   gpc615_5 gpc1826 (
      {stage0_47[358], stage0_47[359], stage0_47[360], stage0_47[361], stage0_47[362]},
      {stage0_48[198]},
      {stage0_49[264], stage0_49[265], stage0_49[266], stage0_49[267], stage0_49[268], stage0_49[269]},
      {stage1_51[44],stage1_50[68],stage1_49[92],stage1_48[123],stage1_47[176]}
   );
   gpc615_5 gpc1827 (
      {stage0_47[363], stage0_47[364], stage0_47[365], stage0_47[366], stage0_47[367]},
      {stage0_48[199]},
      {stage0_49[270], stage0_49[271], stage0_49[272], stage0_49[273], stage0_49[274], stage0_49[275]},
      {stage1_51[45],stage1_50[69],stage1_49[93],stage1_48[124],stage1_47[177]}
   );
   gpc615_5 gpc1828 (
      {stage0_47[368], stage0_47[369], stage0_47[370], stage0_47[371], stage0_47[372]},
      {stage0_48[200]},
      {stage0_49[276], stage0_49[277], stage0_49[278], stage0_49[279], stage0_49[280], stage0_49[281]},
      {stage1_51[46],stage1_50[70],stage1_49[94],stage1_48[125],stage1_47[178]}
   );
   gpc615_5 gpc1829 (
      {stage0_47[373], stage0_47[374], stage0_47[375], stage0_47[376], stage0_47[377]},
      {stage0_48[201]},
      {stage0_49[282], stage0_49[283], stage0_49[284], stage0_49[285], stage0_49[286], stage0_49[287]},
      {stage1_51[47],stage1_50[71],stage1_49[95],stage1_48[126],stage1_47[179]}
   );
   gpc615_5 gpc1830 (
      {stage0_47[378], stage0_47[379], stage0_47[380], stage0_47[381], stage0_47[382]},
      {stage0_48[202]},
      {stage0_49[288], stage0_49[289], stage0_49[290], stage0_49[291], stage0_49[292], stage0_49[293]},
      {stage1_51[48],stage1_50[72],stage1_49[96],stage1_48[127],stage1_47[180]}
   );
   gpc615_5 gpc1831 (
      {stage0_47[383], stage0_47[384], stage0_47[385], stage0_47[386], stage0_47[387]},
      {stage0_48[203]},
      {stage0_49[294], stage0_49[295], stage0_49[296], stage0_49[297], stage0_49[298], stage0_49[299]},
      {stage1_51[49],stage1_50[73],stage1_49[97],stage1_48[128],stage1_47[181]}
   );
   gpc615_5 gpc1832 (
      {stage0_47[388], stage0_47[389], stage0_47[390], stage0_47[391], stage0_47[392]},
      {stage0_48[204]},
      {stage0_49[300], stage0_49[301], stage0_49[302], stage0_49[303], stage0_49[304], stage0_49[305]},
      {stage1_51[50],stage1_50[74],stage1_49[98],stage1_48[129],stage1_47[182]}
   );
   gpc615_5 gpc1833 (
      {stage0_47[393], stage0_47[394], stage0_47[395], stage0_47[396], stage0_47[397]},
      {stage0_48[205]},
      {stage0_49[306], stage0_49[307], stage0_49[308], stage0_49[309], stage0_49[310], stage0_49[311]},
      {stage1_51[51],stage1_50[75],stage1_49[99],stage1_48[130],stage1_47[183]}
   );
   gpc615_5 gpc1834 (
      {stage0_47[398], stage0_47[399], stage0_47[400], stage0_47[401], stage0_47[402]},
      {stage0_48[206]},
      {stage0_49[312], stage0_49[313], stage0_49[314], stage0_49[315], stage0_49[316], stage0_49[317]},
      {stage1_51[52],stage1_50[76],stage1_49[100],stage1_48[131],stage1_47[184]}
   );
   gpc615_5 gpc1835 (
      {stage0_47[403], stage0_47[404], stage0_47[405], stage0_47[406], stage0_47[407]},
      {stage0_48[207]},
      {stage0_49[318], stage0_49[319], stage0_49[320], stage0_49[321], stage0_49[322], stage0_49[323]},
      {stage1_51[53],stage1_50[77],stage1_49[101],stage1_48[132],stage1_47[185]}
   );
   gpc615_5 gpc1836 (
      {stage0_47[408], stage0_47[409], stage0_47[410], stage0_47[411], stage0_47[412]},
      {stage0_48[208]},
      {stage0_49[324], stage0_49[325], stage0_49[326], stage0_49[327], stage0_49[328], stage0_49[329]},
      {stage1_51[54],stage1_50[78],stage1_49[102],stage1_48[133],stage1_47[186]}
   );
   gpc615_5 gpc1837 (
      {stage0_47[413], stage0_47[414], stage0_47[415], stage0_47[416], stage0_47[417]},
      {stage0_48[209]},
      {stage0_49[330], stage0_49[331], stage0_49[332], stage0_49[333], stage0_49[334], stage0_49[335]},
      {stage1_51[55],stage1_50[79],stage1_49[103],stage1_48[134],stage1_47[187]}
   );
   gpc615_5 gpc1838 (
      {stage0_47[418], stage0_47[419], stage0_47[420], stage0_47[421], stage0_47[422]},
      {stage0_48[210]},
      {stage0_49[336], stage0_49[337], stage0_49[338], stage0_49[339], stage0_49[340], stage0_49[341]},
      {stage1_51[56],stage1_50[80],stage1_49[104],stage1_48[135],stage1_47[188]}
   );
   gpc615_5 gpc1839 (
      {stage0_47[423], stage0_47[424], stage0_47[425], stage0_47[426], stage0_47[427]},
      {stage0_48[211]},
      {stage0_49[342], stage0_49[343], stage0_49[344], stage0_49[345], stage0_49[346], stage0_49[347]},
      {stage1_51[57],stage1_50[81],stage1_49[105],stage1_48[136],stage1_47[189]}
   );
   gpc615_5 gpc1840 (
      {stage0_47[428], stage0_47[429], stage0_47[430], stage0_47[431], stage0_47[432]},
      {stage0_48[212]},
      {stage0_49[348], stage0_49[349], stage0_49[350], stage0_49[351], stage0_49[352], stage0_49[353]},
      {stage1_51[58],stage1_50[82],stage1_49[106],stage1_48[137],stage1_47[190]}
   );
   gpc615_5 gpc1841 (
      {stage0_47[433], stage0_47[434], stage0_47[435], stage0_47[436], stage0_47[437]},
      {stage0_48[213]},
      {stage0_49[354], stage0_49[355], stage0_49[356], stage0_49[357], stage0_49[358], stage0_49[359]},
      {stage1_51[59],stage1_50[83],stage1_49[107],stage1_48[138],stage1_47[191]}
   );
   gpc615_5 gpc1842 (
      {stage0_47[438], stage0_47[439], stage0_47[440], stage0_47[441], stage0_47[442]},
      {stage0_48[214]},
      {stage0_49[360], stage0_49[361], stage0_49[362], stage0_49[363], stage0_49[364], stage0_49[365]},
      {stage1_51[60],stage1_50[84],stage1_49[108],stage1_48[139],stage1_47[192]}
   );
   gpc606_5 gpc1843 (
      {stage0_48[215], stage0_48[216], stage0_48[217], stage0_48[218], stage0_48[219], stage0_48[220]},
      {stage0_50[0], stage0_50[1], stage0_50[2], stage0_50[3], stage0_50[4], stage0_50[5]},
      {stage1_52[0],stage1_51[61],stage1_50[85],stage1_49[109],stage1_48[140]}
   );
   gpc606_5 gpc1844 (
      {stage0_48[221], stage0_48[222], stage0_48[223], stage0_48[224], stage0_48[225], stage0_48[226]},
      {stage0_50[6], stage0_50[7], stage0_50[8], stage0_50[9], stage0_50[10], stage0_50[11]},
      {stage1_52[1],stage1_51[62],stage1_50[86],stage1_49[110],stage1_48[141]}
   );
   gpc606_5 gpc1845 (
      {stage0_48[227], stage0_48[228], stage0_48[229], stage0_48[230], stage0_48[231], stage0_48[232]},
      {stage0_50[12], stage0_50[13], stage0_50[14], stage0_50[15], stage0_50[16], stage0_50[17]},
      {stage1_52[2],stage1_51[63],stage1_50[87],stage1_49[111],stage1_48[142]}
   );
   gpc606_5 gpc1846 (
      {stage0_48[233], stage0_48[234], stage0_48[235], stage0_48[236], stage0_48[237], stage0_48[238]},
      {stage0_50[18], stage0_50[19], stage0_50[20], stage0_50[21], stage0_50[22], stage0_50[23]},
      {stage1_52[3],stage1_51[64],stage1_50[88],stage1_49[112],stage1_48[143]}
   );
   gpc606_5 gpc1847 (
      {stage0_48[239], stage0_48[240], stage0_48[241], stage0_48[242], stage0_48[243], stage0_48[244]},
      {stage0_50[24], stage0_50[25], stage0_50[26], stage0_50[27], stage0_50[28], stage0_50[29]},
      {stage1_52[4],stage1_51[65],stage1_50[89],stage1_49[113],stage1_48[144]}
   );
   gpc606_5 gpc1848 (
      {stage0_48[245], stage0_48[246], stage0_48[247], stage0_48[248], stage0_48[249], stage0_48[250]},
      {stage0_50[30], stage0_50[31], stage0_50[32], stage0_50[33], stage0_50[34], stage0_50[35]},
      {stage1_52[5],stage1_51[66],stage1_50[90],stage1_49[114],stage1_48[145]}
   );
   gpc606_5 gpc1849 (
      {stage0_48[251], stage0_48[252], stage0_48[253], stage0_48[254], stage0_48[255], stage0_48[256]},
      {stage0_50[36], stage0_50[37], stage0_50[38], stage0_50[39], stage0_50[40], stage0_50[41]},
      {stage1_52[6],stage1_51[67],stage1_50[91],stage1_49[115],stage1_48[146]}
   );
   gpc606_5 gpc1850 (
      {stage0_48[257], stage0_48[258], stage0_48[259], stage0_48[260], stage0_48[261], stage0_48[262]},
      {stage0_50[42], stage0_50[43], stage0_50[44], stage0_50[45], stage0_50[46], stage0_50[47]},
      {stage1_52[7],stage1_51[68],stage1_50[92],stage1_49[116],stage1_48[147]}
   );
   gpc606_5 gpc1851 (
      {stage0_48[263], stage0_48[264], stage0_48[265], stage0_48[266], stage0_48[267], stage0_48[268]},
      {stage0_50[48], stage0_50[49], stage0_50[50], stage0_50[51], stage0_50[52], stage0_50[53]},
      {stage1_52[8],stage1_51[69],stage1_50[93],stage1_49[117],stage1_48[148]}
   );
   gpc606_5 gpc1852 (
      {stage0_48[269], stage0_48[270], stage0_48[271], stage0_48[272], stage0_48[273], stage0_48[274]},
      {stage0_50[54], stage0_50[55], stage0_50[56], stage0_50[57], stage0_50[58], stage0_50[59]},
      {stage1_52[9],stage1_51[70],stage1_50[94],stage1_49[118],stage1_48[149]}
   );
   gpc606_5 gpc1853 (
      {stage0_48[275], stage0_48[276], stage0_48[277], stage0_48[278], stage0_48[279], stage0_48[280]},
      {stage0_50[60], stage0_50[61], stage0_50[62], stage0_50[63], stage0_50[64], stage0_50[65]},
      {stage1_52[10],stage1_51[71],stage1_50[95],stage1_49[119],stage1_48[150]}
   );
   gpc606_5 gpc1854 (
      {stage0_48[281], stage0_48[282], stage0_48[283], stage0_48[284], stage0_48[285], stage0_48[286]},
      {stage0_50[66], stage0_50[67], stage0_50[68], stage0_50[69], stage0_50[70], stage0_50[71]},
      {stage1_52[11],stage1_51[72],stage1_50[96],stage1_49[120],stage1_48[151]}
   );
   gpc606_5 gpc1855 (
      {stage0_48[287], stage0_48[288], stage0_48[289], stage0_48[290], stage0_48[291], stage0_48[292]},
      {stage0_50[72], stage0_50[73], stage0_50[74], stage0_50[75], stage0_50[76], stage0_50[77]},
      {stage1_52[12],stage1_51[73],stage1_50[97],stage1_49[121],stage1_48[152]}
   );
   gpc615_5 gpc1856 (
      {stage0_48[293], stage0_48[294], stage0_48[295], stage0_48[296], stage0_48[297]},
      {stage0_49[366]},
      {stage0_50[78], stage0_50[79], stage0_50[80], stage0_50[81], stage0_50[82], stage0_50[83]},
      {stage1_52[13],stage1_51[74],stage1_50[98],stage1_49[122],stage1_48[153]}
   );
   gpc615_5 gpc1857 (
      {stage0_48[298], stage0_48[299], stage0_48[300], stage0_48[301], stage0_48[302]},
      {stage0_49[367]},
      {stage0_50[84], stage0_50[85], stage0_50[86], stage0_50[87], stage0_50[88], stage0_50[89]},
      {stage1_52[14],stage1_51[75],stage1_50[99],stage1_49[123],stage1_48[154]}
   );
   gpc615_5 gpc1858 (
      {stage0_48[303], stage0_48[304], stage0_48[305], stage0_48[306], stage0_48[307]},
      {stage0_49[368]},
      {stage0_50[90], stage0_50[91], stage0_50[92], stage0_50[93], stage0_50[94], stage0_50[95]},
      {stage1_52[15],stage1_51[76],stage1_50[100],stage1_49[124],stage1_48[155]}
   );
   gpc615_5 gpc1859 (
      {stage0_48[308], stage0_48[309], stage0_48[310], stage0_48[311], stage0_48[312]},
      {stage0_49[369]},
      {stage0_50[96], stage0_50[97], stage0_50[98], stage0_50[99], stage0_50[100], stage0_50[101]},
      {stage1_52[16],stage1_51[77],stage1_50[101],stage1_49[125],stage1_48[156]}
   );
   gpc615_5 gpc1860 (
      {stage0_48[313], stage0_48[314], stage0_48[315], stage0_48[316], stage0_48[317]},
      {stage0_49[370]},
      {stage0_50[102], stage0_50[103], stage0_50[104], stage0_50[105], stage0_50[106], stage0_50[107]},
      {stage1_52[17],stage1_51[78],stage1_50[102],stage1_49[126],stage1_48[157]}
   );
   gpc615_5 gpc1861 (
      {stage0_48[318], stage0_48[319], stage0_48[320], stage0_48[321], stage0_48[322]},
      {stage0_49[371]},
      {stage0_50[108], stage0_50[109], stage0_50[110], stage0_50[111], stage0_50[112], stage0_50[113]},
      {stage1_52[18],stage1_51[79],stage1_50[103],stage1_49[127],stage1_48[158]}
   );
   gpc615_5 gpc1862 (
      {stage0_48[323], stage0_48[324], stage0_48[325], stage0_48[326], stage0_48[327]},
      {stage0_49[372]},
      {stage0_50[114], stage0_50[115], stage0_50[116], stage0_50[117], stage0_50[118], stage0_50[119]},
      {stage1_52[19],stage1_51[80],stage1_50[104],stage1_49[128],stage1_48[159]}
   );
   gpc615_5 gpc1863 (
      {stage0_48[328], stage0_48[329], stage0_48[330], stage0_48[331], stage0_48[332]},
      {stage0_49[373]},
      {stage0_50[120], stage0_50[121], stage0_50[122], stage0_50[123], stage0_50[124], stage0_50[125]},
      {stage1_52[20],stage1_51[81],stage1_50[105],stage1_49[129],stage1_48[160]}
   );
   gpc615_5 gpc1864 (
      {stage0_48[333], stage0_48[334], stage0_48[335], stage0_48[336], stage0_48[337]},
      {stage0_49[374]},
      {stage0_50[126], stage0_50[127], stage0_50[128], stage0_50[129], stage0_50[130], stage0_50[131]},
      {stage1_52[21],stage1_51[82],stage1_50[106],stage1_49[130],stage1_48[161]}
   );
   gpc615_5 gpc1865 (
      {stage0_48[338], stage0_48[339], stage0_48[340], stage0_48[341], stage0_48[342]},
      {stage0_49[375]},
      {stage0_50[132], stage0_50[133], stage0_50[134], stage0_50[135], stage0_50[136], stage0_50[137]},
      {stage1_52[22],stage1_51[83],stage1_50[107],stage1_49[131],stage1_48[162]}
   );
   gpc615_5 gpc1866 (
      {stage0_48[343], stage0_48[344], stage0_48[345], stage0_48[346], stage0_48[347]},
      {stage0_49[376]},
      {stage0_50[138], stage0_50[139], stage0_50[140], stage0_50[141], stage0_50[142], stage0_50[143]},
      {stage1_52[23],stage1_51[84],stage1_50[108],stage1_49[132],stage1_48[163]}
   );
   gpc615_5 gpc1867 (
      {stage0_48[348], stage0_48[349], stage0_48[350], stage0_48[351], stage0_48[352]},
      {stage0_49[377]},
      {stage0_50[144], stage0_50[145], stage0_50[146], stage0_50[147], stage0_50[148], stage0_50[149]},
      {stage1_52[24],stage1_51[85],stage1_50[109],stage1_49[133],stage1_48[164]}
   );
   gpc615_5 gpc1868 (
      {stage0_48[353], stage0_48[354], stage0_48[355], stage0_48[356], stage0_48[357]},
      {stage0_49[378]},
      {stage0_50[150], stage0_50[151], stage0_50[152], stage0_50[153], stage0_50[154], stage0_50[155]},
      {stage1_52[25],stage1_51[86],stage1_50[110],stage1_49[134],stage1_48[165]}
   );
   gpc615_5 gpc1869 (
      {stage0_48[358], stage0_48[359], stage0_48[360], stage0_48[361], stage0_48[362]},
      {stage0_49[379]},
      {stage0_50[156], stage0_50[157], stage0_50[158], stage0_50[159], stage0_50[160], stage0_50[161]},
      {stage1_52[26],stage1_51[87],stage1_50[111],stage1_49[135],stage1_48[166]}
   );
   gpc615_5 gpc1870 (
      {stage0_48[363], stage0_48[364], stage0_48[365], stage0_48[366], stage0_48[367]},
      {stage0_49[380]},
      {stage0_50[162], stage0_50[163], stage0_50[164], stage0_50[165], stage0_50[166], stage0_50[167]},
      {stage1_52[27],stage1_51[88],stage1_50[112],stage1_49[136],stage1_48[167]}
   );
   gpc615_5 gpc1871 (
      {stage0_48[368], stage0_48[369], stage0_48[370], stage0_48[371], stage0_48[372]},
      {stage0_49[381]},
      {stage0_50[168], stage0_50[169], stage0_50[170], stage0_50[171], stage0_50[172], stage0_50[173]},
      {stage1_52[28],stage1_51[89],stage1_50[113],stage1_49[137],stage1_48[168]}
   );
   gpc615_5 gpc1872 (
      {stage0_48[373], stage0_48[374], stage0_48[375], stage0_48[376], stage0_48[377]},
      {stage0_49[382]},
      {stage0_50[174], stage0_50[175], stage0_50[176], stage0_50[177], stage0_50[178], stage0_50[179]},
      {stage1_52[29],stage1_51[90],stage1_50[114],stage1_49[138],stage1_48[169]}
   );
   gpc615_5 gpc1873 (
      {stage0_48[378], stage0_48[379], stage0_48[380], stage0_48[381], stage0_48[382]},
      {stage0_49[383]},
      {stage0_50[180], stage0_50[181], stage0_50[182], stage0_50[183], stage0_50[184], stage0_50[185]},
      {stage1_52[30],stage1_51[91],stage1_50[115],stage1_49[139],stage1_48[170]}
   );
   gpc615_5 gpc1874 (
      {stage0_48[383], stage0_48[384], stage0_48[385], stage0_48[386], stage0_48[387]},
      {stage0_49[384]},
      {stage0_50[186], stage0_50[187], stage0_50[188], stage0_50[189], stage0_50[190], stage0_50[191]},
      {stage1_52[31],stage1_51[92],stage1_50[116],stage1_49[140],stage1_48[171]}
   );
   gpc615_5 gpc1875 (
      {stage0_48[388], stage0_48[389], stage0_48[390], stage0_48[391], stage0_48[392]},
      {stage0_49[385]},
      {stage0_50[192], stage0_50[193], stage0_50[194], stage0_50[195], stage0_50[196], stage0_50[197]},
      {stage1_52[32],stage1_51[93],stage1_50[117],stage1_49[141],stage1_48[172]}
   );
   gpc615_5 gpc1876 (
      {stage0_48[393], stage0_48[394], stage0_48[395], stage0_48[396], stage0_48[397]},
      {stage0_49[386]},
      {stage0_50[198], stage0_50[199], stage0_50[200], stage0_50[201], stage0_50[202], stage0_50[203]},
      {stage1_52[33],stage1_51[94],stage1_50[118],stage1_49[142],stage1_48[173]}
   );
   gpc615_5 gpc1877 (
      {stage0_48[398], stage0_48[399], stage0_48[400], stage0_48[401], stage0_48[402]},
      {stage0_49[387]},
      {stage0_50[204], stage0_50[205], stage0_50[206], stage0_50[207], stage0_50[208], stage0_50[209]},
      {stage1_52[34],stage1_51[95],stage1_50[119],stage1_49[143],stage1_48[174]}
   );
   gpc615_5 gpc1878 (
      {stage0_48[403], stage0_48[404], stage0_48[405], stage0_48[406], stage0_48[407]},
      {stage0_49[388]},
      {stage0_50[210], stage0_50[211], stage0_50[212], stage0_50[213], stage0_50[214], stage0_50[215]},
      {stage1_52[35],stage1_51[96],stage1_50[120],stage1_49[144],stage1_48[175]}
   );
   gpc615_5 gpc1879 (
      {stage0_48[408], stage0_48[409], stage0_48[410], stage0_48[411], stage0_48[412]},
      {stage0_49[389]},
      {stage0_50[216], stage0_50[217], stage0_50[218], stage0_50[219], stage0_50[220], stage0_50[221]},
      {stage1_52[36],stage1_51[97],stage1_50[121],stage1_49[145],stage1_48[176]}
   );
   gpc615_5 gpc1880 (
      {stage0_48[413], stage0_48[414], stage0_48[415], stage0_48[416], stage0_48[417]},
      {stage0_49[390]},
      {stage0_50[222], stage0_50[223], stage0_50[224], stage0_50[225], stage0_50[226], stage0_50[227]},
      {stage1_52[37],stage1_51[98],stage1_50[122],stage1_49[146],stage1_48[177]}
   );
   gpc615_5 gpc1881 (
      {stage0_48[418], stage0_48[419], stage0_48[420], stage0_48[421], stage0_48[422]},
      {stage0_49[391]},
      {stage0_50[228], stage0_50[229], stage0_50[230], stage0_50[231], stage0_50[232], stage0_50[233]},
      {stage1_52[38],stage1_51[99],stage1_50[123],stage1_49[147],stage1_48[178]}
   );
   gpc615_5 gpc1882 (
      {stage0_48[423], stage0_48[424], stage0_48[425], stage0_48[426], stage0_48[427]},
      {stage0_49[392]},
      {stage0_50[234], stage0_50[235], stage0_50[236], stage0_50[237], stage0_50[238], stage0_50[239]},
      {stage1_52[39],stage1_51[100],stage1_50[124],stage1_49[148],stage1_48[179]}
   );
   gpc615_5 gpc1883 (
      {stage0_48[428], stage0_48[429], stage0_48[430], stage0_48[431], stage0_48[432]},
      {stage0_49[393]},
      {stage0_50[240], stage0_50[241], stage0_50[242], stage0_50[243], stage0_50[244], stage0_50[245]},
      {stage1_52[40],stage1_51[101],stage1_50[125],stage1_49[149],stage1_48[180]}
   );
   gpc615_5 gpc1884 (
      {stage0_48[433], stage0_48[434], stage0_48[435], stage0_48[436], stage0_48[437]},
      {stage0_49[394]},
      {stage0_50[246], stage0_50[247], stage0_50[248], stage0_50[249], stage0_50[250], stage0_50[251]},
      {stage1_52[41],stage1_51[102],stage1_50[126],stage1_49[150],stage1_48[181]}
   );
   gpc615_5 gpc1885 (
      {stage0_48[438], stage0_48[439], stage0_48[440], stage0_48[441], stage0_48[442]},
      {stage0_49[395]},
      {stage0_50[252], stage0_50[253], stage0_50[254], stage0_50[255], stage0_50[256], stage0_50[257]},
      {stage1_52[42],stage1_51[103],stage1_50[127],stage1_49[151],stage1_48[182]}
   );
   gpc615_5 gpc1886 (
      {stage0_48[443], stage0_48[444], stage0_48[445], stage0_48[446], stage0_48[447]},
      {stage0_49[396]},
      {stage0_50[258], stage0_50[259], stage0_50[260], stage0_50[261], stage0_50[262], stage0_50[263]},
      {stage1_52[43],stage1_51[104],stage1_50[128],stage1_49[152],stage1_48[183]}
   );
   gpc615_5 gpc1887 (
      {stage0_48[448], stage0_48[449], stage0_48[450], stage0_48[451], stage0_48[452]},
      {stage0_49[397]},
      {stage0_50[264], stage0_50[265], stage0_50[266], stage0_50[267], stage0_50[268], stage0_50[269]},
      {stage1_52[44],stage1_51[105],stage1_50[129],stage1_49[153],stage1_48[184]}
   );
   gpc615_5 gpc1888 (
      {stage0_48[453], stage0_48[454], stage0_48[455], stage0_48[456], stage0_48[457]},
      {stage0_49[398]},
      {stage0_50[270], stage0_50[271], stage0_50[272], stage0_50[273], stage0_50[274], stage0_50[275]},
      {stage1_52[45],stage1_51[106],stage1_50[130],stage1_49[154],stage1_48[185]}
   );
   gpc615_5 gpc1889 (
      {stage0_48[458], stage0_48[459], stage0_48[460], stage0_48[461], stage0_48[462]},
      {stage0_49[399]},
      {stage0_50[276], stage0_50[277], stage0_50[278], stage0_50[279], stage0_50[280], stage0_50[281]},
      {stage1_52[46],stage1_51[107],stage1_50[131],stage1_49[155],stage1_48[186]}
   );
   gpc615_5 gpc1890 (
      {stage0_48[463], stage0_48[464], stage0_48[465], stage0_48[466], stage0_48[467]},
      {stage0_49[400]},
      {stage0_50[282], stage0_50[283], stage0_50[284], stage0_50[285], stage0_50[286], stage0_50[287]},
      {stage1_52[47],stage1_51[108],stage1_50[132],stage1_49[156],stage1_48[187]}
   );
   gpc615_5 gpc1891 (
      {stage0_48[468], stage0_48[469], stage0_48[470], stage0_48[471], stage0_48[472]},
      {stage0_49[401]},
      {stage0_50[288], stage0_50[289], stage0_50[290], stage0_50[291], stage0_50[292], stage0_50[293]},
      {stage1_52[48],stage1_51[109],stage1_50[133],stage1_49[157],stage1_48[188]}
   );
   gpc615_5 gpc1892 (
      {stage0_48[473], stage0_48[474], stage0_48[475], stage0_48[476], stage0_48[477]},
      {stage0_49[402]},
      {stage0_50[294], stage0_50[295], stage0_50[296], stage0_50[297], stage0_50[298], stage0_50[299]},
      {stage1_52[49],stage1_51[110],stage1_50[134],stage1_49[158],stage1_48[189]}
   );
   gpc606_5 gpc1893 (
      {stage0_49[403], stage0_49[404], stage0_49[405], stage0_49[406], stage0_49[407], stage0_49[408]},
      {stage0_51[0], stage0_51[1], stage0_51[2], stage0_51[3], stage0_51[4], stage0_51[5]},
      {stage1_53[0],stage1_52[50],stage1_51[111],stage1_50[135],stage1_49[159]}
   );
   gpc606_5 gpc1894 (
      {stage0_49[409], stage0_49[410], stage0_49[411], stage0_49[412], stage0_49[413], stage0_49[414]},
      {stage0_51[6], stage0_51[7], stage0_51[8], stage0_51[9], stage0_51[10], stage0_51[11]},
      {stage1_53[1],stage1_52[51],stage1_51[112],stage1_50[136],stage1_49[160]}
   );
   gpc606_5 gpc1895 (
      {stage0_49[415], stage0_49[416], stage0_49[417], stage0_49[418], stage0_49[419], stage0_49[420]},
      {stage0_51[12], stage0_51[13], stage0_51[14], stage0_51[15], stage0_51[16], stage0_51[17]},
      {stage1_53[2],stage1_52[52],stage1_51[113],stage1_50[137],stage1_49[161]}
   );
   gpc606_5 gpc1896 (
      {stage0_49[421], stage0_49[422], stage0_49[423], stage0_49[424], stage0_49[425], stage0_49[426]},
      {stage0_51[18], stage0_51[19], stage0_51[20], stage0_51[21], stage0_51[22], stage0_51[23]},
      {stage1_53[3],stage1_52[53],stage1_51[114],stage1_50[138],stage1_49[162]}
   );
   gpc606_5 gpc1897 (
      {stage0_49[427], stage0_49[428], stage0_49[429], stage0_49[430], stage0_49[431], stage0_49[432]},
      {stage0_51[24], stage0_51[25], stage0_51[26], stage0_51[27], stage0_51[28], stage0_51[29]},
      {stage1_53[4],stage1_52[54],stage1_51[115],stage1_50[139],stage1_49[163]}
   );
   gpc606_5 gpc1898 (
      {stage0_49[433], stage0_49[434], stage0_49[435], stage0_49[436], stage0_49[437], stage0_49[438]},
      {stage0_51[30], stage0_51[31], stage0_51[32], stage0_51[33], stage0_51[34], stage0_51[35]},
      {stage1_53[5],stage1_52[55],stage1_51[116],stage1_50[140],stage1_49[164]}
   );
   gpc606_5 gpc1899 (
      {stage0_49[439], stage0_49[440], stage0_49[441], stage0_49[442], stage0_49[443], stage0_49[444]},
      {stage0_51[36], stage0_51[37], stage0_51[38], stage0_51[39], stage0_51[40], stage0_51[41]},
      {stage1_53[6],stage1_52[56],stage1_51[117],stage1_50[141],stage1_49[165]}
   );
   gpc606_5 gpc1900 (
      {stage0_49[445], stage0_49[446], stage0_49[447], stage0_49[448], stage0_49[449], stage0_49[450]},
      {stage0_51[42], stage0_51[43], stage0_51[44], stage0_51[45], stage0_51[46], stage0_51[47]},
      {stage1_53[7],stage1_52[57],stage1_51[118],stage1_50[142],stage1_49[166]}
   );
   gpc606_5 gpc1901 (
      {stage0_49[451], stage0_49[452], stage0_49[453], stage0_49[454], stage0_49[455], stage0_49[456]},
      {stage0_51[48], stage0_51[49], stage0_51[50], stage0_51[51], stage0_51[52], stage0_51[53]},
      {stage1_53[8],stage1_52[58],stage1_51[119],stage1_50[143],stage1_49[167]}
   );
   gpc606_5 gpc1902 (
      {stage0_49[457], stage0_49[458], stage0_49[459], stage0_49[460], stage0_49[461], stage0_49[462]},
      {stage0_51[54], stage0_51[55], stage0_51[56], stage0_51[57], stage0_51[58], stage0_51[59]},
      {stage1_53[9],stage1_52[59],stage1_51[120],stage1_50[144],stage1_49[168]}
   );
   gpc606_5 gpc1903 (
      {stage0_49[463], stage0_49[464], stage0_49[465], stage0_49[466], stage0_49[467], stage0_49[468]},
      {stage0_51[60], stage0_51[61], stage0_51[62], stage0_51[63], stage0_51[64], stage0_51[65]},
      {stage1_53[10],stage1_52[60],stage1_51[121],stage1_50[145],stage1_49[169]}
   );
   gpc606_5 gpc1904 (
      {stage0_49[469], stage0_49[470], stage0_49[471], stage0_49[472], stage0_49[473], stage0_49[474]},
      {stage0_51[66], stage0_51[67], stage0_51[68], stage0_51[69], stage0_51[70], stage0_51[71]},
      {stage1_53[11],stage1_52[61],stage1_51[122],stage1_50[146],stage1_49[170]}
   );
   gpc606_5 gpc1905 (
      {stage0_49[475], stage0_49[476], stage0_49[477], stage0_49[478], stage0_49[479], stage0_49[480]},
      {stage0_51[72], stage0_51[73], stage0_51[74], stage0_51[75], stage0_51[76], stage0_51[77]},
      {stage1_53[12],stage1_52[62],stage1_51[123],stage1_50[147],stage1_49[171]}
   );
   gpc615_5 gpc1906 (
      {stage0_49[481], stage0_49[482], stage0_49[483], stage0_49[484], stage0_49[485]},
      {stage0_50[300]},
      {stage0_51[78], stage0_51[79], stage0_51[80], stage0_51[81], stage0_51[82], stage0_51[83]},
      {stage1_53[13],stage1_52[63],stage1_51[124],stage1_50[148],stage1_49[172]}
   );
   gpc615_5 gpc1907 (
      {stage0_50[301], stage0_50[302], stage0_50[303], stage0_50[304], stage0_50[305]},
      {stage0_51[84]},
      {stage0_52[0], stage0_52[1], stage0_52[2], stage0_52[3], stage0_52[4], stage0_52[5]},
      {stage1_54[0],stage1_53[14],stage1_52[64],stage1_51[125],stage1_50[149]}
   );
   gpc615_5 gpc1908 (
      {stage0_50[306], stage0_50[307], stage0_50[308], stage0_50[309], stage0_50[310]},
      {stage0_51[85]},
      {stage0_52[6], stage0_52[7], stage0_52[8], stage0_52[9], stage0_52[10], stage0_52[11]},
      {stage1_54[1],stage1_53[15],stage1_52[65],stage1_51[126],stage1_50[150]}
   );
   gpc615_5 gpc1909 (
      {stage0_50[311], stage0_50[312], stage0_50[313], stage0_50[314], stage0_50[315]},
      {stage0_51[86]},
      {stage0_52[12], stage0_52[13], stage0_52[14], stage0_52[15], stage0_52[16], stage0_52[17]},
      {stage1_54[2],stage1_53[16],stage1_52[66],stage1_51[127],stage1_50[151]}
   );
   gpc615_5 gpc1910 (
      {stage0_50[316], stage0_50[317], stage0_50[318], stage0_50[319], stage0_50[320]},
      {stage0_51[87]},
      {stage0_52[18], stage0_52[19], stage0_52[20], stage0_52[21], stage0_52[22], stage0_52[23]},
      {stage1_54[3],stage1_53[17],stage1_52[67],stage1_51[128],stage1_50[152]}
   );
   gpc615_5 gpc1911 (
      {stage0_50[321], stage0_50[322], stage0_50[323], stage0_50[324], stage0_50[325]},
      {stage0_51[88]},
      {stage0_52[24], stage0_52[25], stage0_52[26], stage0_52[27], stage0_52[28], stage0_52[29]},
      {stage1_54[4],stage1_53[18],stage1_52[68],stage1_51[129],stage1_50[153]}
   );
   gpc615_5 gpc1912 (
      {stage0_50[326], stage0_50[327], stage0_50[328], stage0_50[329], stage0_50[330]},
      {stage0_51[89]},
      {stage0_52[30], stage0_52[31], stage0_52[32], stage0_52[33], stage0_52[34], stage0_52[35]},
      {stage1_54[5],stage1_53[19],stage1_52[69],stage1_51[130],stage1_50[154]}
   );
   gpc615_5 gpc1913 (
      {stage0_50[331], stage0_50[332], stage0_50[333], stage0_50[334], stage0_50[335]},
      {stage0_51[90]},
      {stage0_52[36], stage0_52[37], stage0_52[38], stage0_52[39], stage0_52[40], stage0_52[41]},
      {stage1_54[6],stage1_53[20],stage1_52[70],stage1_51[131],stage1_50[155]}
   );
   gpc615_5 gpc1914 (
      {stage0_50[336], stage0_50[337], stage0_50[338], stage0_50[339], stage0_50[340]},
      {stage0_51[91]},
      {stage0_52[42], stage0_52[43], stage0_52[44], stage0_52[45], stage0_52[46], stage0_52[47]},
      {stage1_54[7],stage1_53[21],stage1_52[71],stage1_51[132],stage1_50[156]}
   );
   gpc615_5 gpc1915 (
      {stage0_50[341], stage0_50[342], stage0_50[343], stage0_50[344], stage0_50[345]},
      {stage0_51[92]},
      {stage0_52[48], stage0_52[49], stage0_52[50], stage0_52[51], stage0_52[52], stage0_52[53]},
      {stage1_54[8],stage1_53[22],stage1_52[72],stage1_51[133],stage1_50[157]}
   );
   gpc615_5 gpc1916 (
      {stage0_50[346], stage0_50[347], stage0_50[348], stage0_50[349], stage0_50[350]},
      {stage0_51[93]},
      {stage0_52[54], stage0_52[55], stage0_52[56], stage0_52[57], stage0_52[58], stage0_52[59]},
      {stage1_54[9],stage1_53[23],stage1_52[73],stage1_51[134],stage1_50[158]}
   );
   gpc615_5 gpc1917 (
      {stage0_50[351], stage0_50[352], stage0_50[353], stage0_50[354], stage0_50[355]},
      {stage0_51[94]},
      {stage0_52[60], stage0_52[61], stage0_52[62], stage0_52[63], stage0_52[64], stage0_52[65]},
      {stage1_54[10],stage1_53[24],stage1_52[74],stage1_51[135],stage1_50[159]}
   );
   gpc615_5 gpc1918 (
      {stage0_50[356], stage0_50[357], stage0_50[358], stage0_50[359], stage0_50[360]},
      {stage0_51[95]},
      {stage0_52[66], stage0_52[67], stage0_52[68], stage0_52[69], stage0_52[70], stage0_52[71]},
      {stage1_54[11],stage1_53[25],stage1_52[75],stage1_51[136],stage1_50[160]}
   );
   gpc615_5 gpc1919 (
      {stage0_50[361], stage0_50[362], stage0_50[363], stage0_50[364], stage0_50[365]},
      {stage0_51[96]},
      {stage0_52[72], stage0_52[73], stage0_52[74], stage0_52[75], stage0_52[76], stage0_52[77]},
      {stage1_54[12],stage1_53[26],stage1_52[76],stage1_51[137],stage1_50[161]}
   );
   gpc615_5 gpc1920 (
      {stage0_50[366], stage0_50[367], stage0_50[368], stage0_50[369], stage0_50[370]},
      {stage0_51[97]},
      {stage0_52[78], stage0_52[79], stage0_52[80], stage0_52[81], stage0_52[82], stage0_52[83]},
      {stage1_54[13],stage1_53[27],stage1_52[77],stage1_51[138],stage1_50[162]}
   );
   gpc615_5 gpc1921 (
      {stage0_50[371], stage0_50[372], stage0_50[373], stage0_50[374], stage0_50[375]},
      {stage0_51[98]},
      {stage0_52[84], stage0_52[85], stage0_52[86], stage0_52[87], stage0_52[88], stage0_52[89]},
      {stage1_54[14],stage1_53[28],stage1_52[78],stage1_51[139],stage1_50[163]}
   );
   gpc615_5 gpc1922 (
      {stage0_50[376], stage0_50[377], stage0_50[378], stage0_50[379], stage0_50[380]},
      {stage0_51[99]},
      {stage0_52[90], stage0_52[91], stage0_52[92], stage0_52[93], stage0_52[94], stage0_52[95]},
      {stage1_54[15],stage1_53[29],stage1_52[79],stage1_51[140],stage1_50[164]}
   );
   gpc615_5 gpc1923 (
      {stage0_50[381], stage0_50[382], stage0_50[383], stage0_50[384], stage0_50[385]},
      {stage0_51[100]},
      {stage0_52[96], stage0_52[97], stage0_52[98], stage0_52[99], stage0_52[100], stage0_52[101]},
      {stage1_54[16],stage1_53[30],stage1_52[80],stage1_51[141],stage1_50[165]}
   );
   gpc615_5 gpc1924 (
      {stage0_50[386], stage0_50[387], stage0_50[388], stage0_50[389], stage0_50[390]},
      {stage0_51[101]},
      {stage0_52[102], stage0_52[103], stage0_52[104], stage0_52[105], stage0_52[106], stage0_52[107]},
      {stage1_54[17],stage1_53[31],stage1_52[81],stage1_51[142],stage1_50[166]}
   );
   gpc615_5 gpc1925 (
      {stage0_50[391], stage0_50[392], stage0_50[393], stage0_50[394], stage0_50[395]},
      {stage0_51[102]},
      {stage0_52[108], stage0_52[109], stage0_52[110], stage0_52[111], stage0_52[112], stage0_52[113]},
      {stage1_54[18],stage1_53[32],stage1_52[82],stage1_51[143],stage1_50[167]}
   );
   gpc615_5 gpc1926 (
      {stage0_50[396], stage0_50[397], stage0_50[398], stage0_50[399], stage0_50[400]},
      {stage0_51[103]},
      {stage0_52[114], stage0_52[115], stage0_52[116], stage0_52[117], stage0_52[118], stage0_52[119]},
      {stage1_54[19],stage1_53[33],stage1_52[83],stage1_51[144],stage1_50[168]}
   );
   gpc615_5 gpc1927 (
      {stage0_50[401], stage0_50[402], stage0_50[403], stage0_50[404], stage0_50[405]},
      {stage0_51[104]},
      {stage0_52[120], stage0_52[121], stage0_52[122], stage0_52[123], stage0_52[124], stage0_52[125]},
      {stage1_54[20],stage1_53[34],stage1_52[84],stage1_51[145],stage1_50[169]}
   );
   gpc615_5 gpc1928 (
      {stage0_50[406], stage0_50[407], stage0_50[408], stage0_50[409], stage0_50[410]},
      {stage0_51[105]},
      {stage0_52[126], stage0_52[127], stage0_52[128], stage0_52[129], stage0_52[130], stage0_52[131]},
      {stage1_54[21],stage1_53[35],stage1_52[85],stage1_51[146],stage1_50[170]}
   );
   gpc615_5 gpc1929 (
      {stage0_50[411], stage0_50[412], stage0_50[413], stage0_50[414], stage0_50[415]},
      {stage0_51[106]},
      {stage0_52[132], stage0_52[133], stage0_52[134], stage0_52[135], stage0_52[136], stage0_52[137]},
      {stage1_54[22],stage1_53[36],stage1_52[86],stage1_51[147],stage1_50[171]}
   );
   gpc615_5 gpc1930 (
      {stage0_50[416], stage0_50[417], stage0_50[418], stage0_50[419], stage0_50[420]},
      {stage0_51[107]},
      {stage0_52[138], stage0_52[139], stage0_52[140], stage0_52[141], stage0_52[142], stage0_52[143]},
      {stage1_54[23],stage1_53[37],stage1_52[87],stage1_51[148],stage1_50[172]}
   );
   gpc615_5 gpc1931 (
      {stage0_50[421], stage0_50[422], stage0_50[423], stage0_50[424], stage0_50[425]},
      {stage0_51[108]},
      {stage0_52[144], stage0_52[145], stage0_52[146], stage0_52[147], stage0_52[148], stage0_52[149]},
      {stage1_54[24],stage1_53[38],stage1_52[88],stage1_51[149],stage1_50[173]}
   );
   gpc615_5 gpc1932 (
      {stage0_50[426], stage0_50[427], stage0_50[428], stage0_50[429], stage0_50[430]},
      {stage0_51[109]},
      {stage0_52[150], stage0_52[151], stage0_52[152], stage0_52[153], stage0_52[154], stage0_52[155]},
      {stage1_54[25],stage1_53[39],stage1_52[89],stage1_51[150],stage1_50[174]}
   );
   gpc615_5 gpc1933 (
      {stage0_50[431], stage0_50[432], stage0_50[433], stage0_50[434], stage0_50[435]},
      {stage0_51[110]},
      {stage0_52[156], stage0_52[157], stage0_52[158], stage0_52[159], stage0_52[160], stage0_52[161]},
      {stage1_54[26],stage1_53[40],stage1_52[90],stage1_51[151],stage1_50[175]}
   );
   gpc615_5 gpc1934 (
      {stage0_50[436], stage0_50[437], stage0_50[438], stage0_50[439], stage0_50[440]},
      {stage0_51[111]},
      {stage0_52[162], stage0_52[163], stage0_52[164], stage0_52[165], stage0_52[166], stage0_52[167]},
      {stage1_54[27],stage1_53[41],stage1_52[91],stage1_51[152],stage1_50[176]}
   );
   gpc615_5 gpc1935 (
      {stage0_50[441], stage0_50[442], stage0_50[443], stage0_50[444], stage0_50[445]},
      {stage0_51[112]},
      {stage0_52[168], stage0_52[169], stage0_52[170], stage0_52[171], stage0_52[172], stage0_52[173]},
      {stage1_54[28],stage1_53[42],stage1_52[92],stage1_51[153],stage1_50[177]}
   );
   gpc615_5 gpc1936 (
      {stage0_50[446], stage0_50[447], stage0_50[448], stage0_50[449], stage0_50[450]},
      {stage0_51[113]},
      {stage0_52[174], stage0_52[175], stage0_52[176], stage0_52[177], stage0_52[178], stage0_52[179]},
      {stage1_54[29],stage1_53[43],stage1_52[93],stage1_51[154],stage1_50[178]}
   );
   gpc615_5 gpc1937 (
      {stage0_50[451], stage0_50[452], stage0_50[453], stage0_50[454], stage0_50[455]},
      {stage0_51[114]},
      {stage0_52[180], stage0_52[181], stage0_52[182], stage0_52[183], stage0_52[184], stage0_52[185]},
      {stage1_54[30],stage1_53[44],stage1_52[94],stage1_51[155],stage1_50[179]}
   );
   gpc615_5 gpc1938 (
      {stage0_50[456], stage0_50[457], stage0_50[458], stage0_50[459], stage0_50[460]},
      {stage0_51[115]},
      {stage0_52[186], stage0_52[187], stage0_52[188], stage0_52[189], stage0_52[190], stage0_52[191]},
      {stage1_54[31],stage1_53[45],stage1_52[95],stage1_51[156],stage1_50[180]}
   );
   gpc615_5 gpc1939 (
      {stage0_50[461], stage0_50[462], stage0_50[463], stage0_50[464], stage0_50[465]},
      {stage0_51[116]},
      {stage0_52[192], stage0_52[193], stage0_52[194], stage0_52[195], stage0_52[196], stage0_52[197]},
      {stage1_54[32],stage1_53[46],stage1_52[96],stage1_51[157],stage1_50[181]}
   );
   gpc615_5 gpc1940 (
      {stage0_50[466], stage0_50[467], stage0_50[468], stage0_50[469], stage0_50[470]},
      {stage0_51[117]},
      {stage0_52[198], stage0_52[199], stage0_52[200], stage0_52[201], stage0_52[202], stage0_52[203]},
      {stage1_54[33],stage1_53[47],stage1_52[97],stage1_51[158],stage1_50[182]}
   );
   gpc615_5 gpc1941 (
      {stage0_50[471], stage0_50[472], stage0_50[473], stage0_50[474], stage0_50[475]},
      {stage0_51[118]},
      {stage0_52[204], stage0_52[205], stage0_52[206], stage0_52[207], stage0_52[208], stage0_52[209]},
      {stage1_54[34],stage1_53[48],stage1_52[98],stage1_51[159],stage1_50[183]}
   );
   gpc615_5 gpc1942 (
      {stage0_50[476], stage0_50[477], stage0_50[478], stage0_50[479], stage0_50[480]},
      {stage0_51[119]},
      {stage0_52[210], stage0_52[211], stage0_52[212], stage0_52[213], stage0_52[214], stage0_52[215]},
      {stage1_54[35],stage1_53[49],stage1_52[99],stage1_51[160],stage1_50[184]}
   );
   gpc615_5 gpc1943 (
      {stage0_51[120], stage0_51[121], stage0_51[122], stage0_51[123], stage0_51[124]},
      {stage0_52[216]},
      {stage0_53[0], stage0_53[1], stage0_53[2], stage0_53[3], stage0_53[4], stage0_53[5]},
      {stage1_55[0],stage1_54[36],stage1_53[50],stage1_52[100],stage1_51[161]}
   );
   gpc615_5 gpc1944 (
      {stage0_51[125], stage0_51[126], stage0_51[127], stage0_51[128], stage0_51[129]},
      {stage0_52[217]},
      {stage0_53[6], stage0_53[7], stage0_53[8], stage0_53[9], stage0_53[10], stage0_53[11]},
      {stage1_55[1],stage1_54[37],stage1_53[51],stage1_52[101],stage1_51[162]}
   );
   gpc615_5 gpc1945 (
      {stage0_51[130], stage0_51[131], stage0_51[132], stage0_51[133], stage0_51[134]},
      {stage0_52[218]},
      {stage0_53[12], stage0_53[13], stage0_53[14], stage0_53[15], stage0_53[16], stage0_53[17]},
      {stage1_55[2],stage1_54[38],stage1_53[52],stage1_52[102],stage1_51[163]}
   );
   gpc615_5 gpc1946 (
      {stage0_51[135], stage0_51[136], stage0_51[137], stage0_51[138], stage0_51[139]},
      {stage0_52[219]},
      {stage0_53[18], stage0_53[19], stage0_53[20], stage0_53[21], stage0_53[22], stage0_53[23]},
      {stage1_55[3],stage1_54[39],stage1_53[53],stage1_52[103],stage1_51[164]}
   );
   gpc615_5 gpc1947 (
      {stage0_51[140], stage0_51[141], stage0_51[142], stage0_51[143], stage0_51[144]},
      {stage0_52[220]},
      {stage0_53[24], stage0_53[25], stage0_53[26], stage0_53[27], stage0_53[28], stage0_53[29]},
      {stage1_55[4],stage1_54[40],stage1_53[54],stage1_52[104],stage1_51[165]}
   );
   gpc615_5 gpc1948 (
      {stage0_51[145], stage0_51[146], stage0_51[147], stage0_51[148], stage0_51[149]},
      {stage0_52[221]},
      {stage0_53[30], stage0_53[31], stage0_53[32], stage0_53[33], stage0_53[34], stage0_53[35]},
      {stage1_55[5],stage1_54[41],stage1_53[55],stage1_52[105],stage1_51[166]}
   );
   gpc615_5 gpc1949 (
      {stage0_51[150], stage0_51[151], stage0_51[152], stage0_51[153], stage0_51[154]},
      {stage0_52[222]},
      {stage0_53[36], stage0_53[37], stage0_53[38], stage0_53[39], stage0_53[40], stage0_53[41]},
      {stage1_55[6],stage1_54[42],stage1_53[56],stage1_52[106],stage1_51[167]}
   );
   gpc615_5 gpc1950 (
      {stage0_51[155], stage0_51[156], stage0_51[157], stage0_51[158], stage0_51[159]},
      {stage0_52[223]},
      {stage0_53[42], stage0_53[43], stage0_53[44], stage0_53[45], stage0_53[46], stage0_53[47]},
      {stage1_55[7],stage1_54[43],stage1_53[57],stage1_52[107],stage1_51[168]}
   );
   gpc615_5 gpc1951 (
      {stage0_51[160], stage0_51[161], stage0_51[162], stage0_51[163], stage0_51[164]},
      {stage0_52[224]},
      {stage0_53[48], stage0_53[49], stage0_53[50], stage0_53[51], stage0_53[52], stage0_53[53]},
      {stage1_55[8],stage1_54[44],stage1_53[58],stage1_52[108],stage1_51[169]}
   );
   gpc615_5 gpc1952 (
      {stage0_51[165], stage0_51[166], stage0_51[167], stage0_51[168], stage0_51[169]},
      {stage0_52[225]},
      {stage0_53[54], stage0_53[55], stage0_53[56], stage0_53[57], stage0_53[58], stage0_53[59]},
      {stage1_55[9],stage1_54[45],stage1_53[59],stage1_52[109],stage1_51[170]}
   );
   gpc615_5 gpc1953 (
      {stage0_51[170], stage0_51[171], stage0_51[172], stage0_51[173], stage0_51[174]},
      {stage0_52[226]},
      {stage0_53[60], stage0_53[61], stage0_53[62], stage0_53[63], stage0_53[64], stage0_53[65]},
      {stage1_55[10],stage1_54[46],stage1_53[60],stage1_52[110],stage1_51[171]}
   );
   gpc615_5 gpc1954 (
      {stage0_51[175], stage0_51[176], stage0_51[177], stage0_51[178], stage0_51[179]},
      {stage0_52[227]},
      {stage0_53[66], stage0_53[67], stage0_53[68], stage0_53[69], stage0_53[70], stage0_53[71]},
      {stage1_55[11],stage1_54[47],stage1_53[61],stage1_52[111],stage1_51[172]}
   );
   gpc615_5 gpc1955 (
      {stage0_51[180], stage0_51[181], stage0_51[182], stage0_51[183], stage0_51[184]},
      {stage0_52[228]},
      {stage0_53[72], stage0_53[73], stage0_53[74], stage0_53[75], stage0_53[76], stage0_53[77]},
      {stage1_55[12],stage1_54[48],stage1_53[62],stage1_52[112],stage1_51[173]}
   );
   gpc615_5 gpc1956 (
      {stage0_51[185], stage0_51[186], stage0_51[187], stage0_51[188], stage0_51[189]},
      {stage0_52[229]},
      {stage0_53[78], stage0_53[79], stage0_53[80], stage0_53[81], stage0_53[82], stage0_53[83]},
      {stage1_55[13],stage1_54[49],stage1_53[63],stage1_52[113],stage1_51[174]}
   );
   gpc615_5 gpc1957 (
      {stage0_51[190], stage0_51[191], stage0_51[192], stage0_51[193], stage0_51[194]},
      {stage0_52[230]},
      {stage0_53[84], stage0_53[85], stage0_53[86], stage0_53[87], stage0_53[88], stage0_53[89]},
      {stage1_55[14],stage1_54[50],stage1_53[64],stage1_52[114],stage1_51[175]}
   );
   gpc615_5 gpc1958 (
      {stage0_51[195], stage0_51[196], stage0_51[197], stage0_51[198], stage0_51[199]},
      {stage0_52[231]},
      {stage0_53[90], stage0_53[91], stage0_53[92], stage0_53[93], stage0_53[94], stage0_53[95]},
      {stage1_55[15],stage1_54[51],stage1_53[65],stage1_52[115],stage1_51[176]}
   );
   gpc615_5 gpc1959 (
      {stage0_51[200], stage0_51[201], stage0_51[202], stage0_51[203], stage0_51[204]},
      {stage0_52[232]},
      {stage0_53[96], stage0_53[97], stage0_53[98], stage0_53[99], stage0_53[100], stage0_53[101]},
      {stage1_55[16],stage1_54[52],stage1_53[66],stage1_52[116],stage1_51[177]}
   );
   gpc615_5 gpc1960 (
      {stage0_51[205], stage0_51[206], stage0_51[207], stage0_51[208], stage0_51[209]},
      {stage0_52[233]},
      {stage0_53[102], stage0_53[103], stage0_53[104], stage0_53[105], stage0_53[106], stage0_53[107]},
      {stage1_55[17],stage1_54[53],stage1_53[67],stage1_52[117],stage1_51[178]}
   );
   gpc615_5 gpc1961 (
      {stage0_51[210], stage0_51[211], stage0_51[212], stage0_51[213], stage0_51[214]},
      {stage0_52[234]},
      {stage0_53[108], stage0_53[109], stage0_53[110], stage0_53[111], stage0_53[112], stage0_53[113]},
      {stage1_55[18],stage1_54[54],stage1_53[68],stage1_52[118],stage1_51[179]}
   );
   gpc615_5 gpc1962 (
      {stage0_51[215], stage0_51[216], stage0_51[217], stage0_51[218], stage0_51[219]},
      {stage0_52[235]},
      {stage0_53[114], stage0_53[115], stage0_53[116], stage0_53[117], stage0_53[118], stage0_53[119]},
      {stage1_55[19],stage1_54[55],stage1_53[69],stage1_52[119],stage1_51[180]}
   );
   gpc615_5 gpc1963 (
      {stage0_51[220], stage0_51[221], stage0_51[222], stage0_51[223], stage0_51[224]},
      {stage0_52[236]},
      {stage0_53[120], stage0_53[121], stage0_53[122], stage0_53[123], stage0_53[124], stage0_53[125]},
      {stage1_55[20],stage1_54[56],stage1_53[70],stage1_52[120],stage1_51[181]}
   );
   gpc615_5 gpc1964 (
      {stage0_51[225], stage0_51[226], stage0_51[227], stage0_51[228], stage0_51[229]},
      {stage0_52[237]},
      {stage0_53[126], stage0_53[127], stage0_53[128], stage0_53[129], stage0_53[130], stage0_53[131]},
      {stage1_55[21],stage1_54[57],stage1_53[71],stage1_52[121],stage1_51[182]}
   );
   gpc615_5 gpc1965 (
      {stage0_51[230], stage0_51[231], stage0_51[232], stage0_51[233], stage0_51[234]},
      {stage0_52[238]},
      {stage0_53[132], stage0_53[133], stage0_53[134], stage0_53[135], stage0_53[136], stage0_53[137]},
      {stage1_55[22],stage1_54[58],stage1_53[72],stage1_52[122],stage1_51[183]}
   );
   gpc615_5 gpc1966 (
      {stage0_51[235], stage0_51[236], stage0_51[237], stage0_51[238], stage0_51[239]},
      {stage0_52[239]},
      {stage0_53[138], stage0_53[139], stage0_53[140], stage0_53[141], stage0_53[142], stage0_53[143]},
      {stage1_55[23],stage1_54[59],stage1_53[73],stage1_52[123],stage1_51[184]}
   );
   gpc615_5 gpc1967 (
      {stage0_51[240], stage0_51[241], stage0_51[242], stage0_51[243], stage0_51[244]},
      {stage0_52[240]},
      {stage0_53[144], stage0_53[145], stage0_53[146], stage0_53[147], stage0_53[148], stage0_53[149]},
      {stage1_55[24],stage1_54[60],stage1_53[74],stage1_52[124],stage1_51[185]}
   );
   gpc615_5 gpc1968 (
      {stage0_51[245], stage0_51[246], stage0_51[247], stage0_51[248], stage0_51[249]},
      {stage0_52[241]},
      {stage0_53[150], stage0_53[151], stage0_53[152], stage0_53[153], stage0_53[154], stage0_53[155]},
      {stage1_55[25],stage1_54[61],stage1_53[75],stage1_52[125],stage1_51[186]}
   );
   gpc615_5 gpc1969 (
      {stage0_51[250], stage0_51[251], stage0_51[252], stage0_51[253], stage0_51[254]},
      {stage0_52[242]},
      {stage0_53[156], stage0_53[157], stage0_53[158], stage0_53[159], stage0_53[160], stage0_53[161]},
      {stage1_55[26],stage1_54[62],stage1_53[76],stage1_52[126],stage1_51[187]}
   );
   gpc615_5 gpc1970 (
      {stage0_51[255], stage0_51[256], stage0_51[257], stage0_51[258], stage0_51[259]},
      {stage0_52[243]},
      {stage0_53[162], stage0_53[163], stage0_53[164], stage0_53[165], stage0_53[166], stage0_53[167]},
      {stage1_55[27],stage1_54[63],stage1_53[77],stage1_52[127],stage1_51[188]}
   );
   gpc615_5 gpc1971 (
      {stage0_51[260], stage0_51[261], stage0_51[262], stage0_51[263], stage0_51[264]},
      {stage0_52[244]},
      {stage0_53[168], stage0_53[169], stage0_53[170], stage0_53[171], stage0_53[172], stage0_53[173]},
      {stage1_55[28],stage1_54[64],stage1_53[78],stage1_52[128],stage1_51[189]}
   );
   gpc615_5 gpc1972 (
      {stage0_51[265], stage0_51[266], stage0_51[267], stage0_51[268], stage0_51[269]},
      {stage0_52[245]},
      {stage0_53[174], stage0_53[175], stage0_53[176], stage0_53[177], stage0_53[178], stage0_53[179]},
      {stage1_55[29],stage1_54[65],stage1_53[79],stage1_52[129],stage1_51[190]}
   );
   gpc615_5 gpc1973 (
      {stage0_51[270], stage0_51[271], stage0_51[272], stage0_51[273], stage0_51[274]},
      {stage0_52[246]},
      {stage0_53[180], stage0_53[181], stage0_53[182], stage0_53[183], stage0_53[184], stage0_53[185]},
      {stage1_55[30],stage1_54[66],stage1_53[80],stage1_52[130],stage1_51[191]}
   );
   gpc615_5 gpc1974 (
      {stage0_51[275], stage0_51[276], stage0_51[277], stage0_51[278], stage0_51[279]},
      {stage0_52[247]},
      {stage0_53[186], stage0_53[187], stage0_53[188], stage0_53[189], stage0_53[190], stage0_53[191]},
      {stage1_55[31],stage1_54[67],stage1_53[81],stage1_52[131],stage1_51[192]}
   );
   gpc615_5 gpc1975 (
      {stage0_51[280], stage0_51[281], stage0_51[282], stage0_51[283], stage0_51[284]},
      {stage0_52[248]},
      {stage0_53[192], stage0_53[193], stage0_53[194], stage0_53[195], stage0_53[196], stage0_53[197]},
      {stage1_55[32],stage1_54[68],stage1_53[82],stage1_52[132],stage1_51[193]}
   );
   gpc615_5 gpc1976 (
      {stage0_51[285], stage0_51[286], stage0_51[287], stage0_51[288], stage0_51[289]},
      {stage0_52[249]},
      {stage0_53[198], stage0_53[199], stage0_53[200], stage0_53[201], stage0_53[202], stage0_53[203]},
      {stage1_55[33],stage1_54[69],stage1_53[83],stage1_52[133],stage1_51[194]}
   );
   gpc615_5 gpc1977 (
      {stage0_51[290], stage0_51[291], stage0_51[292], stage0_51[293], stage0_51[294]},
      {stage0_52[250]},
      {stage0_53[204], stage0_53[205], stage0_53[206], stage0_53[207], stage0_53[208], stage0_53[209]},
      {stage1_55[34],stage1_54[70],stage1_53[84],stage1_52[134],stage1_51[195]}
   );
   gpc615_5 gpc1978 (
      {stage0_51[295], stage0_51[296], stage0_51[297], stage0_51[298], stage0_51[299]},
      {stage0_52[251]},
      {stage0_53[210], stage0_53[211], stage0_53[212], stage0_53[213], stage0_53[214], stage0_53[215]},
      {stage1_55[35],stage1_54[71],stage1_53[85],stage1_52[135],stage1_51[196]}
   );
   gpc615_5 gpc1979 (
      {stage0_51[300], stage0_51[301], stage0_51[302], stage0_51[303], stage0_51[304]},
      {stage0_52[252]},
      {stage0_53[216], stage0_53[217], stage0_53[218], stage0_53[219], stage0_53[220], stage0_53[221]},
      {stage1_55[36],stage1_54[72],stage1_53[86],stage1_52[136],stage1_51[197]}
   );
   gpc615_5 gpc1980 (
      {stage0_51[305], stage0_51[306], stage0_51[307], stage0_51[308], stage0_51[309]},
      {stage0_52[253]},
      {stage0_53[222], stage0_53[223], stage0_53[224], stage0_53[225], stage0_53[226], stage0_53[227]},
      {stage1_55[37],stage1_54[73],stage1_53[87],stage1_52[137],stage1_51[198]}
   );
   gpc615_5 gpc1981 (
      {stage0_51[310], stage0_51[311], stage0_51[312], stage0_51[313], stage0_51[314]},
      {stage0_52[254]},
      {stage0_53[228], stage0_53[229], stage0_53[230], stage0_53[231], stage0_53[232], stage0_53[233]},
      {stage1_55[38],stage1_54[74],stage1_53[88],stage1_52[138],stage1_51[199]}
   );
   gpc615_5 gpc1982 (
      {stage0_51[315], stage0_51[316], stage0_51[317], stage0_51[318], stage0_51[319]},
      {stage0_52[255]},
      {stage0_53[234], stage0_53[235], stage0_53[236], stage0_53[237], stage0_53[238], stage0_53[239]},
      {stage1_55[39],stage1_54[75],stage1_53[89],stage1_52[139],stage1_51[200]}
   );
   gpc615_5 gpc1983 (
      {stage0_51[320], stage0_51[321], stage0_51[322], stage0_51[323], stage0_51[324]},
      {stage0_52[256]},
      {stage0_53[240], stage0_53[241], stage0_53[242], stage0_53[243], stage0_53[244], stage0_53[245]},
      {stage1_55[40],stage1_54[76],stage1_53[90],stage1_52[140],stage1_51[201]}
   );
   gpc615_5 gpc1984 (
      {stage0_51[325], stage0_51[326], stage0_51[327], stage0_51[328], stage0_51[329]},
      {stage0_52[257]},
      {stage0_53[246], stage0_53[247], stage0_53[248], stage0_53[249], stage0_53[250], stage0_53[251]},
      {stage1_55[41],stage1_54[77],stage1_53[91],stage1_52[141],stage1_51[202]}
   );
   gpc615_5 gpc1985 (
      {stage0_51[330], stage0_51[331], stage0_51[332], stage0_51[333], stage0_51[334]},
      {stage0_52[258]},
      {stage0_53[252], stage0_53[253], stage0_53[254], stage0_53[255], stage0_53[256], stage0_53[257]},
      {stage1_55[42],stage1_54[78],stage1_53[92],stage1_52[142],stage1_51[203]}
   );
   gpc615_5 gpc1986 (
      {stage0_51[335], stage0_51[336], stage0_51[337], stage0_51[338], stage0_51[339]},
      {stage0_52[259]},
      {stage0_53[258], stage0_53[259], stage0_53[260], stage0_53[261], stage0_53[262], stage0_53[263]},
      {stage1_55[43],stage1_54[79],stage1_53[93],stage1_52[143],stage1_51[204]}
   );
   gpc615_5 gpc1987 (
      {stage0_51[340], stage0_51[341], stage0_51[342], stage0_51[343], stage0_51[344]},
      {stage0_52[260]},
      {stage0_53[264], stage0_53[265], stage0_53[266], stage0_53[267], stage0_53[268], stage0_53[269]},
      {stage1_55[44],stage1_54[80],stage1_53[94],stage1_52[144],stage1_51[205]}
   );
   gpc615_5 gpc1988 (
      {stage0_51[345], stage0_51[346], stage0_51[347], stage0_51[348], stage0_51[349]},
      {stage0_52[261]},
      {stage0_53[270], stage0_53[271], stage0_53[272], stage0_53[273], stage0_53[274], stage0_53[275]},
      {stage1_55[45],stage1_54[81],stage1_53[95],stage1_52[145],stage1_51[206]}
   );
   gpc615_5 gpc1989 (
      {stage0_51[350], stage0_51[351], stage0_51[352], stage0_51[353], stage0_51[354]},
      {stage0_52[262]},
      {stage0_53[276], stage0_53[277], stage0_53[278], stage0_53[279], stage0_53[280], stage0_53[281]},
      {stage1_55[46],stage1_54[82],stage1_53[96],stage1_52[146],stage1_51[207]}
   );
   gpc615_5 gpc1990 (
      {stage0_51[355], stage0_51[356], stage0_51[357], stage0_51[358], stage0_51[359]},
      {stage0_52[263]},
      {stage0_53[282], stage0_53[283], stage0_53[284], stage0_53[285], stage0_53[286], stage0_53[287]},
      {stage1_55[47],stage1_54[83],stage1_53[97],stage1_52[147],stage1_51[208]}
   );
   gpc615_5 gpc1991 (
      {stage0_51[360], stage0_51[361], stage0_51[362], stage0_51[363], stage0_51[364]},
      {stage0_52[264]},
      {stage0_53[288], stage0_53[289], stage0_53[290], stage0_53[291], stage0_53[292], stage0_53[293]},
      {stage1_55[48],stage1_54[84],stage1_53[98],stage1_52[148],stage1_51[209]}
   );
   gpc615_5 gpc1992 (
      {stage0_51[365], stage0_51[366], stage0_51[367], stage0_51[368], stage0_51[369]},
      {stage0_52[265]},
      {stage0_53[294], stage0_53[295], stage0_53[296], stage0_53[297], stage0_53[298], stage0_53[299]},
      {stage1_55[49],stage1_54[85],stage1_53[99],stage1_52[149],stage1_51[210]}
   );
   gpc615_5 gpc1993 (
      {stage0_51[370], stage0_51[371], stage0_51[372], stage0_51[373], stage0_51[374]},
      {stage0_52[266]},
      {stage0_53[300], stage0_53[301], stage0_53[302], stage0_53[303], stage0_53[304], stage0_53[305]},
      {stage1_55[50],stage1_54[86],stage1_53[100],stage1_52[150],stage1_51[211]}
   );
   gpc615_5 gpc1994 (
      {stage0_51[375], stage0_51[376], stage0_51[377], stage0_51[378], stage0_51[379]},
      {stage0_52[267]},
      {stage0_53[306], stage0_53[307], stage0_53[308], stage0_53[309], stage0_53[310], stage0_53[311]},
      {stage1_55[51],stage1_54[87],stage1_53[101],stage1_52[151],stage1_51[212]}
   );
   gpc615_5 gpc1995 (
      {stage0_51[380], stage0_51[381], stage0_51[382], stage0_51[383], stage0_51[384]},
      {stage0_52[268]},
      {stage0_53[312], stage0_53[313], stage0_53[314], stage0_53[315], stage0_53[316], stage0_53[317]},
      {stage1_55[52],stage1_54[88],stage1_53[102],stage1_52[152],stage1_51[213]}
   );
   gpc615_5 gpc1996 (
      {stage0_51[385], stage0_51[386], stage0_51[387], stage0_51[388], stage0_51[389]},
      {stage0_52[269]},
      {stage0_53[318], stage0_53[319], stage0_53[320], stage0_53[321], stage0_53[322], stage0_53[323]},
      {stage1_55[53],stage1_54[89],stage1_53[103],stage1_52[153],stage1_51[214]}
   );
   gpc615_5 gpc1997 (
      {stage0_51[390], stage0_51[391], stage0_51[392], stage0_51[393], stage0_51[394]},
      {stage0_52[270]},
      {stage0_53[324], stage0_53[325], stage0_53[326], stage0_53[327], stage0_53[328], stage0_53[329]},
      {stage1_55[54],stage1_54[90],stage1_53[104],stage1_52[154],stage1_51[215]}
   );
   gpc615_5 gpc1998 (
      {stage0_51[395], stage0_51[396], stage0_51[397], stage0_51[398], stage0_51[399]},
      {stage0_52[271]},
      {stage0_53[330], stage0_53[331], stage0_53[332], stage0_53[333], stage0_53[334], stage0_53[335]},
      {stage1_55[55],stage1_54[91],stage1_53[105],stage1_52[155],stage1_51[216]}
   );
   gpc615_5 gpc1999 (
      {stage0_51[400], stage0_51[401], stage0_51[402], stage0_51[403], stage0_51[404]},
      {stage0_52[272]},
      {stage0_53[336], stage0_53[337], stage0_53[338], stage0_53[339], stage0_53[340], stage0_53[341]},
      {stage1_55[56],stage1_54[92],stage1_53[106],stage1_52[156],stage1_51[217]}
   );
   gpc615_5 gpc2000 (
      {stage0_51[405], stage0_51[406], stage0_51[407], stage0_51[408], stage0_51[409]},
      {stage0_52[273]},
      {stage0_53[342], stage0_53[343], stage0_53[344], stage0_53[345], stage0_53[346], stage0_53[347]},
      {stage1_55[57],stage1_54[93],stage1_53[107],stage1_52[157],stage1_51[218]}
   );
   gpc615_5 gpc2001 (
      {stage0_51[410], stage0_51[411], stage0_51[412], stage0_51[413], stage0_51[414]},
      {stage0_52[274]},
      {stage0_53[348], stage0_53[349], stage0_53[350], stage0_53[351], stage0_53[352], stage0_53[353]},
      {stage1_55[58],stage1_54[94],stage1_53[108],stage1_52[158],stage1_51[219]}
   );
   gpc615_5 gpc2002 (
      {stage0_51[415], stage0_51[416], stage0_51[417], stage0_51[418], stage0_51[419]},
      {stage0_52[275]},
      {stage0_53[354], stage0_53[355], stage0_53[356], stage0_53[357], stage0_53[358], stage0_53[359]},
      {stage1_55[59],stage1_54[95],stage1_53[109],stage1_52[159],stage1_51[220]}
   );
   gpc615_5 gpc2003 (
      {stage0_51[420], stage0_51[421], stage0_51[422], stage0_51[423], stage0_51[424]},
      {stage0_52[276]},
      {stage0_53[360], stage0_53[361], stage0_53[362], stage0_53[363], stage0_53[364], stage0_53[365]},
      {stage1_55[60],stage1_54[96],stage1_53[110],stage1_52[160],stage1_51[221]}
   );
   gpc615_5 gpc2004 (
      {stage0_51[425], stage0_51[426], stage0_51[427], stage0_51[428], stage0_51[429]},
      {stage0_52[277]},
      {stage0_53[366], stage0_53[367], stage0_53[368], stage0_53[369], stage0_53[370], stage0_53[371]},
      {stage1_55[61],stage1_54[97],stage1_53[111],stage1_52[161],stage1_51[222]}
   );
   gpc615_5 gpc2005 (
      {stage0_51[430], stage0_51[431], stage0_51[432], stage0_51[433], stage0_51[434]},
      {stage0_52[278]},
      {stage0_53[372], stage0_53[373], stage0_53[374], stage0_53[375], stage0_53[376], stage0_53[377]},
      {stage1_55[62],stage1_54[98],stage1_53[112],stage1_52[162],stage1_51[223]}
   );
   gpc606_5 gpc2006 (
      {stage0_52[279], stage0_52[280], stage0_52[281], stage0_52[282], stage0_52[283], stage0_52[284]},
      {stage0_54[0], stage0_54[1], stage0_54[2], stage0_54[3], stage0_54[4], stage0_54[5]},
      {stage1_56[0],stage1_55[63],stage1_54[99],stage1_53[113],stage1_52[163]}
   );
   gpc606_5 gpc2007 (
      {stage0_52[285], stage0_52[286], stage0_52[287], stage0_52[288], stage0_52[289], stage0_52[290]},
      {stage0_54[6], stage0_54[7], stage0_54[8], stage0_54[9], stage0_54[10], stage0_54[11]},
      {stage1_56[1],stage1_55[64],stage1_54[100],stage1_53[114],stage1_52[164]}
   );
   gpc606_5 gpc2008 (
      {stage0_52[291], stage0_52[292], stage0_52[293], stage0_52[294], stage0_52[295], stage0_52[296]},
      {stage0_54[12], stage0_54[13], stage0_54[14], stage0_54[15], stage0_54[16], stage0_54[17]},
      {stage1_56[2],stage1_55[65],stage1_54[101],stage1_53[115],stage1_52[165]}
   );
   gpc606_5 gpc2009 (
      {stage0_52[297], stage0_52[298], stage0_52[299], stage0_52[300], stage0_52[301], stage0_52[302]},
      {stage0_54[18], stage0_54[19], stage0_54[20], stage0_54[21], stage0_54[22], stage0_54[23]},
      {stage1_56[3],stage1_55[66],stage1_54[102],stage1_53[116],stage1_52[166]}
   );
   gpc606_5 gpc2010 (
      {stage0_52[303], stage0_52[304], stage0_52[305], stage0_52[306], stage0_52[307], stage0_52[308]},
      {stage0_54[24], stage0_54[25], stage0_54[26], stage0_54[27], stage0_54[28], stage0_54[29]},
      {stage1_56[4],stage1_55[67],stage1_54[103],stage1_53[117],stage1_52[167]}
   );
   gpc606_5 gpc2011 (
      {stage0_52[309], stage0_52[310], stage0_52[311], stage0_52[312], stage0_52[313], stage0_52[314]},
      {stage0_54[30], stage0_54[31], stage0_54[32], stage0_54[33], stage0_54[34], stage0_54[35]},
      {stage1_56[5],stage1_55[68],stage1_54[104],stage1_53[118],stage1_52[168]}
   );
   gpc606_5 gpc2012 (
      {stage0_52[315], stage0_52[316], stage0_52[317], stage0_52[318], stage0_52[319], stage0_52[320]},
      {stage0_54[36], stage0_54[37], stage0_54[38], stage0_54[39], stage0_54[40], stage0_54[41]},
      {stage1_56[6],stage1_55[69],stage1_54[105],stage1_53[119],stage1_52[169]}
   );
   gpc606_5 gpc2013 (
      {stage0_52[321], stage0_52[322], stage0_52[323], stage0_52[324], stage0_52[325], stage0_52[326]},
      {stage0_54[42], stage0_54[43], stage0_54[44], stage0_54[45], stage0_54[46], stage0_54[47]},
      {stage1_56[7],stage1_55[70],stage1_54[106],stage1_53[120],stage1_52[170]}
   );
   gpc606_5 gpc2014 (
      {stage0_52[327], stage0_52[328], stage0_52[329], stage0_52[330], stage0_52[331], stage0_52[332]},
      {stage0_54[48], stage0_54[49], stage0_54[50], stage0_54[51], stage0_54[52], stage0_54[53]},
      {stage1_56[8],stage1_55[71],stage1_54[107],stage1_53[121],stage1_52[171]}
   );
   gpc606_5 gpc2015 (
      {stage0_52[333], stage0_52[334], stage0_52[335], stage0_52[336], stage0_52[337], stage0_52[338]},
      {stage0_54[54], stage0_54[55], stage0_54[56], stage0_54[57], stage0_54[58], stage0_54[59]},
      {stage1_56[9],stage1_55[72],stage1_54[108],stage1_53[122],stage1_52[172]}
   );
   gpc606_5 gpc2016 (
      {stage0_52[339], stage0_52[340], stage0_52[341], stage0_52[342], stage0_52[343], stage0_52[344]},
      {stage0_54[60], stage0_54[61], stage0_54[62], stage0_54[63], stage0_54[64], stage0_54[65]},
      {stage1_56[10],stage1_55[73],stage1_54[109],stage1_53[123],stage1_52[173]}
   );
   gpc606_5 gpc2017 (
      {stage0_52[345], stage0_52[346], stage0_52[347], stage0_52[348], stage0_52[349], stage0_52[350]},
      {stage0_54[66], stage0_54[67], stage0_54[68], stage0_54[69], stage0_54[70], stage0_54[71]},
      {stage1_56[11],stage1_55[74],stage1_54[110],stage1_53[124],stage1_52[174]}
   );
   gpc606_5 gpc2018 (
      {stage0_52[351], stage0_52[352], stage0_52[353], stage0_52[354], stage0_52[355], stage0_52[356]},
      {stage0_54[72], stage0_54[73], stage0_54[74], stage0_54[75], stage0_54[76], stage0_54[77]},
      {stage1_56[12],stage1_55[75],stage1_54[111],stage1_53[125],stage1_52[175]}
   );
   gpc606_5 gpc2019 (
      {stage0_52[357], stage0_52[358], stage0_52[359], stage0_52[360], stage0_52[361], stage0_52[362]},
      {stage0_54[78], stage0_54[79], stage0_54[80], stage0_54[81], stage0_54[82], stage0_54[83]},
      {stage1_56[13],stage1_55[76],stage1_54[112],stage1_53[126],stage1_52[176]}
   );
   gpc606_5 gpc2020 (
      {stage0_52[363], stage0_52[364], stage0_52[365], stage0_52[366], stage0_52[367], stage0_52[368]},
      {stage0_54[84], stage0_54[85], stage0_54[86], stage0_54[87], stage0_54[88], stage0_54[89]},
      {stage1_56[14],stage1_55[77],stage1_54[113],stage1_53[127],stage1_52[177]}
   );
   gpc606_5 gpc2021 (
      {stage0_52[369], stage0_52[370], stage0_52[371], stage0_52[372], stage0_52[373], stage0_52[374]},
      {stage0_54[90], stage0_54[91], stage0_54[92], stage0_54[93], stage0_54[94], stage0_54[95]},
      {stage1_56[15],stage1_55[78],stage1_54[114],stage1_53[128],stage1_52[178]}
   );
   gpc606_5 gpc2022 (
      {stage0_52[375], stage0_52[376], stage0_52[377], stage0_52[378], stage0_52[379], stage0_52[380]},
      {stage0_54[96], stage0_54[97], stage0_54[98], stage0_54[99], stage0_54[100], stage0_54[101]},
      {stage1_56[16],stage1_55[79],stage1_54[115],stage1_53[129],stage1_52[179]}
   );
   gpc606_5 gpc2023 (
      {stage0_52[381], stage0_52[382], stage0_52[383], stage0_52[384], stage0_52[385], stage0_52[386]},
      {stage0_54[102], stage0_54[103], stage0_54[104], stage0_54[105], stage0_54[106], stage0_54[107]},
      {stage1_56[17],stage1_55[80],stage1_54[116],stage1_53[130],stage1_52[180]}
   );
   gpc606_5 gpc2024 (
      {stage0_52[387], stage0_52[388], stage0_52[389], stage0_52[390], stage0_52[391], stage0_52[392]},
      {stage0_54[108], stage0_54[109], stage0_54[110], stage0_54[111], stage0_54[112], stage0_54[113]},
      {stage1_56[18],stage1_55[81],stage1_54[117],stage1_53[131],stage1_52[181]}
   );
   gpc606_5 gpc2025 (
      {stage0_52[393], stage0_52[394], stage0_52[395], stage0_52[396], stage0_52[397], stage0_52[398]},
      {stage0_54[114], stage0_54[115], stage0_54[116], stage0_54[117], stage0_54[118], stage0_54[119]},
      {stage1_56[19],stage1_55[82],stage1_54[118],stage1_53[132],stage1_52[182]}
   );
   gpc606_5 gpc2026 (
      {stage0_52[399], stage0_52[400], stage0_52[401], stage0_52[402], stage0_52[403], stage0_52[404]},
      {stage0_54[120], stage0_54[121], stage0_54[122], stage0_54[123], stage0_54[124], stage0_54[125]},
      {stage1_56[20],stage1_55[83],stage1_54[119],stage1_53[133],stage1_52[183]}
   );
   gpc606_5 gpc2027 (
      {stage0_52[405], stage0_52[406], stage0_52[407], stage0_52[408], stage0_52[409], stage0_52[410]},
      {stage0_54[126], stage0_54[127], stage0_54[128], stage0_54[129], stage0_54[130], stage0_54[131]},
      {stage1_56[21],stage1_55[84],stage1_54[120],stage1_53[134],stage1_52[184]}
   );
   gpc606_5 gpc2028 (
      {stage0_52[411], stage0_52[412], stage0_52[413], stage0_52[414], stage0_52[415], stage0_52[416]},
      {stage0_54[132], stage0_54[133], stage0_54[134], stage0_54[135], stage0_54[136], stage0_54[137]},
      {stage1_56[22],stage1_55[85],stage1_54[121],stage1_53[135],stage1_52[185]}
   );
   gpc606_5 gpc2029 (
      {stage0_52[417], stage0_52[418], stage0_52[419], stage0_52[420], stage0_52[421], stage0_52[422]},
      {stage0_54[138], stage0_54[139], stage0_54[140], stage0_54[141], stage0_54[142], stage0_54[143]},
      {stage1_56[23],stage1_55[86],stage1_54[122],stage1_53[136],stage1_52[186]}
   );
   gpc606_5 gpc2030 (
      {stage0_52[423], stage0_52[424], stage0_52[425], stage0_52[426], stage0_52[427], stage0_52[428]},
      {stage0_54[144], stage0_54[145], stage0_54[146], stage0_54[147], stage0_54[148], stage0_54[149]},
      {stage1_56[24],stage1_55[87],stage1_54[123],stage1_53[137],stage1_52[187]}
   );
   gpc606_5 gpc2031 (
      {stage0_52[429], stage0_52[430], stage0_52[431], stage0_52[432], stage0_52[433], stage0_52[434]},
      {stage0_54[150], stage0_54[151], stage0_54[152], stage0_54[153], stage0_54[154], stage0_54[155]},
      {stage1_56[25],stage1_55[88],stage1_54[124],stage1_53[138],stage1_52[188]}
   );
   gpc606_5 gpc2032 (
      {stage0_52[435], stage0_52[436], stage0_52[437], stage0_52[438], stage0_52[439], stage0_52[440]},
      {stage0_54[156], stage0_54[157], stage0_54[158], stage0_54[159], stage0_54[160], stage0_54[161]},
      {stage1_56[26],stage1_55[89],stage1_54[125],stage1_53[139],stage1_52[189]}
   );
   gpc606_5 gpc2033 (
      {stage0_52[441], stage0_52[442], stage0_52[443], stage0_52[444], stage0_52[445], stage0_52[446]},
      {stage0_54[162], stage0_54[163], stage0_54[164], stage0_54[165], stage0_54[166], stage0_54[167]},
      {stage1_56[27],stage1_55[90],stage1_54[126],stage1_53[140],stage1_52[190]}
   );
   gpc615_5 gpc2034 (
      {stage0_52[447], stage0_52[448], stage0_52[449], stage0_52[450], stage0_52[451]},
      {stage0_53[378]},
      {stage0_54[168], stage0_54[169], stage0_54[170], stage0_54[171], stage0_54[172], stage0_54[173]},
      {stage1_56[28],stage1_55[91],stage1_54[127],stage1_53[141],stage1_52[191]}
   );
   gpc615_5 gpc2035 (
      {stage0_52[452], stage0_52[453], stage0_52[454], stage0_52[455], stage0_52[456]},
      {stage0_53[379]},
      {stage0_54[174], stage0_54[175], stage0_54[176], stage0_54[177], stage0_54[178], stage0_54[179]},
      {stage1_56[29],stage1_55[92],stage1_54[128],stage1_53[142],stage1_52[192]}
   );
   gpc615_5 gpc2036 (
      {stage0_52[457], stage0_52[458], stage0_52[459], stage0_52[460], stage0_52[461]},
      {stage0_53[380]},
      {stage0_54[180], stage0_54[181], stage0_54[182], stage0_54[183], stage0_54[184], stage0_54[185]},
      {stage1_56[30],stage1_55[93],stage1_54[129],stage1_53[143],stage1_52[193]}
   );
   gpc615_5 gpc2037 (
      {stage0_52[462], stage0_52[463], stage0_52[464], stage0_52[465], stage0_52[466]},
      {stage0_53[381]},
      {stage0_54[186], stage0_54[187], stage0_54[188], stage0_54[189], stage0_54[190], stage0_54[191]},
      {stage1_56[31],stage1_55[94],stage1_54[130],stage1_53[144],stage1_52[194]}
   );
   gpc615_5 gpc2038 (
      {stage0_52[467], stage0_52[468], stage0_52[469], stage0_52[470], stage0_52[471]},
      {stage0_53[382]},
      {stage0_54[192], stage0_54[193], stage0_54[194], stage0_54[195], stage0_54[196], stage0_54[197]},
      {stage1_56[32],stage1_55[95],stage1_54[131],stage1_53[145],stage1_52[195]}
   );
   gpc615_5 gpc2039 (
      {stage0_52[472], stage0_52[473], stage0_52[474], stage0_52[475], stage0_52[476]},
      {stage0_53[383]},
      {stage0_54[198], stage0_54[199], stage0_54[200], stage0_54[201], stage0_54[202], stage0_54[203]},
      {stage1_56[33],stage1_55[96],stage1_54[132],stage1_53[146],stage1_52[196]}
   );
   gpc615_5 gpc2040 (
      {stage0_52[477], stage0_52[478], stage0_52[479], stage0_52[480], stage0_52[481]},
      {stage0_53[384]},
      {stage0_54[204], stage0_54[205], stage0_54[206], stage0_54[207], stage0_54[208], stage0_54[209]},
      {stage1_56[34],stage1_55[97],stage1_54[133],stage1_53[147],stage1_52[197]}
   );
   gpc615_5 gpc2041 (
      {stage0_52[482], stage0_52[483], stage0_52[484], stage0_52[485], 1'b0},
      {stage0_53[385]},
      {stage0_54[210], stage0_54[211], stage0_54[212], stage0_54[213], stage0_54[214], stage0_54[215]},
      {stage1_56[35],stage1_55[98],stage1_54[134],stage1_53[148],stage1_52[198]}
   );
   gpc615_5 gpc2042 (
      {stage0_53[386], stage0_53[387], stage0_53[388], stage0_53[389], stage0_53[390]},
      {stage0_54[216]},
      {stage0_55[0], stage0_55[1], stage0_55[2], stage0_55[3], stage0_55[4], stage0_55[5]},
      {stage1_57[0],stage1_56[36],stage1_55[99],stage1_54[135],stage1_53[149]}
   );
   gpc615_5 gpc2043 (
      {stage0_53[391], stage0_53[392], stage0_53[393], stage0_53[394], stage0_53[395]},
      {stage0_54[217]},
      {stage0_55[6], stage0_55[7], stage0_55[8], stage0_55[9], stage0_55[10], stage0_55[11]},
      {stage1_57[1],stage1_56[37],stage1_55[100],stage1_54[136],stage1_53[150]}
   );
   gpc615_5 gpc2044 (
      {stage0_53[396], stage0_53[397], stage0_53[398], stage0_53[399], stage0_53[400]},
      {stage0_54[218]},
      {stage0_55[12], stage0_55[13], stage0_55[14], stage0_55[15], stage0_55[16], stage0_55[17]},
      {stage1_57[2],stage1_56[38],stage1_55[101],stage1_54[137],stage1_53[151]}
   );
   gpc615_5 gpc2045 (
      {stage0_53[401], stage0_53[402], stage0_53[403], stage0_53[404], stage0_53[405]},
      {stage0_54[219]},
      {stage0_55[18], stage0_55[19], stage0_55[20], stage0_55[21], stage0_55[22], stage0_55[23]},
      {stage1_57[3],stage1_56[39],stage1_55[102],stage1_54[138],stage1_53[152]}
   );
   gpc615_5 gpc2046 (
      {stage0_53[406], stage0_53[407], stage0_53[408], stage0_53[409], stage0_53[410]},
      {stage0_54[220]},
      {stage0_55[24], stage0_55[25], stage0_55[26], stage0_55[27], stage0_55[28], stage0_55[29]},
      {stage1_57[4],stage1_56[40],stage1_55[103],stage1_54[139],stage1_53[153]}
   );
   gpc615_5 gpc2047 (
      {stage0_53[411], stage0_53[412], stage0_53[413], stage0_53[414], stage0_53[415]},
      {stage0_54[221]},
      {stage0_55[30], stage0_55[31], stage0_55[32], stage0_55[33], stage0_55[34], stage0_55[35]},
      {stage1_57[5],stage1_56[41],stage1_55[104],stage1_54[140],stage1_53[154]}
   );
   gpc615_5 gpc2048 (
      {stage0_53[416], stage0_53[417], stage0_53[418], stage0_53[419], stage0_53[420]},
      {stage0_54[222]},
      {stage0_55[36], stage0_55[37], stage0_55[38], stage0_55[39], stage0_55[40], stage0_55[41]},
      {stage1_57[6],stage1_56[42],stage1_55[105],stage1_54[141],stage1_53[155]}
   );
   gpc615_5 gpc2049 (
      {stage0_53[421], stage0_53[422], stage0_53[423], stage0_53[424], stage0_53[425]},
      {stage0_54[223]},
      {stage0_55[42], stage0_55[43], stage0_55[44], stage0_55[45], stage0_55[46], stage0_55[47]},
      {stage1_57[7],stage1_56[43],stage1_55[106],stage1_54[142],stage1_53[156]}
   );
   gpc615_5 gpc2050 (
      {stage0_53[426], stage0_53[427], stage0_53[428], stage0_53[429], stage0_53[430]},
      {stage0_54[224]},
      {stage0_55[48], stage0_55[49], stage0_55[50], stage0_55[51], stage0_55[52], stage0_55[53]},
      {stage1_57[8],stage1_56[44],stage1_55[107],stage1_54[143],stage1_53[157]}
   );
   gpc615_5 gpc2051 (
      {stage0_53[431], stage0_53[432], stage0_53[433], stage0_53[434], stage0_53[435]},
      {stage0_54[225]},
      {stage0_55[54], stage0_55[55], stage0_55[56], stage0_55[57], stage0_55[58], stage0_55[59]},
      {stage1_57[9],stage1_56[45],stage1_55[108],stage1_54[144],stage1_53[158]}
   );
   gpc615_5 gpc2052 (
      {stage0_53[436], stage0_53[437], stage0_53[438], stage0_53[439], stage0_53[440]},
      {stage0_54[226]},
      {stage0_55[60], stage0_55[61], stage0_55[62], stage0_55[63], stage0_55[64], stage0_55[65]},
      {stage1_57[10],stage1_56[46],stage1_55[109],stage1_54[145],stage1_53[159]}
   );
   gpc615_5 gpc2053 (
      {stage0_53[441], stage0_53[442], stage0_53[443], stage0_53[444], stage0_53[445]},
      {stage0_54[227]},
      {stage0_55[66], stage0_55[67], stage0_55[68], stage0_55[69], stage0_55[70], stage0_55[71]},
      {stage1_57[11],stage1_56[47],stage1_55[110],stage1_54[146],stage1_53[160]}
   );
   gpc615_5 gpc2054 (
      {stage0_53[446], stage0_53[447], stage0_53[448], stage0_53[449], stage0_53[450]},
      {stage0_54[228]},
      {stage0_55[72], stage0_55[73], stage0_55[74], stage0_55[75], stage0_55[76], stage0_55[77]},
      {stage1_57[12],stage1_56[48],stage1_55[111],stage1_54[147],stage1_53[161]}
   );
   gpc615_5 gpc2055 (
      {stage0_53[451], stage0_53[452], stage0_53[453], stage0_53[454], stage0_53[455]},
      {stage0_54[229]},
      {stage0_55[78], stage0_55[79], stage0_55[80], stage0_55[81], stage0_55[82], stage0_55[83]},
      {stage1_57[13],stage1_56[49],stage1_55[112],stage1_54[148],stage1_53[162]}
   );
   gpc615_5 gpc2056 (
      {stage0_53[456], stage0_53[457], stage0_53[458], stage0_53[459], stage0_53[460]},
      {stage0_54[230]},
      {stage0_55[84], stage0_55[85], stage0_55[86], stage0_55[87], stage0_55[88], stage0_55[89]},
      {stage1_57[14],stage1_56[50],stage1_55[113],stage1_54[149],stage1_53[163]}
   );
   gpc615_5 gpc2057 (
      {stage0_53[461], stage0_53[462], stage0_53[463], stage0_53[464], stage0_53[465]},
      {stage0_54[231]},
      {stage0_55[90], stage0_55[91], stage0_55[92], stage0_55[93], stage0_55[94], stage0_55[95]},
      {stage1_57[15],stage1_56[51],stage1_55[114],stage1_54[150],stage1_53[164]}
   );
   gpc615_5 gpc2058 (
      {stage0_53[466], stage0_53[467], stage0_53[468], stage0_53[469], stage0_53[470]},
      {stage0_54[232]},
      {stage0_55[96], stage0_55[97], stage0_55[98], stage0_55[99], stage0_55[100], stage0_55[101]},
      {stage1_57[16],stage1_56[52],stage1_55[115],stage1_54[151],stage1_53[165]}
   );
   gpc615_5 gpc2059 (
      {stage0_53[471], stage0_53[472], stage0_53[473], stage0_53[474], stage0_53[475]},
      {stage0_54[233]},
      {stage0_55[102], stage0_55[103], stage0_55[104], stage0_55[105], stage0_55[106], stage0_55[107]},
      {stage1_57[17],stage1_56[53],stage1_55[116],stage1_54[152],stage1_53[166]}
   );
   gpc615_5 gpc2060 (
      {stage0_53[476], stage0_53[477], stage0_53[478], stage0_53[479], stage0_53[480]},
      {stage0_54[234]},
      {stage0_55[108], stage0_55[109], stage0_55[110], stage0_55[111], stage0_55[112], stage0_55[113]},
      {stage1_57[18],stage1_56[54],stage1_55[117],stage1_54[153],stage1_53[167]}
   );
   gpc615_5 gpc2061 (
      {stage0_53[481], stage0_53[482], stage0_53[483], stage0_53[484], stage0_53[485]},
      {stage0_54[235]},
      {stage0_55[114], stage0_55[115], stage0_55[116], stage0_55[117], stage0_55[118], stage0_55[119]},
      {stage1_57[19],stage1_56[55],stage1_55[118],stage1_54[154],stage1_53[168]}
   );
   gpc117_4 gpc2062 (
      {stage0_54[236], stage0_54[237], stage0_54[238], stage0_54[239], stage0_54[240], stage0_54[241], stage0_54[242]},
      {stage0_55[120]},
      {stage0_56[0]},
      {stage1_57[20],stage1_56[56],stage1_55[119],stage1_54[155]}
   );
   gpc615_5 gpc2063 (
      {stage0_54[243], stage0_54[244], stage0_54[245], stage0_54[246], stage0_54[247]},
      {stage0_55[121]},
      {stage0_56[1], stage0_56[2], stage0_56[3], stage0_56[4], stage0_56[5], stage0_56[6]},
      {stage1_58[0],stage1_57[21],stage1_56[57],stage1_55[120],stage1_54[156]}
   );
   gpc615_5 gpc2064 (
      {stage0_54[248], stage0_54[249], stage0_54[250], stage0_54[251], stage0_54[252]},
      {stage0_55[122]},
      {stage0_56[7], stage0_56[8], stage0_56[9], stage0_56[10], stage0_56[11], stage0_56[12]},
      {stage1_58[1],stage1_57[22],stage1_56[58],stage1_55[121],stage1_54[157]}
   );
   gpc615_5 gpc2065 (
      {stage0_54[253], stage0_54[254], stage0_54[255], stage0_54[256], stage0_54[257]},
      {stage0_55[123]},
      {stage0_56[13], stage0_56[14], stage0_56[15], stage0_56[16], stage0_56[17], stage0_56[18]},
      {stage1_58[2],stage1_57[23],stage1_56[59],stage1_55[122],stage1_54[158]}
   );
   gpc615_5 gpc2066 (
      {stage0_54[258], stage0_54[259], stage0_54[260], stage0_54[261], stage0_54[262]},
      {stage0_55[124]},
      {stage0_56[19], stage0_56[20], stage0_56[21], stage0_56[22], stage0_56[23], stage0_56[24]},
      {stage1_58[3],stage1_57[24],stage1_56[60],stage1_55[123],stage1_54[159]}
   );
   gpc615_5 gpc2067 (
      {stage0_54[263], stage0_54[264], stage0_54[265], stage0_54[266], stage0_54[267]},
      {stage0_55[125]},
      {stage0_56[25], stage0_56[26], stage0_56[27], stage0_56[28], stage0_56[29], stage0_56[30]},
      {stage1_58[4],stage1_57[25],stage1_56[61],stage1_55[124],stage1_54[160]}
   );
   gpc615_5 gpc2068 (
      {stage0_54[268], stage0_54[269], stage0_54[270], stage0_54[271], stage0_54[272]},
      {stage0_55[126]},
      {stage0_56[31], stage0_56[32], stage0_56[33], stage0_56[34], stage0_56[35], stage0_56[36]},
      {stage1_58[5],stage1_57[26],stage1_56[62],stage1_55[125],stage1_54[161]}
   );
   gpc615_5 gpc2069 (
      {stage0_54[273], stage0_54[274], stage0_54[275], stage0_54[276], stage0_54[277]},
      {stage0_55[127]},
      {stage0_56[37], stage0_56[38], stage0_56[39], stage0_56[40], stage0_56[41], stage0_56[42]},
      {stage1_58[6],stage1_57[27],stage1_56[63],stage1_55[126],stage1_54[162]}
   );
   gpc615_5 gpc2070 (
      {stage0_54[278], stage0_54[279], stage0_54[280], stage0_54[281], stage0_54[282]},
      {stage0_55[128]},
      {stage0_56[43], stage0_56[44], stage0_56[45], stage0_56[46], stage0_56[47], stage0_56[48]},
      {stage1_58[7],stage1_57[28],stage1_56[64],stage1_55[127],stage1_54[163]}
   );
   gpc615_5 gpc2071 (
      {stage0_54[283], stage0_54[284], stage0_54[285], stage0_54[286], stage0_54[287]},
      {stage0_55[129]},
      {stage0_56[49], stage0_56[50], stage0_56[51], stage0_56[52], stage0_56[53], stage0_56[54]},
      {stage1_58[8],stage1_57[29],stage1_56[65],stage1_55[128],stage1_54[164]}
   );
   gpc615_5 gpc2072 (
      {stage0_54[288], stage0_54[289], stage0_54[290], stage0_54[291], stage0_54[292]},
      {stage0_55[130]},
      {stage0_56[55], stage0_56[56], stage0_56[57], stage0_56[58], stage0_56[59], stage0_56[60]},
      {stage1_58[9],stage1_57[30],stage1_56[66],stage1_55[129],stage1_54[165]}
   );
   gpc615_5 gpc2073 (
      {stage0_54[293], stage0_54[294], stage0_54[295], stage0_54[296], stage0_54[297]},
      {stage0_55[131]},
      {stage0_56[61], stage0_56[62], stage0_56[63], stage0_56[64], stage0_56[65], stage0_56[66]},
      {stage1_58[10],stage1_57[31],stage1_56[67],stage1_55[130],stage1_54[166]}
   );
   gpc615_5 gpc2074 (
      {stage0_54[298], stage0_54[299], stage0_54[300], stage0_54[301], stage0_54[302]},
      {stage0_55[132]},
      {stage0_56[67], stage0_56[68], stage0_56[69], stage0_56[70], stage0_56[71], stage0_56[72]},
      {stage1_58[11],stage1_57[32],stage1_56[68],stage1_55[131],stage1_54[167]}
   );
   gpc615_5 gpc2075 (
      {stage0_54[303], stage0_54[304], stage0_54[305], stage0_54[306], stage0_54[307]},
      {stage0_55[133]},
      {stage0_56[73], stage0_56[74], stage0_56[75], stage0_56[76], stage0_56[77], stage0_56[78]},
      {stage1_58[12],stage1_57[33],stage1_56[69],stage1_55[132],stage1_54[168]}
   );
   gpc615_5 gpc2076 (
      {stage0_54[308], stage0_54[309], stage0_54[310], stage0_54[311], stage0_54[312]},
      {stage0_55[134]},
      {stage0_56[79], stage0_56[80], stage0_56[81], stage0_56[82], stage0_56[83], stage0_56[84]},
      {stage1_58[13],stage1_57[34],stage1_56[70],stage1_55[133],stage1_54[169]}
   );
   gpc615_5 gpc2077 (
      {stage0_54[313], stage0_54[314], stage0_54[315], stage0_54[316], stage0_54[317]},
      {stage0_55[135]},
      {stage0_56[85], stage0_56[86], stage0_56[87], stage0_56[88], stage0_56[89], stage0_56[90]},
      {stage1_58[14],stage1_57[35],stage1_56[71],stage1_55[134],stage1_54[170]}
   );
   gpc615_5 gpc2078 (
      {stage0_54[318], stage0_54[319], stage0_54[320], stage0_54[321], stage0_54[322]},
      {stage0_55[136]},
      {stage0_56[91], stage0_56[92], stage0_56[93], stage0_56[94], stage0_56[95], stage0_56[96]},
      {stage1_58[15],stage1_57[36],stage1_56[72],stage1_55[135],stage1_54[171]}
   );
   gpc615_5 gpc2079 (
      {stage0_54[323], stage0_54[324], stage0_54[325], stage0_54[326], stage0_54[327]},
      {stage0_55[137]},
      {stage0_56[97], stage0_56[98], stage0_56[99], stage0_56[100], stage0_56[101], stage0_56[102]},
      {stage1_58[16],stage1_57[37],stage1_56[73],stage1_55[136],stage1_54[172]}
   );
   gpc615_5 gpc2080 (
      {stage0_54[328], stage0_54[329], stage0_54[330], stage0_54[331], stage0_54[332]},
      {stage0_55[138]},
      {stage0_56[103], stage0_56[104], stage0_56[105], stage0_56[106], stage0_56[107], stage0_56[108]},
      {stage1_58[17],stage1_57[38],stage1_56[74],stage1_55[137],stage1_54[173]}
   );
   gpc615_5 gpc2081 (
      {stage0_54[333], stage0_54[334], stage0_54[335], stage0_54[336], stage0_54[337]},
      {stage0_55[139]},
      {stage0_56[109], stage0_56[110], stage0_56[111], stage0_56[112], stage0_56[113], stage0_56[114]},
      {stage1_58[18],stage1_57[39],stage1_56[75],stage1_55[138],stage1_54[174]}
   );
   gpc615_5 gpc2082 (
      {stage0_54[338], stage0_54[339], stage0_54[340], stage0_54[341], stage0_54[342]},
      {stage0_55[140]},
      {stage0_56[115], stage0_56[116], stage0_56[117], stage0_56[118], stage0_56[119], stage0_56[120]},
      {stage1_58[19],stage1_57[40],stage1_56[76],stage1_55[139],stage1_54[175]}
   );
   gpc615_5 gpc2083 (
      {stage0_54[343], stage0_54[344], stage0_54[345], stage0_54[346], stage0_54[347]},
      {stage0_55[141]},
      {stage0_56[121], stage0_56[122], stage0_56[123], stage0_56[124], stage0_56[125], stage0_56[126]},
      {stage1_58[20],stage1_57[41],stage1_56[77],stage1_55[140],stage1_54[176]}
   );
   gpc615_5 gpc2084 (
      {stage0_54[348], stage0_54[349], stage0_54[350], stage0_54[351], stage0_54[352]},
      {stage0_55[142]},
      {stage0_56[127], stage0_56[128], stage0_56[129], stage0_56[130], stage0_56[131], stage0_56[132]},
      {stage1_58[21],stage1_57[42],stage1_56[78],stage1_55[141],stage1_54[177]}
   );
   gpc615_5 gpc2085 (
      {stage0_54[353], stage0_54[354], stage0_54[355], stage0_54[356], stage0_54[357]},
      {stage0_55[143]},
      {stage0_56[133], stage0_56[134], stage0_56[135], stage0_56[136], stage0_56[137], stage0_56[138]},
      {stage1_58[22],stage1_57[43],stage1_56[79],stage1_55[142],stage1_54[178]}
   );
   gpc615_5 gpc2086 (
      {stage0_54[358], stage0_54[359], stage0_54[360], stage0_54[361], stage0_54[362]},
      {stage0_55[144]},
      {stage0_56[139], stage0_56[140], stage0_56[141], stage0_56[142], stage0_56[143], stage0_56[144]},
      {stage1_58[23],stage1_57[44],stage1_56[80],stage1_55[143],stage1_54[179]}
   );
   gpc615_5 gpc2087 (
      {stage0_54[363], stage0_54[364], stage0_54[365], stage0_54[366], stage0_54[367]},
      {stage0_55[145]},
      {stage0_56[145], stage0_56[146], stage0_56[147], stage0_56[148], stage0_56[149], stage0_56[150]},
      {stage1_58[24],stage1_57[45],stage1_56[81],stage1_55[144],stage1_54[180]}
   );
   gpc615_5 gpc2088 (
      {stage0_54[368], stage0_54[369], stage0_54[370], stage0_54[371], stage0_54[372]},
      {stage0_55[146]},
      {stage0_56[151], stage0_56[152], stage0_56[153], stage0_56[154], stage0_56[155], stage0_56[156]},
      {stage1_58[25],stage1_57[46],stage1_56[82],stage1_55[145],stage1_54[181]}
   );
   gpc615_5 gpc2089 (
      {stage0_54[373], stage0_54[374], stage0_54[375], stage0_54[376], stage0_54[377]},
      {stage0_55[147]},
      {stage0_56[157], stage0_56[158], stage0_56[159], stage0_56[160], stage0_56[161], stage0_56[162]},
      {stage1_58[26],stage1_57[47],stage1_56[83],stage1_55[146],stage1_54[182]}
   );
   gpc615_5 gpc2090 (
      {stage0_54[378], stage0_54[379], stage0_54[380], stage0_54[381], stage0_54[382]},
      {stage0_55[148]},
      {stage0_56[163], stage0_56[164], stage0_56[165], stage0_56[166], stage0_56[167], stage0_56[168]},
      {stage1_58[27],stage1_57[48],stage1_56[84],stage1_55[147],stage1_54[183]}
   );
   gpc615_5 gpc2091 (
      {stage0_54[383], stage0_54[384], stage0_54[385], stage0_54[386], stage0_54[387]},
      {stage0_55[149]},
      {stage0_56[169], stage0_56[170], stage0_56[171], stage0_56[172], stage0_56[173], stage0_56[174]},
      {stage1_58[28],stage1_57[49],stage1_56[85],stage1_55[148],stage1_54[184]}
   );
   gpc615_5 gpc2092 (
      {stage0_54[388], stage0_54[389], stage0_54[390], stage0_54[391], stage0_54[392]},
      {stage0_55[150]},
      {stage0_56[175], stage0_56[176], stage0_56[177], stage0_56[178], stage0_56[179], stage0_56[180]},
      {stage1_58[29],stage1_57[50],stage1_56[86],stage1_55[149],stage1_54[185]}
   );
   gpc615_5 gpc2093 (
      {stage0_54[393], stage0_54[394], stage0_54[395], stage0_54[396], stage0_54[397]},
      {stage0_55[151]},
      {stage0_56[181], stage0_56[182], stage0_56[183], stage0_56[184], stage0_56[185], stage0_56[186]},
      {stage1_58[30],stage1_57[51],stage1_56[87],stage1_55[150],stage1_54[186]}
   );
   gpc615_5 gpc2094 (
      {stage0_54[398], stage0_54[399], stage0_54[400], stage0_54[401], stage0_54[402]},
      {stage0_55[152]},
      {stage0_56[187], stage0_56[188], stage0_56[189], stage0_56[190], stage0_56[191], stage0_56[192]},
      {stage1_58[31],stage1_57[52],stage1_56[88],stage1_55[151],stage1_54[187]}
   );
   gpc615_5 gpc2095 (
      {stage0_54[403], stage0_54[404], stage0_54[405], stage0_54[406], stage0_54[407]},
      {stage0_55[153]},
      {stage0_56[193], stage0_56[194], stage0_56[195], stage0_56[196], stage0_56[197], stage0_56[198]},
      {stage1_58[32],stage1_57[53],stage1_56[89],stage1_55[152],stage1_54[188]}
   );
   gpc615_5 gpc2096 (
      {stage0_54[408], stage0_54[409], stage0_54[410], stage0_54[411], stage0_54[412]},
      {stage0_55[154]},
      {stage0_56[199], stage0_56[200], stage0_56[201], stage0_56[202], stage0_56[203], stage0_56[204]},
      {stage1_58[33],stage1_57[54],stage1_56[90],stage1_55[153],stage1_54[189]}
   );
   gpc615_5 gpc2097 (
      {stage0_54[413], stage0_54[414], stage0_54[415], stage0_54[416], stage0_54[417]},
      {stage0_55[155]},
      {stage0_56[205], stage0_56[206], stage0_56[207], stage0_56[208], stage0_56[209], stage0_56[210]},
      {stage1_58[34],stage1_57[55],stage1_56[91],stage1_55[154],stage1_54[190]}
   );
   gpc615_5 gpc2098 (
      {stage0_54[418], stage0_54[419], stage0_54[420], stage0_54[421], stage0_54[422]},
      {stage0_55[156]},
      {stage0_56[211], stage0_56[212], stage0_56[213], stage0_56[214], stage0_56[215], stage0_56[216]},
      {stage1_58[35],stage1_57[56],stage1_56[92],stage1_55[155],stage1_54[191]}
   );
   gpc615_5 gpc2099 (
      {stage0_54[423], stage0_54[424], stage0_54[425], stage0_54[426], stage0_54[427]},
      {stage0_55[157]},
      {stage0_56[217], stage0_56[218], stage0_56[219], stage0_56[220], stage0_56[221], stage0_56[222]},
      {stage1_58[36],stage1_57[57],stage1_56[93],stage1_55[156],stage1_54[192]}
   );
   gpc615_5 gpc2100 (
      {stage0_54[428], stage0_54[429], stage0_54[430], stage0_54[431], stage0_54[432]},
      {stage0_55[158]},
      {stage0_56[223], stage0_56[224], stage0_56[225], stage0_56[226], stage0_56[227], stage0_56[228]},
      {stage1_58[37],stage1_57[58],stage1_56[94],stage1_55[157],stage1_54[193]}
   );
   gpc615_5 gpc2101 (
      {stage0_54[433], stage0_54[434], stage0_54[435], stage0_54[436], stage0_54[437]},
      {stage0_55[159]},
      {stage0_56[229], stage0_56[230], stage0_56[231], stage0_56[232], stage0_56[233], stage0_56[234]},
      {stage1_58[38],stage1_57[59],stage1_56[95],stage1_55[158],stage1_54[194]}
   );
   gpc615_5 gpc2102 (
      {stage0_54[438], stage0_54[439], stage0_54[440], stage0_54[441], stage0_54[442]},
      {stage0_55[160]},
      {stage0_56[235], stage0_56[236], stage0_56[237], stage0_56[238], stage0_56[239], stage0_56[240]},
      {stage1_58[39],stage1_57[60],stage1_56[96],stage1_55[159],stage1_54[195]}
   );
   gpc615_5 gpc2103 (
      {stage0_54[443], stage0_54[444], stage0_54[445], stage0_54[446], stage0_54[447]},
      {stage0_55[161]},
      {stage0_56[241], stage0_56[242], stage0_56[243], stage0_56[244], stage0_56[245], stage0_56[246]},
      {stage1_58[40],stage1_57[61],stage1_56[97],stage1_55[160],stage1_54[196]}
   );
   gpc615_5 gpc2104 (
      {stage0_54[448], stage0_54[449], stage0_54[450], stage0_54[451], stage0_54[452]},
      {stage0_55[162]},
      {stage0_56[247], stage0_56[248], stage0_56[249], stage0_56[250], stage0_56[251], stage0_56[252]},
      {stage1_58[41],stage1_57[62],stage1_56[98],stage1_55[161],stage1_54[197]}
   );
   gpc606_5 gpc2105 (
      {stage0_55[163], stage0_55[164], stage0_55[165], stage0_55[166], stage0_55[167], stage0_55[168]},
      {stage0_57[0], stage0_57[1], stage0_57[2], stage0_57[3], stage0_57[4], stage0_57[5]},
      {stage1_59[0],stage1_58[42],stage1_57[63],stage1_56[99],stage1_55[162]}
   );
   gpc606_5 gpc2106 (
      {stage0_55[169], stage0_55[170], stage0_55[171], stage0_55[172], stage0_55[173], stage0_55[174]},
      {stage0_57[6], stage0_57[7], stage0_57[8], stage0_57[9], stage0_57[10], stage0_57[11]},
      {stage1_59[1],stage1_58[43],stage1_57[64],stage1_56[100],stage1_55[163]}
   );
   gpc606_5 gpc2107 (
      {stage0_55[175], stage0_55[176], stage0_55[177], stage0_55[178], stage0_55[179], stage0_55[180]},
      {stage0_57[12], stage0_57[13], stage0_57[14], stage0_57[15], stage0_57[16], stage0_57[17]},
      {stage1_59[2],stage1_58[44],stage1_57[65],stage1_56[101],stage1_55[164]}
   );
   gpc606_5 gpc2108 (
      {stage0_55[181], stage0_55[182], stage0_55[183], stage0_55[184], stage0_55[185], stage0_55[186]},
      {stage0_57[18], stage0_57[19], stage0_57[20], stage0_57[21], stage0_57[22], stage0_57[23]},
      {stage1_59[3],stage1_58[45],stage1_57[66],stage1_56[102],stage1_55[165]}
   );
   gpc606_5 gpc2109 (
      {stage0_55[187], stage0_55[188], stage0_55[189], stage0_55[190], stage0_55[191], stage0_55[192]},
      {stage0_57[24], stage0_57[25], stage0_57[26], stage0_57[27], stage0_57[28], stage0_57[29]},
      {stage1_59[4],stage1_58[46],stage1_57[67],stage1_56[103],stage1_55[166]}
   );
   gpc606_5 gpc2110 (
      {stage0_55[193], stage0_55[194], stage0_55[195], stage0_55[196], stage0_55[197], stage0_55[198]},
      {stage0_57[30], stage0_57[31], stage0_57[32], stage0_57[33], stage0_57[34], stage0_57[35]},
      {stage1_59[5],stage1_58[47],stage1_57[68],stage1_56[104],stage1_55[167]}
   );
   gpc606_5 gpc2111 (
      {stage0_55[199], stage0_55[200], stage0_55[201], stage0_55[202], stage0_55[203], stage0_55[204]},
      {stage0_57[36], stage0_57[37], stage0_57[38], stage0_57[39], stage0_57[40], stage0_57[41]},
      {stage1_59[6],stage1_58[48],stage1_57[69],stage1_56[105],stage1_55[168]}
   );
   gpc606_5 gpc2112 (
      {stage0_55[205], stage0_55[206], stage0_55[207], stage0_55[208], stage0_55[209], stage0_55[210]},
      {stage0_57[42], stage0_57[43], stage0_57[44], stage0_57[45], stage0_57[46], stage0_57[47]},
      {stage1_59[7],stage1_58[49],stage1_57[70],stage1_56[106],stage1_55[169]}
   );
   gpc606_5 gpc2113 (
      {stage0_55[211], stage0_55[212], stage0_55[213], stage0_55[214], stage0_55[215], stage0_55[216]},
      {stage0_57[48], stage0_57[49], stage0_57[50], stage0_57[51], stage0_57[52], stage0_57[53]},
      {stage1_59[8],stage1_58[50],stage1_57[71],stage1_56[107],stage1_55[170]}
   );
   gpc606_5 gpc2114 (
      {stage0_55[217], stage0_55[218], stage0_55[219], stage0_55[220], stage0_55[221], stage0_55[222]},
      {stage0_57[54], stage0_57[55], stage0_57[56], stage0_57[57], stage0_57[58], stage0_57[59]},
      {stage1_59[9],stage1_58[51],stage1_57[72],stage1_56[108],stage1_55[171]}
   );
   gpc606_5 gpc2115 (
      {stage0_55[223], stage0_55[224], stage0_55[225], stage0_55[226], stage0_55[227], stage0_55[228]},
      {stage0_57[60], stage0_57[61], stage0_57[62], stage0_57[63], stage0_57[64], stage0_57[65]},
      {stage1_59[10],stage1_58[52],stage1_57[73],stage1_56[109],stage1_55[172]}
   );
   gpc606_5 gpc2116 (
      {stage0_55[229], stage0_55[230], stage0_55[231], stage0_55[232], stage0_55[233], stage0_55[234]},
      {stage0_57[66], stage0_57[67], stage0_57[68], stage0_57[69], stage0_57[70], stage0_57[71]},
      {stage1_59[11],stage1_58[53],stage1_57[74],stage1_56[110],stage1_55[173]}
   );
   gpc606_5 gpc2117 (
      {stage0_55[235], stage0_55[236], stage0_55[237], stage0_55[238], stage0_55[239], stage0_55[240]},
      {stage0_57[72], stage0_57[73], stage0_57[74], stage0_57[75], stage0_57[76], stage0_57[77]},
      {stage1_59[12],stage1_58[54],stage1_57[75],stage1_56[111],stage1_55[174]}
   );
   gpc606_5 gpc2118 (
      {stage0_55[241], stage0_55[242], stage0_55[243], stage0_55[244], stage0_55[245], stage0_55[246]},
      {stage0_57[78], stage0_57[79], stage0_57[80], stage0_57[81], stage0_57[82], stage0_57[83]},
      {stage1_59[13],stage1_58[55],stage1_57[76],stage1_56[112],stage1_55[175]}
   );
   gpc606_5 gpc2119 (
      {stage0_55[247], stage0_55[248], stage0_55[249], stage0_55[250], stage0_55[251], stage0_55[252]},
      {stage0_57[84], stage0_57[85], stage0_57[86], stage0_57[87], stage0_57[88], stage0_57[89]},
      {stage1_59[14],stage1_58[56],stage1_57[77],stage1_56[113],stage1_55[176]}
   );
   gpc606_5 gpc2120 (
      {stage0_55[253], stage0_55[254], stage0_55[255], stage0_55[256], stage0_55[257], stage0_55[258]},
      {stage0_57[90], stage0_57[91], stage0_57[92], stage0_57[93], stage0_57[94], stage0_57[95]},
      {stage1_59[15],stage1_58[57],stage1_57[78],stage1_56[114],stage1_55[177]}
   );
   gpc606_5 gpc2121 (
      {stage0_55[259], stage0_55[260], stage0_55[261], stage0_55[262], stage0_55[263], stage0_55[264]},
      {stage0_57[96], stage0_57[97], stage0_57[98], stage0_57[99], stage0_57[100], stage0_57[101]},
      {stage1_59[16],stage1_58[58],stage1_57[79],stage1_56[115],stage1_55[178]}
   );
   gpc606_5 gpc2122 (
      {stage0_55[265], stage0_55[266], stage0_55[267], stage0_55[268], stage0_55[269], stage0_55[270]},
      {stage0_57[102], stage0_57[103], stage0_57[104], stage0_57[105], stage0_57[106], stage0_57[107]},
      {stage1_59[17],stage1_58[59],stage1_57[80],stage1_56[116],stage1_55[179]}
   );
   gpc606_5 gpc2123 (
      {stage0_55[271], stage0_55[272], stage0_55[273], stage0_55[274], stage0_55[275], stage0_55[276]},
      {stage0_57[108], stage0_57[109], stage0_57[110], stage0_57[111], stage0_57[112], stage0_57[113]},
      {stage1_59[18],stage1_58[60],stage1_57[81],stage1_56[117],stage1_55[180]}
   );
   gpc606_5 gpc2124 (
      {stage0_55[277], stage0_55[278], stage0_55[279], stage0_55[280], stage0_55[281], stage0_55[282]},
      {stage0_57[114], stage0_57[115], stage0_57[116], stage0_57[117], stage0_57[118], stage0_57[119]},
      {stage1_59[19],stage1_58[61],stage1_57[82],stage1_56[118],stage1_55[181]}
   );
   gpc606_5 gpc2125 (
      {stage0_55[283], stage0_55[284], stage0_55[285], stage0_55[286], stage0_55[287], stage0_55[288]},
      {stage0_57[120], stage0_57[121], stage0_57[122], stage0_57[123], stage0_57[124], stage0_57[125]},
      {stage1_59[20],stage1_58[62],stage1_57[83],stage1_56[119],stage1_55[182]}
   );
   gpc606_5 gpc2126 (
      {stage0_55[289], stage0_55[290], stage0_55[291], stage0_55[292], stage0_55[293], stage0_55[294]},
      {stage0_57[126], stage0_57[127], stage0_57[128], stage0_57[129], stage0_57[130], stage0_57[131]},
      {stage1_59[21],stage1_58[63],stage1_57[84],stage1_56[120],stage1_55[183]}
   );
   gpc606_5 gpc2127 (
      {stage0_55[295], stage0_55[296], stage0_55[297], stage0_55[298], stage0_55[299], stage0_55[300]},
      {stage0_57[132], stage0_57[133], stage0_57[134], stage0_57[135], stage0_57[136], stage0_57[137]},
      {stage1_59[22],stage1_58[64],stage1_57[85],stage1_56[121],stage1_55[184]}
   );
   gpc606_5 gpc2128 (
      {stage0_55[301], stage0_55[302], stage0_55[303], stage0_55[304], stage0_55[305], stage0_55[306]},
      {stage0_57[138], stage0_57[139], stage0_57[140], stage0_57[141], stage0_57[142], stage0_57[143]},
      {stage1_59[23],stage1_58[65],stage1_57[86],stage1_56[122],stage1_55[185]}
   );
   gpc606_5 gpc2129 (
      {stage0_55[307], stage0_55[308], stage0_55[309], stage0_55[310], stage0_55[311], stage0_55[312]},
      {stage0_57[144], stage0_57[145], stage0_57[146], stage0_57[147], stage0_57[148], stage0_57[149]},
      {stage1_59[24],stage1_58[66],stage1_57[87],stage1_56[123],stage1_55[186]}
   );
   gpc606_5 gpc2130 (
      {stage0_55[313], stage0_55[314], stage0_55[315], stage0_55[316], stage0_55[317], stage0_55[318]},
      {stage0_57[150], stage0_57[151], stage0_57[152], stage0_57[153], stage0_57[154], stage0_57[155]},
      {stage1_59[25],stage1_58[67],stage1_57[88],stage1_56[124],stage1_55[187]}
   );
   gpc606_5 gpc2131 (
      {stage0_55[319], stage0_55[320], stage0_55[321], stage0_55[322], stage0_55[323], stage0_55[324]},
      {stage0_57[156], stage0_57[157], stage0_57[158], stage0_57[159], stage0_57[160], stage0_57[161]},
      {stage1_59[26],stage1_58[68],stage1_57[89],stage1_56[125],stage1_55[188]}
   );
   gpc606_5 gpc2132 (
      {stage0_55[325], stage0_55[326], stage0_55[327], stage0_55[328], stage0_55[329], stage0_55[330]},
      {stage0_57[162], stage0_57[163], stage0_57[164], stage0_57[165], stage0_57[166], stage0_57[167]},
      {stage1_59[27],stage1_58[69],stage1_57[90],stage1_56[126],stage1_55[189]}
   );
   gpc606_5 gpc2133 (
      {stage0_55[331], stage0_55[332], stage0_55[333], stage0_55[334], stage0_55[335], stage0_55[336]},
      {stage0_57[168], stage0_57[169], stage0_57[170], stage0_57[171], stage0_57[172], stage0_57[173]},
      {stage1_59[28],stage1_58[70],stage1_57[91],stage1_56[127],stage1_55[190]}
   );
   gpc606_5 gpc2134 (
      {stage0_55[337], stage0_55[338], stage0_55[339], stage0_55[340], stage0_55[341], stage0_55[342]},
      {stage0_57[174], stage0_57[175], stage0_57[176], stage0_57[177], stage0_57[178], stage0_57[179]},
      {stage1_59[29],stage1_58[71],stage1_57[92],stage1_56[128],stage1_55[191]}
   );
   gpc606_5 gpc2135 (
      {stage0_55[343], stage0_55[344], stage0_55[345], stage0_55[346], stage0_55[347], stage0_55[348]},
      {stage0_57[180], stage0_57[181], stage0_57[182], stage0_57[183], stage0_57[184], stage0_57[185]},
      {stage1_59[30],stage1_58[72],stage1_57[93],stage1_56[129],stage1_55[192]}
   );
   gpc606_5 gpc2136 (
      {stage0_55[349], stage0_55[350], stage0_55[351], stage0_55[352], stage0_55[353], stage0_55[354]},
      {stage0_57[186], stage0_57[187], stage0_57[188], stage0_57[189], stage0_57[190], stage0_57[191]},
      {stage1_59[31],stage1_58[73],stage1_57[94],stage1_56[130],stage1_55[193]}
   );
   gpc606_5 gpc2137 (
      {stage0_55[355], stage0_55[356], stage0_55[357], stage0_55[358], stage0_55[359], stage0_55[360]},
      {stage0_57[192], stage0_57[193], stage0_57[194], stage0_57[195], stage0_57[196], stage0_57[197]},
      {stage1_59[32],stage1_58[74],stage1_57[95],stage1_56[131],stage1_55[194]}
   );
   gpc606_5 gpc2138 (
      {stage0_55[361], stage0_55[362], stage0_55[363], stage0_55[364], stage0_55[365], stage0_55[366]},
      {stage0_57[198], stage0_57[199], stage0_57[200], stage0_57[201], stage0_57[202], stage0_57[203]},
      {stage1_59[33],stage1_58[75],stage1_57[96],stage1_56[132],stage1_55[195]}
   );
   gpc606_5 gpc2139 (
      {stage0_55[367], stage0_55[368], stage0_55[369], stage0_55[370], stage0_55[371], stage0_55[372]},
      {stage0_57[204], stage0_57[205], stage0_57[206], stage0_57[207], stage0_57[208], stage0_57[209]},
      {stage1_59[34],stage1_58[76],stage1_57[97],stage1_56[133],stage1_55[196]}
   );
   gpc606_5 gpc2140 (
      {stage0_55[373], stage0_55[374], stage0_55[375], stage0_55[376], stage0_55[377], stage0_55[378]},
      {stage0_57[210], stage0_57[211], stage0_57[212], stage0_57[213], stage0_57[214], stage0_57[215]},
      {stage1_59[35],stage1_58[77],stage1_57[98],stage1_56[134],stage1_55[197]}
   );
   gpc606_5 gpc2141 (
      {stage0_55[379], stage0_55[380], stage0_55[381], stage0_55[382], stage0_55[383], stage0_55[384]},
      {stage0_57[216], stage0_57[217], stage0_57[218], stage0_57[219], stage0_57[220], stage0_57[221]},
      {stage1_59[36],stage1_58[78],stage1_57[99],stage1_56[135],stage1_55[198]}
   );
   gpc606_5 gpc2142 (
      {stage0_55[385], stage0_55[386], stage0_55[387], stage0_55[388], stage0_55[389], stage0_55[390]},
      {stage0_57[222], stage0_57[223], stage0_57[224], stage0_57[225], stage0_57[226], stage0_57[227]},
      {stage1_59[37],stage1_58[79],stage1_57[100],stage1_56[136],stage1_55[199]}
   );
   gpc606_5 gpc2143 (
      {stage0_55[391], stage0_55[392], stage0_55[393], stage0_55[394], stage0_55[395], stage0_55[396]},
      {stage0_57[228], stage0_57[229], stage0_57[230], stage0_57[231], stage0_57[232], stage0_57[233]},
      {stage1_59[38],stage1_58[80],stage1_57[101],stage1_56[137],stage1_55[200]}
   );
   gpc606_5 gpc2144 (
      {stage0_55[397], stage0_55[398], stage0_55[399], stage0_55[400], stage0_55[401], stage0_55[402]},
      {stage0_57[234], stage0_57[235], stage0_57[236], stage0_57[237], stage0_57[238], stage0_57[239]},
      {stage1_59[39],stage1_58[81],stage1_57[102],stage1_56[138],stage1_55[201]}
   );
   gpc606_5 gpc2145 (
      {stage0_55[403], stage0_55[404], stage0_55[405], stage0_55[406], stage0_55[407], stage0_55[408]},
      {stage0_57[240], stage0_57[241], stage0_57[242], stage0_57[243], stage0_57[244], stage0_57[245]},
      {stage1_59[40],stage1_58[82],stage1_57[103],stage1_56[139],stage1_55[202]}
   );
   gpc606_5 gpc2146 (
      {stage0_55[409], stage0_55[410], stage0_55[411], stage0_55[412], stage0_55[413], stage0_55[414]},
      {stage0_57[246], stage0_57[247], stage0_57[248], stage0_57[249], stage0_57[250], stage0_57[251]},
      {stage1_59[41],stage1_58[83],stage1_57[104],stage1_56[140],stage1_55[203]}
   );
   gpc615_5 gpc2147 (
      {stage0_55[415], stage0_55[416], stage0_55[417], stage0_55[418], stage0_55[419]},
      {stage0_56[253]},
      {stage0_57[252], stage0_57[253], stage0_57[254], stage0_57[255], stage0_57[256], stage0_57[257]},
      {stage1_59[42],stage1_58[84],stage1_57[105],stage1_56[141],stage1_55[204]}
   );
   gpc615_5 gpc2148 (
      {stage0_55[420], stage0_55[421], stage0_55[422], stage0_55[423], stage0_55[424]},
      {stage0_56[254]},
      {stage0_57[258], stage0_57[259], stage0_57[260], stage0_57[261], stage0_57[262], stage0_57[263]},
      {stage1_59[43],stage1_58[85],stage1_57[106],stage1_56[142],stage1_55[205]}
   );
   gpc606_5 gpc2149 (
      {stage0_56[255], stage0_56[256], stage0_56[257], stage0_56[258], stage0_56[259], stage0_56[260]},
      {stage0_58[0], stage0_58[1], stage0_58[2], stage0_58[3], stage0_58[4], stage0_58[5]},
      {stage1_60[0],stage1_59[44],stage1_58[86],stage1_57[107],stage1_56[143]}
   );
   gpc606_5 gpc2150 (
      {stage0_56[261], stage0_56[262], stage0_56[263], stage0_56[264], stage0_56[265], stage0_56[266]},
      {stage0_58[6], stage0_58[7], stage0_58[8], stage0_58[9], stage0_58[10], stage0_58[11]},
      {stage1_60[1],stage1_59[45],stage1_58[87],stage1_57[108],stage1_56[144]}
   );
   gpc606_5 gpc2151 (
      {stage0_56[267], stage0_56[268], stage0_56[269], stage0_56[270], stage0_56[271], stage0_56[272]},
      {stage0_58[12], stage0_58[13], stage0_58[14], stage0_58[15], stage0_58[16], stage0_58[17]},
      {stage1_60[2],stage1_59[46],stage1_58[88],stage1_57[109],stage1_56[145]}
   );
   gpc606_5 gpc2152 (
      {stage0_56[273], stage0_56[274], stage0_56[275], stage0_56[276], stage0_56[277], stage0_56[278]},
      {stage0_58[18], stage0_58[19], stage0_58[20], stage0_58[21], stage0_58[22], stage0_58[23]},
      {stage1_60[3],stage1_59[47],stage1_58[89],stage1_57[110],stage1_56[146]}
   );
   gpc606_5 gpc2153 (
      {stage0_56[279], stage0_56[280], stage0_56[281], stage0_56[282], stage0_56[283], stage0_56[284]},
      {stage0_58[24], stage0_58[25], stage0_58[26], stage0_58[27], stage0_58[28], stage0_58[29]},
      {stage1_60[4],stage1_59[48],stage1_58[90],stage1_57[111],stage1_56[147]}
   );
   gpc606_5 gpc2154 (
      {stage0_56[285], stage0_56[286], stage0_56[287], stage0_56[288], stage0_56[289], stage0_56[290]},
      {stage0_58[30], stage0_58[31], stage0_58[32], stage0_58[33], stage0_58[34], stage0_58[35]},
      {stage1_60[5],stage1_59[49],stage1_58[91],stage1_57[112],stage1_56[148]}
   );
   gpc606_5 gpc2155 (
      {stage0_56[291], stage0_56[292], stage0_56[293], stage0_56[294], stage0_56[295], stage0_56[296]},
      {stage0_58[36], stage0_58[37], stage0_58[38], stage0_58[39], stage0_58[40], stage0_58[41]},
      {stage1_60[6],stage1_59[50],stage1_58[92],stage1_57[113],stage1_56[149]}
   );
   gpc606_5 gpc2156 (
      {stage0_56[297], stage0_56[298], stage0_56[299], stage0_56[300], stage0_56[301], stage0_56[302]},
      {stage0_58[42], stage0_58[43], stage0_58[44], stage0_58[45], stage0_58[46], stage0_58[47]},
      {stage1_60[7],stage1_59[51],stage1_58[93],stage1_57[114],stage1_56[150]}
   );
   gpc606_5 gpc2157 (
      {stage0_56[303], stage0_56[304], stage0_56[305], stage0_56[306], stage0_56[307], stage0_56[308]},
      {stage0_58[48], stage0_58[49], stage0_58[50], stage0_58[51], stage0_58[52], stage0_58[53]},
      {stage1_60[8],stage1_59[52],stage1_58[94],stage1_57[115],stage1_56[151]}
   );
   gpc606_5 gpc2158 (
      {stage0_56[309], stage0_56[310], stage0_56[311], stage0_56[312], stage0_56[313], stage0_56[314]},
      {stage0_58[54], stage0_58[55], stage0_58[56], stage0_58[57], stage0_58[58], stage0_58[59]},
      {stage1_60[9],stage1_59[53],stage1_58[95],stage1_57[116],stage1_56[152]}
   );
   gpc606_5 gpc2159 (
      {stage0_56[315], stage0_56[316], stage0_56[317], stage0_56[318], stage0_56[319], stage0_56[320]},
      {stage0_58[60], stage0_58[61], stage0_58[62], stage0_58[63], stage0_58[64], stage0_58[65]},
      {stage1_60[10],stage1_59[54],stage1_58[96],stage1_57[117],stage1_56[153]}
   );
   gpc615_5 gpc2160 (
      {stage0_56[321], stage0_56[322], stage0_56[323], stage0_56[324], stage0_56[325]},
      {stage0_57[264]},
      {stage0_58[66], stage0_58[67], stage0_58[68], stage0_58[69], stage0_58[70], stage0_58[71]},
      {stage1_60[11],stage1_59[55],stage1_58[97],stage1_57[118],stage1_56[154]}
   );
   gpc615_5 gpc2161 (
      {stage0_56[326], stage0_56[327], stage0_56[328], stage0_56[329], stage0_56[330]},
      {stage0_57[265]},
      {stage0_58[72], stage0_58[73], stage0_58[74], stage0_58[75], stage0_58[76], stage0_58[77]},
      {stage1_60[12],stage1_59[56],stage1_58[98],stage1_57[119],stage1_56[155]}
   );
   gpc615_5 gpc2162 (
      {stage0_56[331], stage0_56[332], stage0_56[333], stage0_56[334], stage0_56[335]},
      {stage0_57[266]},
      {stage0_58[78], stage0_58[79], stage0_58[80], stage0_58[81], stage0_58[82], stage0_58[83]},
      {stage1_60[13],stage1_59[57],stage1_58[99],stage1_57[120],stage1_56[156]}
   );
   gpc615_5 gpc2163 (
      {stage0_56[336], stage0_56[337], stage0_56[338], stage0_56[339], stage0_56[340]},
      {stage0_57[267]},
      {stage0_58[84], stage0_58[85], stage0_58[86], stage0_58[87], stage0_58[88], stage0_58[89]},
      {stage1_60[14],stage1_59[58],stage1_58[100],stage1_57[121],stage1_56[157]}
   );
   gpc615_5 gpc2164 (
      {stage0_56[341], stage0_56[342], stage0_56[343], stage0_56[344], stage0_56[345]},
      {stage0_57[268]},
      {stage0_58[90], stage0_58[91], stage0_58[92], stage0_58[93], stage0_58[94], stage0_58[95]},
      {stage1_60[15],stage1_59[59],stage1_58[101],stage1_57[122],stage1_56[158]}
   );
   gpc615_5 gpc2165 (
      {stage0_56[346], stage0_56[347], stage0_56[348], stage0_56[349], stage0_56[350]},
      {stage0_57[269]},
      {stage0_58[96], stage0_58[97], stage0_58[98], stage0_58[99], stage0_58[100], stage0_58[101]},
      {stage1_60[16],stage1_59[60],stage1_58[102],stage1_57[123],stage1_56[159]}
   );
   gpc615_5 gpc2166 (
      {stage0_56[351], stage0_56[352], stage0_56[353], stage0_56[354], stage0_56[355]},
      {stage0_57[270]},
      {stage0_58[102], stage0_58[103], stage0_58[104], stage0_58[105], stage0_58[106], stage0_58[107]},
      {stage1_60[17],stage1_59[61],stage1_58[103],stage1_57[124],stage1_56[160]}
   );
   gpc615_5 gpc2167 (
      {stage0_56[356], stage0_56[357], stage0_56[358], stage0_56[359], stage0_56[360]},
      {stage0_57[271]},
      {stage0_58[108], stage0_58[109], stage0_58[110], stage0_58[111], stage0_58[112], stage0_58[113]},
      {stage1_60[18],stage1_59[62],stage1_58[104],stage1_57[125],stage1_56[161]}
   );
   gpc615_5 gpc2168 (
      {stage0_56[361], stage0_56[362], stage0_56[363], stage0_56[364], stage0_56[365]},
      {stage0_57[272]},
      {stage0_58[114], stage0_58[115], stage0_58[116], stage0_58[117], stage0_58[118], stage0_58[119]},
      {stage1_60[19],stage1_59[63],stage1_58[105],stage1_57[126],stage1_56[162]}
   );
   gpc615_5 gpc2169 (
      {stage0_56[366], stage0_56[367], stage0_56[368], stage0_56[369], stage0_56[370]},
      {stage0_57[273]},
      {stage0_58[120], stage0_58[121], stage0_58[122], stage0_58[123], stage0_58[124], stage0_58[125]},
      {stage1_60[20],stage1_59[64],stage1_58[106],stage1_57[127],stage1_56[163]}
   );
   gpc615_5 gpc2170 (
      {stage0_56[371], stage0_56[372], stage0_56[373], stage0_56[374], stage0_56[375]},
      {stage0_57[274]},
      {stage0_58[126], stage0_58[127], stage0_58[128], stage0_58[129], stage0_58[130], stage0_58[131]},
      {stage1_60[21],stage1_59[65],stage1_58[107],stage1_57[128],stage1_56[164]}
   );
   gpc615_5 gpc2171 (
      {stage0_56[376], stage0_56[377], stage0_56[378], stage0_56[379], stage0_56[380]},
      {stage0_57[275]},
      {stage0_58[132], stage0_58[133], stage0_58[134], stage0_58[135], stage0_58[136], stage0_58[137]},
      {stage1_60[22],stage1_59[66],stage1_58[108],stage1_57[129],stage1_56[165]}
   );
   gpc615_5 gpc2172 (
      {stage0_56[381], stage0_56[382], stage0_56[383], stage0_56[384], stage0_56[385]},
      {stage0_57[276]},
      {stage0_58[138], stage0_58[139], stage0_58[140], stage0_58[141], stage0_58[142], stage0_58[143]},
      {stage1_60[23],stage1_59[67],stage1_58[109],stage1_57[130],stage1_56[166]}
   );
   gpc615_5 gpc2173 (
      {stage0_56[386], stage0_56[387], stage0_56[388], stage0_56[389], stage0_56[390]},
      {stage0_57[277]},
      {stage0_58[144], stage0_58[145], stage0_58[146], stage0_58[147], stage0_58[148], stage0_58[149]},
      {stage1_60[24],stage1_59[68],stage1_58[110],stage1_57[131],stage1_56[167]}
   );
   gpc615_5 gpc2174 (
      {stage0_56[391], stage0_56[392], stage0_56[393], stage0_56[394], stage0_56[395]},
      {stage0_57[278]},
      {stage0_58[150], stage0_58[151], stage0_58[152], stage0_58[153], stage0_58[154], stage0_58[155]},
      {stage1_60[25],stage1_59[69],stage1_58[111],stage1_57[132],stage1_56[168]}
   );
   gpc615_5 gpc2175 (
      {stage0_56[396], stage0_56[397], stage0_56[398], stage0_56[399], stage0_56[400]},
      {stage0_57[279]},
      {stage0_58[156], stage0_58[157], stage0_58[158], stage0_58[159], stage0_58[160], stage0_58[161]},
      {stage1_60[26],stage1_59[70],stage1_58[112],stage1_57[133],stage1_56[169]}
   );
   gpc615_5 gpc2176 (
      {stage0_56[401], stage0_56[402], stage0_56[403], stage0_56[404], stage0_56[405]},
      {stage0_57[280]},
      {stage0_58[162], stage0_58[163], stage0_58[164], stage0_58[165], stage0_58[166], stage0_58[167]},
      {stage1_60[27],stage1_59[71],stage1_58[113],stage1_57[134],stage1_56[170]}
   );
   gpc615_5 gpc2177 (
      {stage0_56[406], stage0_56[407], stage0_56[408], stage0_56[409], stage0_56[410]},
      {stage0_57[281]},
      {stage0_58[168], stage0_58[169], stage0_58[170], stage0_58[171], stage0_58[172], stage0_58[173]},
      {stage1_60[28],stage1_59[72],stage1_58[114],stage1_57[135],stage1_56[171]}
   );
   gpc615_5 gpc2178 (
      {stage0_56[411], stage0_56[412], stage0_56[413], stage0_56[414], stage0_56[415]},
      {stage0_57[282]},
      {stage0_58[174], stage0_58[175], stage0_58[176], stage0_58[177], stage0_58[178], stage0_58[179]},
      {stage1_60[29],stage1_59[73],stage1_58[115],stage1_57[136],stage1_56[172]}
   );
   gpc615_5 gpc2179 (
      {stage0_56[416], stage0_56[417], stage0_56[418], stage0_56[419], stage0_56[420]},
      {stage0_57[283]},
      {stage0_58[180], stage0_58[181], stage0_58[182], stage0_58[183], stage0_58[184], stage0_58[185]},
      {stage1_60[30],stage1_59[74],stage1_58[116],stage1_57[137],stage1_56[173]}
   );
   gpc615_5 gpc2180 (
      {stage0_56[421], stage0_56[422], stage0_56[423], stage0_56[424], stage0_56[425]},
      {stage0_57[284]},
      {stage0_58[186], stage0_58[187], stage0_58[188], stage0_58[189], stage0_58[190], stage0_58[191]},
      {stage1_60[31],stage1_59[75],stage1_58[117],stage1_57[138],stage1_56[174]}
   );
   gpc615_5 gpc2181 (
      {stage0_56[426], stage0_56[427], stage0_56[428], stage0_56[429], stage0_56[430]},
      {stage0_57[285]},
      {stage0_58[192], stage0_58[193], stage0_58[194], stage0_58[195], stage0_58[196], stage0_58[197]},
      {stage1_60[32],stage1_59[76],stage1_58[118],stage1_57[139],stage1_56[175]}
   );
   gpc615_5 gpc2182 (
      {stage0_56[431], stage0_56[432], stage0_56[433], stage0_56[434], stage0_56[435]},
      {stage0_57[286]},
      {stage0_58[198], stage0_58[199], stage0_58[200], stage0_58[201], stage0_58[202], stage0_58[203]},
      {stage1_60[33],stage1_59[77],stage1_58[119],stage1_57[140],stage1_56[176]}
   );
   gpc615_5 gpc2183 (
      {stage0_56[436], stage0_56[437], stage0_56[438], stage0_56[439], stage0_56[440]},
      {stage0_57[287]},
      {stage0_58[204], stage0_58[205], stage0_58[206], stage0_58[207], stage0_58[208], stage0_58[209]},
      {stage1_60[34],stage1_59[78],stage1_58[120],stage1_57[141],stage1_56[177]}
   );
   gpc615_5 gpc2184 (
      {stage0_56[441], stage0_56[442], stage0_56[443], stage0_56[444], stage0_56[445]},
      {stage0_57[288]},
      {stage0_58[210], stage0_58[211], stage0_58[212], stage0_58[213], stage0_58[214], stage0_58[215]},
      {stage1_60[35],stage1_59[79],stage1_58[121],stage1_57[142],stage1_56[178]}
   );
   gpc615_5 gpc2185 (
      {stage0_56[446], stage0_56[447], stage0_56[448], stage0_56[449], stage0_56[450]},
      {stage0_57[289]},
      {stage0_58[216], stage0_58[217], stage0_58[218], stage0_58[219], stage0_58[220], stage0_58[221]},
      {stage1_60[36],stage1_59[80],stage1_58[122],stage1_57[143],stage1_56[179]}
   );
   gpc615_5 gpc2186 (
      {stage0_56[451], stage0_56[452], stage0_56[453], stage0_56[454], stage0_56[455]},
      {stage0_57[290]},
      {stage0_58[222], stage0_58[223], stage0_58[224], stage0_58[225], stage0_58[226], stage0_58[227]},
      {stage1_60[37],stage1_59[81],stage1_58[123],stage1_57[144],stage1_56[180]}
   );
   gpc615_5 gpc2187 (
      {stage0_56[456], stage0_56[457], stage0_56[458], stage0_56[459], stage0_56[460]},
      {stage0_57[291]},
      {stage0_58[228], stage0_58[229], stage0_58[230], stage0_58[231], stage0_58[232], stage0_58[233]},
      {stage1_60[38],stage1_59[82],stage1_58[124],stage1_57[145],stage1_56[181]}
   );
   gpc615_5 gpc2188 (
      {stage0_56[461], stage0_56[462], stage0_56[463], stage0_56[464], stage0_56[465]},
      {stage0_57[292]},
      {stage0_58[234], stage0_58[235], stage0_58[236], stage0_58[237], stage0_58[238], stage0_58[239]},
      {stage1_60[39],stage1_59[83],stage1_58[125],stage1_57[146],stage1_56[182]}
   );
   gpc615_5 gpc2189 (
      {stage0_56[466], stage0_56[467], stage0_56[468], stage0_56[469], stage0_56[470]},
      {stage0_57[293]},
      {stage0_58[240], stage0_58[241], stage0_58[242], stage0_58[243], stage0_58[244], stage0_58[245]},
      {stage1_60[40],stage1_59[84],stage1_58[126],stage1_57[147],stage1_56[183]}
   );
   gpc615_5 gpc2190 (
      {stage0_56[471], stage0_56[472], stage0_56[473], stage0_56[474], stage0_56[475]},
      {stage0_57[294]},
      {stage0_58[246], stage0_58[247], stage0_58[248], stage0_58[249], stage0_58[250], stage0_58[251]},
      {stage1_60[41],stage1_59[85],stage1_58[127],stage1_57[148],stage1_56[184]}
   );
   gpc615_5 gpc2191 (
      {stage0_56[476], stage0_56[477], stage0_56[478], stage0_56[479], stage0_56[480]},
      {stage0_57[295]},
      {stage0_58[252], stage0_58[253], stage0_58[254], stage0_58[255], stage0_58[256], stage0_58[257]},
      {stage1_60[42],stage1_59[86],stage1_58[128],stage1_57[149],stage1_56[185]}
   );
   gpc615_5 gpc2192 (
      {stage0_56[481], stage0_56[482], stage0_56[483], stage0_56[484], stage0_56[485]},
      {stage0_57[296]},
      {stage0_58[258], stage0_58[259], stage0_58[260], stage0_58[261], stage0_58[262], stage0_58[263]},
      {stage1_60[43],stage1_59[87],stage1_58[129],stage1_57[150],stage1_56[186]}
   );
   gpc615_5 gpc2193 (
      {stage0_57[297], stage0_57[298], stage0_57[299], stage0_57[300], stage0_57[301]},
      {stage0_58[264]},
      {stage0_59[0], stage0_59[1], stage0_59[2], stage0_59[3], stage0_59[4], stage0_59[5]},
      {stage1_61[0],stage1_60[44],stage1_59[88],stage1_58[130],stage1_57[151]}
   );
   gpc615_5 gpc2194 (
      {stage0_57[302], stage0_57[303], stage0_57[304], stage0_57[305], stage0_57[306]},
      {stage0_58[265]},
      {stage0_59[6], stage0_59[7], stage0_59[8], stage0_59[9], stage0_59[10], stage0_59[11]},
      {stage1_61[1],stage1_60[45],stage1_59[89],stage1_58[131],stage1_57[152]}
   );
   gpc615_5 gpc2195 (
      {stage0_57[307], stage0_57[308], stage0_57[309], stage0_57[310], stage0_57[311]},
      {stage0_58[266]},
      {stage0_59[12], stage0_59[13], stage0_59[14], stage0_59[15], stage0_59[16], stage0_59[17]},
      {stage1_61[2],stage1_60[46],stage1_59[90],stage1_58[132],stage1_57[153]}
   );
   gpc615_5 gpc2196 (
      {stage0_57[312], stage0_57[313], stage0_57[314], stage0_57[315], stage0_57[316]},
      {stage0_58[267]},
      {stage0_59[18], stage0_59[19], stage0_59[20], stage0_59[21], stage0_59[22], stage0_59[23]},
      {stage1_61[3],stage1_60[47],stage1_59[91],stage1_58[133],stage1_57[154]}
   );
   gpc615_5 gpc2197 (
      {stage0_57[317], stage0_57[318], stage0_57[319], stage0_57[320], stage0_57[321]},
      {stage0_58[268]},
      {stage0_59[24], stage0_59[25], stage0_59[26], stage0_59[27], stage0_59[28], stage0_59[29]},
      {stage1_61[4],stage1_60[48],stage1_59[92],stage1_58[134],stage1_57[155]}
   );
   gpc615_5 gpc2198 (
      {stage0_57[322], stage0_57[323], stage0_57[324], stage0_57[325], stage0_57[326]},
      {stage0_58[269]},
      {stage0_59[30], stage0_59[31], stage0_59[32], stage0_59[33], stage0_59[34], stage0_59[35]},
      {stage1_61[5],stage1_60[49],stage1_59[93],stage1_58[135],stage1_57[156]}
   );
   gpc615_5 gpc2199 (
      {stage0_57[327], stage0_57[328], stage0_57[329], stage0_57[330], stage0_57[331]},
      {stage0_58[270]},
      {stage0_59[36], stage0_59[37], stage0_59[38], stage0_59[39], stage0_59[40], stage0_59[41]},
      {stage1_61[6],stage1_60[50],stage1_59[94],stage1_58[136],stage1_57[157]}
   );
   gpc615_5 gpc2200 (
      {stage0_57[332], stage0_57[333], stage0_57[334], stage0_57[335], stage0_57[336]},
      {stage0_58[271]},
      {stage0_59[42], stage0_59[43], stage0_59[44], stage0_59[45], stage0_59[46], stage0_59[47]},
      {stage1_61[7],stage1_60[51],stage1_59[95],stage1_58[137],stage1_57[158]}
   );
   gpc615_5 gpc2201 (
      {stage0_57[337], stage0_57[338], stage0_57[339], stage0_57[340], stage0_57[341]},
      {stage0_58[272]},
      {stage0_59[48], stage0_59[49], stage0_59[50], stage0_59[51], stage0_59[52], stage0_59[53]},
      {stage1_61[8],stage1_60[52],stage1_59[96],stage1_58[138],stage1_57[159]}
   );
   gpc615_5 gpc2202 (
      {stage0_57[342], stage0_57[343], stage0_57[344], stage0_57[345], stage0_57[346]},
      {stage0_58[273]},
      {stage0_59[54], stage0_59[55], stage0_59[56], stage0_59[57], stage0_59[58], stage0_59[59]},
      {stage1_61[9],stage1_60[53],stage1_59[97],stage1_58[139],stage1_57[160]}
   );
   gpc615_5 gpc2203 (
      {stage0_57[347], stage0_57[348], stage0_57[349], stage0_57[350], stage0_57[351]},
      {stage0_58[274]},
      {stage0_59[60], stage0_59[61], stage0_59[62], stage0_59[63], stage0_59[64], stage0_59[65]},
      {stage1_61[10],stage1_60[54],stage1_59[98],stage1_58[140],stage1_57[161]}
   );
   gpc615_5 gpc2204 (
      {stage0_57[352], stage0_57[353], stage0_57[354], stage0_57[355], stage0_57[356]},
      {stage0_58[275]},
      {stage0_59[66], stage0_59[67], stage0_59[68], stage0_59[69], stage0_59[70], stage0_59[71]},
      {stage1_61[11],stage1_60[55],stage1_59[99],stage1_58[141],stage1_57[162]}
   );
   gpc615_5 gpc2205 (
      {stage0_57[357], stage0_57[358], stage0_57[359], stage0_57[360], stage0_57[361]},
      {stage0_58[276]},
      {stage0_59[72], stage0_59[73], stage0_59[74], stage0_59[75], stage0_59[76], stage0_59[77]},
      {stage1_61[12],stage1_60[56],stage1_59[100],stage1_58[142],stage1_57[163]}
   );
   gpc615_5 gpc2206 (
      {stage0_57[362], stage0_57[363], stage0_57[364], stage0_57[365], stage0_57[366]},
      {stage0_58[277]},
      {stage0_59[78], stage0_59[79], stage0_59[80], stage0_59[81], stage0_59[82], stage0_59[83]},
      {stage1_61[13],stage1_60[57],stage1_59[101],stage1_58[143],stage1_57[164]}
   );
   gpc615_5 gpc2207 (
      {stage0_57[367], stage0_57[368], stage0_57[369], stage0_57[370], stage0_57[371]},
      {stage0_58[278]},
      {stage0_59[84], stage0_59[85], stage0_59[86], stage0_59[87], stage0_59[88], stage0_59[89]},
      {stage1_61[14],stage1_60[58],stage1_59[102],stage1_58[144],stage1_57[165]}
   );
   gpc615_5 gpc2208 (
      {stage0_57[372], stage0_57[373], stage0_57[374], stage0_57[375], stage0_57[376]},
      {stage0_58[279]},
      {stage0_59[90], stage0_59[91], stage0_59[92], stage0_59[93], stage0_59[94], stage0_59[95]},
      {stage1_61[15],stage1_60[59],stage1_59[103],stage1_58[145],stage1_57[166]}
   );
   gpc615_5 gpc2209 (
      {stage0_57[377], stage0_57[378], stage0_57[379], stage0_57[380], stage0_57[381]},
      {stage0_58[280]},
      {stage0_59[96], stage0_59[97], stage0_59[98], stage0_59[99], stage0_59[100], stage0_59[101]},
      {stage1_61[16],stage1_60[60],stage1_59[104],stage1_58[146],stage1_57[167]}
   );
   gpc615_5 gpc2210 (
      {stage0_57[382], stage0_57[383], stage0_57[384], stage0_57[385], stage0_57[386]},
      {stage0_58[281]},
      {stage0_59[102], stage0_59[103], stage0_59[104], stage0_59[105], stage0_59[106], stage0_59[107]},
      {stage1_61[17],stage1_60[61],stage1_59[105],stage1_58[147],stage1_57[168]}
   );
   gpc615_5 gpc2211 (
      {stage0_57[387], stage0_57[388], stage0_57[389], stage0_57[390], stage0_57[391]},
      {stage0_58[282]},
      {stage0_59[108], stage0_59[109], stage0_59[110], stage0_59[111], stage0_59[112], stage0_59[113]},
      {stage1_61[18],stage1_60[62],stage1_59[106],stage1_58[148],stage1_57[169]}
   );
   gpc615_5 gpc2212 (
      {stage0_57[392], stage0_57[393], stage0_57[394], stage0_57[395], stage0_57[396]},
      {stage0_58[283]},
      {stage0_59[114], stage0_59[115], stage0_59[116], stage0_59[117], stage0_59[118], stage0_59[119]},
      {stage1_61[19],stage1_60[63],stage1_59[107],stage1_58[149],stage1_57[170]}
   );
   gpc615_5 gpc2213 (
      {stage0_57[397], stage0_57[398], stage0_57[399], stage0_57[400], stage0_57[401]},
      {stage0_58[284]},
      {stage0_59[120], stage0_59[121], stage0_59[122], stage0_59[123], stage0_59[124], stage0_59[125]},
      {stage1_61[20],stage1_60[64],stage1_59[108],stage1_58[150],stage1_57[171]}
   );
   gpc615_5 gpc2214 (
      {stage0_57[402], stage0_57[403], stage0_57[404], stage0_57[405], stage0_57[406]},
      {stage0_58[285]},
      {stage0_59[126], stage0_59[127], stage0_59[128], stage0_59[129], stage0_59[130], stage0_59[131]},
      {stage1_61[21],stage1_60[65],stage1_59[109],stage1_58[151],stage1_57[172]}
   );
   gpc615_5 gpc2215 (
      {stage0_57[407], stage0_57[408], stage0_57[409], stage0_57[410], stage0_57[411]},
      {stage0_58[286]},
      {stage0_59[132], stage0_59[133], stage0_59[134], stage0_59[135], stage0_59[136], stage0_59[137]},
      {stage1_61[22],stage1_60[66],stage1_59[110],stage1_58[152],stage1_57[173]}
   );
   gpc615_5 gpc2216 (
      {stage0_57[412], stage0_57[413], stage0_57[414], stage0_57[415], stage0_57[416]},
      {stage0_58[287]},
      {stage0_59[138], stage0_59[139], stage0_59[140], stage0_59[141], stage0_59[142], stage0_59[143]},
      {stage1_61[23],stage1_60[67],stage1_59[111],stage1_58[153],stage1_57[174]}
   );
   gpc615_5 gpc2217 (
      {stage0_57[417], stage0_57[418], stage0_57[419], stage0_57[420], stage0_57[421]},
      {stage0_58[288]},
      {stage0_59[144], stage0_59[145], stage0_59[146], stage0_59[147], stage0_59[148], stage0_59[149]},
      {stage1_61[24],stage1_60[68],stage1_59[112],stage1_58[154],stage1_57[175]}
   );
   gpc615_5 gpc2218 (
      {stage0_57[422], stage0_57[423], stage0_57[424], stage0_57[425], stage0_57[426]},
      {stage0_58[289]},
      {stage0_59[150], stage0_59[151], stage0_59[152], stage0_59[153], stage0_59[154], stage0_59[155]},
      {stage1_61[25],stage1_60[69],stage1_59[113],stage1_58[155],stage1_57[176]}
   );
   gpc615_5 gpc2219 (
      {stage0_57[427], stage0_57[428], stage0_57[429], stage0_57[430], stage0_57[431]},
      {stage0_58[290]},
      {stage0_59[156], stage0_59[157], stage0_59[158], stage0_59[159], stage0_59[160], stage0_59[161]},
      {stage1_61[26],stage1_60[70],stage1_59[114],stage1_58[156],stage1_57[177]}
   );
   gpc615_5 gpc2220 (
      {stage0_57[432], stage0_57[433], stage0_57[434], stage0_57[435], stage0_57[436]},
      {stage0_58[291]},
      {stage0_59[162], stage0_59[163], stage0_59[164], stage0_59[165], stage0_59[166], stage0_59[167]},
      {stage1_61[27],stage1_60[71],stage1_59[115],stage1_58[157],stage1_57[178]}
   );
   gpc615_5 gpc2221 (
      {stage0_57[437], stage0_57[438], stage0_57[439], stage0_57[440], stage0_57[441]},
      {stage0_58[292]},
      {stage0_59[168], stage0_59[169], stage0_59[170], stage0_59[171], stage0_59[172], stage0_59[173]},
      {stage1_61[28],stage1_60[72],stage1_59[116],stage1_58[158],stage1_57[179]}
   );
   gpc615_5 gpc2222 (
      {stage0_57[442], stage0_57[443], stage0_57[444], stage0_57[445], stage0_57[446]},
      {stage0_58[293]},
      {stage0_59[174], stage0_59[175], stage0_59[176], stage0_59[177], stage0_59[178], stage0_59[179]},
      {stage1_61[29],stage1_60[73],stage1_59[117],stage1_58[159],stage1_57[180]}
   );
   gpc615_5 gpc2223 (
      {stage0_57[447], stage0_57[448], stage0_57[449], stage0_57[450], stage0_57[451]},
      {stage0_58[294]},
      {stage0_59[180], stage0_59[181], stage0_59[182], stage0_59[183], stage0_59[184], stage0_59[185]},
      {stage1_61[30],stage1_60[74],stage1_59[118],stage1_58[160],stage1_57[181]}
   );
   gpc615_5 gpc2224 (
      {stage0_57[452], stage0_57[453], stage0_57[454], stage0_57[455], stage0_57[456]},
      {stage0_58[295]},
      {stage0_59[186], stage0_59[187], stage0_59[188], stage0_59[189], stage0_59[190], stage0_59[191]},
      {stage1_61[31],stage1_60[75],stage1_59[119],stage1_58[161],stage1_57[182]}
   );
   gpc615_5 gpc2225 (
      {stage0_57[457], stage0_57[458], stage0_57[459], stage0_57[460], stage0_57[461]},
      {stage0_58[296]},
      {stage0_59[192], stage0_59[193], stage0_59[194], stage0_59[195], stage0_59[196], stage0_59[197]},
      {stage1_61[32],stage1_60[76],stage1_59[120],stage1_58[162],stage1_57[183]}
   );
   gpc615_5 gpc2226 (
      {stage0_57[462], stage0_57[463], stage0_57[464], stage0_57[465], stage0_57[466]},
      {stage0_58[297]},
      {stage0_59[198], stage0_59[199], stage0_59[200], stage0_59[201], stage0_59[202], stage0_59[203]},
      {stage1_61[33],stage1_60[77],stage1_59[121],stage1_58[163],stage1_57[184]}
   );
   gpc615_5 gpc2227 (
      {stage0_57[467], stage0_57[468], stage0_57[469], stage0_57[470], stage0_57[471]},
      {stage0_58[298]},
      {stage0_59[204], stage0_59[205], stage0_59[206], stage0_59[207], stage0_59[208], stage0_59[209]},
      {stage1_61[34],stage1_60[78],stage1_59[122],stage1_58[164],stage1_57[185]}
   );
   gpc615_5 gpc2228 (
      {stage0_57[472], stage0_57[473], stage0_57[474], stage0_57[475], stage0_57[476]},
      {stage0_58[299]},
      {stage0_59[210], stage0_59[211], stage0_59[212], stage0_59[213], stage0_59[214], stage0_59[215]},
      {stage1_61[35],stage1_60[79],stage1_59[123],stage1_58[165],stage1_57[186]}
   );
   gpc615_5 gpc2229 (
      {stage0_57[477], stage0_57[478], stage0_57[479], stage0_57[480], stage0_57[481]},
      {stage0_58[300]},
      {stage0_59[216], stage0_59[217], stage0_59[218], stage0_59[219], stage0_59[220], stage0_59[221]},
      {stage1_61[36],stage1_60[80],stage1_59[124],stage1_58[166],stage1_57[187]}
   );
   gpc615_5 gpc2230 (
      {stage0_57[482], stage0_57[483], stage0_57[484], stage0_57[485], 1'b0},
      {stage0_58[301]},
      {stage0_59[222], stage0_59[223], stage0_59[224], stage0_59[225], stage0_59[226], stage0_59[227]},
      {stage1_61[37],stage1_60[81],stage1_59[125],stage1_58[167],stage1_57[188]}
   );
   gpc7_3 gpc2231 (
      {stage0_58[302], stage0_58[303], stage0_58[304], stage0_58[305], stage0_58[306], stage0_58[307], stage0_58[308]},
      {stage1_60[82],stage1_59[126],stage1_58[168]}
   );
   gpc7_3 gpc2232 (
      {stage0_58[309], stage0_58[310], stage0_58[311], stage0_58[312], stage0_58[313], stage0_58[314], stage0_58[315]},
      {stage1_60[83],stage1_59[127],stage1_58[169]}
   );
   gpc7_3 gpc2233 (
      {stage0_58[316], stage0_58[317], stage0_58[318], stage0_58[319], stage0_58[320], stage0_58[321], stage0_58[322]},
      {stage1_60[84],stage1_59[128],stage1_58[170]}
   );
   gpc7_3 gpc2234 (
      {stage0_58[323], stage0_58[324], stage0_58[325], stage0_58[326], stage0_58[327], stage0_58[328], stage0_58[329]},
      {stage1_60[85],stage1_59[129],stage1_58[171]}
   );
   gpc7_3 gpc2235 (
      {stage0_58[330], stage0_58[331], stage0_58[332], stage0_58[333], stage0_58[334], stage0_58[335], stage0_58[336]},
      {stage1_60[86],stage1_59[130],stage1_58[172]}
   );
   gpc7_3 gpc2236 (
      {stage0_58[337], stage0_58[338], stage0_58[339], stage0_58[340], stage0_58[341], stage0_58[342], stage0_58[343]},
      {stage1_60[87],stage1_59[131],stage1_58[173]}
   );
   gpc606_5 gpc2237 (
      {stage0_58[344], stage0_58[345], stage0_58[346], stage0_58[347], stage0_58[348], stage0_58[349]},
      {stage0_60[0], stage0_60[1], stage0_60[2], stage0_60[3], stage0_60[4], stage0_60[5]},
      {stage1_62[0],stage1_61[38],stage1_60[88],stage1_59[132],stage1_58[174]}
   );
   gpc606_5 gpc2238 (
      {stage0_58[350], stage0_58[351], stage0_58[352], stage0_58[353], stage0_58[354], stage0_58[355]},
      {stage0_60[6], stage0_60[7], stage0_60[8], stage0_60[9], stage0_60[10], stage0_60[11]},
      {stage1_62[1],stage1_61[39],stage1_60[89],stage1_59[133],stage1_58[175]}
   );
   gpc606_5 gpc2239 (
      {stage0_58[356], stage0_58[357], stage0_58[358], stage0_58[359], stage0_58[360], stage0_58[361]},
      {stage0_60[12], stage0_60[13], stage0_60[14], stage0_60[15], stage0_60[16], stage0_60[17]},
      {stage1_62[2],stage1_61[40],stage1_60[90],stage1_59[134],stage1_58[176]}
   );
   gpc606_5 gpc2240 (
      {stage0_58[362], stage0_58[363], stage0_58[364], stage0_58[365], stage0_58[366], stage0_58[367]},
      {stage0_60[18], stage0_60[19], stage0_60[20], stage0_60[21], stage0_60[22], stage0_60[23]},
      {stage1_62[3],stage1_61[41],stage1_60[91],stage1_59[135],stage1_58[177]}
   );
   gpc606_5 gpc2241 (
      {stage0_58[368], stage0_58[369], stage0_58[370], stage0_58[371], stage0_58[372], stage0_58[373]},
      {stage0_60[24], stage0_60[25], stage0_60[26], stage0_60[27], stage0_60[28], stage0_60[29]},
      {stage1_62[4],stage1_61[42],stage1_60[92],stage1_59[136],stage1_58[178]}
   );
   gpc606_5 gpc2242 (
      {stage0_58[374], stage0_58[375], stage0_58[376], stage0_58[377], stage0_58[378], stage0_58[379]},
      {stage0_60[30], stage0_60[31], stage0_60[32], stage0_60[33], stage0_60[34], stage0_60[35]},
      {stage1_62[5],stage1_61[43],stage1_60[93],stage1_59[137],stage1_58[179]}
   );
   gpc606_5 gpc2243 (
      {stage0_58[380], stage0_58[381], stage0_58[382], stage0_58[383], stage0_58[384], stage0_58[385]},
      {stage0_60[36], stage0_60[37], stage0_60[38], stage0_60[39], stage0_60[40], stage0_60[41]},
      {stage1_62[6],stage1_61[44],stage1_60[94],stage1_59[138],stage1_58[180]}
   );
   gpc606_5 gpc2244 (
      {stage0_58[386], stage0_58[387], stage0_58[388], stage0_58[389], stage0_58[390], stage0_58[391]},
      {stage0_60[42], stage0_60[43], stage0_60[44], stage0_60[45], stage0_60[46], stage0_60[47]},
      {stage1_62[7],stage1_61[45],stage1_60[95],stage1_59[139],stage1_58[181]}
   );
   gpc606_5 gpc2245 (
      {stage0_58[392], stage0_58[393], stage0_58[394], stage0_58[395], stage0_58[396], stage0_58[397]},
      {stage0_60[48], stage0_60[49], stage0_60[50], stage0_60[51], stage0_60[52], stage0_60[53]},
      {stage1_62[8],stage1_61[46],stage1_60[96],stage1_59[140],stage1_58[182]}
   );
   gpc606_5 gpc2246 (
      {stage0_58[398], stage0_58[399], stage0_58[400], stage0_58[401], stage0_58[402], stage0_58[403]},
      {stage0_60[54], stage0_60[55], stage0_60[56], stage0_60[57], stage0_60[58], stage0_60[59]},
      {stage1_62[9],stage1_61[47],stage1_60[97],stage1_59[141],stage1_58[183]}
   );
   gpc606_5 gpc2247 (
      {stage0_58[404], stage0_58[405], stage0_58[406], stage0_58[407], stage0_58[408], stage0_58[409]},
      {stage0_60[60], stage0_60[61], stage0_60[62], stage0_60[63], stage0_60[64], stage0_60[65]},
      {stage1_62[10],stage1_61[48],stage1_60[98],stage1_59[142],stage1_58[184]}
   );
   gpc606_5 gpc2248 (
      {stage0_58[410], stage0_58[411], stage0_58[412], stage0_58[413], stage0_58[414], stage0_58[415]},
      {stage0_60[66], stage0_60[67], stage0_60[68], stage0_60[69], stage0_60[70], stage0_60[71]},
      {stage1_62[11],stage1_61[49],stage1_60[99],stage1_59[143],stage1_58[185]}
   );
   gpc606_5 gpc2249 (
      {stage0_58[416], stage0_58[417], stage0_58[418], stage0_58[419], stage0_58[420], stage0_58[421]},
      {stage0_60[72], stage0_60[73], stage0_60[74], stage0_60[75], stage0_60[76], stage0_60[77]},
      {stage1_62[12],stage1_61[50],stage1_60[100],stage1_59[144],stage1_58[186]}
   );
   gpc606_5 gpc2250 (
      {stage0_58[422], stage0_58[423], stage0_58[424], stage0_58[425], stage0_58[426], stage0_58[427]},
      {stage0_60[78], stage0_60[79], stage0_60[80], stage0_60[81], stage0_60[82], stage0_60[83]},
      {stage1_62[13],stage1_61[51],stage1_60[101],stage1_59[145],stage1_58[187]}
   );
   gpc606_5 gpc2251 (
      {stage0_58[428], stage0_58[429], stage0_58[430], stage0_58[431], stage0_58[432], stage0_58[433]},
      {stage0_60[84], stage0_60[85], stage0_60[86], stage0_60[87], stage0_60[88], stage0_60[89]},
      {stage1_62[14],stage1_61[52],stage1_60[102],stage1_59[146],stage1_58[188]}
   );
   gpc606_5 gpc2252 (
      {stage0_58[434], stage0_58[435], stage0_58[436], stage0_58[437], stage0_58[438], stage0_58[439]},
      {stage0_60[90], stage0_60[91], stage0_60[92], stage0_60[93], stage0_60[94], stage0_60[95]},
      {stage1_62[15],stage1_61[53],stage1_60[103],stage1_59[147],stage1_58[189]}
   );
   gpc615_5 gpc2253 (
      {stage0_58[440], stage0_58[441], stage0_58[442], stage0_58[443], stage0_58[444]},
      {stage0_59[228]},
      {stage0_60[96], stage0_60[97], stage0_60[98], stage0_60[99], stage0_60[100], stage0_60[101]},
      {stage1_62[16],stage1_61[54],stage1_60[104],stage1_59[148],stage1_58[190]}
   );
   gpc615_5 gpc2254 (
      {stage0_58[445], stage0_58[446], stage0_58[447], stage0_58[448], stage0_58[449]},
      {stage0_59[229]},
      {stage0_60[102], stage0_60[103], stage0_60[104], stage0_60[105], stage0_60[106], stage0_60[107]},
      {stage1_62[17],stage1_61[55],stage1_60[105],stage1_59[149],stage1_58[191]}
   );
   gpc615_5 gpc2255 (
      {stage0_58[450], stage0_58[451], stage0_58[452], stage0_58[453], stage0_58[454]},
      {stage0_59[230]},
      {stage0_60[108], stage0_60[109], stage0_60[110], stage0_60[111], stage0_60[112], stage0_60[113]},
      {stage1_62[18],stage1_61[56],stage1_60[106],stage1_59[150],stage1_58[192]}
   );
   gpc615_5 gpc2256 (
      {stage0_58[455], stage0_58[456], stage0_58[457], stage0_58[458], stage0_58[459]},
      {stage0_59[231]},
      {stage0_60[114], stage0_60[115], stage0_60[116], stage0_60[117], stage0_60[118], stage0_60[119]},
      {stage1_62[19],stage1_61[57],stage1_60[107],stage1_59[151],stage1_58[193]}
   );
   gpc117_4 gpc2257 (
      {stage0_59[232], stage0_59[233], stage0_59[234], stage0_59[235], stage0_59[236], stage0_59[237], stage0_59[238]},
      {stage0_60[120]},
      {stage0_61[0]},
      {stage1_62[20],stage1_61[58],stage1_60[108],stage1_59[152]}
   );
   gpc117_4 gpc2258 (
      {stage0_59[239], stage0_59[240], stage0_59[241], stage0_59[242], stage0_59[243], stage0_59[244], stage0_59[245]},
      {stage0_60[121]},
      {stage0_61[1]},
      {stage1_62[21],stage1_61[59],stage1_60[109],stage1_59[153]}
   );
   gpc117_4 gpc2259 (
      {stage0_59[246], stage0_59[247], stage0_59[248], stage0_59[249], stage0_59[250], stage0_59[251], stage0_59[252]},
      {stage0_60[122]},
      {stage0_61[2]},
      {stage1_62[22],stage1_61[60],stage1_60[110],stage1_59[154]}
   );
   gpc117_4 gpc2260 (
      {stage0_59[253], stage0_59[254], stage0_59[255], stage0_59[256], stage0_59[257], stage0_59[258], stage0_59[259]},
      {stage0_60[123]},
      {stage0_61[3]},
      {stage1_62[23],stage1_61[61],stage1_60[111],stage1_59[155]}
   );
   gpc117_4 gpc2261 (
      {stage0_59[260], stage0_59[261], stage0_59[262], stage0_59[263], stage0_59[264], stage0_59[265], stage0_59[266]},
      {stage0_60[124]},
      {stage0_61[4]},
      {stage1_62[24],stage1_61[62],stage1_60[112],stage1_59[156]}
   );
   gpc117_4 gpc2262 (
      {stage0_59[267], stage0_59[268], stage0_59[269], stage0_59[270], stage0_59[271], stage0_59[272], stage0_59[273]},
      {stage0_60[125]},
      {stage0_61[5]},
      {stage1_62[25],stage1_61[63],stage1_60[113],stage1_59[157]}
   );
   gpc117_4 gpc2263 (
      {stage0_59[274], stage0_59[275], stage0_59[276], stage0_59[277], stage0_59[278], stage0_59[279], stage0_59[280]},
      {stage0_60[126]},
      {stage0_61[6]},
      {stage1_62[26],stage1_61[64],stage1_60[114],stage1_59[158]}
   );
   gpc117_4 gpc2264 (
      {stage0_59[281], stage0_59[282], stage0_59[283], stage0_59[284], stage0_59[285], stage0_59[286], stage0_59[287]},
      {stage0_60[127]},
      {stage0_61[7]},
      {stage1_62[27],stage1_61[65],stage1_60[115],stage1_59[159]}
   );
   gpc117_4 gpc2265 (
      {stage0_59[288], stage0_59[289], stage0_59[290], stage0_59[291], stage0_59[292], stage0_59[293], stage0_59[294]},
      {stage0_60[128]},
      {stage0_61[8]},
      {stage1_62[28],stage1_61[66],stage1_60[116],stage1_59[160]}
   );
   gpc117_4 gpc2266 (
      {stage0_59[295], stage0_59[296], stage0_59[297], stage0_59[298], stage0_59[299], stage0_59[300], stage0_59[301]},
      {stage0_60[129]},
      {stage0_61[9]},
      {stage1_62[29],stage1_61[67],stage1_60[117],stage1_59[161]}
   );
   gpc117_4 gpc2267 (
      {stage0_59[302], stage0_59[303], stage0_59[304], stage0_59[305], stage0_59[306], stage0_59[307], stage0_59[308]},
      {stage0_60[130]},
      {stage0_61[10]},
      {stage1_62[30],stage1_61[68],stage1_60[118],stage1_59[162]}
   );
   gpc117_4 gpc2268 (
      {stage0_59[309], stage0_59[310], stage0_59[311], stage0_59[312], stage0_59[313], stage0_59[314], stage0_59[315]},
      {stage0_60[131]},
      {stage0_61[11]},
      {stage1_62[31],stage1_61[69],stage1_60[119],stage1_59[163]}
   );
   gpc117_4 gpc2269 (
      {stage0_59[316], stage0_59[317], stage0_59[318], stage0_59[319], stage0_59[320], stage0_59[321], stage0_59[322]},
      {stage0_60[132]},
      {stage0_61[12]},
      {stage1_62[32],stage1_61[70],stage1_60[120],stage1_59[164]}
   );
   gpc117_4 gpc2270 (
      {stage0_59[323], stage0_59[324], stage0_59[325], stage0_59[326], stage0_59[327], stage0_59[328], stage0_59[329]},
      {stage0_60[133]},
      {stage0_61[13]},
      {stage1_62[33],stage1_61[71],stage1_60[121],stage1_59[165]}
   );
   gpc117_4 gpc2271 (
      {stage0_59[330], stage0_59[331], stage0_59[332], stage0_59[333], stage0_59[334], stage0_59[335], stage0_59[336]},
      {stage0_60[134]},
      {stage0_61[14]},
      {stage1_62[34],stage1_61[72],stage1_60[122],stage1_59[166]}
   );
   gpc606_5 gpc2272 (
      {stage0_59[337], stage0_59[338], stage0_59[339], stage0_59[340], stage0_59[341], stage0_59[342]},
      {stage0_61[15], stage0_61[16], stage0_61[17], stage0_61[18], stage0_61[19], stage0_61[20]},
      {stage1_63[0],stage1_62[35],stage1_61[73],stage1_60[123],stage1_59[167]}
   );
   gpc606_5 gpc2273 (
      {stage0_59[343], stage0_59[344], stage0_59[345], stage0_59[346], stage0_59[347], stage0_59[348]},
      {stage0_61[21], stage0_61[22], stage0_61[23], stage0_61[24], stage0_61[25], stage0_61[26]},
      {stage1_63[1],stage1_62[36],stage1_61[74],stage1_60[124],stage1_59[168]}
   );
   gpc606_5 gpc2274 (
      {stage0_59[349], stage0_59[350], stage0_59[351], stage0_59[352], stage0_59[353], stage0_59[354]},
      {stage0_61[27], stage0_61[28], stage0_61[29], stage0_61[30], stage0_61[31], stage0_61[32]},
      {stage1_63[2],stage1_62[37],stage1_61[75],stage1_60[125],stage1_59[169]}
   );
   gpc606_5 gpc2275 (
      {stage0_59[355], stage0_59[356], stage0_59[357], stage0_59[358], stage0_59[359], stage0_59[360]},
      {stage0_61[33], stage0_61[34], stage0_61[35], stage0_61[36], stage0_61[37], stage0_61[38]},
      {stage1_63[3],stage1_62[38],stage1_61[76],stage1_60[126],stage1_59[170]}
   );
   gpc606_5 gpc2276 (
      {stage0_59[361], stage0_59[362], stage0_59[363], stage0_59[364], stage0_59[365], stage0_59[366]},
      {stage0_61[39], stage0_61[40], stage0_61[41], stage0_61[42], stage0_61[43], stage0_61[44]},
      {stage1_63[4],stage1_62[39],stage1_61[77],stage1_60[127],stage1_59[171]}
   );
   gpc606_5 gpc2277 (
      {stage0_59[367], stage0_59[368], stage0_59[369], stage0_59[370], stage0_59[371], stage0_59[372]},
      {stage0_61[45], stage0_61[46], stage0_61[47], stage0_61[48], stage0_61[49], stage0_61[50]},
      {stage1_63[5],stage1_62[40],stage1_61[78],stage1_60[128],stage1_59[172]}
   );
   gpc606_5 gpc2278 (
      {stage0_59[373], stage0_59[374], stage0_59[375], stage0_59[376], stage0_59[377], stage0_59[378]},
      {stage0_61[51], stage0_61[52], stage0_61[53], stage0_61[54], stage0_61[55], stage0_61[56]},
      {stage1_63[6],stage1_62[41],stage1_61[79],stage1_60[129],stage1_59[173]}
   );
   gpc606_5 gpc2279 (
      {stage0_59[379], stage0_59[380], stage0_59[381], stage0_59[382], stage0_59[383], stage0_59[384]},
      {stage0_61[57], stage0_61[58], stage0_61[59], stage0_61[60], stage0_61[61], stage0_61[62]},
      {stage1_63[7],stage1_62[42],stage1_61[80],stage1_60[130],stage1_59[174]}
   );
   gpc606_5 gpc2280 (
      {stage0_59[385], stage0_59[386], stage0_59[387], stage0_59[388], stage0_59[389], stage0_59[390]},
      {stage0_61[63], stage0_61[64], stage0_61[65], stage0_61[66], stage0_61[67], stage0_61[68]},
      {stage1_63[8],stage1_62[43],stage1_61[81],stage1_60[131],stage1_59[175]}
   );
   gpc606_5 gpc2281 (
      {stage0_59[391], stage0_59[392], stage0_59[393], stage0_59[394], stage0_59[395], stage0_59[396]},
      {stage0_61[69], stage0_61[70], stage0_61[71], stage0_61[72], stage0_61[73], stage0_61[74]},
      {stage1_63[9],stage1_62[44],stage1_61[82],stage1_60[132],stage1_59[176]}
   );
   gpc606_5 gpc2282 (
      {stage0_59[397], stage0_59[398], stage0_59[399], stage0_59[400], stage0_59[401], stage0_59[402]},
      {stage0_61[75], stage0_61[76], stage0_61[77], stage0_61[78], stage0_61[79], stage0_61[80]},
      {stage1_63[10],stage1_62[45],stage1_61[83],stage1_60[133],stage1_59[177]}
   );
   gpc606_5 gpc2283 (
      {stage0_59[403], stage0_59[404], stage0_59[405], stage0_59[406], stage0_59[407], stage0_59[408]},
      {stage0_61[81], stage0_61[82], stage0_61[83], stage0_61[84], stage0_61[85], stage0_61[86]},
      {stage1_63[11],stage1_62[46],stage1_61[84],stage1_60[134],stage1_59[178]}
   );
   gpc606_5 gpc2284 (
      {stage0_59[409], stage0_59[410], stage0_59[411], stage0_59[412], stage0_59[413], stage0_59[414]},
      {stage0_61[87], stage0_61[88], stage0_61[89], stage0_61[90], stage0_61[91], stage0_61[92]},
      {stage1_63[12],stage1_62[47],stage1_61[85],stage1_60[135],stage1_59[179]}
   );
   gpc606_5 gpc2285 (
      {stage0_59[415], stage0_59[416], stage0_59[417], stage0_59[418], stage0_59[419], stage0_59[420]},
      {stage0_61[93], stage0_61[94], stage0_61[95], stage0_61[96], stage0_61[97], stage0_61[98]},
      {stage1_63[13],stage1_62[48],stage1_61[86],stage1_60[136],stage1_59[180]}
   );
   gpc606_5 gpc2286 (
      {stage0_59[421], stage0_59[422], stage0_59[423], stage0_59[424], stage0_59[425], stage0_59[426]},
      {stage0_61[99], stage0_61[100], stage0_61[101], stage0_61[102], stage0_61[103], stage0_61[104]},
      {stage1_63[14],stage1_62[49],stage1_61[87],stage1_60[137],stage1_59[181]}
   );
   gpc606_5 gpc2287 (
      {stage0_59[427], stage0_59[428], stage0_59[429], stage0_59[430], stage0_59[431], stage0_59[432]},
      {stage0_61[105], stage0_61[106], stage0_61[107], stage0_61[108], stage0_61[109], stage0_61[110]},
      {stage1_63[15],stage1_62[50],stage1_61[88],stage1_60[138],stage1_59[182]}
   );
   gpc606_5 gpc2288 (
      {stage0_59[433], stage0_59[434], stage0_59[435], stage0_59[436], stage0_59[437], stage0_59[438]},
      {stage0_61[111], stage0_61[112], stage0_61[113], stage0_61[114], stage0_61[115], stage0_61[116]},
      {stage1_63[16],stage1_62[51],stage1_61[89],stage1_60[139],stage1_59[183]}
   );
   gpc606_5 gpc2289 (
      {stage0_59[439], stage0_59[440], stage0_59[441], stage0_59[442], stage0_59[443], stage0_59[444]},
      {stage0_61[117], stage0_61[118], stage0_61[119], stage0_61[120], stage0_61[121], stage0_61[122]},
      {stage1_63[17],stage1_62[52],stage1_61[90],stage1_60[140],stage1_59[184]}
   );
   gpc606_5 gpc2290 (
      {stage0_59[445], stage0_59[446], stage0_59[447], stage0_59[448], stage0_59[449], stage0_59[450]},
      {stage0_61[123], stage0_61[124], stage0_61[125], stage0_61[126], stage0_61[127], stage0_61[128]},
      {stage1_63[18],stage1_62[53],stage1_61[91],stage1_60[141],stage1_59[185]}
   );
   gpc606_5 gpc2291 (
      {stage0_59[451], stage0_59[452], stage0_59[453], stage0_59[454], stage0_59[455], stage0_59[456]},
      {stage0_61[129], stage0_61[130], stage0_61[131], stage0_61[132], stage0_61[133], stage0_61[134]},
      {stage1_63[19],stage1_62[54],stage1_61[92],stage1_60[142],stage1_59[186]}
   );
   gpc606_5 gpc2292 (
      {stage0_59[457], stage0_59[458], stage0_59[459], stage0_59[460], stage0_59[461], stage0_59[462]},
      {stage0_61[135], stage0_61[136], stage0_61[137], stage0_61[138], stage0_61[139], stage0_61[140]},
      {stage1_63[20],stage1_62[55],stage1_61[93],stage1_60[143],stage1_59[187]}
   );
   gpc606_5 gpc2293 (
      {stage0_59[463], stage0_59[464], stage0_59[465], stage0_59[466], stage0_59[467], stage0_59[468]},
      {stage0_61[141], stage0_61[142], stage0_61[143], stage0_61[144], stage0_61[145], stage0_61[146]},
      {stage1_63[21],stage1_62[56],stage1_61[94],stage1_60[144],stage1_59[188]}
   );
   gpc606_5 gpc2294 (
      {stage0_60[135], stage0_60[136], stage0_60[137], stage0_60[138], stage0_60[139], stage0_60[140]},
      {stage0_62[0], stage0_62[1], stage0_62[2], stage0_62[3], stage0_62[4], stage0_62[5]},
      {stage1_64[0],stage1_63[22],stage1_62[57],stage1_61[95],stage1_60[145]}
   );
   gpc615_5 gpc2295 (
      {stage0_60[141], stage0_60[142], stage0_60[143], stage0_60[144], stage0_60[145]},
      {stage0_61[147]},
      {stage0_62[6], stage0_62[7], stage0_62[8], stage0_62[9], stage0_62[10], stage0_62[11]},
      {stage1_64[1],stage1_63[23],stage1_62[58],stage1_61[96],stage1_60[146]}
   );
   gpc615_5 gpc2296 (
      {stage0_60[146], stage0_60[147], stage0_60[148], stage0_60[149], stage0_60[150]},
      {stage0_61[148]},
      {stage0_62[12], stage0_62[13], stage0_62[14], stage0_62[15], stage0_62[16], stage0_62[17]},
      {stage1_64[2],stage1_63[24],stage1_62[59],stage1_61[97],stage1_60[147]}
   );
   gpc615_5 gpc2297 (
      {stage0_60[151], stage0_60[152], stage0_60[153], stage0_60[154], stage0_60[155]},
      {stage0_61[149]},
      {stage0_62[18], stage0_62[19], stage0_62[20], stage0_62[21], stage0_62[22], stage0_62[23]},
      {stage1_64[3],stage1_63[25],stage1_62[60],stage1_61[98],stage1_60[148]}
   );
   gpc615_5 gpc2298 (
      {stage0_60[156], stage0_60[157], stage0_60[158], stage0_60[159], stage0_60[160]},
      {stage0_61[150]},
      {stage0_62[24], stage0_62[25], stage0_62[26], stage0_62[27], stage0_62[28], stage0_62[29]},
      {stage1_64[4],stage1_63[26],stage1_62[61],stage1_61[99],stage1_60[149]}
   );
   gpc615_5 gpc2299 (
      {stage0_60[161], stage0_60[162], stage0_60[163], stage0_60[164], stage0_60[165]},
      {stage0_61[151]},
      {stage0_62[30], stage0_62[31], stage0_62[32], stage0_62[33], stage0_62[34], stage0_62[35]},
      {stage1_64[5],stage1_63[27],stage1_62[62],stage1_61[100],stage1_60[150]}
   );
   gpc615_5 gpc2300 (
      {stage0_60[166], stage0_60[167], stage0_60[168], stage0_60[169], stage0_60[170]},
      {stage0_61[152]},
      {stage0_62[36], stage0_62[37], stage0_62[38], stage0_62[39], stage0_62[40], stage0_62[41]},
      {stage1_64[6],stage1_63[28],stage1_62[63],stage1_61[101],stage1_60[151]}
   );
   gpc615_5 gpc2301 (
      {stage0_60[171], stage0_60[172], stage0_60[173], stage0_60[174], stage0_60[175]},
      {stage0_61[153]},
      {stage0_62[42], stage0_62[43], stage0_62[44], stage0_62[45], stage0_62[46], stage0_62[47]},
      {stage1_64[7],stage1_63[29],stage1_62[64],stage1_61[102],stage1_60[152]}
   );
   gpc615_5 gpc2302 (
      {stage0_60[176], stage0_60[177], stage0_60[178], stage0_60[179], stage0_60[180]},
      {stage0_61[154]},
      {stage0_62[48], stage0_62[49], stage0_62[50], stage0_62[51], stage0_62[52], stage0_62[53]},
      {stage1_64[8],stage1_63[30],stage1_62[65],stage1_61[103],stage1_60[153]}
   );
   gpc615_5 gpc2303 (
      {stage0_60[181], stage0_60[182], stage0_60[183], stage0_60[184], stage0_60[185]},
      {stage0_61[155]},
      {stage0_62[54], stage0_62[55], stage0_62[56], stage0_62[57], stage0_62[58], stage0_62[59]},
      {stage1_64[9],stage1_63[31],stage1_62[66],stage1_61[104],stage1_60[154]}
   );
   gpc615_5 gpc2304 (
      {stage0_60[186], stage0_60[187], stage0_60[188], stage0_60[189], stage0_60[190]},
      {stage0_61[156]},
      {stage0_62[60], stage0_62[61], stage0_62[62], stage0_62[63], stage0_62[64], stage0_62[65]},
      {stage1_64[10],stage1_63[32],stage1_62[67],stage1_61[105],stage1_60[155]}
   );
   gpc615_5 gpc2305 (
      {stage0_60[191], stage0_60[192], stage0_60[193], stage0_60[194], stage0_60[195]},
      {stage0_61[157]},
      {stage0_62[66], stage0_62[67], stage0_62[68], stage0_62[69], stage0_62[70], stage0_62[71]},
      {stage1_64[11],stage1_63[33],stage1_62[68],stage1_61[106],stage1_60[156]}
   );
   gpc615_5 gpc2306 (
      {stage0_60[196], stage0_60[197], stage0_60[198], stage0_60[199], stage0_60[200]},
      {stage0_61[158]},
      {stage0_62[72], stage0_62[73], stage0_62[74], stage0_62[75], stage0_62[76], stage0_62[77]},
      {stage1_64[12],stage1_63[34],stage1_62[69],stage1_61[107],stage1_60[157]}
   );
   gpc615_5 gpc2307 (
      {stage0_60[201], stage0_60[202], stage0_60[203], stage0_60[204], stage0_60[205]},
      {stage0_61[159]},
      {stage0_62[78], stage0_62[79], stage0_62[80], stage0_62[81], stage0_62[82], stage0_62[83]},
      {stage1_64[13],stage1_63[35],stage1_62[70],stage1_61[108],stage1_60[158]}
   );
   gpc615_5 gpc2308 (
      {stage0_60[206], stage0_60[207], stage0_60[208], stage0_60[209], stage0_60[210]},
      {stage0_61[160]},
      {stage0_62[84], stage0_62[85], stage0_62[86], stage0_62[87], stage0_62[88], stage0_62[89]},
      {stage1_64[14],stage1_63[36],stage1_62[71],stage1_61[109],stage1_60[159]}
   );
   gpc615_5 gpc2309 (
      {stage0_60[211], stage0_60[212], stage0_60[213], stage0_60[214], stage0_60[215]},
      {stage0_61[161]},
      {stage0_62[90], stage0_62[91], stage0_62[92], stage0_62[93], stage0_62[94], stage0_62[95]},
      {stage1_64[15],stage1_63[37],stage1_62[72],stage1_61[110],stage1_60[160]}
   );
   gpc615_5 gpc2310 (
      {stage0_60[216], stage0_60[217], stage0_60[218], stage0_60[219], stage0_60[220]},
      {stage0_61[162]},
      {stage0_62[96], stage0_62[97], stage0_62[98], stage0_62[99], stage0_62[100], stage0_62[101]},
      {stage1_64[16],stage1_63[38],stage1_62[73],stage1_61[111],stage1_60[161]}
   );
   gpc615_5 gpc2311 (
      {stage0_60[221], stage0_60[222], stage0_60[223], stage0_60[224], stage0_60[225]},
      {stage0_61[163]},
      {stage0_62[102], stage0_62[103], stage0_62[104], stage0_62[105], stage0_62[106], stage0_62[107]},
      {stage1_64[17],stage1_63[39],stage1_62[74],stage1_61[112],stage1_60[162]}
   );
   gpc615_5 gpc2312 (
      {stage0_60[226], stage0_60[227], stage0_60[228], stage0_60[229], stage0_60[230]},
      {stage0_61[164]},
      {stage0_62[108], stage0_62[109], stage0_62[110], stage0_62[111], stage0_62[112], stage0_62[113]},
      {stage1_64[18],stage1_63[40],stage1_62[75],stage1_61[113],stage1_60[163]}
   );
   gpc615_5 gpc2313 (
      {stage0_60[231], stage0_60[232], stage0_60[233], stage0_60[234], stage0_60[235]},
      {stage0_61[165]},
      {stage0_62[114], stage0_62[115], stage0_62[116], stage0_62[117], stage0_62[118], stage0_62[119]},
      {stage1_64[19],stage1_63[41],stage1_62[76],stage1_61[114],stage1_60[164]}
   );
   gpc615_5 gpc2314 (
      {stage0_60[236], stage0_60[237], stage0_60[238], stage0_60[239], stage0_60[240]},
      {stage0_61[166]},
      {stage0_62[120], stage0_62[121], stage0_62[122], stage0_62[123], stage0_62[124], stage0_62[125]},
      {stage1_64[20],stage1_63[42],stage1_62[77],stage1_61[115],stage1_60[165]}
   );
   gpc615_5 gpc2315 (
      {stage0_60[241], stage0_60[242], stage0_60[243], stage0_60[244], stage0_60[245]},
      {stage0_61[167]},
      {stage0_62[126], stage0_62[127], stage0_62[128], stage0_62[129], stage0_62[130], stage0_62[131]},
      {stage1_64[21],stage1_63[43],stage1_62[78],stage1_61[116],stage1_60[166]}
   );
   gpc615_5 gpc2316 (
      {stage0_60[246], stage0_60[247], stage0_60[248], stage0_60[249], stage0_60[250]},
      {stage0_61[168]},
      {stage0_62[132], stage0_62[133], stage0_62[134], stage0_62[135], stage0_62[136], stage0_62[137]},
      {stage1_64[22],stage1_63[44],stage1_62[79],stage1_61[117],stage1_60[167]}
   );
   gpc615_5 gpc2317 (
      {stage0_60[251], stage0_60[252], stage0_60[253], stage0_60[254], stage0_60[255]},
      {stage0_61[169]},
      {stage0_62[138], stage0_62[139], stage0_62[140], stage0_62[141], stage0_62[142], stage0_62[143]},
      {stage1_64[23],stage1_63[45],stage1_62[80],stage1_61[118],stage1_60[168]}
   );
   gpc615_5 gpc2318 (
      {stage0_60[256], stage0_60[257], stage0_60[258], stage0_60[259], stage0_60[260]},
      {stage0_61[170]},
      {stage0_62[144], stage0_62[145], stage0_62[146], stage0_62[147], stage0_62[148], stage0_62[149]},
      {stage1_64[24],stage1_63[46],stage1_62[81],stage1_61[119],stage1_60[169]}
   );
   gpc615_5 gpc2319 (
      {stage0_60[261], stage0_60[262], stage0_60[263], stage0_60[264], stage0_60[265]},
      {stage0_61[171]},
      {stage0_62[150], stage0_62[151], stage0_62[152], stage0_62[153], stage0_62[154], stage0_62[155]},
      {stage1_64[25],stage1_63[47],stage1_62[82],stage1_61[120],stage1_60[170]}
   );
   gpc615_5 gpc2320 (
      {stage0_60[266], stage0_60[267], stage0_60[268], stage0_60[269], stage0_60[270]},
      {stage0_61[172]},
      {stage0_62[156], stage0_62[157], stage0_62[158], stage0_62[159], stage0_62[160], stage0_62[161]},
      {stage1_64[26],stage1_63[48],stage1_62[83],stage1_61[121],stage1_60[171]}
   );
   gpc615_5 gpc2321 (
      {stage0_60[271], stage0_60[272], stage0_60[273], stage0_60[274], stage0_60[275]},
      {stage0_61[173]},
      {stage0_62[162], stage0_62[163], stage0_62[164], stage0_62[165], stage0_62[166], stage0_62[167]},
      {stage1_64[27],stage1_63[49],stage1_62[84],stage1_61[122],stage1_60[172]}
   );
   gpc615_5 gpc2322 (
      {stage0_60[276], stage0_60[277], stage0_60[278], stage0_60[279], stage0_60[280]},
      {stage0_61[174]},
      {stage0_62[168], stage0_62[169], stage0_62[170], stage0_62[171], stage0_62[172], stage0_62[173]},
      {stage1_64[28],stage1_63[50],stage1_62[85],stage1_61[123],stage1_60[173]}
   );
   gpc615_5 gpc2323 (
      {stage0_60[281], stage0_60[282], stage0_60[283], stage0_60[284], stage0_60[285]},
      {stage0_61[175]},
      {stage0_62[174], stage0_62[175], stage0_62[176], stage0_62[177], stage0_62[178], stage0_62[179]},
      {stage1_64[29],stage1_63[51],stage1_62[86],stage1_61[124],stage1_60[174]}
   );
   gpc615_5 gpc2324 (
      {stage0_60[286], stage0_60[287], stage0_60[288], stage0_60[289], stage0_60[290]},
      {stage0_61[176]},
      {stage0_62[180], stage0_62[181], stage0_62[182], stage0_62[183], stage0_62[184], stage0_62[185]},
      {stage1_64[30],stage1_63[52],stage1_62[87],stage1_61[125],stage1_60[175]}
   );
   gpc615_5 gpc2325 (
      {stage0_60[291], stage0_60[292], stage0_60[293], stage0_60[294], stage0_60[295]},
      {stage0_61[177]},
      {stage0_62[186], stage0_62[187], stage0_62[188], stage0_62[189], stage0_62[190], stage0_62[191]},
      {stage1_64[31],stage1_63[53],stage1_62[88],stage1_61[126],stage1_60[176]}
   );
   gpc615_5 gpc2326 (
      {stage0_60[296], stage0_60[297], stage0_60[298], stage0_60[299], stage0_60[300]},
      {stage0_61[178]},
      {stage0_62[192], stage0_62[193], stage0_62[194], stage0_62[195], stage0_62[196], stage0_62[197]},
      {stage1_64[32],stage1_63[54],stage1_62[89],stage1_61[127],stage1_60[177]}
   );
   gpc615_5 gpc2327 (
      {stage0_60[301], stage0_60[302], stage0_60[303], stage0_60[304], stage0_60[305]},
      {stage0_61[179]},
      {stage0_62[198], stage0_62[199], stage0_62[200], stage0_62[201], stage0_62[202], stage0_62[203]},
      {stage1_64[33],stage1_63[55],stage1_62[90],stage1_61[128],stage1_60[178]}
   );
   gpc615_5 gpc2328 (
      {stage0_60[306], stage0_60[307], stage0_60[308], stage0_60[309], stage0_60[310]},
      {stage0_61[180]},
      {stage0_62[204], stage0_62[205], stage0_62[206], stage0_62[207], stage0_62[208], stage0_62[209]},
      {stage1_64[34],stage1_63[56],stage1_62[91],stage1_61[129],stage1_60[179]}
   );
   gpc615_5 gpc2329 (
      {stage0_60[311], stage0_60[312], stage0_60[313], stage0_60[314], stage0_60[315]},
      {stage0_61[181]},
      {stage0_62[210], stage0_62[211], stage0_62[212], stage0_62[213], stage0_62[214], stage0_62[215]},
      {stage1_64[35],stage1_63[57],stage1_62[92],stage1_61[130],stage1_60[180]}
   );
   gpc615_5 gpc2330 (
      {stage0_60[316], stage0_60[317], stage0_60[318], stage0_60[319], stage0_60[320]},
      {stage0_61[182]},
      {stage0_62[216], stage0_62[217], stage0_62[218], stage0_62[219], stage0_62[220], stage0_62[221]},
      {stage1_64[36],stage1_63[58],stage1_62[93],stage1_61[131],stage1_60[181]}
   );
   gpc615_5 gpc2331 (
      {stage0_60[321], stage0_60[322], stage0_60[323], stage0_60[324], stage0_60[325]},
      {stage0_61[183]},
      {stage0_62[222], stage0_62[223], stage0_62[224], stage0_62[225], stage0_62[226], stage0_62[227]},
      {stage1_64[37],stage1_63[59],stage1_62[94],stage1_61[132],stage1_60[182]}
   );
   gpc615_5 gpc2332 (
      {stage0_60[326], stage0_60[327], stage0_60[328], stage0_60[329], stage0_60[330]},
      {stage0_61[184]},
      {stage0_62[228], stage0_62[229], stage0_62[230], stage0_62[231], stage0_62[232], stage0_62[233]},
      {stage1_64[38],stage1_63[60],stage1_62[95],stage1_61[133],stage1_60[183]}
   );
   gpc615_5 gpc2333 (
      {stage0_60[331], stage0_60[332], stage0_60[333], stage0_60[334], stage0_60[335]},
      {stage0_61[185]},
      {stage0_62[234], stage0_62[235], stage0_62[236], stage0_62[237], stage0_62[238], stage0_62[239]},
      {stage1_64[39],stage1_63[61],stage1_62[96],stage1_61[134],stage1_60[184]}
   );
   gpc615_5 gpc2334 (
      {stage0_60[336], stage0_60[337], stage0_60[338], stage0_60[339], stage0_60[340]},
      {stage0_61[186]},
      {stage0_62[240], stage0_62[241], stage0_62[242], stage0_62[243], stage0_62[244], stage0_62[245]},
      {stage1_64[40],stage1_63[62],stage1_62[97],stage1_61[135],stage1_60[185]}
   );
   gpc615_5 gpc2335 (
      {stage0_60[341], stage0_60[342], stage0_60[343], stage0_60[344], stage0_60[345]},
      {stage0_61[187]},
      {stage0_62[246], stage0_62[247], stage0_62[248], stage0_62[249], stage0_62[250], stage0_62[251]},
      {stage1_64[41],stage1_63[63],stage1_62[98],stage1_61[136],stage1_60[186]}
   );
   gpc615_5 gpc2336 (
      {stage0_60[346], stage0_60[347], stage0_60[348], stage0_60[349], stage0_60[350]},
      {stage0_61[188]},
      {stage0_62[252], stage0_62[253], stage0_62[254], stage0_62[255], stage0_62[256], stage0_62[257]},
      {stage1_64[42],stage1_63[64],stage1_62[99],stage1_61[137],stage1_60[187]}
   );
   gpc615_5 gpc2337 (
      {stage0_60[351], stage0_60[352], stage0_60[353], stage0_60[354], stage0_60[355]},
      {stage0_61[189]},
      {stage0_62[258], stage0_62[259], stage0_62[260], stage0_62[261], stage0_62[262], stage0_62[263]},
      {stage1_64[43],stage1_63[65],stage1_62[100],stage1_61[138],stage1_60[188]}
   );
   gpc615_5 gpc2338 (
      {stage0_60[356], stage0_60[357], stage0_60[358], stage0_60[359], stage0_60[360]},
      {stage0_61[190]},
      {stage0_62[264], stage0_62[265], stage0_62[266], stage0_62[267], stage0_62[268], stage0_62[269]},
      {stage1_64[44],stage1_63[66],stage1_62[101],stage1_61[139],stage1_60[189]}
   );
   gpc615_5 gpc2339 (
      {stage0_60[361], stage0_60[362], stage0_60[363], stage0_60[364], stage0_60[365]},
      {stage0_61[191]},
      {stage0_62[270], stage0_62[271], stage0_62[272], stage0_62[273], stage0_62[274], stage0_62[275]},
      {stage1_64[45],stage1_63[67],stage1_62[102],stage1_61[140],stage1_60[190]}
   );
   gpc615_5 gpc2340 (
      {stage0_60[366], stage0_60[367], stage0_60[368], stage0_60[369], stage0_60[370]},
      {stage0_61[192]},
      {stage0_62[276], stage0_62[277], stage0_62[278], stage0_62[279], stage0_62[280], stage0_62[281]},
      {stage1_64[46],stage1_63[68],stage1_62[103],stage1_61[141],stage1_60[191]}
   );
   gpc615_5 gpc2341 (
      {stage0_60[371], stage0_60[372], stage0_60[373], stage0_60[374], stage0_60[375]},
      {stage0_61[193]},
      {stage0_62[282], stage0_62[283], stage0_62[284], stage0_62[285], stage0_62[286], stage0_62[287]},
      {stage1_64[47],stage1_63[69],stage1_62[104],stage1_61[142],stage1_60[192]}
   );
   gpc615_5 gpc2342 (
      {stage0_60[376], stage0_60[377], stage0_60[378], stage0_60[379], stage0_60[380]},
      {stage0_61[194]},
      {stage0_62[288], stage0_62[289], stage0_62[290], stage0_62[291], stage0_62[292], stage0_62[293]},
      {stage1_64[48],stage1_63[70],stage1_62[105],stage1_61[143],stage1_60[193]}
   );
   gpc615_5 gpc2343 (
      {stage0_60[381], stage0_60[382], stage0_60[383], stage0_60[384], stage0_60[385]},
      {stage0_61[195]},
      {stage0_62[294], stage0_62[295], stage0_62[296], stage0_62[297], stage0_62[298], stage0_62[299]},
      {stage1_64[49],stage1_63[71],stage1_62[106],stage1_61[144],stage1_60[194]}
   );
   gpc615_5 gpc2344 (
      {stage0_60[386], stage0_60[387], stage0_60[388], stage0_60[389], stage0_60[390]},
      {stage0_61[196]},
      {stage0_62[300], stage0_62[301], stage0_62[302], stage0_62[303], stage0_62[304], stage0_62[305]},
      {stage1_64[50],stage1_63[72],stage1_62[107],stage1_61[145],stage1_60[195]}
   );
   gpc615_5 gpc2345 (
      {stage0_60[391], stage0_60[392], stage0_60[393], stage0_60[394], stage0_60[395]},
      {stage0_61[197]},
      {stage0_62[306], stage0_62[307], stage0_62[308], stage0_62[309], stage0_62[310], stage0_62[311]},
      {stage1_64[51],stage1_63[73],stage1_62[108],stage1_61[146],stage1_60[196]}
   );
   gpc615_5 gpc2346 (
      {stage0_60[396], stage0_60[397], stage0_60[398], stage0_60[399], stage0_60[400]},
      {stage0_61[198]},
      {stage0_62[312], stage0_62[313], stage0_62[314], stage0_62[315], stage0_62[316], stage0_62[317]},
      {stage1_64[52],stage1_63[74],stage1_62[109],stage1_61[147],stage1_60[197]}
   );
   gpc615_5 gpc2347 (
      {stage0_60[401], stage0_60[402], stage0_60[403], stage0_60[404], stage0_60[405]},
      {stage0_61[199]},
      {stage0_62[318], stage0_62[319], stage0_62[320], stage0_62[321], stage0_62[322], stage0_62[323]},
      {stage1_64[53],stage1_63[75],stage1_62[110],stage1_61[148],stage1_60[198]}
   );
   gpc615_5 gpc2348 (
      {stage0_60[406], stage0_60[407], stage0_60[408], stage0_60[409], stage0_60[410]},
      {stage0_61[200]},
      {stage0_62[324], stage0_62[325], stage0_62[326], stage0_62[327], stage0_62[328], stage0_62[329]},
      {stage1_64[54],stage1_63[76],stage1_62[111],stage1_61[149],stage1_60[199]}
   );
   gpc615_5 gpc2349 (
      {stage0_60[411], stage0_60[412], stage0_60[413], stage0_60[414], stage0_60[415]},
      {stage0_61[201]},
      {stage0_62[330], stage0_62[331], stage0_62[332], stage0_62[333], stage0_62[334], stage0_62[335]},
      {stage1_64[55],stage1_63[77],stage1_62[112],stage1_61[150],stage1_60[200]}
   );
   gpc615_5 gpc2350 (
      {stage0_60[416], stage0_60[417], stage0_60[418], stage0_60[419], stage0_60[420]},
      {stage0_61[202]},
      {stage0_62[336], stage0_62[337], stage0_62[338], stage0_62[339], stage0_62[340], stage0_62[341]},
      {stage1_64[56],stage1_63[78],stage1_62[113],stage1_61[151],stage1_60[201]}
   );
   gpc615_5 gpc2351 (
      {stage0_60[421], stage0_60[422], stage0_60[423], stage0_60[424], stage0_60[425]},
      {stage0_61[203]},
      {stage0_62[342], stage0_62[343], stage0_62[344], stage0_62[345], stage0_62[346], stage0_62[347]},
      {stage1_64[57],stage1_63[79],stage1_62[114],stage1_61[152],stage1_60[202]}
   );
   gpc615_5 gpc2352 (
      {stage0_60[426], stage0_60[427], stage0_60[428], stage0_60[429], stage0_60[430]},
      {stage0_61[204]},
      {stage0_62[348], stage0_62[349], stage0_62[350], stage0_62[351], stage0_62[352], stage0_62[353]},
      {stage1_64[58],stage1_63[80],stage1_62[115],stage1_61[153],stage1_60[203]}
   );
   gpc615_5 gpc2353 (
      {stage0_60[431], stage0_60[432], stage0_60[433], stage0_60[434], stage0_60[435]},
      {stage0_61[205]},
      {stage0_62[354], stage0_62[355], stage0_62[356], stage0_62[357], stage0_62[358], stage0_62[359]},
      {stage1_64[59],stage1_63[81],stage1_62[116],stage1_61[154],stage1_60[204]}
   );
   gpc615_5 gpc2354 (
      {stage0_60[436], stage0_60[437], stage0_60[438], stage0_60[439], stage0_60[440]},
      {stage0_61[206]},
      {stage0_62[360], stage0_62[361], stage0_62[362], stage0_62[363], stage0_62[364], stage0_62[365]},
      {stage1_64[60],stage1_63[82],stage1_62[117],stage1_61[155],stage1_60[205]}
   );
   gpc615_5 gpc2355 (
      {stage0_60[441], stage0_60[442], stage0_60[443], stage0_60[444], stage0_60[445]},
      {stage0_61[207]},
      {stage0_62[366], stage0_62[367], stage0_62[368], stage0_62[369], stage0_62[370], stage0_62[371]},
      {stage1_64[61],stage1_63[83],stage1_62[118],stage1_61[156],stage1_60[206]}
   );
   gpc615_5 gpc2356 (
      {stage0_60[446], stage0_60[447], stage0_60[448], stage0_60[449], stage0_60[450]},
      {stage0_61[208]},
      {stage0_62[372], stage0_62[373], stage0_62[374], stage0_62[375], stage0_62[376], stage0_62[377]},
      {stage1_64[62],stage1_63[84],stage1_62[119],stage1_61[157],stage1_60[207]}
   );
   gpc615_5 gpc2357 (
      {stage0_60[451], stage0_60[452], stage0_60[453], stage0_60[454], stage0_60[455]},
      {stage0_61[209]},
      {stage0_62[378], stage0_62[379], stage0_62[380], stage0_62[381], stage0_62[382], stage0_62[383]},
      {stage1_64[63],stage1_63[85],stage1_62[120],stage1_61[158],stage1_60[208]}
   );
   gpc615_5 gpc2358 (
      {stage0_60[456], stage0_60[457], stage0_60[458], stage0_60[459], stage0_60[460]},
      {stage0_61[210]},
      {stage0_62[384], stage0_62[385], stage0_62[386], stage0_62[387], stage0_62[388], stage0_62[389]},
      {stage1_64[64],stage1_63[86],stage1_62[121],stage1_61[159],stage1_60[209]}
   );
   gpc615_5 gpc2359 (
      {stage0_60[461], stage0_60[462], stage0_60[463], stage0_60[464], stage0_60[465]},
      {stage0_61[211]},
      {stage0_62[390], stage0_62[391], stage0_62[392], stage0_62[393], stage0_62[394], stage0_62[395]},
      {stage1_64[65],stage1_63[87],stage1_62[122],stage1_61[160],stage1_60[210]}
   );
   gpc615_5 gpc2360 (
      {stage0_60[466], stage0_60[467], stage0_60[468], stage0_60[469], stage0_60[470]},
      {stage0_61[212]},
      {stage0_62[396], stage0_62[397], stage0_62[398], stage0_62[399], stage0_62[400], stage0_62[401]},
      {stage1_64[66],stage1_63[88],stage1_62[123],stage1_61[161],stage1_60[211]}
   );
   gpc615_5 gpc2361 (
      {stage0_60[471], stage0_60[472], stage0_60[473], stage0_60[474], stage0_60[475]},
      {stage0_61[213]},
      {stage0_62[402], stage0_62[403], stage0_62[404], stage0_62[405], stage0_62[406], stage0_62[407]},
      {stage1_64[67],stage1_63[89],stage1_62[124],stage1_61[162],stage1_60[212]}
   );
   gpc615_5 gpc2362 (
      {stage0_60[476], stage0_60[477], stage0_60[478], stage0_60[479], stage0_60[480]},
      {stage0_61[214]},
      {stage0_62[408], stage0_62[409], stage0_62[410], stage0_62[411], stage0_62[412], stage0_62[413]},
      {stage1_64[68],stage1_63[90],stage1_62[125],stage1_61[163],stage1_60[213]}
   );
   gpc615_5 gpc2363 (
      {stage0_60[481], stage0_60[482], stage0_60[483], stage0_60[484], stage0_60[485]},
      {stage0_61[215]},
      {stage0_62[414], stage0_62[415], stage0_62[416], stage0_62[417], stage0_62[418], stage0_62[419]},
      {stage1_64[69],stage1_63[91],stage1_62[126],stage1_61[164],stage1_60[214]}
   );
   gpc615_5 gpc2364 (
      {stage0_61[216], stage0_61[217], stage0_61[218], stage0_61[219], stage0_61[220]},
      {stage0_62[420]},
      {stage0_63[0], stage0_63[1], stage0_63[2], stage0_63[3], stage0_63[4], stage0_63[5]},
      {stage1_65[0],stage1_64[70],stage1_63[92],stage1_62[127],stage1_61[165]}
   );
   gpc615_5 gpc2365 (
      {stage0_61[221], stage0_61[222], stage0_61[223], stage0_61[224], stage0_61[225]},
      {stage0_62[421]},
      {stage0_63[6], stage0_63[7], stage0_63[8], stage0_63[9], stage0_63[10], stage0_63[11]},
      {stage1_65[1],stage1_64[71],stage1_63[93],stage1_62[128],stage1_61[166]}
   );
   gpc615_5 gpc2366 (
      {stage0_61[226], stage0_61[227], stage0_61[228], stage0_61[229], stage0_61[230]},
      {stage0_62[422]},
      {stage0_63[12], stage0_63[13], stage0_63[14], stage0_63[15], stage0_63[16], stage0_63[17]},
      {stage1_65[2],stage1_64[72],stage1_63[94],stage1_62[129],stage1_61[167]}
   );
   gpc615_5 gpc2367 (
      {stage0_61[231], stage0_61[232], stage0_61[233], stage0_61[234], stage0_61[235]},
      {stage0_62[423]},
      {stage0_63[18], stage0_63[19], stage0_63[20], stage0_63[21], stage0_63[22], stage0_63[23]},
      {stage1_65[3],stage1_64[73],stage1_63[95],stage1_62[130],stage1_61[168]}
   );
   gpc615_5 gpc2368 (
      {stage0_61[236], stage0_61[237], stage0_61[238], stage0_61[239], stage0_61[240]},
      {stage0_62[424]},
      {stage0_63[24], stage0_63[25], stage0_63[26], stage0_63[27], stage0_63[28], stage0_63[29]},
      {stage1_65[4],stage1_64[74],stage1_63[96],stage1_62[131],stage1_61[169]}
   );
   gpc615_5 gpc2369 (
      {stage0_61[241], stage0_61[242], stage0_61[243], stage0_61[244], stage0_61[245]},
      {stage0_62[425]},
      {stage0_63[30], stage0_63[31], stage0_63[32], stage0_63[33], stage0_63[34], stage0_63[35]},
      {stage1_65[5],stage1_64[75],stage1_63[97],stage1_62[132],stage1_61[170]}
   );
   gpc615_5 gpc2370 (
      {stage0_61[246], stage0_61[247], stage0_61[248], stage0_61[249], stage0_61[250]},
      {stage0_62[426]},
      {stage0_63[36], stage0_63[37], stage0_63[38], stage0_63[39], stage0_63[40], stage0_63[41]},
      {stage1_65[6],stage1_64[76],stage1_63[98],stage1_62[133],stage1_61[171]}
   );
   gpc615_5 gpc2371 (
      {stage0_61[251], stage0_61[252], stage0_61[253], stage0_61[254], stage0_61[255]},
      {stage0_62[427]},
      {stage0_63[42], stage0_63[43], stage0_63[44], stage0_63[45], stage0_63[46], stage0_63[47]},
      {stage1_65[7],stage1_64[77],stage1_63[99],stage1_62[134],stage1_61[172]}
   );
   gpc615_5 gpc2372 (
      {stage0_61[256], stage0_61[257], stage0_61[258], stage0_61[259], stage0_61[260]},
      {stage0_62[428]},
      {stage0_63[48], stage0_63[49], stage0_63[50], stage0_63[51], stage0_63[52], stage0_63[53]},
      {stage1_65[8],stage1_64[78],stage1_63[100],stage1_62[135],stage1_61[173]}
   );
   gpc615_5 gpc2373 (
      {stage0_61[261], stage0_61[262], stage0_61[263], stage0_61[264], stage0_61[265]},
      {stage0_62[429]},
      {stage0_63[54], stage0_63[55], stage0_63[56], stage0_63[57], stage0_63[58], stage0_63[59]},
      {stage1_65[9],stage1_64[79],stage1_63[101],stage1_62[136],stage1_61[174]}
   );
   gpc615_5 gpc2374 (
      {stage0_61[266], stage0_61[267], stage0_61[268], stage0_61[269], stage0_61[270]},
      {stage0_62[430]},
      {stage0_63[60], stage0_63[61], stage0_63[62], stage0_63[63], stage0_63[64], stage0_63[65]},
      {stage1_65[10],stage1_64[80],stage1_63[102],stage1_62[137],stage1_61[175]}
   );
   gpc615_5 gpc2375 (
      {stage0_61[271], stage0_61[272], stage0_61[273], stage0_61[274], stage0_61[275]},
      {stage0_62[431]},
      {stage0_63[66], stage0_63[67], stage0_63[68], stage0_63[69], stage0_63[70], stage0_63[71]},
      {stage1_65[11],stage1_64[81],stage1_63[103],stage1_62[138],stage1_61[176]}
   );
   gpc615_5 gpc2376 (
      {stage0_61[276], stage0_61[277], stage0_61[278], stage0_61[279], stage0_61[280]},
      {stage0_62[432]},
      {stage0_63[72], stage0_63[73], stage0_63[74], stage0_63[75], stage0_63[76], stage0_63[77]},
      {stage1_65[12],stage1_64[82],stage1_63[104],stage1_62[139],stage1_61[177]}
   );
   gpc615_5 gpc2377 (
      {stage0_61[281], stage0_61[282], stage0_61[283], stage0_61[284], stage0_61[285]},
      {stage0_62[433]},
      {stage0_63[78], stage0_63[79], stage0_63[80], stage0_63[81], stage0_63[82], stage0_63[83]},
      {stage1_65[13],stage1_64[83],stage1_63[105],stage1_62[140],stage1_61[178]}
   );
   gpc615_5 gpc2378 (
      {stage0_61[286], stage0_61[287], stage0_61[288], stage0_61[289], stage0_61[290]},
      {stage0_62[434]},
      {stage0_63[84], stage0_63[85], stage0_63[86], stage0_63[87], stage0_63[88], stage0_63[89]},
      {stage1_65[14],stage1_64[84],stage1_63[106],stage1_62[141],stage1_61[179]}
   );
   gpc615_5 gpc2379 (
      {stage0_61[291], stage0_61[292], stage0_61[293], stage0_61[294], stage0_61[295]},
      {stage0_62[435]},
      {stage0_63[90], stage0_63[91], stage0_63[92], stage0_63[93], stage0_63[94], stage0_63[95]},
      {stage1_65[15],stage1_64[85],stage1_63[107],stage1_62[142],stage1_61[180]}
   );
   gpc615_5 gpc2380 (
      {stage0_61[296], stage0_61[297], stage0_61[298], stage0_61[299], stage0_61[300]},
      {stage0_62[436]},
      {stage0_63[96], stage0_63[97], stage0_63[98], stage0_63[99], stage0_63[100], stage0_63[101]},
      {stage1_65[16],stage1_64[86],stage1_63[108],stage1_62[143],stage1_61[181]}
   );
   gpc615_5 gpc2381 (
      {stage0_61[301], stage0_61[302], stage0_61[303], stage0_61[304], stage0_61[305]},
      {stage0_62[437]},
      {stage0_63[102], stage0_63[103], stage0_63[104], stage0_63[105], stage0_63[106], stage0_63[107]},
      {stage1_65[17],stage1_64[87],stage1_63[109],stage1_62[144],stage1_61[182]}
   );
   gpc615_5 gpc2382 (
      {stage0_61[306], stage0_61[307], stage0_61[308], stage0_61[309], stage0_61[310]},
      {stage0_62[438]},
      {stage0_63[108], stage0_63[109], stage0_63[110], stage0_63[111], stage0_63[112], stage0_63[113]},
      {stage1_65[18],stage1_64[88],stage1_63[110],stage1_62[145],stage1_61[183]}
   );
   gpc615_5 gpc2383 (
      {stage0_61[311], stage0_61[312], stage0_61[313], stage0_61[314], stage0_61[315]},
      {stage0_62[439]},
      {stage0_63[114], stage0_63[115], stage0_63[116], stage0_63[117], stage0_63[118], stage0_63[119]},
      {stage1_65[19],stage1_64[89],stage1_63[111],stage1_62[146],stage1_61[184]}
   );
   gpc615_5 gpc2384 (
      {stage0_61[316], stage0_61[317], stage0_61[318], stage0_61[319], stage0_61[320]},
      {stage0_62[440]},
      {stage0_63[120], stage0_63[121], stage0_63[122], stage0_63[123], stage0_63[124], stage0_63[125]},
      {stage1_65[20],stage1_64[90],stage1_63[112],stage1_62[147],stage1_61[185]}
   );
   gpc615_5 gpc2385 (
      {stage0_61[321], stage0_61[322], stage0_61[323], stage0_61[324], stage0_61[325]},
      {stage0_62[441]},
      {stage0_63[126], stage0_63[127], stage0_63[128], stage0_63[129], stage0_63[130], stage0_63[131]},
      {stage1_65[21],stage1_64[91],stage1_63[113],stage1_62[148],stage1_61[186]}
   );
   gpc615_5 gpc2386 (
      {stage0_61[326], stage0_61[327], stage0_61[328], stage0_61[329], stage0_61[330]},
      {stage0_62[442]},
      {stage0_63[132], stage0_63[133], stage0_63[134], stage0_63[135], stage0_63[136], stage0_63[137]},
      {stage1_65[22],stage1_64[92],stage1_63[114],stage1_62[149],stage1_61[187]}
   );
   gpc615_5 gpc2387 (
      {stage0_61[331], stage0_61[332], stage0_61[333], stage0_61[334], stage0_61[335]},
      {stage0_62[443]},
      {stage0_63[138], stage0_63[139], stage0_63[140], stage0_63[141], stage0_63[142], stage0_63[143]},
      {stage1_65[23],stage1_64[93],stage1_63[115],stage1_62[150],stage1_61[188]}
   );
   gpc615_5 gpc2388 (
      {stage0_61[336], stage0_61[337], stage0_61[338], stage0_61[339], stage0_61[340]},
      {stage0_62[444]},
      {stage0_63[144], stage0_63[145], stage0_63[146], stage0_63[147], stage0_63[148], stage0_63[149]},
      {stage1_65[24],stage1_64[94],stage1_63[116],stage1_62[151],stage1_61[189]}
   );
   gpc615_5 gpc2389 (
      {stage0_61[341], stage0_61[342], stage0_61[343], stage0_61[344], stage0_61[345]},
      {stage0_62[445]},
      {stage0_63[150], stage0_63[151], stage0_63[152], stage0_63[153], stage0_63[154], stage0_63[155]},
      {stage1_65[25],stage1_64[95],stage1_63[117],stage1_62[152],stage1_61[190]}
   );
   gpc615_5 gpc2390 (
      {stage0_61[346], stage0_61[347], stage0_61[348], stage0_61[349], stage0_61[350]},
      {stage0_62[446]},
      {stage0_63[156], stage0_63[157], stage0_63[158], stage0_63[159], stage0_63[160], stage0_63[161]},
      {stage1_65[26],stage1_64[96],stage1_63[118],stage1_62[153],stage1_61[191]}
   );
   gpc615_5 gpc2391 (
      {stage0_61[351], stage0_61[352], stage0_61[353], stage0_61[354], stage0_61[355]},
      {stage0_62[447]},
      {stage0_63[162], stage0_63[163], stage0_63[164], stage0_63[165], stage0_63[166], stage0_63[167]},
      {stage1_65[27],stage1_64[97],stage1_63[119],stage1_62[154],stage1_61[192]}
   );
   gpc615_5 gpc2392 (
      {stage0_61[356], stage0_61[357], stage0_61[358], stage0_61[359], stage0_61[360]},
      {stage0_62[448]},
      {stage0_63[168], stage0_63[169], stage0_63[170], stage0_63[171], stage0_63[172], stage0_63[173]},
      {stage1_65[28],stage1_64[98],stage1_63[120],stage1_62[155],stage1_61[193]}
   );
   gpc615_5 gpc2393 (
      {stage0_61[361], stage0_61[362], stage0_61[363], stage0_61[364], stage0_61[365]},
      {stage0_62[449]},
      {stage0_63[174], stage0_63[175], stage0_63[176], stage0_63[177], stage0_63[178], stage0_63[179]},
      {stage1_65[29],stage1_64[99],stage1_63[121],stage1_62[156],stage1_61[194]}
   );
   gpc615_5 gpc2394 (
      {stage0_61[366], stage0_61[367], stage0_61[368], stage0_61[369], stage0_61[370]},
      {stage0_62[450]},
      {stage0_63[180], stage0_63[181], stage0_63[182], stage0_63[183], stage0_63[184], stage0_63[185]},
      {stage1_65[30],stage1_64[100],stage1_63[122],stage1_62[157],stage1_61[195]}
   );
   gpc615_5 gpc2395 (
      {stage0_61[371], stage0_61[372], stage0_61[373], stage0_61[374], stage0_61[375]},
      {stage0_62[451]},
      {stage0_63[186], stage0_63[187], stage0_63[188], stage0_63[189], stage0_63[190], stage0_63[191]},
      {stage1_65[31],stage1_64[101],stage1_63[123],stage1_62[158],stage1_61[196]}
   );
   gpc615_5 gpc2396 (
      {stage0_61[376], stage0_61[377], stage0_61[378], stage0_61[379], stage0_61[380]},
      {stage0_62[452]},
      {stage0_63[192], stage0_63[193], stage0_63[194], stage0_63[195], stage0_63[196], stage0_63[197]},
      {stage1_65[32],stage1_64[102],stage1_63[124],stage1_62[159],stage1_61[197]}
   );
   gpc615_5 gpc2397 (
      {stage0_61[381], stage0_61[382], stage0_61[383], stage0_61[384], stage0_61[385]},
      {stage0_62[453]},
      {stage0_63[198], stage0_63[199], stage0_63[200], stage0_63[201], stage0_63[202], stage0_63[203]},
      {stage1_65[33],stage1_64[103],stage1_63[125],stage1_62[160],stage1_61[198]}
   );
   gpc615_5 gpc2398 (
      {stage0_61[386], stage0_61[387], stage0_61[388], stage0_61[389], stage0_61[390]},
      {stage0_62[454]},
      {stage0_63[204], stage0_63[205], stage0_63[206], stage0_63[207], stage0_63[208], stage0_63[209]},
      {stage1_65[34],stage1_64[104],stage1_63[126],stage1_62[161],stage1_61[199]}
   );
   gpc615_5 gpc2399 (
      {stage0_61[391], stage0_61[392], stage0_61[393], stage0_61[394], stage0_61[395]},
      {stage0_62[455]},
      {stage0_63[210], stage0_63[211], stage0_63[212], stage0_63[213], stage0_63[214], stage0_63[215]},
      {stage1_65[35],stage1_64[105],stage1_63[127],stage1_62[162],stage1_61[200]}
   );
   gpc615_5 gpc2400 (
      {stage0_61[396], stage0_61[397], stage0_61[398], stage0_61[399], stage0_61[400]},
      {stage0_62[456]},
      {stage0_63[216], stage0_63[217], stage0_63[218], stage0_63[219], stage0_63[220], stage0_63[221]},
      {stage1_65[36],stage1_64[106],stage1_63[128],stage1_62[163],stage1_61[201]}
   );
   gpc615_5 gpc2401 (
      {stage0_61[401], stage0_61[402], stage0_61[403], stage0_61[404], stage0_61[405]},
      {stage0_62[457]},
      {stage0_63[222], stage0_63[223], stage0_63[224], stage0_63[225], stage0_63[226], stage0_63[227]},
      {stage1_65[37],stage1_64[107],stage1_63[129],stage1_62[164],stage1_61[202]}
   );
   gpc615_5 gpc2402 (
      {stage0_61[406], stage0_61[407], stage0_61[408], stage0_61[409], stage0_61[410]},
      {stage0_62[458]},
      {stage0_63[228], stage0_63[229], stage0_63[230], stage0_63[231], stage0_63[232], stage0_63[233]},
      {stage1_65[38],stage1_64[108],stage1_63[130],stage1_62[165],stage1_61[203]}
   );
   gpc615_5 gpc2403 (
      {stage0_61[411], stage0_61[412], stage0_61[413], stage0_61[414], stage0_61[415]},
      {stage0_62[459]},
      {stage0_63[234], stage0_63[235], stage0_63[236], stage0_63[237], stage0_63[238], stage0_63[239]},
      {stage1_65[39],stage1_64[109],stage1_63[131],stage1_62[166],stage1_61[204]}
   );
   gpc615_5 gpc2404 (
      {stage0_61[416], stage0_61[417], stage0_61[418], stage0_61[419], stage0_61[420]},
      {stage0_62[460]},
      {stage0_63[240], stage0_63[241], stage0_63[242], stage0_63[243], stage0_63[244], stage0_63[245]},
      {stage1_65[40],stage1_64[110],stage1_63[132],stage1_62[167],stage1_61[205]}
   );
   gpc615_5 gpc2405 (
      {stage0_61[421], stage0_61[422], stage0_61[423], stage0_61[424], stage0_61[425]},
      {stage0_62[461]},
      {stage0_63[246], stage0_63[247], stage0_63[248], stage0_63[249], stage0_63[250], stage0_63[251]},
      {stage1_65[41],stage1_64[111],stage1_63[133],stage1_62[168],stage1_61[206]}
   );
   gpc615_5 gpc2406 (
      {stage0_61[426], stage0_61[427], stage0_61[428], stage0_61[429], stage0_61[430]},
      {stage0_62[462]},
      {stage0_63[252], stage0_63[253], stage0_63[254], stage0_63[255], stage0_63[256], stage0_63[257]},
      {stage1_65[42],stage1_64[112],stage1_63[134],stage1_62[169],stage1_61[207]}
   );
   gpc615_5 gpc2407 (
      {stage0_61[431], stage0_61[432], stage0_61[433], stage0_61[434], stage0_61[435]},
      {stage0_62[463]},
      {stage0_63[258], stage0_63[259], stage0_63[260], stage0_63[261], stage0_63[262], stage0_63[263]},
      {stage1_65[43],stage1_64[113],stage1_63[135],stage1_62[170],stage1_61[208]}
   );
   gpc615_5 gpc2408 (
      {stage0_61[436], stage0_61[437], stage0_61[438], stage0_61[439], stage0_61[440]},
      {stage0_62[464]},
      {stage0_63[264], stage0_63[265], stage0_63[266], stage0_63[267], stage0_63[268], stage0_63[269]},
      {stage1_65[44],stage1_64[114],stage1_63[136],stage1_62[171],stage1_61[209]}
   );
   gpc615_5 gpc2409 (
      {stage0_61[441], stage0_61[442], stage0_61[443], stage0_61[444], stage0_61[445]},
      {stage0_62[465]},
      {stage0_63[270], stage0_63[271], stage0_63[272], stage0_63[273], stage0_63[274], stage0_63[275]},
      {stage1_65[45],stage1_64[115],stage1_63[137],stage1_62[172],stage1_61[210]}
   );
   gpc615_5 gpc2410 (
      {stage0_61[446], stage0_61[447], stage0_61[448], stage0_61[449], stage0_61[450]},
      {stage0_62[466]},
      {stage0_63[276], stage0_63[277], stage0_63[278], stage0_63[279], stage0_63[280], stage0_63[281]},
      {stage1_65[46],stage1_64[116],stage1_63[138],stage1_62[173],stage1_61[211]}
   );
   gpc615_5 gpc2411 (
      {stage0_61[451], stage0_61[452], stage0_61[453], stage0_61[454], stage0_61[455]},
      {stage0_62[467]},
      {stage0_63[282], stage0_63[283], stage0_63[284], stage0_63[285], stage0_63[286], stage0_63[287]},
      {stage1_65[47],stage1_64[117],stage1_63[139],stage1_62[174],stage1_61[212]}
   );
   gpc615_5 gpc2412 (
      {stage0_61[456], stage0_61[457], stage0_61[458], stage0_61[459], stage0_61[460]},
      {stage0_62[468]},
      {stage0_63[288], stage0_63[289], stage0_63[290], stage0_63[291], stage0_63[292], stage0_63[293]},
      {stage1_65[48],stage1_64[118],stage1_63[140],stage1_62[175],stage1_61[213]}
   );
   gpc615_5 gpc2413 (
      {stage0_61[461], stage0_61[462], stage0_61[463], stage0_61[464], stage0_61[465]},
      {stage0_62[469]},
      {stage0_63[294], stage0_63[295], stage0_63[296], stage0_63[297], stage0_63[298], stage0_63[299]},
      {stage1_65[49],stage1_64[119],stage1_63[141],stage1_62[176],stage1_61[214]}
   );
   gpc615_5 gpc2414 (
      {stage0_61[466], stage0_61[467], stage0_61[468], stage0_61[469], stage0_61[470]},
      {stage0_62[470]},
      {stage0_63[300], stage0_63[301], stage0_63[302], stage0_63[303], stage0_63[304], stage0_63[305]},
      {stage1_65[50],stage1_64[120],stage1_63[142],stage1_62[177],stage1_61[215]}
   );
   gpc615_5 gpc2415 (
      {stage0_61[471], stage0_61[472], stage0_61[473], stage0_61[474], stage0_61[475]},
      {stage0_62[471]},
      {stage0_63[306], stage0_63[307], stage0_63[308], stage0_63[309], stage0_63[310], stage0_63[311]},
      {stage1_65[51],stage1_64[121],stage1_63[143],stage1_62[178],stage1_61[216]}
   );
   gpc615_5 gpc2416 (
      {stage0_61[476], stage0_61[477], stage0_61[478], stage0_61[479], stage0_61[480]},
      {stage0_62[472]},
      {stage0_63[312], stage0_63[313], stage0_63[314], stage0_63[315], stage0_63[316], stage0_63[317]},
      {stage1_65[52],stage1_64[122],stage1_63[144],stage1_62[179],stage1_61[217]}
   );
   gpc615_5 gpc2417 (
      {stage0_61[481], stage0_61[482], stage0_61[483], stage0_61[484], stage0_61[485]},
      {stage0_62[473]},
      {stage0_63[318], stage0_63[319], stage0_63[320], stage0_63[321], stage0_63[322], stage0_63[323]},
      {stage1_65[53],stage1_64[123],stage1_63[145],stage1_62[180],stage1_61[218]}
   );
   gpc1_1 gpc2418 (
      {stage0_0[448]},
      {stage1_0[87]}
   );
   gpc1_1 gpc2419 (
      {stage0_0[449]},
      {stage1_0[88]}
   );
   gpc1_1 gpc2420 (
      {stage0_0[450]},
      {stage1_0[89]}
   );
   gpc1_1 gpc2421 (
      {stage0_0[451]},
      {stage1_0[90]}
   );
   gpc1_1 gpc2422 (
      {stage0_0[452]},
      {stage1_0[91]}
   );
   gpc1_1 gpc2423 (
      {stage0_0[453]},
      {stage1_0[92]}
   );
   gpc1_1 gpc2424 (
      {stage0_0[454]},
      {stage1_0[93]}
   );
   gpc1_1 gpc2425 (
      {stage0_0[455]},
      {stage1_0[94]}
   );
   gpc1_1 gpc2426 (
      {stage0_0[456]},
      {stage1_0[95]}
   );
   gpc1_1 gpc2427 (
      {stage0_0[457]},
      {stage1_0[96]}
   );
   gpc1_1 gpc2428 (
      {stage0_0[458]},
      {stage1_0[97]}
   );
   gpc1_1 gpc2429 (
      {stage0_0[459]},
      {stage1_0[98]}
   );
   gpc1_1 gpc2430 (
      {stage0_0[460]},
      {stage1_0[99]}
   );
   gpc1_1 gpc2431 (
      {stage0_0[461]},
      {stage1_0[100]}
   );
   gpc1_1 gpc2432 (
      {stage0_0[462]},
      {stage1_0[101]}
   );
   gpc1_1 gpc2433 (
      {stage0_0[463]},
      {stage1_0[102]}
   );
   gpc1_1 gpc2434 (
      {stage0_0[464]},
      {stage1_0[103]}
   );
   gpc1_1 gpc2435 (
      {stage0_0[465]},
      {stage1_0[104]}
   );
   gpc1_1 gpc2436 (
      {stage0_0[466]},
      {stage1_0[105]}
   );
   gpc1_1 gpc2437 (
      {stage0_0[467]},
      {stage1_0[106]}
   );
   gpc1_1 gpc2438 (
      {stage0_0[468]},
      {stage1_0[107]}
   );
   gpc1_1 gpc2439 (
      {stage0_0[469]},
      {stage1_0[108]}
   );
   gpc1_1 gpc2440 (
      {stage0_0[470]},
      {stage1_0[109]}
   );
   gpc1_1 gpc2441 (
      {stage0_0[471]},
      {stage1_0[110]}
   );
   gpc1_1 gpc2442 (
      {stage0_0[472]},
      {stage1_0[111]}
   );
   gpc1_1 gpc2443 (
      {stage0_0[473]},
      {stage1_0[112]}
   );
   gpc1_1 gpc2444 (
      {stage0_0[474]},
      {stage1_0[113]}
   );
   gpc1_1 gpc2445 (
      {stage0_0[475]},
      {stage1_0[114]}
   );
   gpc1_1 gpc2446 (
      {stage0_0[476]},
      {stage1_0[115]}
   );
   gpc1_1 gpc2447 (
      {stage0_0[477]},
      {stage1_0[116]}
   );
   gpc1_1 gpc2448 (
      {stage0_0[478]},
      {stage1_0[117]}
   );
   gpc1_1 gpc2449 (
      {stage0_0[479]},
      {stage1_0[118]}
   );
   gpc1_1 gpc2450 (
      {stage0_0[480]},
      {stage1_0[119]}
   );
   gpc1_1 gpc2451 (
      {stage0_0[481]},
      {stage1_0[120]}
   );
   gpc1_1 gpc2452 (
      {stage0_0[482]},
      {stage1_0[121]}
   );
   gpc1_1 gpc2453 (
      {stage0_0[483]},
      {stage1_0[122]}
   );
   gpc1_1 gpc2454 (
      {stage0_0[484]},
      {stage1_0[123]}
   );
   gpc1_1 gpc2455 (
      {stage0_0[485]},
      {stage1_0[124]}
   );
   gpc1_1 gpc2456 (
      {stage0_1[439]},
      {stage1_1[129]}
   );
   gpc1_1 gpc2457 (
      {stage0_1[440]},
      {stage1_1[130]}
   );
   gpc1_1 gpc2458 (
      {stage0_1[441]},
      {stage1_1[131]}
   );
   gpc1_1 gpc2459 (
      {stage0_1[442]},
      {stage1_1[132]}
   );
   gpc1_1 gpc2460 (
      {stage0_1[443]},
      {stage1_1[133]}
   );
   gpc1_1 gpc2461 (
      {stage0_1[444]},
      {stage1_1[134]}
   );
   gpc1_1 gpc2462 (
      {stage0_1[445]},
      {stage1_1[135]}
   );
   gpc1_1 gpc2463 (
      {stage0_1[446]},
      {stage1_1[136]}
   );
   gpc1_1 gpc2464 (
      {stage0_1[447]},
      {stage1_1[137]}
   );
   gpc1_1 gpc2465 (
      {stage0_1[448]},
      {stage1_1[138]}
   );
   gpc1_1 gpc2466 (
      {stage0_1[449]},
      {stage1_1[139]}
   );
   gpc1_1 gpc2467 (
      {stage0_1[450]},
      {stage1_1[140]}
   );
   gpc1_1 gpc2468 (
      {stage0_1[451]},
      {stage1_1[141]}
   );
   gpc1_1 gpc2469 (
      {stage0_1[452]},
      {stage1_1[142]}
   );
   gpc1_1 gpc2470 (
      {stage0_1[453]},
      {stage1_1[143]}
   );
   gpc1_1 gpc2471 (
      {stage0_1[454]},
      {stage1_1[144]}
   );
   gpc1_1 gpc2472 (
      {stage0_1[455]},
      {stage1_1[145]}
   );
   gpc1_1 gpc2473 (
      {stage0_1[456]},
      {stage1_1[146]}
   );
   gpc1_1 gpc2474 (
      {stage0_1[457]},
      {stage1_1[147]}
   );
   gpc1_1 gpc2475 (
      {stage0_1[458]},
      {stage1_1[148]}
   );
   gpc1_1 gpc2476 (
      {stage0_1[459]},
      {stage1_1[149]}
   );
   gpc1_1 gpc2477 (
      {stage0_1[460]},
      {stage1_1[150]}
   );
   gpc1_1 gpc2478 (
      {stage0_1[461]},
      {stage1_1[151]}
   );
   gpc1_1 gpc2479 (
      {stage0_1[462]},
      {stage1_1[152]}
   );
   gpc1_1 gpc2480 (
      {stage0_1[463]},
      {stage1_1[153]}
   );
   gpc1_1 gpc2481 (
      {stage0_1[464]},
      {stage1_1[154]}
   );
   gpc1_1 gpc2482 (
      {stage0_1[465]},
      {stage1_1[155]}
   );
   gpc1_1 gpc2483 (
      {stage0_1[466]},
      {stage1_1[156]}
   );
   gpc1_1 gpc2484 (
      {stage0_1[467]},
      {stage1_1[157]}
   );
   gpc1_1 gpc2485 (
      {stage0_1[468]},
      {stage1_1[158]}
   );
   gpc1_1 gpc2486 (
      {stage0_1[469]},
      {stage1_1[159]}
   );
   gpc1_1 gpc2487 (
      {stage0_1[470]},
      {stage1_1[160]}
   );
   gpc1_1 gpc2488 (
      {stage0_1[471]},
      {stage1_1[161]}
   );
   gpc1_1 gpc2489 (
      {stage0_1[472]},
      {stage1_1[162]}
   );
   gpc1_1 gpc2490 (
      {stage0_1[473]},
      {stage1_1[163]}
   );
   gpc1_1 gpc2491 (
      {stage0_1[474]},
      {stage1_1[164]}
   );
   gpc1_1 gpc2492 (
      {stage0_1[475]},
      {stage1_1[165]}
   );
   gpc1_1 gpc2493 (
      {stage0_1[476]},
      {stage1_1[166]}
   );
   gpc1_1 gpc2494 (
      {stage0_1[477]},
      {stage1_1[167]}
   );
   gpc1_1 gpc2495 (
      {stage0_1[478]},
      {stage1_1[168]}
   );
   gpc1_1 gpc2496 (
      {stage0_1[479]},
      {stage1_1[169]}
   );
   gpc1_1 gpc2497 (
      {stage0_1[480]},
      {stage1_1[170]}
   );
   gpc1_1 gpc2498 (
      {stage0_1[481]},
      {stage1_1[171]}
   );
   gpc1_1 gpc2499 (
      {stage0_1[482]},
      {stage1_1[172]}
   );
   gpc1_1 gpc2500 (
      {stage0_1[483]},
      {stage1_1[173]}
   );
   gpc1_1 gpc2501 (
      {stage0_1[484]},
      {stage1_1[174]}
   );
   gpc1_1 gpc2502 (
      {stage0_1[485]},
      {stage1_1[175]}
   );
   gpc1_1 gpc2503 (
      {stage0_3[466]},
      {stage1_3[195]}
   );
   gpc1_1 gpc2504 (
      {stage0_3[467]},
      {stage1_3[196]}
   );
   gpc1_1 gpc2505 (
      {stage0_3[468]},
      {stage1_3[197]}
   );
   gpc1_1 gpc2506 (
      {stage0_3[469]},
      {stage1_3[198]}
   );
   gpc1_1 gpc2507 (
      {stage0_3[470]},
      {stage1_3[199]}
   );
   gpc1_1 gpc2508 (
      {stage0_3[471]},
      {stage1_3[200]}
   );
   gpc1_1 gpc2509 (
      {stage0_3[472]},
      {stage1_3[201]}
   );
   gpc1_1 gpc2510 (
      {stage0_3[473]},
      {stage1_3[202]}
   );
   gpc1_1 gpc2511 (
      {stage0_3[474]},
      {stage1_3[203]}
   );
   gpc1_1 gpc2512 (
      {stage0_3[475]},
      {stage1_3[204]}
   );
   gpc1_1 gpc2513 (
      {stage0_3[476]},
      {stage1_3[205]}
   );
   gpc1_1 gpc2514 (
      {stage0_3[477]},
      {stage1_3[206]}
   );
   gpc1_1 gpc2515 (
      {stage0_3[478]},
      {stage1_3[207]}
   );
   gpc1_1 gpc2516 (
      {stage0_3[479]},
      {stage1_3[208]}
   );
   gpc1_1 gpc2517 (
      {stage0_3[480]},
      {stage1_3[209]}
   );
   gpc1_1 gpc2518 (
      {stage0_3[481]},
      {stage1_3[210]}
   );
   gpc1_1 gpc2519 (
      {stage0_3[482]},
      {stage1_3[211]}
   );
   gpc1_1 gpc2520 (
      {stage0_3[483]},
      {stage1_3[212]}
   );
   gpc1_1 gpc2521 (
      {stage0_3[484]},
      {stage1_3[213]}
   );
   gpc1_1 gpc2522 (
      {stage0_3[485]},
      {stage1_3[214]}
   );
   gpc1_1 gpc2523 (
      {stage0_6[466]},
      {stage1_6[194]}
   );
   gpc1_1 gpc2524 (
      {stage0_6[467]},
      {stage1_6[195]}
   );
   gpc1_1 gpc2525 (
      {stage0_6[468]},
      {stage1_6[196]}
   );
   gpc1_1 gpc2526 (
      {stage0_6[469]},
      {stage1_6[197]}
   );
   gpc1_1 gpc2527 (
      {stage0_6[470]},
      {stage1_6[198]}
   );
   gpc1_1 gpc2528 (
      {stage0_6[471]},
      {stage1_6[199]}
   );
   gpc1_1 gpc2529 (
      {stage0_6[472]},
      {stage1_6[200]}
   );
   gpc1_1 gpc2530 (
      {stage0_6[473]},
      {stage1_6[201]}
   );
   gpc1_1 gpc2531 (
      {stage0_6[474]},
      {stage1_6[202]}
   );
   gpc1_1 gpc2532 (
      {stage0_6[475]},
      {stage1_6[203]}
   );
   gpc1_1 gpc2533 (
      {stage0_6[476]},
      {stage1_6[204]}
   );
   gpc1_1 gpc2534 (
      {stage0_6[477]},
      {stage1_6[205]}
   );
   gpc1_1 gpc2535 (
      {stage0_6[478]},
      {stage1_6[206]}
   );
   gpc1_1 gpc2536 (
      {stage0_6[479]},
      {stage1_6[207]}
   );
   gpc1_1 gpc2537 (
      {stage0_6[480]},
      {stage1_6[208]}
   );
   gpc1_1 gpc2538 (
      {stage0_6[481]},
      {stage1_6[209]}
   );
   gpc1_1 gpc2539 (
      {stage0_6[482]},
      {stage1_6[210]}
   );
   gpc1_1 gpc2540 (
      {stage0_6[483]},
      {stage1_6[211]}
   );
   gpc1_1 gpc2541 (
      {stage0_6[484]},
      {stage1_6[212]}
   );
   gpc1_1 gpc2542 (
      {stage0_6[485]},
      {stage1_6[213]}
   );
   gpc1_1 gpc2543 (
      {stage0_7[462]},
      {stage1_7[197]}
   );
   gpc1_1 gpc2544 (
      {stage0_7[463]},
      {stage1_7[198]}
   );
   gpc1_1 gpc2545 (
      {stage0_7[464]},
      {stage1_7[199]}
   );
   gpc1_1 gpc2546 (
      {stage0_7[465]},
      {stage1_7[200]}
   );
   gpc1_1 gpc2547 (
      {stage0_7[466]},
      {stage1_7[201]}
   );
   gpc1_1 gpc2548 (
      {stage0_7[467]},
      {stage1_7[202]}
   );
   gpc1_1 gpc2549 (
      {stage0_7[468]},
      {stage1_7[203]}
   );
   gpc1_1 gpc2550 (
      {stage0_7[469]},
      {stage1_7[204]}
   );
   gpc1_1 gpc2551 (
      {stage0_7[470]},
      {stage1_7[205]}
   );
   gpc1_1 gpc2552 (
      {stage0_7[471]},
      {stage1_7[206]}
   );
   gpc1_1 gpc2553 (
      {stage0_7[472]},
      {stage1_7[207]}
   );
   gpc1_1 gpc2554 (
      {stage0_7[473]},
      {stage1_7[208]}
   );
   gpc1_1 gpc2555 (
      {stage0_7[474]},
      {stage1_7[209]}
   );
   gpc1_1 gpc2556 (
      {stage0_7[475]},
      {stage1_7[210]}
   );
   gpc1_1 gpc2557 (
      {stage0_7[476]},
      {stage1_7[211]}
   );
   gpc1_1 gpc2558 (
      {stage0_7[477]},
      {stage1_7[212]}
   );
   gpc1_1 gpc2559 (
      {stage0_7[478]},
      {stage1_7[213]}
   );
   gpc1_1 gpc2560 (
      {stage0_7[479]},
      {stage1_7[214]}
   );
   gpc1_1 gpc2561 (
      {stage0_7[480]},
      {stage1_7[215]}
   );
   gpc1_1 gpc2562 (
      {stage0_7[481]},
      {stage1_7[216]}
   );
   gpc1_1 gpc2563 (
      {stage0_7[482]},
      {stage1_7[217]}
   );
   gpc1_1 gpc2564 (
      {stage0_7[483]},
      {stage1_7[218]}
   );
   gpc1_1 gpc2565 (
      {stage0_7[484]},
      {stage1_7[219]}
   );
   gpc1_1 gpc2566 (
      {stage0_7[485]},
      {stage1_7[220]}
   );
   gpc1_1 gpc2567 (
      {stage0_8[476]},
      {stage1_8[196]}
   );
   gpc1_1 gpc2568 (
      {stage0_8[477]},
      {stage1_8[197]}
   );
   gpc1_1 gpc2569 (
      {stage0_8[478]},
      {stage1_8[198]}
   );
   gpc1_1 gpc2570 (
      {stage0_8[479]},
      {stage1_8[199]}
   );
   gpc1_1 gpc2571 (
      {stage0_8[480]},
      {stage1_8[200]}
   );
   gpc1_1 gpc2572 (
      {stage0_8[481]},
      {stage1_8[201]}
   );
   gpc1_1 gpc2573 (
      {stage0_8[482]},
      {stage1_8[202]}
   );
   gpc1_1 gpc2574 (
      {stage0_8[483]},
      {stage1_8[203]}
   );
   gpc1_1 gpc2575 (
      {stage0_8[484]},
      {stage1_8[204]}
   );
   gpc1_1 gpc2576 (
      {stage0_8[485]},
      {stage1_8[205]}
   );
   gpc1_1 gpc2577 (
      {stage0_9[468]},
      {stage1_9[196]}
   );
   gpc1_1 gpc2578 (
      {stage0_9[469]},
      {stage1_9[197]}
   );
   gpc1_1 gpc2579 (
      {stage0_9[470]},
      {stage1_9[198]}
   );
   gpc1_1 gpc2580 (
      {stage0_9[471]},
      {stage1_9[199]}
   );
   gpc1_1 gpc2581 (
      {stage0_9[472]},
      {stage1_9[200]}
   );
   gpc1_1 gpc2582 (
      {stage0_9[473]},
      {stage1_9[201]}
   );
   gpc1_1 gpc2583 (
      {stage0_9[474]},
      {stage1_9[202]}
   );
   gpc1_1 gpc2584 (
      {stage0_9[475]},
      {stage1_9[203]}
   );
   gpc1_1 gpc2585 (
      {stage0_9[476]},
      {stage1_9[204]}
   );
   gpc1_1 gpc2586 (
      {stage0_9[477]},
      {stage1_9[205]}
   );
   gpc1_1 gpc2587 (
      {stage0_9[478]},
      {stage1_9[206]}
   );
   gpc1_1 gpc2588 (
      {stage0_9[479]},
      {stage1_9[207]}
   );
   gpc1_1 gpc2589 (
      {stage0_9[480]},
      {stage1_9[208]}
   );
   gpc1_1 gpc2590 (
      {stage0_9[481]},
      {stage1_9[209]}
   );
   gpc1_1 gpc2591 (
      {stage0_9[482]},
      {stage1_9[210]}
   );
   gpc1_1 gpc2592 (
      {stage0_9[483]},
      {stage1_9[211]}
   );
   gpc1_1 gpc2593 (
      {stage0_9[484]},
      {stage1_9[212]}
   );
   gpc1_1 gpc2594 (
      {stage0_9[485]},
      {stage1_9[213]}
   );
   gpc1_1 gpc2595 (
      {stage0_10[384]},
      {stage1_10[183]}
   );
   gpc1_1 gpc2596 (
      {stage0_10[385]},
      {stage1_10[184]}
   );
   gpc1_1 gpc2597 (
      {stage0_10[386]},
      {stage1_10[185]}
   );
   gpc1_1 gpc2598 (
      {stage0_10[387]},
      {stage1_10[186]}
   );
   gpc1_1 gpc2599 (
      {stage0_10[388]},
      {stage1_10[187]}
   );
   gpc1_1 gpc2600 (
      {stage0_10[389]},
      {stage1_10[188]}
   );
   gpc1_1 gpc2601 (
      {stage0_10[390]},
      {stage1_10[189]}
   );
   gpc1_1 gpc2602 (
      {stage0_10[391]},
      {stage1_10[190]}
   );
   gpc1_1 gpc2603 (
      {stage0_10[392]},
      {stage1_10[191]}
   );
   gpc1_1 gpc2604 (
      {stage0_10[393]},
      {stage1_10[192]}
   );
   gpc1_1 gpc2605 (
      {stage0_10[394]},
      {stage1_10[193]}
   );
   gpc1_1 gpc2606 (
      {stage0_10[395]},
      {stage1_10[194]}
   );
   gpc1_1 gpc2607 (
      {stage0_10[396]},
      {stage1_10[195]}
   );
   gpc1_1 gpc2608 (
      {stage0_10[397]},
      {stage1_10[196]}
   );
   gpc1_1 gpc2609 (
      {stage0_10[398]},
      {stage1_10[197]}
   );
   gpc1_1 gpc2610 (
      {stage0_10[399]},
      {stage1_10[198]}
   );
   gpc1_1 gpc2611 (
      {stage0_10[400]},
      {stage1_10[199]}
   );
   gpc1_1 gpc2612 (
      {stage0_10[401]},
      {stage1_10[200]}
   );
   gpc1_1 gpc2613 (
      {stage0_10[402]},
      {stage1_10[201]}
   );
   gpc1_1 gpc2614 (
      {stage0_10[403]},
      {stage1_10[202]}
   );
   gpc1_1 gpc2615 (
      {stage0_10[404]},
      {stage1_10[203]}
   );
   gpc1_1 gpc2616 (
      {stage0_10[405]},
      {stage1_10[204]}
   );
   gpc1_1 gpc2617 (
      {stage0_10[406]},
      {stage1_10[205]}
   );
   gpc1_1 gpc2618 (
      {stage0_10[407]},
      {stage1_10[206]}
   );
   gpc1_1 gpc2619 (
      {stage0_10[408]},
      {stage1_10[207]}
   );
   gpc1_1 gpc2620 (
      {stage0_10[409]},
      {stage1_10[208]}
   );
   gpc1_1 gpc2621 (
      {stage0_10[410]},
      {stage1_10[209]}
   );
   gpc1_1 gpc2622 (
      {stage0_10[411]},
      {stage1_10[210]}
   );
   gpc1_1 gpc2623 (
      {stage0_10[412]},
      {stage1_10[211]}
   );
   gpc1_1 gpc2624 (
      {stage0_10[413]},
      {stage1_10[212]}
   );
   gpc1_1 gpc2625 (
      {stage0_10[414]},
      {stage1_10[213]}
   );
   gpc1_1 gpc2626 (
      {stage0_10[415]},
      {stage1_10[214]}
   );
   gpc1_1 gpc2627 (
      {stage0_10[416]},
      {stage1_10[215]}
   );
   gpc1_1 gpc2628 (
      {stage0_10[417]},
      {stage1_10[216]}
   );
   gpc1_1 gpc2629 (
      {stage0_10[418]},
      {stage1_10[217]}
   );
   gpc1_1 gpc2630 (
      {stage0_10[419]},
      {stage1_10[218]}
   );
   gpc1_1 gpc2631 (
      {stage0_10[420]},
      {stage1_10[219]}
   );
   gpc1_1 gpc2632 (
      {stage0_10[421]},
      {stage1_10[220]}
   );
   gpc1_1 gpc2633 (
      {stage0_10[422]},
      {stage1_10[221]}
   );
   gpc1_1 gpc2634 (
      {stage0_10[423]},
      {stage1_10[222]}
   );
   gpc1_1 gpc2635 (
      {stage0_10[424]},
      {stage1_10[223]}
   );
   gpc1_1 gpc2636 (
      {stage0_10[425]},
      {stage1_10[224]}
   );
   gpc1_1 gpc2637 (
      {stage0_10[426]},
      {stage1_10[225]}
   );
   gpc1_1 gpc2638 (
      {stage0_10[427]},
      {stage1_10[226]}
   );
   gpc1_1 gpc2639 (
      {stage0_10[428]},
      {stage1_10[227]}
   );
   gpc1_1 gpc2640 (
      {stage0_10[429]},
      {stage1_10[228]}
   );
   gpc1_1 gpc2641 (
      {stage0_10[430]},
      {stage1_10[229]}
   );
   gpc1_1 gpc2642 (
      {stage0_10[431]},
      {stage1_10[230]}
   );
   gpc1_1 gpc2643 (
      {stage0_10[432]},
      {stage1_10[231]}
   );
   gpc1_1 gpc2644 (
      {stage0_10[433]},
      {stage1_10[232]}
   );
   gpc1_1 gpc2645 (
      {stage0_10[434]},
      {stage1_10[233]}
   );
   gpc1_1 gpc2646 (
      {stage0_10[435]},
      {stage1_10[234]}
   );
   gpc1_1 gpc2647 (
      {stage0_10[436]},
      {stage1_10[235]}
   );
   gpc1_1 gpc2648 (
      {stage0_10[437]},
      {stage1_10[236]}
   );
   gpc1_1 gpc2649 (
      {stage0_10[438]},
      {stage1_10[237]}
   );
   gpc1_1 gpc2650 (
      {stage0_10[439]},
      {stage1_10[238]}
   );
   gpc1_1 gpc2651 (
      {stage0_10[440]},
      {stage1_10[239]}
   );
   gpc1_1 gpc2652 (
      {stage0_10[441]},
      {stage1_10[240]}
   );
   gpc1_1 gpc2653 (
      {stage0_10[442]},
      {stage1_10[241]}
   );
   gpc1_1 gpc2654 (
      {stage0_10[443]},
      {stage1_10[242]}
   );
   gpc1_1 gpc2655 (
      {stage0_10[444]},
      {stage1_10[243]}
   );
   gpc1_1 gpc2656 (
      {stage0_10[445]},
      {stage1_10[244]}
   );
   gpc1_1 gpc2657 (
      {stage0_10[446]},
      {stage1_10[245]}
   );
   gpc1_1 gpc2658 (
      {stage0_10[447]},
      {stage1_10[246]}
   );
   gpc1_1 gpc2659 (
      {stage0_10[448]},
      {stage1_10[247]}
   );
   gpc1_1 gpc2660 (
      {stage0_10[449]},
      {stage1_10[248]}
   );
   gpc1_1 gpc2661 (
      {stage0_10[450]},
      {stage1_10[249]}
   );
   gpc1_1 gpc2662 (
      {stage0_10[451]},
      {stage1_10[250]}
   );
   gpc1_1 gpc2663 (
      {stage0_10[452]},
      {stage1_10[251]}
   );
   gpc1_1 gpc2664 (
      {stage0_10[453]},
      {stage1_10[252]}
   );
   gpc1_1 gpc2665 (
      {stage0_10[454]},
      {stage1_10[253]}
   );
   gpc1_1 gpc2666 (
      {stage0_10[455]},
      {stage1_10[254]}
   );
   gpc1_1 gpc2667 (
      {stage0_10[456]},
      {stage1_10[255]}
   );
   gpc1_1 gpc2668 (
      {stage0_10[457]},
      {stage1_10[256]}
   );
   gpc1_1 gpc2669 (
      {stage0_10[458]},
      {stage1_10[257]}
   );
   gpc1_1 gpc2670 (
      {stage0_10[459]},
      {stage1_10[258]}
   );
   gpc1_1 gpc2671 (
      {stage0_10[460]},
      {stage1_10[259]}
   );
   gpc1_1 gpc2672 (
      {stage0_10[461]},
      {stage1_10[260]}
   );
   gpc1_1 gpc2673 (
      {stage0_10[462]},
      {stage1_10[261]}
   );
   gpc1_1 gpc2674 (
      {stage0_10[463]},
      {stage1_10[262]}
   );
   gpc1_1 gpc2675 (
      {stage0_10[464]},
      {stage1_10[263]}
   );
   gpc1_1 gpc2676 (
      {stage0_10[465]},
      {stage1_10[264]}
   );
   gpc1_1 gpc2677 (
      {stage0_10[466]},
      {stage1_10[265]}
   );
   gpc1_1 gpc2678 (
      {stage0_10[467]},
      {stage1_10[266]}
   );
   gpc1_1 gpc2679 (
      {stage0_10[468]},
      {stage1_10[267]}
   );
   gpc1_1 gpc2680 (
      {stage0_10[469]},
      {stage1_10[268]}
   );
   gpc1_1 gpc2681 (
      {stage0_10[470]},
      {stage1_10[269]}
   );
   gpc1_1 gpc2682 (
      {stage0_10[471]},
      {stage1_10[270]}
   );
   gpc1_1 gpc2683 (
      {stage0_10[472]},
      {stage1_10[271]}
   );
   gpc1_1 gpc2684 (
      {stage0_10[473]},
      {stage1_10[272]}
   );
   gpc1_1 gpc2685 (
      {stage0_10[474]},
      {stage1_10[273]}
   );
   gpc1_1 gpc2686 (
      {stage0_10[475]},
      {stage1_10[274]}
   );
   gpc1_1 gpc2687 (
      {stage0_10[476]},
      {stage1_10[275]}
   );
   gpc1_1 gpc2688 (
      {stage0_10[477]},
      {stage1_10[276]}
   );
   gpc1_1 gpc2689 (
      {stage0_10[478]},
      {stage1_10[277]}
   );
   gpc1_1 gpc2690 (
      {stage0_10[479]},
      {stage1_10[278]}
   );
   gpc1_1 gpc2691 (
      {stage0_10[480]},
      {stage1_10[279]}
   );
   gpc1_1 gpc2692 (
      {stage0_10[481]},
      {stage1_10[280]}
   );
   gpc1_1 gpc2693 (
      {stage0_10[482]},
      {stage1_10[281]}
   );
   gpc1_1 gpc2694 (
      {stage0_10[483]},
      {stage1_10[282]}
   );
   gpc1_1 gpc2695 (
      {stage0_10[484]},
      {stage1_10[283]}
   );
   gpc1_1 gpc2696 (
      {stage0_10[485]},
      {stage1_10[284]}
   );
   gpc1_1 gpc2697 (
      {stage0_11[367]},
      {stage1_11[158]}
   );
   gpc1_1 gpc2698 (
      {stage0_11[368]},
      {stage1_11[159]}
   );
   gpc1_1 gpc2699 (
      {stage0_11[369]},
      {stage1_11[160]}
   );
   gpc1_1 gpc2700 (
      {stage0_11[370]},
      {stage1_11[161]}
   );
   gpc1_1 gpc2701 (
      {stage0_11[371]},
      {stage1_11[162]}
   );
   gpc1_1 gpc2702 (
      {stage0_11[372]},
      {stage1_11[163]}
   );
   gpc1_1 gpc2703 (
      {stage0_11[373]},
      {stage1_11[164]}
   );
   gpc1_1 gpc2704 (
      {stage0_11[374]},
      {stage1_11[165]}
   );
   gpc1_1 gpc2705 (
      {stage0_11[375]},
      {stage1_11[166]}
   );
   gpc1_1 gpc2706 (
      {stage0_11[376]},
      {stage1_11[167]}
   );
   gpc1_1 gpc2707 (
      {stage0_11[377]},
      {stage1_11[168]}
   );
   gpc1_1 gpc2708 (
      {stage0_11[378]},
      {stage1_11[169]}
   );
   gpc1_1 gpc2709 (
      {stage0_11[379]},
      {stage1_11[170]}
   );
   gpc1_1 gpc2710 (
      {stage0_11[380]},
      {stage1_11[171]}
   );
   gpc1_1 gpc2711 (
      {stage0_11[381]},
      {stage1_11[172]}
   );
   gpc1_1 gpc2712 (
      {stage0_11[382]},
      {stage1_11[173]}
   );
   gpc1_1 gpc2713 (
      {stage0_11[383]},
      {stage1_11[174]}
   );
   gpc1_1 gpc2714 (
      {stage0_11[384]},
      {stage1_11[175]}
   );
   gpc1_1 gpc2715 (
      {stage0_11[385]},
      {stage1_11[176]}
   );
   gpc1_1 gpc2716 (
      {stage0_11[386]},
      {stage1_11[177]}
   );
   gpc1_1 gpc2717 (
      {stage0_11[387]},
      {stage1_11[178]}
   );
   gpc1_1 gpc2718 (
      {stage0_11[388]},
      {stage1_11[179]}
   );
   gpc1_1 gpc2719 (
      {stage0_11[389]},
      {stage1_11[180]}
   );
   gpc1_1 gpc2720 (
      {stage0_11[390]},
      {stage1_11[181]}
   );
   gpc1_1 gpc2721 (
      {stage0_11[391]},
      {stage1_11[182]}
   );
   gpc1_1 gpc2722 (
      {stage0_11[392]},
      {stage1_11[183]}
   );
   gpc1_1 gpc2723 (
      {stage0_11[393]},
      {stage1_11[184]}
   );
   gpc1_1 gpc2724 (
      {stage0_11[394]},
      {stage1_11[185]}
   );
   gpc1_1 gpc2725 (
      {stage0_11[395]},
      {stage1_11[186]}
   );
   gpc1_1 gpc2726 (
      {stage0_11[396]},
      {stage1_11[187]}
   );
   gpc1_1 gpc2727 (
      {stage0_11[397]},
      {stage1_11[188]}
   );
   gpc1_1 gpc2728 (
      {stage0_11[398]},
      {stage1_11[189]}
   );
   gpc1_1 gpc2729 (
      {stage0_11[399]},
      {stage1_11[190]}
   );
   gpc1_1 gpc2730 (
      {stage0_11[400]},
      {stage1_11[191]}
   );
   gpc1_1 gpc2731 (
      {stage0_11[401]},
      {stage1_11[192]}
   );
   gpc1_1 gpc2732 (
      {stage0_11[402]},
      {stage1_11[193]}
   );
   gpc1_1 gpc2733 (
      {stage0_11[403]},
      {stage1_11[194]}
   );
   gpc1_1 gpc2734 (
      {stage0_11[404]},
      {stage1_11[195]}
   );
   gpc1_1 gpc2735 (
      {stage0_11[405]},
      {stage1_11[196]}
   );
   gpc1_1 gpc2736 (
      {stage0_11[406]},
      {stage1_11[197]}
   );
   gpc1_1 gpc2737 (
      {stage0_11[407]},
      {stage1_11[198]}
   );
   gpc1_1 gpc2738 (
      {stage0_11[408]},
      {stage1_11[199]}
   );
   gpc1_1 gpc2739 (
      {stage0_11[409]},
      {stage1_11[200]}
   );
   gpc1_1 gpc2740 (
      {stage0_11[410]},
      {stage1_11[201]}
   );
   gpc1_1 gpc2741 (
      {stage0_11[411]},
      {stage1_11[202]}
   );
   gpc1_1 gpc2742 (
      {stage0_11[412]},
      {stage1_11[203]}
   );
   gpc1_1 gpc2743 (
      {stage0_11[413]},
      {stage1_11[204]}
   );
   gpc1_1 gpc2744 (
      {stage0_11[414]},
      {stage1_11[205]}
   );
   gpc1_1 gpc2745 (
      {stage0_11[415]},
      {stage1_11[206]}
   );
   gpc1_1 gpc2746 (
      {stage0_11[416]},
      {stage1_11[207]}
   );
   gpc1_1 gpc2747 (
      {stage0_11[417]},
      {stage1_11[208]}
   );
   gpc1_1 gpc2748 (
      {stage0_11[418]},
      {stage1_11[209]}
   );
   gpc1_1 gpc2749 (
      {stage0_11[419]},
      {stage1_11[210]}
   );
   gpc1_1 gpc2750 (
      {stage0_11[420]},
      {stage1_11[211]}
   );
   gpc1_1 gpc2751 (
      {stage0_11[421]},
      {stage1_11[212]}
   );
   gpc1_1 gpc2752 (
      {stage0_11[422]},
      {stage1_11[213]}
   );
   gpc1_1 gpc2753 (
      {stage0_11[423]},
      {stage1_11[214]}
   );
   gpc1_1 gpc2754 (
      {stage0_11[424]},
      {stage1_11[215]}
   );
   gpc1_1 gpc2755 (
      {stage0_11[425]},
      {stage1_11[216]}
   );
   gpc1_1 gpc2756 (
      {stage0_11[426]},
      {stage1_11[217]}
   );
   gpc1_1 gpc2757 (
      {stage0_11[427]},
      {stage1_11[218]}
   );
   gpc1_1 gpc2758 (
      {stage0_11[428]},
      {stage1_11[219]}
   );
   gpc1_1 gpc2759 (
      {stage0_11[429]},
      {stage1_11[220]}
   );
   gpc1_1 gpc2760 (
      {stage0_11[430]},
      {stage1_11[221]}
   );
   gpc1_1 gpc2761 (
      {stage0_11[431]},
      {stage1_11[222]}
   );
   gpc1_1 gpc2762 (
      {stage0_11[432]},
      {stage1_11[223]}
   );
   gpc1_1 gpc2763 (
      {stage0_11[433]},
      {stage1_11[224]}
   );
   gpc1_1 gpc2764 (
      {stage0_11[434]},
      {stage1_11[225]}
   );
   gpc1_1 gpc2765 (
      {stage0_11[435]},
      {stage1_11[226]}
   );
   gpc1_1 gpc2766 (
      {stage0_11[436]},
      {stage1_11[227]}
   );
   gpc1_1 gpc2767 (
      {stage0_11[437]},
      {stage1_11[228]}
   );
   gpc1_1 gpc2768 (
      {stage0_11[438]},
      {stage1_11[229]}
   );
   gpc1_1 gpc2769 (
      {stage0_11[439]},
      {stage1_11[230]}
   );
   gpc1_1 gpc2770 (
      {stage0_11[440]},
      {stage1_11[231]}
   );
   gpc1_1 gpc2771 (
      {stage0_11[441]},
      {stage1_11[232]}
   );
   gpc1_1 gpc2772 (
      {stage0_11[442]},
      {stage1_11[233]}
   );
   gpc1_1 gpc2773 (
      {stage0_11[443]},
      {stage1_11[234]}
   );
   gpc1_1 gpc2774 (
      {stage0_11[444]},
      {stage1_11[235]}
   );
   gpc1_1 gpc2775 (
      {stage0_11[445]},
      {stage1_11[236]}
   );
   gpc1_1 gpc2776 (
      {stage0_11[446]},
      {stage1_11[237]}
   );
   gpc1_1 gpc2777 (
      {stage0_11[447]},
      {stage1_11[238]}
   );
   gpc1_1 gpc2778 (
      {stage0_11[448]},
      {stage1_11[239]}
   );
   gpc1_1 gpc2779 (
      {stage0_11[449]},
      {stage1_11[240]}
   );
   gpc1_1 gpc2780 (
      {stage0_11[450]},
      {stage1_11[241]}
   );
   gpc1_1 gpc2781 (
      {stage0_11[451]},
      {stage1_11[242]}
   );
   gpc1_1 gpc2782 (
      {stage0_11[452]},
      {stage1_11[243]}
   );
   gpc1_1 gpc2783 (
      {stage0_11[453]},
      {stage1_11[244]}
   );
   gpc1_1 gpc2784 (
      {stage0_11[454]},
      {stage1_11[245]}
   );
   gpc1_1 gpc2785 (
      {stage0_11[455]},
      {stage1_11[246]}
   );
   gpc1_1 gpc2786 (
      {stage0_11[456]},
      {stage1_11[247]}
   );
   gpc1_1 gpc2787 (
      {stage0_11[457]},
      {stage1_11[248]}
   );
   gpc1_1 gpc2788 (
      {stage0_11[458]},
      {stage1_11[249]}
   );
   gpc1_1 gpc2789 (
      {stage0_11[459]},
      {stage1_11[250]}
   );
   gpc1_1 gpc2790 (
      {stage0_11[460]},
      {stage1_11[251]}
   );
   gpc1_1 gpc2791 (
      {stage0_11[461]},
      {stage1_11[252]}
   );
   gpc1_1 gpc2792 (
      {stage0_11[462]},
      {stage1_11[253]}
   );
   gpc1_1 gpc2793 (
      {stage0_11[463]},
      {stage1_11[254]}
   );
   gpc1_1 gpc2794 (
      {stage0_11[464]},
      {stage1_11[255]}
   );
   gpc1_1 gpc2795 (
      {stage0_11[465]},
      {stage1_11[256]}
   );
   gpc1_1 gpc2796 (
      {stage0_11[466]},
      {stage1_11[257]}
   );
   gpc1_1 gpc2797 (
      {stage0_11[467]},
      {stage1_11[258]}
   );
   gpc1_1 gpc2798 (
      {stage0_11[468]},
      {stage1_11[259]}
   );
   gpc1_1 gpc2799 (
      {stage0_11[469]},
      {stage1_11[260]}
   );
   gpc1_1 gpc2800 (
      {stage0_11[470]},
      {stage1_11[261]}
   );
   gpc1_1 gpc2801 (
      {stage0_11[471]},
      {stage1_11[262]}
   );
   gpc1_1 gpc2802 (
      {stage0_11[472]},
      {stage1_11[263]}
   );
   gpc1_1 gpc2803 (
      {stage0_11[473]},
      {stage1_11[264]}
   );
   gpc1_1 gpc2804 (
      {stage0_11[474]},
      {stage1_11[265]}
   );
   gpc1_1 gpc2805 (
      {stage0_11[475]},
      {stage1_11[266]}
   );
   gpc1_1 gpc2806 (
      {stage0_11[476]},
      {stage1_11[267]}
   );
   gpc1_1 gpc2807 (
      {stage0_11[477]},
      {stage1_11[268]}
   );
   gpc1_1 gpc2808 (
      {stage0_11[478]},
      {stage1_11[269]}
   );
   gpc1_1 gpc2809 (
      {stage0_11[479]},
      {stage1_11[270]}
   );
   gpc1_1 gpc2810 (
      {stage0_11[480]},
      {stage1_11[271]}
   );
   gpc1_1 gpc2811 (
      {stage0_11[481]},
      {stage1_11[272]}
   );
   gpc1_1 gpc2812 (
      {stage0_11[482]},
      {stage1_11[273]}
   );
   gpc1_1 gpc2813 (
      {stage0_11[483]},
      {stage1_11[274]}
   );
   gpc1_1 gpc2814 (
      {stage0_11[484]},
      {stage1_11[275]}
   );
   gpc1_1 gpc2815 (
      {stage0_11[485]},
      {stage1_11[276]}
   );
   gpc1_1 gpc2816 (
      {stage0_12[484]},
      {stage1_12[187]}
   );
   gpc1_1 gpc2817 (
      {stage0_12[485]},
      {stage1_12[188]}
   );
   gpc1_1 gpc2818 (
      {stage0_13[376]},
      {stage1_13[195]}
   );
   gpc1_1 gpc2819 (
      {stage0_13[377]},
      {stage1_13[196]}
   );
   gpc1_1 gpc2820 (
      {stage0_13[378]},
      {stage1_13[197]}
   );
   gpc1_1 gpc2821 (
      {stage0_13[379]},
      {stage1_13[198]}
   );
   gpc1_1 gpc2822 (
      {stage0_13[380]},
      {stage1_13[199]}
   );
   gpc1_1 gpc2823 (
      {stage0_13[381]},
      {stage1_13[200]}
   );
   gpc1_1 gpc2824 (
      {stage0_13[382]},
      {stage1_13[201]}
   );
   gpc1_1 gpc2825 (
      {stage0_13[383]},
      {stage1_13[202]}
   );
   gpc1_1 gpc2826 (
      {stage0_13[384]},
      {stage1_13[203]}
   );
   gpc1_1 gpc2827 (
      {stage0_13[385]},
      {stage1_13[204]}
   );
   gpc1_1 gpc2828 (
      {stage0_13[386]},
      {stage1_13[205]}
   );
   gpc1_1 gpc2829 (
      {stage0_13[387]},
      {stage1_13[206]}
   );
   gpc1_1 gpc2830 (
      {stage0_13[388]},
      {stage1_13[207]}
   );
   gpc1_1 gpc2831 (
      {stage0_13[389]},
      {stage1_13[208]}
   );
   gpc1_1 gpc2832 (
      {stage0_13[390]},
      {stage1_13[209]}
   );
   gpc1_1 gpc2833 (
      {stage0_13[391]},
      {stage1_13[210]}
   );
   gpc1_1 gpc2834 (
      {stage0_13[392]},
      {stage1_13[211]}
   );
   gpc1_1 gpc2835 (
      {stage0_13[393]},
      {stage1_13[212]}
   );
   gpc1_1 gpc2836 (
      {stage0_13[394]},
      {stage1_13[213]}
   );
   gpc1_1 gpc2837 (
      {stage0_13[395]},
      {stage1_13[214]}
   );
   gpc1_1 gpc2838 (
      {stage0_13[396]},
      {stage1_13[215]}
   );
   gpc1_1 gpc2839 (
      {stage0_13[397]},
      {stage1_13[216]}
   );
   gpc1_1 gpc2840 (
      {stage0_13[398]},
      {stage1_13[217]}
   );
   gpc1_1 gpc2841 (
      {stage0_13[399]},
      {stage1_13[218]}
   );
   gpc1_1 gpc2842 (
      {stage0_13[400]},
      {stage1_13[219]}
   );
   gpc1_1 gpc2843 (
      {stage0_13[401]},
      {stage1_13[220]}
   );
   gpc1_1 gpc2844 (
      {stage0_13[402]},
      {stage1_13[221]}
   );
   gpc1_1 gpc2845 (
      {stage0_13[403]},
      {stage1_13[222]}
   );
   gpc1_1 gpc2846 (
      {stage0_13[404]},
      {stage1_13[223]}
   );
   gpc1_1 gpc2847 (
      {stage0_13[405]},
      {stage1_13[224]}
   );
   gpc1_1 gpc2848 (
      {stage0_13[406]},
      {stage1_13[225]}
   );
   gpc1_1 gpc2849 (
      {stage0_13[407]},
      {stage1_13[226]}
   );
   gpc1_1 gpc2850 (
      {stage0_13[408]},
      {stage1_13[227]}
   );
   gpc1_1 gpc2851 (
      {stage0_13[409]},
      {stage1_13[228]}
   );
   gpc1_1 gpc2852 (
      {stage0_13[410]},
      {stage1_13[229]}
   );
   gpc1_1 gpc2853 (
      {stage0_13[411]},
      {stage1_13[230]}
   );
   gpc1_1 gpc2854 (
      {stage0_13[412]},
      {stage1_13[231]}
   );
   gpc1_1 gpc2855 (
      {stage0_13[413]},
      {stage1_13[232]}
   );
   gpc1_1 gpc2856 (
      {stage0_13[414]},
      {stage1_13[233]}
   );
   gpc1_1 gpc2857 (
      {stage0_13[415]},
      {stage1_13[234]}
   );
   gpc1_1 gpc2858 (
      {stage0_13[416]},
      {stage1_13[235]}
   );
   gpc1_1 gpc2859 (
      {stage0_13[417]},
      {stage1_13[236]}
   );
   gpc1_1 gpc2860 (
      {stage0_13[418]},
      {stage1_13[237]}
   );
   gpc1_1 gpc2861 (
      {stage0_13[419]},
      {stage1_13[238]}
   );
   gpc1_1 gpc2862 (
      {stage0_13[420]},
      {stage1_13[239]}
   );
   gpc1_1 gpc2863 (
      {stage0_13[421]},
      {stage1_13[240]}
   );
   gpc1_1 gpc2864 (
      {stage0_13[422]},
      {stage1_13[241]}
   );
   gpc1_1 gpc2865 (
      {stage0_13[423]},
      {stage1_13[242]}
   );
   gpc1_1 gpc2866 (
      {stage0_13[424]},
      {stage1_13[243]}
   );
   gpc1_1 gpc2867 (
      {stage0_13[425]},
      {stage1_13[244]}
   );
   gpc1_1 gpc2868 (
      {stage0_13[426]},
      {stage1_13[245]}
   );
   gpc1_1 gpc2869 (
      {stage0_13[427]},
      {stage1_13[246]}
   );
   gpc1_1 gpc2870 (
      {stage0_13[428]},
      {stage1_13[247]}
   );
   gpc1_1 gpc2871 (
      {stage0_13[429]},
      {stage1_13[248]}
   );
   gpc1_1 gpc2872 (
      {stage0_13[430]},
      {stage1_13[249]}
   );
   gpc1_1 gpc2873 (
      {stage0_13[431]},
      {stage1_13[250]}
   );
   gpc1_1 gpc2874 (
      {stage0_13[432]},
      {stage1_13[251]}
   );
   gpc1_1 gpc2875 (
      {stage0_13[433]},
      {stage1_13[252]}
   );
   gpc1_1 gpc2876 (
      {stage0_13[434]},
      {stage1_13[253]}
   );
   gpc1_1 gpc2877 (
      {stage0_13[435]},
      {stage1_13[254]}
   );
   gpc1_1 gpc2878 (
      {stage0_13[436]},
      {stage1_13[255]}
   );
   gpc1_1 gpc2879 (
      {stage0_13[437]},
      {stage1_13[256]}
   );
   gpc1_1 gpc2880 (
      {stage0_13[438]},
      {stage1_13[257]}
   );
   gpc1_1 gpc2881 (
      {stage0_13[439]},
      {stage1_13[258]}
   );
   gpc1_1 gpc2882 (
      {stage0_13[440]},
      {stage1_13[259]}
   );
   gpc1_1 gpc2883 (
      {stage0_13[441]},
      {stage1_13[260]}
   );
   gpc1_1 gpc2884 (
      {stage0_13[442]},
      {stage1_13[261]}
   );
   gpc1_1 gpc2885 (
      {stage0_13[443]},
      {stage1_13[262]}
   );
   gpc1_1 gpc2886 (
      {stage0_13[444]},
      {stage1_13[263]}
   );
   gpc1_1 gpc2887 (
      {stage0_13[445]},
      {stage1_13[264]}
   );
   gpc1_1 gpc2888 (
      {stage0_13[446]},
      {stage1_13[265]}
   );
   gpc1_1 gpc2889 (
      {stage0_13[447]},
      {stage1_13[266]}
   );
   gpc1_1 gpc2890 (
      {stage0_13[448]},
      {stage1_13[267]}
   );
   gpc1_1 gpc2891 (
      {stage0_13[449]},
      {stage1_13[268]}
   );
   gpc1_1 gpc2892 (
      {stage0_13[450]},
      {stage1_13[269]}
   );
   gpc1_1 gpc2893 (
      {stage0_13[451]},
      {stage1_13[270]}
   );
   gpc1_1 gpc2894 (
      {stage0_13[452]},
      {stage1_13[271]}
   );
   gpc1_1 gpc2895 (
      {stage0_13[453]},
      {stage1_13[272]}
   );
   gpc1_1 gpc2896 (
      {stage0_13[454]},
      {stage1_13[273]}
   );
   gpc1_1 gpc2897 (
      {stage0_13[455]},
      {stage1_13[274]}
   );
   gpc1_1 gpc2898 (
      {stage0_13[456]},
      {stage1_13[275]}
   );
   gpc1_1 gpc2899 (
      {stage0_13[457]},
      {stage1_13[276]}
   );
   gpc1_1 gpc2900 (
      {stage0_13[458]},
      {stage1_13[277]}
   );
   gpc1_1 gpc2901 (
      {stage0_13[459]},
      {stage1_13[278]}
   );
   gpc1_1 gpc2902 (
      {stage0_13[460]},
      {stage1_13[279]}
   );
   gpc1_1 gpc2903 (
      {stage0_13[461]},
      {stage1_13[280]}
   );
   gpc1_1 gpc2904 (
      {stage0_13[462]},
      {stage1_13[281]}
   );
   gpc1_1 gpc2905 (
      {stage0_13[463]},
      {stage1_13[282]}
   );
   gpc1_1 gpc2906 (
      {stage0_13[464]},
      {stage1_13[283]}
   );
   gpc1_1 gpc2907 (
      {stage0_13[465]},
      {stage1_13[284]}
   );
   gpc1_1 gpc2908 (
      {stage0_13[466]},
      {stage1_13[285]}
   );
   gpc1_1 gpc2909 (
      {stage0_13[467]},
      {stage1_13[286]}
   );
   gpc1_1 gpc2910 (
      {stage0_13[468]},
      {stage1_13[287]}
   );
   gpc1_1 gpc2911 (
      {stage0_13[469]},
      {stage1_13[288]}
   );
   gpc1_1 gpc2912 (
      {stage0_13[470]},
      {stage1_13[289]}
   );
   gpc1_1 gpc2913 (
      {stage0_13[471]},
      {stage1_13[290]}
   );
   gpc1_1 gpc2914 (
      {stage0_13[472]},
      {stage1_13[291]}
   );
   gpc1_1 gpc2915 (
      {stage0_13[473]},
      {stage1_13[292]}
   );
   gpc1_1 gpc2916 (
      {stage0_13[474]},
      {stage1_13[293]}
   );
   gpc1_1 gpc2917 (
      {stage0_13[475]},
      {stage1_13[294]}
   );
   gpc1_1 gpc2918 (
      {stage0_13[476]},
      {stage1_13[295]}
   );
   gpc1_1 gpc2919 (
      {stage0_13[477]},
      {stage1_13[296]}
   );
   gpc1_1 gpc2920 (
      {stage0_13[478]},
      {stage1_13[297]}
   );
   gpc1_1 gpc2921 (
      {stage0_13[479]},
      {stage1_13[298]}
   );
   gpc1_1 gpc2922 (
      {stage0_13[480]},
      {stage1_13[299]}
   );
   gpc1_1 gpc2923 (
      {stage0_13[481]},
      {stage1_13[300]}
   );
   gpc1_1 gpc2924 (
      {stage0_13[482]},
      {stage1_13[301]}
   );
   gpc1_1 gpc2925 (
      {stage0_13[483]},
      {stage1_13[302]}
   );
   gpc1_1 gpc2926 (
      {stage0_13[484]},
      {stage1_13[303]}
   );
   gpc1_1 gpc2927 (
      {stage0_13[485]},
      {stage1_13[304]}
   );
   gpc1_1 gpc2928 (
      {stage0_14[419]},
      {stage1_14[152]}
   );
   gpc1_1 gpc2929 (
      {stage0_14[420]},
      {stage1_14[153]}
   );
   gpc1_1 gpc2930 (
      {stage0_14[421]},
      {stage1_14[154]}
   );
   gpc1_1 gpc2931 (
      {stage0_14[422]},
      {stage1_14[155]}
   );
   gpc1_1 gpc2932 (
      {stage0_14[423]},
      {stage1_14[156]}
   );
   gpc1_1 gpc2933 (
      {stage0_14[424]},
      {stage1_14[157]}
   );
   gpc1_1 gpc2934 (
      {stage0_14[425]},
      {stage1_14[158]}
   );
   gpc1_1 gpc2935 (
      {stage0_14[426]},
      {stage1_14[159]}
   );
   gpc1_1 gpc2936 (
      {stage0_14[427]},
      {stage1_14[160]}
   );
   gpc1_1 gpc2937 (
      {stage0_14[428]},
      {stage1_14[161]}
   );
   gpc1_1 gpc2938 (
      {stage0_14[429]},
      {stage1_14[162]}
   );
   gpc1_1 gpc2939 (
      {stage0_14[430]},
      {stage1_14[163]}
   );
   gpc1_1 gpc2940 (
      {stage0_14[431]},
      {stage1_14[164]}
   );
   gpc1_1 gpc2941 (
      {stage0_14[432]},
      {stage1_14[165]}
   );
   gpc1_1 gpc2942 (
      {stage0_14[433]},
      {stage1_14[166]}
   );
   gpc1_1 gpc2943 (
      {stage0_14[434]},
      {stage1_14[167]}
   );
   gpc1_1 gpc2944 (
      {stage0_14[435]},
      {stage1_14[168]}
   );
   gpc1_1 gpc2945 (
      {stage0_14[436]},
      {stage1_14[169]}
   );
   gpc1_1 gpc2946 (
      {stage0_14[437]},
      {stage1_14[170]}
   );
   gpc1_1 gpc2947 (
      {stage0_14[438]},
      {stage1_14[171]}
   );
   gpc1_1 gpc2948 (
      {stage0_14[439]},
      {stage1_14[172]}
   );
   gpc1_1 gpc2949 (
      {stage0_14[440]},
      {stage1_14[173]}
   );
   gpc1_1 gpc2950 (
      {stage0_14[441]},
      {stage1_14[174]}
   );
   gpc1_1 gpc2951 (
      {stage0_14[442]},
      {stage1_14[175]}
   );
   gpc1_1 gpc2952 (
      {stage0_14[443]},
      {stage1_14[176]}
   );
   gpc1_1 gpc2953 (
      {stage0_14[444]},
      {stage1_14[177]}
   );
   gpc1_1 gpc2954 (
      {stage0_14[445]},
      {stage1_14[178]}
   );
   gpc1_1 gpc2955 (
      {stage0_14[446]},
      {stage1_14[179]}
   );
   gpc1_1 gpc2956 (
      {stage0_14[447]},
      {stage1_14[180]}
   );
   gpc1_1 gpc2957 (
      {stage0_14[448]},
      {stage1_14[181]}
   );
   gpc1_1 gpc2958 (
      {stage0_14[449]},
      {stage1_14[182]}
   );
   gpc1_1 gpc2959 (
      {stage0_14[450]},
      {stage1_14[183]}
   );
   gpc1_1 gpc2960 (
      {stage0_14[451]},
      {stage1_14[184]}
   );
   gpc1_1 gpc2961 (
      {stage0_14[452]},
      {stage1_14[185]}
   );
   gpc1_1 gpc2962 (
      {stage0_14[453]},
      {stage1_14[186]}
   );
   gpc1_1 gpc2963 (
      {stage0_14[454]},
      {stage1_14[187]}
   );
   gpc1_1 gpc2964 (
      {stage0_14[455]},
      {stage1_14[188]}
   );
   gpc1_1 gpc2965 (
      {stage0_14[456]},
      {stage1_14[189]}
   );
   gpc1_1 gpc2966 (
      {stage0_14[457]},
      {stage1_14[190]}
   );
   gpc1_1 gpc2967 (
      {stage0_14[458]},
      {stage1_14[191]}
   );
   gpc1_1 gpc2968 (
      {stage0_14[459]},
      {stage1_14[192]}
   );
   gpc1_1 gpc2969 (
      {stage0_14[460]},
      {stage1_14[193]}
   );
   gpc1_1 gpc2970 (
      {stage0_14[461]},
      {stage1_14[194]}
   );
   gpc1_1 gpc2971 (
      {stage0_14[462]},
      {stage1_14[195]}
   );
   gpc1_1 gpc2972 (
      {stage0_14[463]},
      {stage1_14[196]}
   );
   gpc1_1 gpc2973 (
      {stage0_14[464]},
      {stage1_14[197]}
   );
   gpc1_1 gpc2974 (
      {stage0_14[465]},
      {stage1_14[198]}
   );
   gpc1_1 gpc2975 (
      {stage0_14[466]},
      {stage1_14[199]}
   );
   gpc1_1 gpc2976 (
      {stage0_14[467]},
      {stage1_14[200]}
   );
   gpc1_1 gpc2977 (
      {stage0_14[468]},
      {stage1_14[201]}
   );
   gpc1_1 gpc2978 (
      {stage0_14[469]},
      {stage1_14[202]}
   );
   gpc1_1 gpc2979 (
      {stage0_14[470]},
      {stage1_14[203]}
   );
   gpc1_1 gpc2980 (
      {stage0_14[471]},
      {stage1_14[204]}
   );
   gpc1_1 gpc2981 (
      {stage0_14[472]},
      {stage1_14[205]}
   );
   gpc1_1 gpc2982 (
      {stage0_14[473]},
      {stage1_14[206]}
   );
   gpc1_1 gpc2983 (
      {stage0_14[474]},
      {stage1_14[207]}
   );
   gpc1_1 gpc2984 (
      {stage0_14[475]},
      {stage1_14[208]}
   );
   gpc1_1 gpc2985 (
      {stage0_14[476]},
      {stage1_14[209]}
   );
   gpc1_1 gpc2986 (
      {stage0_14[477]},
      {stage1_14[210]}
   );
   gpc1_1 gpc2987 (
      {stage0_14[478]},
      {stage1_14[211]}
   );
   gpc1_1 gpc2988 (
      {stage0_14[479]},
      {stage1_14[212]}
   );
   gpc1_1 gpc2989 (
      {stage0_14[480]},
      {stage1_14[213]}
   );
   gpc1_1 gpc2990 (
      {stage0_14[481]},
      {stage1_14[214]}
   );
   gpc1_1 gpc2991 (
      {stage0_14[482]},
      {stage1_14[215]}
   );
   gpc1_1 gpc2992 (
      {stage0_14[483]},
      {stage1_14[216]}
   );
   gpc1_1 gpc2993 (
      {stage0_14[484]},
      {stage1_14[217]}
   );
   gpc1_1 gpc2994 (
      {stage0_14[485]},
      {stage1_14[218]}
   );
   gpc1_1 gpc2995 (
      {stage0_15[479]},
      {stage1_15[164]}
   );
   gpc1_1 gpc2996 (
      {stage0_15[480]},
      {stage1_15[165]}
   );
   gpc1_1 gpc2997 (
      {stage0_15[481]},
      {stage1_15[166]}
   );
   gpc1_1 gpc2998 (
      {stage0_15[482]},
      {stage1_15[167]}
   );
   gpc1_1 gpc2999 (
      {stage0_15[483]},
      {stage1_15[168]}
   );
   gpc1_1 gpc3000 (
      {stage0_15[484]},
      {stage1_15[169]}
   );
   gpc1_1 gpc3001 (
      {stage0_15[485]},
      {stage1_15[170]}
   );
   gpc1_1 gpc3002 (
      {stage0_17[450]},
      {stage1_17[193]}
   );
   gpc1_1 gpc3003 (
      {stage0_17[451]},
      {stage1_17[194]}
   );
   gpc1_1 gpc3004 (
      {stage0_17[452]},
      {stage1_17[195]}
   );
   gpc1_1 gpc3005 (
      {stage0_17[453]},
      {stage1_17[196]}
   );
   gpc1_1 gpc3006 (
      {stage0_17[454]},
      {stage1_17[197]}
   );
   gpc1_1 gpc3007 (
      {stage0_17[455]},
      {stage1_17[198]}
   );
   gpc1_1 gpc3008 (
      {stage0_17[456]},
      {stage1_17[199]}
   );
   gpc1_1 gpc3009 (
      {stage0_17[457]},
      {stage1_17[200]}
   );
   gpc1_1 gpc3010 (
      {stage0_17[458]},
      {stage1_17[201]}
   );
   gpc1_1 gpc3011 (
      {stage0_17[459]},
      {stage1_17[202]}
   );
   gpc1_1 gpc3012 (
      {stage0_17[460]},
      {stage1_17[203]}
   );
   gpc1_1 gpc3013 (
      {stage0_17[461]},
      {stage1_17[204]}
   );
   gpc1_1 gpc3014 (
      {stage0_17[462]},
      {stage1_17[205]}
   );
   gpc1_1 gpc3015 (
      {stage0_17[463]},
      {stage1_17[206]}
   );
   gpc1_1 gpc3016 (
      {stage0_17[464]},
      {stage1_17[207]}
   );
   gpc1_1 gpc3017 (
      {stage0_17[465]},
      {stage1_17[208]}
   );
   gpc1_1 gpc3018 (
      {stage0_17[466]},
      {stage1_17[209]}
   );
   gpc1_1 gpc3019 (
      {stage0_17[467]},
      {stage1_17[210]}
   );
   gpc1_1 gpc3020 (
      {stage0_17[468]},
      {stage1_17[211]}
   );
   gpc1_1 gpc3021 (
      {stage0_17[469]},
      {stage1_17[212]}
   );
   gpc1_1 gpc3022 (
      {stage0_17[470]},
      {stage1_17[213]}
   );
   gpc1_1 gpc3023 (
      {stage0_17[471]},
      {stage1_17[214]}
   );
   gpc1_1 gpc3024 (
      {stage0_17[472]},
      {stage1_17[215]}
   );
   gpc1_1 gpc3025 (
      {stage0_17[473]},
      {stage1_17[216]}
   );
   gpc1_1 gpc3026 (
      {stage0_17[474]},
      {stage1_17[217]}
   );
   gpc1_1 gpc3027 (
      {stage0_17[475]},
      {stage1_17[218]}
   );
   gpc1_1 gpc3028 (
      {stage0_17[476]},
      {stage1_17[219]}
   );
   gpc1_1 gpc3029 (
      {stage0_17[477]},
      {stage1_17[220]}
   );
   gpc1_1 gpc3030 (
      {stage0_17[478]},
      {stage1_17[221]}
   );
   gpc1_1 gpc3031 (
      {stage0_17[479]},
      {stage1_17[222]}
   );
   gpc1_1 gpc3032 (
      {stage0_17[480]},
      {stage1_17[223]}
   );
   gpc1_1 gpc3033 (
      {stage0_17[481]},
      {stage1_17[224]}
   );
   gpc1_1 gpc3034 (
      {stage0_17[482]},
      {stage1_17[225]}
   );
   gpc1_1 gpc3035 (
      {stage0_17[483]},
      {stage1_17[226]}
   );
   gpc1_1 gpc3036 (
      {stage0_17[484]},
      {stage1_17[227]}
   );
   gpc1_1 gpc3037 (
      {stage0_17[485]},
      {stage1_17[228]}
   );
   gpc1_1 gpc3038 (
      {stage0_18[426]},
      {stage1_18[149]}
   );
   gpc1_1 gpc3039 (
      {stage0_18[427]},
      {stage1_18[150]}
   );
   gpc1_1 gpc3040 (
      {stage0_18[428]},
      {stage1_18[151]}
   );
   gpc1_1 gpc3041 (
      {stage0_18[429]},
      {stage1_18[152]}
   );
   gpc1_1 gpc3042 (
      {stage0_18[430]},
      {stage1_18[153]}
   );
   gpc1_1 gpc3043 (
      {stage0_18[431]},
      {stage1_18[154]}
   );
   gpc1_1 gpc3044 (
      {stage0_18[432]},
      {stage1_18[155]}
   );
   gpc1_1 gpc3045 (
      {stage0_18[433]},
      {stage1_18[156]}
   );
   gpc1_1 gpc3046 (
      {stage0_18[434]},
      {stage1_18[157]}
   );
   gpc1_1 gpc3047 (
      {stage0_18[435]},
      {stage1_18[158]}
   );
   gpc1_1 gpc3048 (
      {stage0_18[436]},
      {stage1_18[159]}
   );
   gpc1_1 gpc3049 (
      {stage0_18[437]},
      {stage1_18[160]}
   );
   gpc1_1 gpc3050 (
      {stage0_18[438]},
      {stage1_18[161]}
   );
   gpc1_1 gpc3051 (
      {stage0_18[439]},
      {stage1_18[162]}
   );
   gpc1_1 gpc3052 (
      {stage0_18[440]},
      {stage1_18[163]}
   );
   gpc1_1 gpc3053 (
      {stage0_18[441]},
      {stage1_18[164]}
   );
   gpc1_1 gpc3054 (
      {stage0_18[442]},
      {stage1_18[165]}
   );
   gpc1_1 gpc3055 (
      {stage0_18[443]},
      {stage1_18[166]}
   );
   gpc1_1 gpc3056 (
      {stage0_18[444]},
      {stage1_18[167]}
   );
   gpc1_1 gpc3057 (
      {stage0_18[445]},
      {stage1_18[168]}
   );
   gpc1_1 gpc3058 (
      {stage0_18[446]},
      {stage1_18[169]}
   );
   gpc1_1 gpc3059 (
      {stage0_18[447]},
      {stage1_18[170]}
   );
   gpc1_1 gpc3060 (
      {stage0_18[448]},
      {stage1_18[171]}
   );
   gpc1_1 gpc3061 (
      {stage0_18[449]},
      {stage1_18[172]}
   );
   gpc1_1 gpc3062 (
      {stage0_18[450]},
      {stage1_18[173]}
   );
   gpc1_1 gpc3063 (
      {stage0_18[451]},
      {stage1_18[174]}
   );
   gpc1_1 gpc3064 (
      {stage0_18[452]},
      {stage1_18[175]}
   );
   gpc1_1 gpc3065 (
      {stage0_18[453]},
      {stage1_18[176]}
   );
   gpc1_1 gpc3066 (
      {stage0_18[454]},
      {stage1_18[177]}
   );
   gpc1_1 gpc3067 (
      {stage0_18[455]},
      {stage1_18[178]}
   );
   gpc1_1 gpc3068 (
      {stage0_18[456]},
      {stage1_18[179]}
   );
   gpc1_1 gpc3069 (
      {stage0_18[457]},
      {stage1_18[180]}
   );
   gpc1_1 gpc3070 (
      {stage0_18[458]},
      {stage1_18[181]}
   );
   gpc1_1 gpc3071 (
      {stage0_18[459]},
      {stage1_18[182]}
   );
   gpc1_1 gpc3072 (
      {stage0_18[460]},
      {stage1_18[183]}
   );
   gpc1_1 gpc3073 (
      {stage0_18[461]},
      {stage1_18[184]}
   );
   gpc1_1 gpc3074 (
      {stage0_18[462]},
      {stage1_18[185]}
   );
   gpc1_1 gpc3075 (
      {stage0_18[463]},
      {stage1_18[186]}
   );
   gpc1_1 gpc3076 (
      {stage0_18[464]},
      {stage1_18[187]}
   );
   gpc1_1 gpc3077 (
      {stage0_18[465]},
      {stage1_18[188]}
   );
   gpc1_1 gpc3078 (
      {stage0_18[466]},
      {stage1_18[189]}
   );
   gpc1_1 gpc3079 (
      {stage0_18[467]},
      {stage1_18[190]}
   );
   gpc1_1 gpc3080 (
      {stage0_18[468]},
      {stage1_18[191]}
   );
   gpc1_1 gpc3081 (
      {stage0_18[469]},
      {stage1_18[192]}
   );
   gpc1_1 gpc3082 (
      {stage0_18[470]},
      {stage1_18[193]}
   );
   gpc1_1 gpc3083 (
      {stage0_18[471]},
      {stage1_18[194]}
   );
   gpc1_1 gpc3084 (
      {stage0_18[472]},
      {stage1_18[195]}
   );
   gpc1_1 gpc3085 (
      {stage0_18[473]},
      {stage1_18[196]}
   );
   gpc1_1 gpc3086 (
      {stage0_18[474]},
      {stage1_18[197]}
   );
   gpc1_1 gpc3087 (
      {stage0_18[475]},
      {stage1_18[198]}
   );
   gpc1_1 gpc3088 (
      {stage0_18[476]},
      {stage1_18[199]}
   );
   gpc1_1 gpc3089 (
      {stage0_18[477]},
      {stage1_18[200]}
   );
   gpc1_1 gpc3090 (
      {stage0_18[478]},
      {stage1_18[201]}
   );
   gpc1_1 gpc3091 (
      {stage0_18[479]},
      {stage1_18[202]}
   );
   gpc1_1 gpc3092 (
      {stage0_18[480]},
      {stage1_18[203]}
   );
   gpc1_1 gpc3093 (
      {stage0_18[481]},
      {stage1_18[204]}
   );
   gpc1_1 gpc3094 (
      {stage0_18[482]},
      {stage1_18[205]}
   );
   gpc1_1 gpc3095 (
      {stage0_18[483]},
      {stage1_18[206]}
   );
   gpc1_1 gpc3096 (
      {stage0_18[484]},
      {stage1_18[207]}
   );
   gpc1_1 gpc3097 (
      {stage0_18[485]},
      {stage1_18[208]}
   );
   gpc1_1 gpc3098 (
      {stage0_19[397]},
      {stage1_19[187]}
   );
   gpc1_1 gpc3099 (
      {stage0_19[398]},
      {stage1_19[188]}
   );
   gpc1_1 gpc3100 (
      {stage0_19[399]},
      {stage1_19[189]}
   );
   gpc1_1 gpc3101 (
      {stage0_19[400]},
      {stage1_19[190]}
   );
   gpc1_1 gpc3102 (
      {stage0_19[401]},
      {stage1_19[191]}
   );
   gpc1_1 gpc3103 (
      {stage0_19[402]},
      {stage1_19[192]}
   );
   gpc1_1 gpc3104 (
      {stage0_19[403]},
      {stage1_19[193]}
   );
   gpc1_1 gpc3105 (
      {stage0_19[404]},
      {stage1_19[194]}
   );
   gpc1_1 gpc3106 (
      {stage0_19[405]},
      {stage1_19[195]}
   );
   gpc1_1 gpc3107 (
      {stage0_19[406]},
      {stage1_19[196]}
   );
   gpc1_1 gpc3108 (
      {stage0_19[407]},
      {stage1_19[197]}
   );
   gpc1_1 gpc3109 (
      {stage0_19[408]},
      {stage1_19[198]}
   );
   gpc1_1 gpc3110 (
      {stage0_19[409]},
      {stage1_19[199]}
   );
   gpc1_1 gpc3111 (
      {stage0_19[410]},
      {stage1_19[200]}
   );
   gpc1_1 gpc3112 (
      {stage0_19[411]},
      {stage1_19[201]}
   );
   gpc1_1 gpc3113 (
      {stage0_19[412]},
      {stage1_19[202]}
   );
   gpc1_1 gpc3114 (
      {stage0_19[413]},
      {stage1_19[203]}
   );
   gpc1_1 gpc3115 (
      {stage0_19[414]},
      {stage1_19[204]}
   );
   gpc1_1 gpc3116 (
      {stage0_19[415]},
      {stage1_19[205]}
   );
   gpc1_1 gpc3117 (
      {stage0_19[416]},
      {stage1_19[206]}
   );
   gpc1_1 gpc3118 (
      {stage0_19[417]},
      {stage1_19[207]}
   );
   gpc1_1 gpc3119 (
      {stage0_19[418]},
      {stage1_19[208]}
   );
   gpc1_1 gpc3120 (
      {stage0_19[419]},
      {stage1_19[209]}
   );
   gpc1_1 gpc3121 (
      {stage0_19[420]},
      {stage1_19[210]}
   );
   gpc1_1 gpc3122 (
      {stage0_19[421]},
      {stage1_19[211]}
   );
   gpc1_1 gpc3123 (
      {stage0_19[422]},
      {stage1_19[212]}
   );
   gpc1_1 gpc3124 (
      {stage0_19[423]},
      {stage1_19[213]}
   );
   gpc1_1 gpc3125 (
      {stage0_19[424]},
      {stage1_19[214]}
   );
   gpc1_1 gpc3126 (
      {stage0_19[425]},
      {stage1_19[215]}
   );
   gpc1_1 gpc3127 (
      {stage0_19[426]},
      {stage1_19[216]}
   );
   gpc1_1 gpc3128 (
      {stage0_19[427]},
      {stage1_19[217]}
   );
   gpc1_1 gpc3129 (
      {stage0_19[428]},
      {stage1_19[218]}
   );
   gpc1_1 gpc3130 (
      {stage0_19[429]},
      {stage1_19[219]}
   );
   gpc1_1 gpc3131 (
      {stage0_19[430]},
      {stage1_19[220]}
   );
   gpc1_1 gpc3132 (
      {stage0_19[431]},
      {stage1_19[221]}
   );
   gpc1_1 gpc3133 (
      {stage0_19[432]},
      {stage1_19[222]}
   );
   gpc1_1 gpc3134 (
      {stage0_19[433]},
      {stage1_19[223]}
   );
   gpc1_1 gpc3135 (
      {stage0_19[434]},
      {stage1_19[224]}
   );
   gpc1_1 gpc3136 (
      {stage0_19[435]},
      {stage1_19[225]}
   );
   gpc1_1 gpc3137 (
      {stage0_19[436]},
      {stage1_19[226]}
   );
   gpc1_1 gpc3138 (
      {stage0_19[437]},
      {stage1_19[227]}
   );
   gpc1_1 gpc3139 (
      {stage0_19[438]},
      {stage1_19[228]}
   );
   gpc1_1 gpc3140 (
      {stage0_19[439]},
      {stage1_19[229]}
   );
   gpc1_1 gpc3141 (
      {stage0_19[440]},
      {stage1_19[230]}
   );
   gpc1_1 gpc3142 (
      {stage0_19[441]},
      {stage1_19[231]}
   );
   gpc1_1 gpc3143 (
      {stage0_19[442]},
      {stage1_19[232]}
   );
   gpc1_1 gpc3144 (
      {stage0_19[443]},
      {stage1_19[233]}
   );
   gpc1_1 gpc3145 (
      {stage0_19[444]},
      {stage1_19[234]}
   );
   gpc1_1 gpc3146 (
      {stage0_19[445]},
      {stage1_19[235]}
   );
   gpc1_1 gpc3147 (
      {stage0_19[446]},
      {stage1_19[236]}
   );
   gpc1_1 gpc3148 (
      {stage0_19[447]},
      {stage1_19[237]}
   );
   gpc1_1 gpc3149 (
      {stage0_19[448]},
      {stage1_19[238]}
   );
   gpc1_1 gpc3150 (
      {stage0_19[449]},
      {stage1_19[239]}
   );
   gpc1_1 gpc3151 (
      {stage0_19[450]},
      {stage1_19[240]}
   );
   gpc1_1 gpc3152 (
      {stage0_19[451]},
      {stage1_19[241]}
   );
   gpc1_1 gpc3153 (
      {stage0_19[452]},
      {stage1_19[242]}
   );
   gpc1_1 gpc3154 (
      {stage0_19[453]},
      {stage1_19[243]}
   );
   gpc1_1 gpc3155 (
      {stage0_19[454]},
      {stage1_19[244]}
   );
   gpc1_1 gpc3156 (
      {stage0_19[455]},
      {stage1_19[245]}
   );
   gpc1_1 gpc3157 (
      {stage0_19[456]},
      {stage1_19[246]}
   );
   gpc1_1 gpc3158 (
      {stage0_19[457]},
      {stage1_19[247]}
   );
   gpc1_1 gpc3159 (
      {stage0_19[458]},
      {stage1_19[248]}
   );
   gpc1_1 gpc3160 (
      {stage0_19[459]},
      {stage1_19[249]}
   );
   gpc1_1 gpc3161 (
      {stage0_19[460]},
      {stage1_19[250]}
   );
   gpc1_1 gpc3162 (
      {stage0_19[461]},
      {stage1_19[251]}
   );
   gpc1_1 gpc3163 (
      {stage0_19[462]},
      {stage1_19[252]}
   );
   gpc1_1 gpc3164 (
      {stage0_19[463]},
      {stage1_19[253]}
   );
   gpc1_1 gpc3165 (
      {stage0_19[464]},
      {stage1_19[254]}
   );
   gpc1_1 gpc3166 (
      {stage0_19[465]},
      {stage1_19[255]}
   );
   gpc1_1 gpc3167 (
      {stage0_19[466]},
      {stage1_19[256]}
   );
   gpc1_1 gpc3168 (
      {stage0_19[467]},
      {stage1_19[257]}
   );
   gpc1_1 gpc3169 (
      {stage0_19[468]},
      {stage1_19[258]}
   );
   gpc1_1 gpc3170 (
      {stage0_19[469]},
      {stage1_19[259]}
   );
   gpc1_1 gpc3171 (
      {stage0_19[470]},
      {stage1_19[260]}
   );
   gpc1_1 gpc3172 (
      {stage0_19[471]},
      {stage1_19[261]}
   );
   gpc1_1 gpc3173 (
      {stage0_19[472]},
      {stage1_19[262]}
   );
   gpc1_1 gpc3174 (
      {stage0_19[473]},
      {stage1_19[263]}
   );
   gpc1_1 gpc3175 (
      {stage0_19[474]},
      {stage1_19[264]}
   );
   gpc1_1 gpc3176 (
      {stage0_19[475]},
      {stage1_19[265]}
   );
   gpc1_1 gpc3177 (
      {stage0_19[476]},
      {stage1_19[266]}
   );
   gpc1_1 gpc3178 (
      {stage0_19[477]},
      {stage1_19[267]}
   );
   gpc1_1 gpc3179 (
      {stage0_19[478]},
      {stage1_19[268]}
   );
   gpc1_1 gpc3180 (
      {stage0_19[479]},
      {stage1_19[269]}
   );
   gpc1_1 gpc3181 (
      {stage0_19[480]},
      {stage1_19[270]}
   );
   gpc1_1 gpc3182 (
      {stage0_19[481]},
      {stage1_19[271]}
   );
   gpc1_1 gpc3183 (
      {stage0_19[482]},
      {stage1_19[272]}
   );
   gpc1_1 gpc3184 (
      {stage0_19[483]},
      {stage1_19[273]}
   );
   gpc1_1 gpc3185 (
      {stage0_19[484]},
      {stage1_19[274]}
   );
   gpc1_1 gpc3186 (
      {stage0_19[485]},
      {stage1_19[275]}
   );
   gpc1_1 gpc3187 (
      {stage0_20[432]},
      {stage1_20[214]}
   );
   gpc1_1 gpc3188 (
      {stage0_20[433]},
      {stage1_20[215]}
   );
   gpc1_1 gpc3189 (
      {stage0_20[434]},
      {stage1_20[216]}
   );
   gpc1_1 gpc3190 (
      {stage0_20[435]},
      {stage1_20[217]}
   );
   gpc1_1 gpc3191 (
      {stage0_20[436]},
      {stage1_20[218]}
   );
   gpc1_1 gpc3192 (
      {stage0_20[437]},
      {stage1_20[219]}
   );
   gpc1_1 gpc3193 (
      {stage0_20[438]},
      {stage1_20[220]}
   );
   gpc1_1 gpc3194 (
      {stage0_20[439]},
      {stage1_20[221]}
   );
   gpc1_1 gpc3195 (
      {stage0_20[440]},
      {stage1_20[222]}
   );
   gpc1_1 gpc3196 (
      {stage0_20[441]},
      {stage1_20[223]}
   );
   gpc1_1 gpc3197 (
      {stage0_20[442]},
      {stage1_20[224]}
   );
   gpc1_1 gpc3198 (
      {stage0_20[443]},
      {stage1_20[225]}
   );
   gpc1_1 gpc3199 (
      {stage0_20[444]},
      {stage1_20[226]}
   );
   gpc1_1 gpc3200 (
      {stage0_20[445]},
      {stage1_20[227]}
   );
   gpc1_1 gpc3201 (
      {stage0_20[446]},
      {stage1_20[228]}
   );
   gpc1_1 gpc3202 (
      {stage0_20[447]},
      {stage1_20[229]}
   );
   gpc1_1 gpc3203 (
      {stage0_20[448]},
      {stage1_20[230]}
   );
   gpc1_1 gpc3204 (
      {stage0_20[449]},
      {stage1_20[231]}
   );
   gpc1_1 gpc3205 (
      {stage0_20[450]},
      {stage1_20[232]}
   );
   gpc1_1 gpc3206 (
      {stage0_20[451]},
      {stage1_20[233]}
   );
   gpc1_1 gpc3207 (
      {stage0_20[452]},
      {stage1_20[234]}
   );
   gpc1_1 gpc3208 (
      {stage0_20[453]},
      {stage1_20[235]}
   );
   gpc1_1 gpc3209 (
      {stage0_20[454]},
      {stage1_20[236]}
   );
   gpc1_1 gpc3210 (
      {stage0_20[455]},
      {stage1_20[237]}
   );
   gpc1_1 gpc3211 (
      {stage0_20[456]},
      {stage1_20[238]}
   );
   gpc1_1 gpc3212 (
      {stage0_20[457]},
      {stage1_20[239]}
   );
   gpc1_1 gpc3213 (
      {stage0_20[458]},
      {stage1_20[240]}
   );
   gpc1_1 gpc3214 (
      {stage0_20[459]},
      {stage1_20[241]}
   );
   gpc1_1 gpc3215 (
      {stage0_20[460]},
      {stage1_20[242]}
   );
   gpc1_1 gpc3216 (
      {stage0_20[461]},
      {stage1_20[243]}
   );
   gpc1_1 gpc3217 (
      {stage0_20[462]},
      {stage1_20[244]}
   );
   gpc1_1 gpc3218 (
      {stage0_20[463]},
      {stage1_20[245]}
   );
   gpc1_1 gpc3219 (
      {stage0_20[464]},
      {stage1_20[246]}
   );
   gpc1_1 gpc3220 (
      {stage0_20[465]},
      {stage1_20[247]}
   );
   gpc1_1 gpc3221 (
      {stage0_20[466]},
      {stage1_20[248]}
   );
   gpc1_1 gpc3222 (
      {stage0_20[467]},
      {stage1_20[249]}
   );
   gpc1_1 gpc3223 (
      {stage0_20[468]},
      {stage1_20[250]}
   );
   gpc1_1 gpc3224 (
      {stage0_20[469]},
      {stage1_20[251]}
   );
   gpc1_1 gpc3225 (
      {stage0_20[470]},
      {stage1_20[252]}
   );
   gpc1_1 gpc3226 (
      {stage0_20[471]},
      {stage1_20[253]}
   );
   gpc1_1 gpc3227 (
      {stage0_20[472]},
      {stage1_20[254]}
   );
   gpc1_1 gpc3228 (
      {stage0_20[473]},
      {stage1_20[255]}
   );
   gpc1_1 gpc3229 (
      {stage0_20[474]},
      {stage1_20[256]}
   );
   gpc1_1 gpc3230 (
      {stage0_20[475]},
      {stage1_20[257]}
   );
   gpc1_1 gpc3231 (
      {stage0_20[476]},
      {stage1_20[258]}
   );
   gpc1_1 gpc3232 (
      {stage0_20[477]},
      {stage1_20[259]}
   );
   gpc1_1 gpc3233 (
      {stage0_20[478]},
      {stage1_20[260]}
   );
   gpc1_1 gpc3234 (
      {stage0_20[479]},
      {stage1_20[261]}
   );
   gpc1_1 gpc3235 (
      {stage0_20[480]},
      {stage1_20[262]}
   );
   gpc1_1 gpc3236 (
      {stage0_20[481]},
      {stage1_20[263]}
   );
   gpc1_1 gpc3237 (
      {stage0_20[482]},
      {stage1_20[264]}
   );
   gpc1_1 gpc3238 (
      {stage0_20[483]},
      {stage1_20[265]}
   );
   gpc1_1 gpc3239 (
      {stage0_20[484]},
      {stage1_20[266]}
   );
   gpc1_1 gpc3240 (
      {stage0_20[485]},
      {stage1_20[267]}
   );
   gpc1_1 gpc3241 (
      {stage0_21[468]},
      {stage1_21[172]}
   );
   gpc1_1 gpc3242 (
      {stage0_21[469]},
      {stage1_21[173]}
   );
   gpc1_1 gpc3243 (
      {stage0_21[470]},
      {stage1_21[174]}
   );
   gpc1_1 gpc3244 (
      {stage0_21[471]},
      {stage1_21[175]}
   );
   gpc1_1 gpc3245 (
      {stage0_21[472]},
      {stage1_21[176]}
   );
   gpc1_1 gpc3246 (
      {stage0_21[473]},
      {stage1_21[177]}
   );
   gpc1_1 gpc3247 (
      {stage0_21[474]},
      {stage1_21[178]}
   );
   gpc1_1 gpc3248 (
      {stage0_21[475]},
      {stage1_21[179]}
   );
   gpc1_1 gpc3249 (
      {stage0_21[476]},
      {stage1_21[180]}
   );
   gpc1_1 gpc3250 (
      {stage0_21[477]},
      {stage1_21[181]}
   );
   gpc1_1 gpc3251 (
      {stage0_21[478]},
      {stage1_21[182]}
   );
   gpc1_1 gpc3252 (
      {stage0_21[479]},
      {stage1_21[183]}
   );
   gpc1_1 gpc3253 (
      {stage0_21[480]},
      {stage1_21[184]}
   );
   gpc1_1 gpc3254 (
      {stage0_21[481]},
      {stage1_21[185]}
   );
   gpc1_1 gpc3255 (
      {stage0_21[482]},
      {stage1_21[186]}
   );
   gpc1_1 gpc3256 (
      {stage0_21[483]},
      {stage1_21[187]}
   );
   gpc1_1 gpc3257 (
      {stage0_21[484]},
      {stage1_21[188]}
   );
   gpc1_1 gpc3258 (
      {stage0_21[485]},
      {stage1_21[189]}
   );
   gpc1_1 gpc3259 (
      {stage0_22[472]},
      {stage1_22[157]}
   );
   gpc1_1 gpc3260 (
      {stage0_22[473]},
      {stage1_22[158]}
   );
   gpc1_1 gpc3261 (
      {stage0_22[474]},
      {stage1_22[159]}
   );
   gpc1_1 gpc3262 (
      {stage0_22[475]},
      {stage1_22[160]}
   );
   gpc1_1 gpc3263 (
      {stage0_22[476]},
      {stage1_22[161]}
   );
   gpc1_1 gpc3264 (
      {stage0_22[477]},
      {stage1_22[162]}
   );
   gpc1_1 gpc3265 (
      {stage0_22[478]},
      {stage1_22[163]}
   );
   gpc1_1 gpc3266 (
      {stage0_22[479]},
      {stage1_22[164]}
   );
   gpc1_1 gpc3267 (
      {stage0_22[480]},
      {stage1_22[165]}
   );
   gpc1_1 gpc3268 (
      {stage0_22[481]},
      {stage1_22[166]}
   );
   gpc1_1 gpc3269 (
      {stage0_22[482]},
      {stage1_22[167]}
   );
   gpc1_1 gpc3270 (
      {stage0_22[483]},
      {stage1_22[168]}
   );
   gpc1_1 gpc3271 (
      {stage0_22[484]},
      {stage1_22[169]}
   );
   gpc1_1 gpc3272 (
      {stage0_22[485]},
      {stage1_22[170]}
   );
   gpc1_1 gpc3273 (
      {stage0_23[396]},
      {stage1_23[197]}
   );
   gpc1_1 gpc3274 (
      {stage0_23[397]},
      {stage1_23[198]}
   );
   gpc1_1 gpc3275 (
      {stage0_23[398]},
      {stage1_23[199]}
   );
   gpc1_1 gpc3276 (
      {stage0_23[399]},
      {stage1_23[200]}
   );
   gpc1_1 gpc3277 (
      {stage0_23[400]},
      {stage1_23[201]}
   );
   gpc1_1 gpc3278 (
      {stage0_23[401]},
      {stage1_23[202]}
   );
   gpc1_1 gpc3279 (
      {stage0_23[402]},
      {stage1_23[203]}
   );
   gpc1_1 gpc3280 (
      {stage0_23[403]},
      {stage1_23[204]}
   );
   gpc1_1 gpc3281 (
      {stage0_23[404]},
      {stage1_23[205]}
   );
   gpc1_1 gpc3282 (
      {stage0_23[405]},
      {stage1_23[206]}
   );
   gpc1_1 gpc3283 (
      {stage0_23[406]},
      {stage1_23[207]}
   );
   gpc1_1 gpc3284 (
      {stage0_23[407]},
      {stage1_23[208]}
   );
   gpc1_1 gpc3285 (
      {stage0_23[408]},
      {stage1_23[209]}
   );
   gpc1_1 gpc3286 (
      {stage0_23[409]},
      {stage1_23[210]}
   );
   gpc1_1 gpc3287 (
      {stage0_23[410]},
      {stage1_23[211]}
   );
   gpc1_1 gpc3288 (
      {stage0_23[411]},
      {stage1_23[212]}
   );
   gpc1_1 gpc3289 (
      {stage0_23[412]},
      {stage1_23[213]}
   );
   gpc1_1 gpc3290 (
      {stage0_23[413]},
      {stage1_23[214]}
   );
   gpc1_1 gpc3291 (
      {stage0_23[414]},
      {stage1_23[215]}
   );
   gpc1_1 gpc3292 (
      {stage0_23[415]},
      {stage1_23[216]}
   );
   gpc1_1 gpc3293 (
      {stage0_23[416]},
      {stage1_23[217]}
   );
   gpc1_1 gpc3294 (
      {stage0_23[417]},
      {stage1_23[218]}
   );
   gpc1_1 gpc3295 (
      {stage0_23[418]},
      {stage1_23[219]}
   );
   gpc1_1 gpc3296 (
      {stage0_23[419]},
      {stage1_23[220]}
   );
   gpc1_1 gpc3297 (
      {stage0_23[420]},
      {stage1_23[221]}
   );
   gpc1_1 gpc3298 (
      {stage0_23[421]},
      {stage1_23[222]}
   );
   gpc1_1 gpc3299 (
      {stage0_23[422]},
      {stage1_23[223]}
   );
   gpc1_1 gpc3300 (
      {stage0_23[423]},
      {stage1_23[224]}
   );
   gpc1_1 gpc3301 (
      {stage0_23[424]},
      {stage1_23[225]}
   );
   gpc1_1 gpc3302 (
      {stage0_23[425]},
      {stage1_23[226]}
   );
   gpc1_1 gpc3303 (
      {stage0_23[426]},
      {stage1_23[227]}
   );
   gpc1_1 gpc3304 (
      {stage0_23[427]},
      {stage1_23[228]}
   );
   gpc1_1 gpc3305 (
      {stage0_23[428]},
      {stage1_23[229]}
   );
   gpc1_1 gpc3306 (
      {stage0_23[429]},
      {stage1_23[230]}
   );
   gpc1_1 gpc3307 (
      {stage0_23[430]},
      {stage1_23[231]}
   );
   gpc1_1 gpc3308 (
      {stage0_23[431]},
      {stage1_23[232]}
   );
   gpc1_1 gpc3309 (
      {stage0_23[432]},
      {stage1_23[233]}
   );
   gpc1_1 gpc3310 (
      {stage0_23[433]},
      {stage1_23[234]}
   );
   gpc1_1 gpc3311 (
      {stage0_23[434]},
      {stage1_23[235]}
   );
   gpc1_1 gpc3312 (
      {stage0_23[435]},
      {stage1_23[236]}
   );
   gpc1_1 gpc3313 (
      {stage0_23[436]},
      {stage1_23[237]}
   );
   gpc1_1 gpc3314 (
      {stage0_23[437]},
      {stage1_23[238]}
   );
   gpc1_1 gpc3315 (
      {stage0_23[438]},
      {stage1_23[239]}
   );
   gpc1_1 gpc3316 (
      {stage0_23[439]},
      {stage1_23[240]}
   );
   gpc1_1 gpc3317 (
      {stage0_23[440]},
      {stage1_23[241]}
   );
   gpc1_1 gpc3318 (
      {stage0_23[441]},
      {stage1_23[242]}
   );
   gpc1_1 gpc3319 (
      {stage0_23[442]},
      {stage1_23[243]}
   );
   gpc1_1 gpc3320 (
      {stage0_23[443]},
      {stage1_23[244]}
   );
   gpc1_1 gpc3321 (
      {stage0_23[444]},
      {stage1_23[245]}
   );
   gpc1_1 gpc3322 (
      {stage0_23[445]},
      {stage1_23[246]}
   );
   gpc1_1 gpc3323 (
      {stage0_23[446]},
      {stage1_23[247]}
   );
   gpc1_1 gpc3324 (
      {stage0_23[447]},
      {stage1_23[248]}
   );
   gpc1_1 gpc3325 (
      {stage0_23[448]},
      {stage1_23[249]}
   );
   gpc1_1 gpc3326 (
      {stage0_23[449]},
      {stage1_23[250]}
   );
   gpc1_1 gpc3327 (
      {stage0_23[450]},
      {stage1_23[251]}
   );
   gpc1_1 gpc3328 (
      {stage0_23[451]},
      {stage1_23[252]}
   );
   gpc1_1 gpc3329 (
      {stage0_23[452]},
      {stage1_23[253]}
   );
   gpc1_1 gpc3330 (
      {stage0_23[453]},
      {stage1_23[254]}
   );
   gpc1_1 gpc3331 (
      {stage0_23[454]},
      {stage1_23[255]}
   );
   gpc1_1 gpc3332 (
      {stage0_23[455]},
      {stage1_23[256]}
   );
   gpc1_1 gpc3333 (
      {stage0_23[456]},
      {stage1_23[257]}
   );
   gpc1_1 gpc3334 (
      {stage0_23[457]},
      {stage1_23[258]}
   );
   gpc1_1 gpc3335 (
      {stage0_23[458]},
      {stage1_23[259]}
   );
   gpc1_1 gpc3336 (
      {stage0_23[459]},
      {stage1_23[260]}
   );
   gpc1_1 gpc3337 (
      {stage0_23[460]},
      {stage1_23[261]}
   );
   gpc1_1 gpc3338 (
      {stage0_23[461]},
      {stage1_23[262]}
   );
   gpc1_1 gpc3339 (
      {stage0_23[462]},
      {stage1_23[263]}
   );
   gpc1_1 gpc3340 (
      {stage0_23[463]},
      {stage1_23[264]}
   );
   gpc1_1 gpc3341 (
      {stage0_23[464]},
      {stage1_23[265]}
   );
   gpc1_1 gpc3342 (
      {stage0_23[465]},
      {stage1_23[266]}
   );
   gpc1_1 gpc3343 (
      {stage0_23[466]},
      {stage1_23[267]}
   );
   gpc1_1 gpc3344 (
      {stage0_23[467]},
      {stage1_23[268]}
   );
   gpc1_1 gpc3345 (
      {stage0_23[468]},
      {stage1_23[269]}
   );
   gpc1_1 gpc3346 (
      {stage0_23[469]},
      {stage1_23[270]}
   );
   gpc1_1 gpc3347 (
      {stage0_23[470]},
      {stage1_23[271]}
   );
   gpc1_1 gpc3348 (
      {stage0_23[471]},
      {stage1_23[272]}
   );
   gpc1_1 gpc3349 (
      {stage0_23[472]},
      {stage1_23[273]}
   );
   gpc1_1 gpc3350 (
      {stage0_23[473]},
      {stage1_23[274]}
   );
   gpc1_1 gpc3351 (
      {stage0_23[474]},
      {stage1_23[275]}
   );
   gpc1_1 gpc3352 (
      {stage0_23[475]},
      {stage1_23[276]}
   );
   gpc1_1 gpc3353 (
      {stage0_23[476]},
      {stage1_23[277]}
   );
   gpc1_1 gpc3354 (
      {stage0_23[477]},
      {stage1_23[278]}
   );
   gpc1_1 gpc3355 (
      {stage0_23[478]},
      {stage1_23[279]}
   );
   gpc1_1 gpc3356 (
      {stage0_23[479]},
      {stage1_23[280]}
   );
   gpc1_1 gpc3357 (
      {stage0_23[480]},
      {stage1_23[281]}
   );
   gpc1_1 gpc3358 (
      {stage0_23[481]},
      {stage1_23[282]}
   );
   gpc1_1 gpc3359 (
      {stage0_23[482]},
      {stage1_23[283]}
   );
   gpc1_1 gpc3360 (
      {stage0_23[483]},
      {stage1_23[284]}
   );
   gpc1_1 gpc3361 (
      {stage0_23[484]},
      {stage1_23[285]}
   );
   gpc1_1 gpc3362 (
      {stage0_23[485]},
      {stage1_23[286]}
   );
   gpc1_1 gpc3363 (
      {stage0_24[485]},
      {stage1_24[213]}
   );
   gpc1_1 gpc3364 (
      {stage0_26[402]},
      {stage1_26[167]}
   );
   gpc1_1 gpc3365 (
      {stage0_26[403]},
      {stage1_26[168]}
   );
   gpc1_1 gpc3366 (
      {stage0_26[404]},
      {stage1_26[169]}
   );
   gpc1_1 gpc3367 (
      {stage0_26[405]},
      {stage1_26[170]}
   );
   gpc1_1 gpc3368 (
      {stage0_26[406]},
      {stage1_26[171]}
   );
   gpc1_1 gpc3369 (
      {stage0_26[407]},
      {stage1_26[172]}
   );
   gpc1_1 gpc3370 (
      {stage0_26[408]},
      {stage1_26[173]}
   );
   gpc1_1 gpc3371 (
      {stage0_26[409]},
      {stage1_26[174]}
   );
   gpc1_1 gpc3372 (
      {stage0_26[410]},
      {stage1_26[175]}
   );
   gpc1_1 gpc3373 (
      {stage0_26[411]},
      {stage1_26[176]}
   );
   gpc1_1 gpc3374 (
      {stage0_26[412]},
      {stage1_26[177]}
   );
   gpc1_1 gpc3375 (
      {stage0_26[413]},
      {stage1_26[178]}
   );
   gpc1_1 gpc3376 (
      {stage0_26[414]},
      {stage1_26[179]}
   );
   gpc1_1 gpc3377 (
      {stage0_26[415]},
      {stage1_26[180]}
   );
   gpc1_1 gpc3378 (
      {stage0_26[416]},
      {stage1_26[181]}
   );
   gpc1_1 gpc3379 (
      {stage0_26[417]},
      {stage1_26[182]}
   );
   gpc1_1 gpc3380 (
      {stage0_26[418]},
      {stage1_26[183]}
   );
   gpc1_1 gpc3381 (
      {stage0_26[419]},
      {stage1_26[184]}
   );
   gpc1_1 gpc3382 (
      {stage0_26[420]},
      {stage1_26[185]}
   );
   gpc1_1 gpc3383 (
      {stage0_26[421]},
      {stage1_26[186]}
   );
   gpc1_1 gpc3384 (
      {stage0_26[422]},
      {stage1_26[187]}
   );
   gpc1_1 gpc3385 (
      {stage0_26[423]},
      {stage1_26[188]}
   );
   gpc1_1 gpc3386 (
      {stage0_26[424]},
      {stage1_26[189]}
   );
   gpc1_1 gpc3387 (
      {stage0_26[425]},
      {stage1_26[190]}
   );
   gpc1_1 gpc3388 (
      {stage0_26[426]},
      {stage1_26[191]}
   );
   gpc1_1 gpc3389 (
      {stage0_26[427]},
      {stage1_26[192]}
   );
   gpc1_1 gpc3390 (
      {stage0_26[428]},
      {stage1_26[193]}
   );
   gpc1_1 gpc3391 (
      {stage0_26[429]},
      {stage1_26[194]}
   );
   gpc1_1 gpc3392 (
      {stage0_26[430]},
      {stage1_26[195]}
   );
   gpc1_1 gpc3393 (
      {stage0_26[431]},
      {stage1_26[196]}
   );
   gpc1_1 gpc3394 (
      {stage0_26[432]},
      {stage1_26[197]}
   );
   gpc1_1 gpc3395 (
      {stage0_26[433]},
      {stage1_26[198]}
   );
   gpc1_1 gpc3396 (
      {stage0_26[434]},
      {stage1_26[199]}
   );
   gpc1_1 gpc3397 (
      {stage0_26[435]},
      {stage1_26[200]}
   );
   gpc1_1 gpc3398 (
      {stage0_26[436]},
      {stage1_26[201]}
   );
   gpc1_1 gpc3399 (
      {stage0_26[437]},
      {stage1_26[202]}
   );
   gpc1_1 gpc3400 (
      {stage0_26[438]},
      {stage1_26[203]}
   );
   gpc1_1 gpc3401 (
      {stage0_26[439]},
      {stage1_26[204]}
   );
   gpc1_1 gpc3402 (
      {stage0_26[440]},
      {stage1_26[205]}
   );
   gpc1_1 gpc3403 (
      {stage0_26[441]},
      {stage1_26[206]}
   );
   gpc1_1 gpc3404 (
      {stage0_26[442]},
      {stage1_26[207]}
   );
   gpc1_1 gpc3405 (
      {stage0_26[443]},
      {stage1_26[208]}
   );
   gpc1_1 gpc3406 (
      {stage0_26[444]},
      {stage1_26[209]}
   );
   gpc1_1 gpc3407 (
      {stage0_26[445]},
      {stage1_26[210]}
   );
   gpc1_1 gpc3408 (
      {stage0_26[446]},
      {stage1_26[211]}
   );
   gpc1_1 gpc3409 (
      {stage0_26[447]},
      {stage1_26[212]}
   );
   gpc1_1 gpc3410 (
      {stage0_26[448]},
      {stage1_26[213]}
   );
   gpc1_1 gpc3411 (
      {stage0_26[449]},
      {stage1_26[214]}
   );
   gpc1_1 gpc3412 (
      {stage0_26[450]},
      {stage1_26[215]}
   );
   gpc1_1 gpc3413 (
      {stage0_26[451]},
      {stage1_26[216]}
   );
   gpc1_1 gpc3414 (
      {stage0_26[452]},
      {stage1_26[217]}
   );
   gpc1_1 gpc3415 (
      {stage0_26[453]},
      {stage1_26[218]}
   );
   gpc1_1 gpc3416 (
      {stage0_26[454]},
      {stage1_26[219]}
   );
   gpc1_1 gpc3417 (
      {stage0_26[455]},
      {stage1_26[220]}
   );
   gpc1_1 gpc3418 (
      {stage0_26[456]},
      {stage1_26[221]}
   );
   gpc1_1 gpc3419 (
      {stage0_26[457]},
      {stage1_26[222]}
   );
   gpc1_1 gpc3420 (
      {stage0_26[458]},
      {stage1_26[223]}
   );
   gpc1_1 gpc3421 (
      {stage0_26[459]},
      {stage1_26[224]}
   );
   gpc1_1 gpc3422 (
      {stage0_26[460]},
      {stage1_26[225]}
   );
   gpc1_1 gpc3423 (
      {stage0_26[461]},
      {stage1_26[226]}
   );
   gpc1_1 gpc3424 (
      {stage0_26[462]},
      {stage1_26[227]}
   );
   gpc1_1 gpc3425 (
      {stage0_26[463]},
      {stage1_26[228]}
   );
   gpc1_1 gpc3426 (
      {stage0_26[464]},
      {stage1_26[229]}
   );
   gpc1_1 gpc3427 (
      {stage0_26[465]},
      {stage1_26[230]}
   );
   gpc1_1 gpc3428 (
      {stage0_26[466]},
      {stage1_26[231]}
   );
   gpc1_1 gpc3429 (
      {stage0_26[467]},
      {stage1_26[232]}
   );
   gpc1_1 gpc3430 (
      {stage0_26[468]},
      {stage1_26[233]}
   );
   gpc1_1 gpc3431 (
      {stage0_26[469]},
      {stage1_26[234]}
   );
   gpc1_1 gpc3432 (
      {stage0_26[470]},
      {stage1_26[235]}
   );
   gpc1_1 gpc3433 (
      {stage0_26[471]},
      {stage1_26[236]}
   );
   gpc1_1 gpc3434 (
      {stage0_26[472]},
      {stage1_26[237]}
   );
   gpc1_1 gpc3435 (
      {stage0_26[473]},
      {stage1_26[238]}
   );
   gpc1_1 gpc3436 (
      {stage0_26[474]},
      {stage1_26[239]}
   );
   gpc1_1 gpc3437 (
      {stage0_26[475]},
      {stage1_26[240]}
   );
   gpc1_1 gpc3438 (
      {stage0_26[476]},
      {stage1_26[241]}
   );
   gpc1_1 gpc3439 (
      {stage0_26[477]},
      {stage1_26[242]}
   );
   gpc1_1 gpc3440 (
      {stage0_26[478]},
      {stage1_26[243]}
   );
   gpc1_1 gpc3441 (
      {stage0_26[479]},
      {stage1_26[244]}
   );
   gpc1_1 gpc3442 (
      {stage0_26[480]},
      {stage1_26[245]}
   );
   gpc1_1 gpc3443 (
      {stage0_26[481]},
      {stage1_26[246]}
   );
   gpc1_1 gpc3444 (
      {stage0_26[482]},
      {stage1_26[247]}
   );
   gpc1_1 gpc3445 (
      {stage0_26[483]},
      {stage1_26[248]}
   );
   gpc1_1 gpc3446 (
      {stage0_26[484]},
      {stage1_26[249]}
   );
   gpc1_1 gpc3447 (
      {stage0_26[485]},
      {stage1_26[250]}
   );
   gpc1_1 gpc3448 (
      {stage0_27[473]},
      {stage1_27[193]}
   );
   gpc1_1 gpc3449 (
      {stage0_27[474]},
      {stage1_27[194]}
   );
   gpc1_1 gpc3450 (
      {stage0_27[475]},
      {stage1_27[195]}
   );
   gpc1_1 gpc3451 (
      {stage0_27[476]},
      {stage1_27[196]}
   );
   gpc1_1 gpc3452 (
      {stage0_27[477]},
      {stage1_27[197]}
   );
   gpc1_1 gpc3453 (
      {stage0_27[478]},
      {stage1_27[198]}
   );
   gpc1_1 gpc3454 (
      {stage0_27[479]},
      {stage1_27[199]}
   );
   gpc1_1 gpc3455 (
      {stage0_27[480]},
      {stage1_27[200]}
   );
   gpc1_1 gpc3456 (
      {stage0_27[481]},
      {stage1_27[201]}
   );
   gpc1_1 gpc3457 (
      {stage0_27[482]},
      {stage1_27[202]}
   );
   gpc1_1 gpc3458 (
      {stage0_27[483]},
      {stage1_27[203]}
   );
   gpc1_1 gpc3459 (
      {stage0_27[484]},
      {stage1_27[204]}
   );
   gpc1_1 gpc3460 (
      {stage0_27[485]},
      {stage1_27[205]}
   );
   gpc1_1 gpc3461 (
      {stage0_28[475]},
      {stage1_28[213]}
   );
   gpc1_1 gpc3462 (
      {stage0_28[476]},
      {stage1_28[214]}
   );
   gpc1_1 gpc3463 (
      {stage0_28[477]},
      {stage1_28[215]}
   );
   gpc1_1 gpc3464 (
      {stage0_28[478]},
      {stage1_28[216]}
   );
   gpc1_1 gpc3465 (
      {stage0_28[479]},
      {stage1_28[217]}
   );
   gpc1_1 gpc3466 (
      {stage0_28[480]},
      {stage1_28[218]}
   );
   gpc1_1 gpc3467 (
      {stage0_28[481]},
      {stage1_28[219]}
   );
   gpc1_1 gpc3468 (
      {stage0_28[482]},
      {stage1_28[220]}
   );
   gpc1_1 gpc3469 (
      {stage0_28[483]},
      {stage1_28[221]}
   );
   gpc1_1 gpc3470 (
      {stage0_28[484]},
      {stage1_28[222]}
   );
   gpc1_1 gpc3471 (
      {stage0_28[485]},
      {stage1_28[223]}
   );
   gpc1_1 gpc3472 (
      {stage0_29[444]},
      {stage1_29[187]}
   );
   gpc1_1 gpc3473 (
      {stage0_29[445]},
      {stage1_29[188]}
   );
   gpc1_1 gpc3474 (
      {stage0_29[446]},
      {stage1_29[189]}
   );
   gpc1_1 gpc3475 (
      {stage0_29[447]},
      {stage1_29[190]}
   );
   gpc1_1 gpc3476 (
      {stage0_29[448]},
      {stage1_29[191]}
   );
   gpc1_1 gpc3477 (
      {stage0_29[449]},
      {stage1_29[192]}
   );
   gpc1_1 gpc3478 (
      {stage0_29[450]},
      {stage1_29[193]}
   );
   gpc1_1 gpc3479 (
      {stage0_29[451]},
      {stage1_29[194]}
   );
   gpc1_1 gpc3480 (
      {stage0_29[452]},
      {stage1_29[195]}
   );
   gpc1_1 gpc3481 (
      {stage0_29[453]},
      {stage1_29[196]}
   );
   gpc1_1 gpc3482 (
      {stage0_29[454]},
      {stage1_29[197]}
   );
   gpc1_1 gpc3483 (
      {stage0_29[455]},
      {stage1_29[198]}
   );
   gpc1_1 gpc3484 (
      {stage0_29[456]},
      {stage1_29[199]}
   );
   gpc1_1 gpc3485 (
      {stage0_29[457]},
      {stage1_29[200]}
   );
   gpc1_1 gpc3486 (
      {stage0_29[458]},
      {stage1_29[201]}
   );
   gpc1_1 gpc3487 (
      {stage0_29[459]},
      {stage1_29[202]}
   );
   gpc1_1 gpc3488 (
      {stage0_29[460]},
      {stage1_29[203]}
   );
   gpc1_1 gpc3489 (
      {stage0_29[461]},
      {stage1_29[204]}
   );
   gpc1_1 gpc3490 (
      {stage0_29[462]},
      {stage1_29[205]}
   );
   gpc1_1 gpc3491 (
      {stage0_29[463]},
      {stage1_29[206]}
   );
   gpc1_1 gpc3492 (
      {stage0_29[464]},
      {stage1_29[207]}
   );
   gpc1_1 gpc3493 (
      {stage0_29[465]},
      {stage1_29[208]}
   );
   gpc1_1 gpc3494 (
      {stage0_29[466]},
      {stage1_29[209]}
   );
   gpc1_1 gpc3495 (
      {stage0_29[467]},
      {stage1_29[210]}
   );
   gpc1_1 gpc3496 (
      {stage0_29[468]},
      {stage1_29[211]}
   );
   gpc1_1 gpc3497 (
      {stage0_29[469]},
      {stage1_29[212]}
   );
   gpc1_1 gpc3498 (
      {stage0_29[470]},
      {stage1_29[213]}
   );
   gpc1_1 gpc3499 (
      {stage0_29[471]},
      {stage1_29[214]}
   );
   gpc1_1 gpc3500 (
      {stage0_29[472]},
      {stage1_29[215]}
   );
   gpc1_1 gpc3501 (
      {stage0_29[473]},
      {stage1_29[216]}
   );
   gpc1_1 gpc3502 (
      {stage0_29[474]},
      {stage1_29[217]}
   );
   gpc1_1 gpc3503 (
      {stage0_29[475]},
      {stage1_29[218]}
   );
   gpc1_1 gpc3504 (
      {stage0_29[476]},
      {stage1_29[219]}
   );
   gpc1_1 gpc3505 (
      {stage0_29[477]},
      {stage1_29[220]}
   );
   gpc1_1 gpc3506 (
      {stage0_29[478]},
      {stage1_29[221]}
   );
   gpc1_1 gpc3507 (
      {stage0_29[479]},
      {stage1_29[222]}
   );
   gpc1_1 gpc3508 (
      {stage0_29[480]},
      {stage1_29[223]}
   );
   gpc1_1 gpc3509 (
      {stage0_29[481]},
      {stage1_29[224]}
   );
   gpc1_1 gpc3510 (
      {stage0_29[482]},
      {stage1_29[225]}
   );
   gpc1_1 gpc3511 (
      {stage0_29[483]},
      {stage1_29[226]}
   );
   gpc1_1 gpc3512 (
      {stage0_29[484]},
      {stage1_29[227]}
   );
   gpc1_1 gpc3513 (
      {stage0_29[485]},
      {stage1_29[228]}
   );
   gpc1_1 gpc3514 (
      {stage0_30[460]},
      {stage1_30[166]}
   );
   gpc1_1 gpc3515 (
      {stage0_30[461]},
      {stage1_30[167]}
   );
   gpc1_1 gpc3516 (
      {stage0_30[462]},
      {stage1_30[168]}
   );
   gpc1_1 gpc3517 (
      {stage0_30[463]},
      {stage1_30[169]}
   );
   gpc1_1 gpc3518 (
      {stage0_30[464]},
      {stage1_30[170]}
   );
   gpc1_1 gpc3519 (
      {stage0_30[465]},
      {stage1_30[171]}
   );
   gpc1_1 gpc3520 (
      {stage0_30[466]},
      {stage1_30[172]}
   );
   gpc1_1 gpc3521 (
      {stage0_30[467]},
      {stage1_30[173]}
   );
   gpc1_1 gpc3522 (
      {stage0_30[468]},
      {stage1_30[174]}
   );
   gpc1_1 gpc3523 (
      {stage0_30[469]},
      {stage1_30[175]}
   );
   gpc1_1 gpc3524 (
      {stage0_30[470]},
      {stage1_30[176]}
   );
   gpc1_1 gpc3525 (
      {stage0_30[471]},
      {stage1_30[177]}
   );
   gpc1_1 gpc3526 (
      {stage0_30[472]},
      {stage1_30[178]}
   );
   gpc1_1 gpc3527 (
      {stage0_30[473]},
      {stage1_30[179]}
   );
   gpc1_1 gpc3528 (
      {stage0_30[474]},
      {stage1_30[180]}
   );
   gpc1_1 gpc3529 (
      {stage0_30[475]},
      {stage1_30[181]}
   );
   gpc1_1 gpc3530 (
      {stage0_30[476]},
      {stage1_30[182]}
   );
   gpc1_1 gpc3531 (
      {stage0_30[477]},
      {stage1_30[183]}
   );
   gpc1_1 gpc3532 (
      {stage0_30[478]},
      {stage1_30[184]}
   );
   gpc1_1 gpc3533 (
      {stage0_30[479]},
      {stage1_30[185]}
   );
   gpc1_1 gpc3534 (
      {stage0_30[480]},
      {stage1_30[186]}
   );
   gpc1_1 gpc3535 (
      {stage0_30[481]},
      {stage1_30[187]}
   );
   gpc1_1 gpc3536 (
      {stage0_30[482]},
      {stage1_30[188]}
   );
   gpc1_1 gpc3537 (
      {stage0_30[483]},
      {stage1_30[189]}
   );
   gpc1_1 gpc3538 (
      {stage0_30[484]},
      {stage1_30[190]}
   );
   gpc1_1 gpc3539 (
      {stage0_30[485]},
      {stage1_30[191]}
   );
   gpc1_1 gpc3540 (
      {stage0_31[476]},
      {stage1_31[208]}
   );
   gpc1_1 gpc3541 (
      {stage0_31[477]},
      {stage1_31[209]}
   );
   gpc1_1 gpc3542 (
      {stage0_31[478]},
      {stage1_31[210]}
   );
   gpc1_1 gpc3543 (
      {stage0_31[479]},
      {stage1_31[211]}
   );
   gpc1_1 gpc3544 (
      {stage0_31[480]},
      {stage1_31[212]}
   );
   gpc1_1 gpc3545 (
      {stage0_31[481]},
      {stage1_31[213]}
   );
   gpc1_1 gpc3546 (
      {stage0_31[482]},
      {stage1_31[214]}
   );
   gpc1_1 gpc3547 (
      {stage0_31[483]},
      {stage1_31[215]}
   );
   gpc1_1 gpc3548 (
      {stage0_31[484]},
      {stage1_31[216]}
   );
   gpc1_1 gpc3549 (
      {stage0_31[485]},
      {stage1_31[217]}
   );
   gpc1_1 gpc3550 (
      {stage0_33[396]},
      {stage1_33[169]}
   );
   gpc1_1 gpc3551 (
      {stage0_33[397]},
      {stage1_33[170]}
   );
   gpc1_1 gpc3552 (
      {stage0_33[398]},
      {stage1_33[171]}
   );
   gpc1_1 gpc3553 (
      {stage0_33[399]},
      {stage1_33[172]}
   );
   gpc1_1 gpc3554 (
      {stage0_33[400]},
      {stage1_33[173]}
   );
   gpc1_1 gpc3555 (
      {stage0_33[401]},
      {stage1_33[174]}
   );
   gpc1_1 gpc3556 (
      {stage0_33[402]},
      {stage1_33[175]}
   );
   gpc1_1 gpc3557 (
      {stage0_33[403]},
      {stage1_33[176]}
   );
   gpc1_1 gpc3558 (
      {stage0_33[404]},
      {stage1_33[177]}
   );
   gpc1_1 gpc3559 (
      {stage0_33[405]},
      {stage1_33[178]}
   );
   gpc1_1 gpc3560 (
      {stage0_33[406]},
      {stage1_33[179]}
   );
   gpc1_1 gpc3561 (
      {stage0_33[407]},
      {stage1_33[180]}
   );
   gpc1_1 gpc3562 (
      {stage0_33[408]},
      {stage1_33[181]}
   );
   gpc1_1 gpc3563 (
      {stage0_33[409]},
      {stage1_33[182]}
   );
   gpc1_1 gpc3564 (
      {stage0_33[410]},
      {stage1_33[183]}
   );
   gpc1_1 gpc3565 (
      {stage0_33[411]},
      {stage1_33[184]}
   );
   gpc1_1 gpc3566 (
      {stage0_33[412]},
      {stage1_33[185]}
   );
   gpc1_1 gpc3567 (
      {stage0_33[413]},
      {stage1_33[186]}
   );
   gpc1_1 gpc3568 (
      {stage0_33[414]},
      {stage1_33[187]}
   );
   gpc1_1 gpc3569 (
      {stage0_33[415]},
      {stage1_33[188]}
   );
   gpc1_1 gpc3570 (
      {stage0_33[416]},
      {stage1_33[189]}
   );
   gpc1_1 gpc3571 (
      {stage0_33[417]},
      {stage1_33[190]}
   );
   gpc1_1 gpc3572 (
      {stage0_33[418]},
      {stage1_33[191]}
   );
   gpc1_1 gpc3573 (
      {stage0_33[419]},
      {stage1_33[192]}
   );
   gpc1_1 gpc3574 (
      {stage0_33[420]},
      {stage1_33[193]}
   );
   gpc1_1 gpc3575 (
      {stage0_33[421]},
      {stage1_33[194]}
   );
   gpc1_1 gpc3576 (
      {stage0_33[422]},
      {stage1_33[195]}
   );
   gpc1_1 gpc3577 (
      {stage0_33[423]},
      {stage1_33[196]}
   );
   gpc1_1 gpc3578 (
      {stage0_33[424]},
      {stage1_33[197]}
   );
   gpc1_1 gpc3579 (
      {stage0_33[425]},
      {stage1_33[198]}
   );
   gpc1_1 gpc3580 (
      {stage0_33[426]},
      {stage1_33[199]}
   );
   gpc1_1 gpc3581 (
      {stage0_33[427]},
      {stage1_33[200]}
   );
   gpc1_1 gpc3582 (
      {stage0_33[428]},
      {stage1_33[201]}
   );
   gpc1_1 gpc3583 (
      {stage0_33[429]},
      {stage1_33[202]}
   );
   gpc1_1 gpc3584 (
      {stage0_33[430]},
      {stage1_33[203]}
   );
   gpc1_1 gpc3585 (
      {stage0_33[431]},
      {stage1_33[204]}
   );
   gpc1_1 gpc3586 (
      {stage0_33[432]},
      {stage1_33[205]}
   );
   gpc1_1 gpc3587 (
      {stage0_33[433]},
      {stage1_33[206]}
   );
   gpc1_1 gpc3588 (
      {stage0_33[434]},
      {stage1_33[207]}
   );
   gpc1_1 gpc3589 (
      {stage0_33[435]},
      {stage1_33[208]}
   );
   gpc1_1 gpc3590 (
      {stage0_33[436]},
      {stage1_33[209]}
   );
   gpc1_1 gpc3591 (
      {stage0_33[437]},
      {stage1_33[210]}
   );
   gpc1_1 gpc3592 (
      {stage0_33[438]},
      {stage1_33[211]}
   );
   gpc1_1 gpc3593 (
      {stage0_33[439]},
      {stage1_33[212]}
   );
   gpc1_1 gpc3594 (
      {stage0_33[440]},
      {stage1_33[213]}
   );
   gpc1_1 gpc3595 (
      {stage0_33[441]},
      {stage1_33[214]}
   );
   gpc1_1 gpc3596 (
      {stage0_33[442]},
      {stage1_33[215]}
   );
   gpc1_1 gpc3597 (
      {stage0_33[443]},
      {stage1_33[216]}
   );
   gpc1_1 gpc3598 (
      {stage0_33[444]},
      {stage1_33[217]}
   );
   gpc1_1 gpc3599 (
      {stage0_33[445]},
      {stage1_33[218]}
   );
   gpc1_1 gpc3600 (
      {stage0_33[446]},
      {stage1_33[219]}
   );
   gpc1_1 gpc3601 (
      {stage0_33[447]},
      {stage1_33[220]}
   );
   gpc1_1 gpc3602 (
      {stage0_33[448]},
      {stage1_33[221]}
   );
   gpc1_1 gpc3603 (
      {stage0_33[449]},
      {stage1_33[222]}
   );
   gpc1_1 gpc3604 (
      {stage0_33[450]},
      {stage1_33[223]}
   );
   gpc1_1 gpc3605 (
      {stage0_33[451]},
      {stage1_33[224]}
   );
   gpc1_1 gpc3606 (
      {stage0_33[452]},
      {stage1_33[225]}
   );
   gpc1_1 gpc3607 (
      {stage0_33[453]},
      {stage1_33[226]}
   );
   gpc1_1 gpc3608 (
      {stage0_33[454]},
      {stage1_33[227]}
   );
   gpc1_1 gpc3609 (
      {stage0_33[455]},
      {stage1_33[228]}
   );
   gpc1_1 gpc3610 (
      {stage0_33[456]},
      {stage1_33[229]}
   );
   gpc1_1 gpc3611 (
      {stage0_33[457]},
      {stage1_33[230]}
   );
   gpc1_1 gpc3612 (
      {stage0_33[458]},
      {stage1_33[231]}
   );
   gpc1_1 gpc3613 (
      {stage0_33[459]},
      {stage1_33[232]}
   );
   gpc1_1 gpc3614 (
      {stage0_33[460]},
      {stage1_33[233]}
   );
   gpc1_1 gpc3615 (
      {stage0_33[461]},
      {stage1_33[234]}
   );
   gpc1_1 gpc3616 (
      {stage0_33[462]},
      {stage1_33[235]}
   );
   gpc1_1 gpc3617 (
      {stage0_33[463]},
      {stage1_33[236]}
   );
   gpc1_1 gpc3618 (
      {stage0_33[464]},
      {stage1_33[237]}
   );
   gpc1_1 gpc3619 (
      {stage0_33[465]},
      {stage1_33[238]}
   );
   gpc1_1 gpc3620 (
      {stage0_33[466]},
      {stage1_33[239]}
   );
   gpc1_1 gpc3621 (
      {stage0_33[467]},
      {stage1_33[240]}
   );
   gpc1_1 gpc3622 (
      {stage0_33[468]},
      {stage1_33[241]}
   );
   gpc1_1 gpc3623 (
      {stage0_33[469]},
      {stage1_33[242]}
   );
   gpc1_1 gpc3624 (
      {stage0_33[470]},
      {stage1_33[243]}
   );
   gpc1_1 gpc3625 (
      {stage0_33[471]},
      {stage1_33[244]}
   );
   gpc1_1 gpc3626 (
      {stage0_33[472]},
      {stage1_33[245]}
   );
   gpc1_1 gpc3627 (
      {stage0_33[473]},
      {stage1_33[246]}
   );
   gpc1_1 gpc3628 (
      {stage0_33[474]},
      {stage1_33[247]}
   );
   gpc1_1 gpc3629 (
      {stage0_33[475]},
      {stage1_33[248]}
   );
   gpc1_1 gpc3630 (
      {stage0_33[476]},
      {stage1_33[249]}
   );
   gpc1_1 gpc3631 (
      {stage0_33[477]},
      {stage1_33[250]}
   );
   gpc1_1 gpc3632 (
      {stage0_33[478]},
      {stage1_33[251]}
   );
   gpc1_1 gpc3633 (
      {stage0_33[479]},
      {stage1_33[252]}
   );
   gpc1_1 gpc3634 (
      {stage0_33[480]},
      {stage1_33[253]}
   );
   gpc1_1 gpc3635 (
      {stage0_33[481]},
      {stage1_33[254]}
   );
   gpc1_1 gpc3636 (
      {stage0_33[482]},
      {stage1_33[255]}
   );
   gpc1_1 gpc3637 (
      {stage0_33[483]},
      {stage1_33[256]}
   );
   gpc1_1 gpc3638 (
      {stage0_33[484]},
      {stage1_33[257]}
   );
   gpc1_1 gpc3639 (
      {stage0_33[485]},
      {stage1_33[258]}
   );
   gpc1_1 gpc3640 (
      {stage0_35[464]},
      {stage1_35[195]}
   );
   gpc1_1 gpc3641 (
      {stage0_35[465]},
      {stage1_35[196]}
   );
   gpc1_1 gpc3642 (
      {stage0_35[466]},
      {stage1_35[197]}
   );
   gpc1_1 gpc3643 (
      {stage0_35[467]},
      {stage1_35[198]}
   );
   gpc1_1 gpc3644 (
      {stage0_35[468]},
      {stage1_35[199]}
   );
   gpc1_1 gpc3645 (
      {stage0_35[469]},
      {stage1_35[200]}
   );
   gpc1_1 gpc3646 (
      {stage0_35[470]},
      {stage1_35[201]}
   );
   gpc1_1 gpc3647 (
      {stage0_35[471]},
      {stage1_35[202]}
   );
   gpc1_1 gpc3648 (
      {stage0_35[472]},
      {stage1_35[203]}
   );
   gpc1_1 gpc3649 (
      {stage0_35[473]},
      {stage1_35[204]}
   );
   gpc1_1 gpc3650 (
      {stage0_35[474]},
      {stage1_35[205]}
   );
   gpc1_1 gpc3651 (
      {stage0_35[475]},
      {stage1_35[206]}
   );
   gpc1_1 gpc3652 (
      {stage0_35[476]},
      {stage1_35[207]}
   );
   gpc1_1 gpc3653 (
      {stage0_35[477]},
      {stage1_35[208]}
   );
   gpc1_1 gpc3654 (
      {stage0_35[478]},
      {stage1_35[209]}
   );
   gpc1_1 gpc3655 (
      {stage0_35[479]},
      {stage1_35[210]}
   );
   gpc1_1 gpc3656 (
      {stage0_35[480]},
      {stage1_35[211]}
   );
   gpc1_1 gpc3657 (
      {stage0_35[481]},
      {stage1_35[212]}
   );
   gpc1_1 gpc3658 (
      {stage0_35[482]},
      {stage1_35[213]}
   );
   gpc1_1 gpc3659 (
      {stage0_35[483]},
      {stage1_35[214]}
   );
   gpc1_1 gpc3660 (
      {stage0_35[484]},
      {stage1_35[215]}
   );
   gpc1_1 gpc3661 (
      {stage0_35[485]},
      {stage1_35[216]}
   );
   gpc1_1 gpc3662 (
      {stage0_37[355]},
      {stage1_37[177]}
   );
   gpc1_1 gpc3663 (
      {stage0_37[356]},
      {stage1_37[178]}
   );
   gpc1_1 gpc3664 (
      {stage0_37[357]},
      {stage1_37[179]}
   );
   gpc1_1 gpc3665 (
      {stage0_37[358]},
      {stage1_37[180]}
   );
   gpc1_1 gpc3666 (
      {stage0_37[359]},
      {stage1_37[181]}
   );
   gpc1_1 gpc3667 (
      {stage0_37[360]},
      {stage1_37[182]}
   );
   gpc1_1 gpc3668 (
      {stage0_37[361]},
      {stage1_37[183]}
   );
   gpc1_1 gpc3669 (
      {stage0_37[362]},
      {stage1_37[184]}
   );
   gpc1_1 gpc3670 (
      {stage0_37[363]},
      {stage1_37[185]}
   );
   gpc1_1 gpc3671 (
      {stage0_37[364]},
      {stage1_37[186]}
   );
   gpc1_1 gpc3672 (
      {stage0_37[365]},
      {stage1_37[187]}
   );
   gpc1_1 gpc3673 (
      {stage0_37[366]},
      {stage1_37[188]}
   );
   gpc1_1 gpc3674 (
      {stage0_37[367]},
      {stage1_37[189]}
   );
   gpc1_1 gpc3675 (
      {stage0_37[368]},
      {stage1_37[190]}
   );
   gpc1_1 gpc3676 (
      {stage0_37[369]},
      {stage1_37[191]}
   );
   gpc1_1 gpc3677 (
      {stage0_37[370]},
      {stage1_37[192]}
   );
   gpc1_1 gpc3678 (
      {stage0_37[371]},
      {stage1_37[193]}
   );
   gpc1_1 gpc3679 (
      {stage0_37[372]},
      {stage1_37[194]}
   );
   gpc1_1 gpc3680 (
      {stage0_37[373]},
      {stage1_37[195]}
   );
   gpc1_1 gpc3681 (
      {stage0_37[374]},
      {stage1_37[196]}
   );
   gpc1_1 gpc3682 (
      {stage0_37[375]},
      {stage1_37[197]}
   );
   gpc1_1 gpc3683 (
      {stage0_37[376]},
      {stage1_37[198]}
   );
   gpc1_1 gpc3684 (
      {stage0_37[377]},
      {stage1_37[199]}
   );
   gpc1_1 gpc3685 (
      {stage0_37[378]},
      {stage1_37[200]}
   );
   gpc1_1 gpc3686 (
      {stage0_37[379]},
      {stage1_37[201]}
   );
   gpc1_1 gpc3687 (
      {stage0_37[380]},
      {stage1_37[202]}
   );
   gpc1_1 gpc3688 (
      {stage0_37[381]},
      {stage1_37[203]}
   );
   gpc1_1 gpc3689 (
      {stage0_37[382]},
      {stage1_37[204]}
   );
   gpc1_1 gpc3690 (
      {stage0_37[383]},
      {stage1_37[205]}
   );
   gpc1_1 gpc3691 (
      {stage0_37[384]},
      {stage1_37[206]}
   );
   gpc1_1 gpc3692 (
      {stage0_37[385]},
      {stage1_37[207]}
   );
   gpc1_1 gpc3693 (
      {stage0_37[386]},
      {stage1_37[208]}
   );
   gpc1_1 gpc3694 (
      {stage0_37[387]},
      {stage1_37[209]}
   );
   gpc1_1 gpc3695 (
      {stage0_37[388]},
      {stage1_37[210]}
   );
   gpc1_1 gpc3696 (
      {stage0_37[389]},
      {stage1_37[211]}
   );
   gpc1_1 gpc3697 (
      {stage0_37[390]},
      {stage1_37[212]}
   );
   gpc1_1 gpc3698 (
      {stage0_37[391]},
      {stage1_37[213]}
   );
   gpc1_1 gpc3699 (
      {stage0_37[392]},
      {stage1_37[214]}
   );
   gpc1_1 gpc3700 (
      {stage0_37[393]},
      {stage1_37[215]}
   );
   gpc1_1 gpc3701 (
      {stage0_37[394]},
      {stage1_37[216]}
   );
   gpc1_1 gpc3702 (
      {stage0_37[395]},
      {stage1_37[217]}
   );
   gpc1_1 gpc3703 (
      {stage0_37[396]},
      {stage1_37[218]}
   );
   gpc1_1 gpc3704 (
      {stage0_37[397]},
      {stage1_37[219]}
   );
   gpc1_1 gpc3705 (
      {stage0_37[398]},
      {stage1_37[220]}
   );
   gpc1_1 gpc3706 (
      {stage0_37[399]},
      {stage1_37[221]}
   );
   gpc1_1 gpc3707 (
      {stage0_37[400]},
      {stage1_37[222]}
   );
   gpc1_1 gpc3708 (
      {stage0_37[401]},
      {stage1_37[223]}
   );
   gpc1_1 gpc3709 (
      {stage0_37[402]},
      {stage1_37[224]}
   );
   gpc1_1 gpc3710 (
      {stage0_37[403]},
      {stage1_37[225]}
   );
   gpc1_1 gpc3711 (
      {stage0_37[404]},
      {stage1_37[226]}
   );
   gpc1_1 gpc3712 (
      {stage0_37[405]},
      {stage1_37[227]}
   );
   gpc1_1 gpc3713 (
      {stage0_37[406]},
      {stage1_37[228]}
   );
   gpc1_1 gpc3714 (
      {stage0_37[407]},
      {stage1_37[229]}
   );
   gpc1_1 gpc3715 (
      {stage0_37[408]},
      {stage1_37[230]}
   );
   gpc1_1 gpc3716 (
      {stage0_37[409]},
      {stage1_37[231]}
   );
   gpc1_1 gpc3717 (
      {stage0_37[410]},
      {stage1_37[232]}
   );
   gpc1_1 gpc3718 (
      {stage0_37[411]},
      {stage1_37[233]}
   );
   gpc1_1 gpc3719 (
      {stage0_37[412]},
      {stage1_37[234]}
   );
   gpc1_1 gpc3720 (
      {stage0_37[413]},
      {stage1_37[235]}
   );
   gpc1_1 gpc3721 (
      {stage0_37[414]},
      {stage1_37[236]}
   );
   gpc1_1 gpc3722 (
      {stage0_37[415]},
      {stage1_37[237]}
   );
   gpc1_1 gpc3723 (
      {stage0_37[416]},
      {stage1_37[238]}
   );
   gpc1_1 gpc3724 (
      {stage0_37[417]},
      {stage1_37[239]}
   );
   gpc1_1 gpc3725 (
      {stage0_37[418]},
      {stage1_37[240]}
   );
   gpc1_1 gpc3726 (
      {stage0_37[419]},
      {stage1_37[241]}
   );
   gpc1_1 gpc3727 (
      {stage0_37[420]},
      {stage1_37[242]}
   );
   gpc1_1 gpc3728 (
      {stage0_37[421]},
      {stage1_37[243]}
   );
   gpc1_1 gpc3729 (
      {stage0_37[422]},
      {stage1_37[244]}
   );
   gpc1_1 gpc3730 (
      {stage0_37[423]},
      {stage1_37[245]}
   );
   gpc1_1 gpc3731 (
      {stage0_37[424]},
      {stage1_37[246]}
   );
   gpc1_1 gpc3732 (
      {stage0_37[425]},
      {stage1_37[247]}
   );
   gpc1_1 gpc3733 (
      {stage0_37[426]},
      {stage1_37[248]}
   );
   gpc1_1 gpc3734 (
      {stage0_37[427]},
      {stage1_37[249]}
   );
   gpc1_1 gpc3735 (
      {stage0_37[428]},
      {stage1_37[250]}
   );
   gpc1_1 gpc3736 (
      {stage0_37[429]},
      {stage1_37[251]}
   );
   gpc1_1 gpc3737 (
      {stage0_37[430]},
      {stage1_37[252]}
   );
   gpc1_1 gpc3738 (
      {stage0_37[431]},
      {stage1_37[253]}
   );
   gpc1_1 gpc3739 (
      {stage0_37[432]},
      {stage1_37[254]}
   );
   gpc1_1 gpc3740 (
      {stage0_37[433]},
      {stage1_37[255]}
   );
   gpc1_1 gpc3741 (
      {stage0_37[434]},
      {stage1_37[256]}
   );
   gpc1_1 gpc3742 (
      {stage0_37[435]},
      {stage1_37[257]}
   );
   gpc1_1 gpc3743 (
      {stage0_37[436]},
      {stage1_37[258]}
   );
   gpc1_1 gpc3744 (
      {stage0_37[437]},
      {stage1_37[259]}
   );
   gpc1_1 gpc3745 (
      {stage0_37[438]},
      {stage1_37[260]}
   );
   gpc1_1 gpc3746 (
      {stage0_37[439]},
      {stage1_37[261]}
   );
   gpc1_1 gpc3747 (
      {stage0_37[440]},
      {stage1_37[262]}
   );
   gpc1_1 gpc3748 (
      {stage0_37[441]},
      {stage1_37[263]}
   );
   gpc1_1 gpc3749 (
      {stage0_37[442]},
      {stage1_37[264]}
   );
   gpc1_1 gpc3750 (
      {stage0_37[443]},
      {stage1_37[265]}
   );
   gpc1_1 gpc3751 (
      {stage0_37[444]},
      {stage1_37[266]}
   );
   gpc1_1 gpc3752 (
      {stage0_37[445]},
      {stage1_37[267]}
   );
   gpc1_1 gpc3753 (
      {stage0_37[446]},
      {stage1_37[268]}
   );
   gpc1_1 gpc3754 (
      {stage0_37[447]},
      {stage1_37[269]}
   );
   gpc1_1 gpc3755 (
      {stage0_37[448]},
      {stage1_37[270]}
   );
   gpc1_1 gpc3756 (
      {stage0_37[449]},
      {stage1_37[271]}
   );
   gpc1_1 gpc3757 (
      {stage0_37[450]},
      {stage1_37[272]}
   );
   gpc1_1 gpc3758 (
      {stage0_37[451]},
      {stage1_37[273]}
   );
   gpc1_1 gpc3759 (
      {stage0_37[452]},
      {stage1_37[274]}
   );
   gpc1_1 gpc3760 (
      {stage0_37[453]},
      {stage1_37[275]}
   );
   gpc1_1 gpc3761 (
      {stage0_37[454]},
      {stage1_37[276]}
   );
   gpc1_1 gpc3762 (
      {stage0_37[455]},
      {stage1_37[277]}
   );
   gpc1_1 gpc3763 (
      {stage0_37[456]},
      {stage1_37[278]}
   );
   gpc1_1 gpc3764 (
      {stage0_37[457]},
      {stage1_37[279]}
   );
   gpc1_1 gpc3765 (
      {stage0_37[458]},
      {stage1_37[280]}
   );
   gpc1_1 gpc3766 (
      {stage0_37[459]},
      {stage1_37[281]}
   );
   gpc1_1 gpc3767 (
      {stage0_37[460]},
      {stage1_37[282]}
   );
   gpc1_1 gpc3768 (
      {stage0_37[461]},
      {stage1_37[283]}
   );
   gpc1_1 gpc3769 (
      {stage0_37[462]},
      {stage1_37[284]}
   );
   gpc1_1 gpc3770 (
      {stage0_37[463]},
      {stage1_37[285]}
   );
   gpc1_1 gpc3771 (
      {stage0_37[464]},
      {stage1_37[286]}
   );
   gpc1_1 gpc3772 (
      {stage0_37[465]},
      {stage1_37[287]}
   );
   gpc1_1 gpc3773 (
      {stage0_37[466]},
      {stage1_37[288]}
   );
   gpc1_1 gpc3774 (
      {stage0_37[467]},
      {stage1_37[289]}
   );
   gpc1_1 gpc3775 (
      {stage0_37[468]},
      {stage1_37[290]}
   );
   gpc1_1 gpc3776 (
      {stage0_37[469]},
      {stage1_37[291]}
   );
   gpc1_1 gpc3777 (
      {stage0_37[470]},
      {stage1_37[292]}
   );
   gpc1_1 gpc3778 (
      {stage0_37[471]},
      {stage1_37[293]}
   );
   gpc1_1 gpc3779 (
      {stage0_37[472]},
      {stage1_37[294]}
   );
   gpc1_1 gpc3780 (
      {stage0_37[473]},
      {stage1_37[295]}
   );
   gpc1_1 gpc3781 (
      {stage0_37[474]},
      {stage1_37[296]}
   );
   gpc1_1 gpc3782 (
      {stage0_37[475]},
      {stage1_37[297]}
   );
   gpc1_1 gpc3783 (
      {stage0_37[476]},
      {stage1_37[298]}
   );
   gpc1_1 gpc3784 (
      {stage0_37[477]},
      {stage1_37[299]}
   );
   gpc1_1 gpc3785 (
      {stage0_37[478]},
      {stage1_37[300]}
   );
   gpc1_1 gpc3786 (
      {stage0_37[479]},
      {stage1_37[301]}
   );
   gpc1_1 gpc3787 (
      {stage0_37[480]},
      {stage1_37[302]}
   );
   gpc1_1 gpc3788 (
      {stage0_37[481]},
      {stage1_37[303]}
   );
   gpc1_1 gpc3789 (
      {stage0_37[482]},
      {stage1_37[304]}
   );
   gpc1_1 gpc3790 (
      {stage0_37[483]},
      {stage1_37[305]}
   );
   gpc1_1 gpc3791 (
      {stage0_37[484]},
      {stage1_37[306]}
   );
   gpc1_1 gpc3792 (
      {stage0_37[485]},
      {stage1_37[307]}
   );
   gpc1_1 gpc3793 (
      {stage0_38[391]},
      {stage1_38[170]}
   );
   gpc1_1 gpc3794 (
      {stage0_38[392]},
      {stage1_38[171]}
   );
   gpc1_1 gpc3795 (
      {stage0_38[393]},
      {stage1_38[172]}
   );
   gpc1_1 gpc3796 (
      {stage0_38[394]},
      {stage1_38[173]}
   );
   gpc1_1 gpc3797 (
      {stage0_38[395]},
      {stage1_38[174]}
   );
   gpc1_1 gpc3798 (
      {stage0_38[396]},
      {stage1_38[175]}
   );
   gpc1_1 gpc3799 (
      {stage0_38[397]},
      {stage1_38[176]}
   );
   gpc1_1 gpc3800 (
      {stage0_38[398]},
      {stage1_38[177]}
   );
   gpc1_1 gpc3801 (
      {stage0_38[399]},
      {stage1_38[178]}
   );
   gpc1_1 gpc3802 (
      {stage0_38[400]},
      {stage1_38[179]}
   );
   gpc1_1 gpc3803 (
      {stage0_38[401]},
      {stage1_38[180]}
   );
   gpc1_1 gpc3804 (
      {stage0_38[402]},
      {stage1_38[181]}
   );
   gpc1_1 gpc3805 (
      {stage0_38[403]},
      {stage1_38[182]}
   );
   gpc1_1 gpc3806 (
      {stage0_38[404]},
      {stage1_38[183]}
   );
   gpc1_1 gpc3807 (
      {stage0_38[405]},
      {stage1_38[184]}
   );
   gpc1_1 gpc3808 (
      {stage0_38[406]},
      {stage1_38[185]}
   );
   gpc1_1 gpc3809 (
      {stage0_38[407]},
      {stage1_38[186]}
   );
   gpc1_1 gpc3810 (
      {stage0_38[408]},
      {stage1_38[187]}
   );
   gpc1_1 gpc3811 (
      {stage0_38[409]},
      {stage1_38[188]}
   );
   gpc1_1 gpc3812 (
      {stage0_38[410]},
      {stage1_38[189]}
   );
   gpc1_1 gpc3813 (
      {stage0_38[411]},
      {stage1_38[190]}
   );
   gpc1_1 gpc3814 (
      {stage0_38[412]},
      {stage1_38[191]}
   );
   gpc1_1 gpc3815 (
      {stage0_38[413]},
      {stage1_38[192]}
   );
   gpc1_1 gpc3816 (
      {stage0_38[414]},
      {stage1_38[193]}
   );
   gpc1_1 gpc3817 (
      {stage0_38[415]},
      {stage1_38[194]}
   );
   gpc1_1 gpc3818 (
      {stage0_38[416]},
      {stage1_38[195]}
   );
   gpc1_1 gpc3819 (
      {stage0_38[417]},
      {stage1_38[196]}
   );
   gpc1_1 gpc3820 (
      {stage0_38[418]},
      {stage1_38[197]}
   );
   gpc1_1 gpc3821 (
      {stage0_38[419]},
      {stage1_38[198]}
   );
   gpc1_1 gpc3822 (
      {stage0_38[420]},
      {stage1_38[199]}
   );
   gpc1_1 gpc3823 (
      {stage0_38[421]},
      {stage1_38[200]}
   );
   gpc1_1 gpc3824 (
      {stage0_38[422]},
      {stage1_38[201]}
   );
   gpc1_1 gpc3825 (
      {stage0_38[423]},
      {stage1_38[202]}
   );
   gpc1_1 gpc3826 (
      {stage0_38[424]},
      {stage1_38[203]}
   );
   gpc1_1 gpc3827 (
      {stage0_38[425]},
      {stage1_38[204]}
   );
   gpc1_1 gpc3828 (
      {stage0_38[426]},
      {stage1_38[205]}
   );
   gpc1_1 gpc3829 (
      {stage0_38[427]},
      {stage1_38[206]}
   );
   gpc1_1 gpc3830 (
      {stage0_38[428]},
      {stage1_38[207]}
   );
   gpc1_1 gpc3831 (
      {stage0_38[429]},
      {stage1_38[208]}
   );
   gpc1_1 gpc3832 (
      {stage0_38[430]},
      {stage1_38[209]}
   );
   gpc1_1 gpc3833 (
      {stage0_38[431]},
      {stage1_38[210]}
   );
   gpc1_1 gpc3834 (
      {stage0_38[432]},
      {stage1_38[211]}
   );
   gpc1_1 gpc3835 (
      {stage0_38[433]},
      {stage1_38[212]}
   );
   gpc1_1 gpc3836 (
      {stage0_38[434]},
      {stage1_38[213]}
   );
   gpc1_1 gpc3837 (
      {stage0_38[435]},
      {stage1_38[214]}
   );
   gpc1_1 gpc3838 (
      {stage0_38[436]},
      {stage1_38[215]}
   );
   gpc1_1 gpc3839 (
      {stage0_38[437]},
      {stage1_38[216]}
   );
   gpc1_1 gpc3840 (
      {stage0_38[438]},
      {stage1_38[217]}
   );
   gpc1_1 gpc3841 (
      {stage0_38[439]},
      {stage1_38[218]}
   );
   gpc1_1 gpc3842 (
      {stage0_38[440]},
      {stage1_38[219]}
   );
   gpc1_1 gpc3843 (
      {stage0_38[441]},
      {stage1_38[220]}
   );
   gpc1_1 gpc3844 (
      {stage0_38[442]},
      {stage1_38[221]}
   );
   gpc1_1 gpc3845 (
      {stage0_38[443]},
      {stage1_38[222]}
   );
   gpc1_1 gpc3846 (
      {stage0_38[444]},
      {stage1_38[223]}
   );
   gpc1_1 gpc3847 (
      {stage0_38[445]},
      {stage1_38[224]}
   );
   gpc1_1 gpc3848 (
      {stage0_38[446]},
      {stage1_38[225]}
   );
   gpc1_1 gpc3849 (
      {stage0_38[447]},
      {stage1_38[226]}
   );
   gpc1_1 gpc3850 (
      {stage0_38[448]},
      {stage1_38[227]}
   );
   gpc1_1 gpc3851 (
      {stage0_38[449]},
      {stage1_38[228]}
   );
   gpc1_1 gpc3852 (
      {stage0_38[450]},
      {stage1_38[229]}
   );
   gpc1_1 gpc3853 (
      {stage0_38[451]},
      {stage1_38[230]}
   );
   gpc1_1 gpc3854 (
      {stage0_38[452]},
      {stage1_38[231]}
   );
   gpc1_1 gpc3855 (
      {stage0_38[453]},
      {stage1_38[232]}
   );
   gpc1_1 gpc3856 (
      {stage0_38[454]},
      {stage1_38[233]}
   );
   gpc1_1 gpc3857 (
      {stage0_38[455]},
      {stage1_38[234]}
   );
   gpc1_1 gpc3858 (
      {stage0_38[456]},
      {stage1_38[235]}
   );
   gpc1_1 gpc3859 (
      {stage0_38[457]},
      {stage1_38[236]}
   );
   gpc1_1 gpc3860 (
      {stage0_38[458]},
      {stage1_38[237]}
   );
   gpc1_1 gpc3861 (
      {stage0_38[459]},
      {stage1_38[238]}
   );
   gpc1_1 gpc3862 (
      {stage0_38[460]},
      {stage1_38[239]}
   );
   gpc1_1 gpc3863 (
      {stage0_38[461]},
      {stage1_38[240]}
   );
   gpc1_1 gpc3864 (
      {stage0_38[462]},
      {stage1_38[241]}
   );
   gpc1_1 gpc3865 (
      {stage0_38[463]},
      {stage1_38[242]}
   );
   gpc1_1 gpc3866 (
      {stage0_38[464]},
      {stage1_38[243]}
   );
   gpc1_1 gpc3867 (
      {stage0_38[465]},
      {stage1_38[244]}
   );
   gpc1_1 gpc3868 (
      {stage0_38[466]},
      {stage1_38[245]}
   );
   gpc1_1 gpc3869 (
      {stage0_38[467]},
      {stage1_38[246]}
   );
   gpc1_1 gpc3870 (
      {stage0_38[468]},
      {stage1_38[247]}
   );
   gpc1_1 gpc3871 (
      {stage0_38[469]},
      {stage1_38[248]}
   );
   gpc1_1 gpc3872 (
      {stage0_38[470]},
      {stage1_38[249]}
   );
   gpc1_1 gpc3873 (
      {stage0_38[471]},
      {stage1_38[250]}
   );
   gpc1_1 gpc3874 (
      {stage0_38[472]},
      {stage1_38[251]}
   );
   gpc1_1 gpc3875 (
      {stage0_38[473]},
      {stage1_38[252]}
   );
   gpc1_1 gpc3876 (
      {stage0_38[474]},
      {stage1_38[253]}
   );
   gpc1_1 gpc3877 (
      {stage0_38[475]},
      {stage1_38[254]}
   );
   gpc1_1 gpc3878 (
      {stage0_38[476]},
      {stage1_38[255]}
   );
   gpc1_1 gpc3879 (
      {stage0_38[477]},
      {stage1_38[256]}
   );
   gpc1_1 gpc3880 (
      {stage0_38[478]},
      {stage1_38[257]}
   );
   gpc1_1 gpc3881 (
      {stage0_38[479]},
      {stage1_38[258]}
   );
   gpc1_1 gpc3882 (
      {stage0_38[480]},
      {stage1_38[259]}
   );
   gpc1_1 gpc3883 (
      {stage0_38[481]},
      {stage1_38[260]}
   );
   gpc1_1 gpc3884 (
      {stage0_38[482]},
      {stage1_38[261]}
   );
   gpc1_1 gpc3885 (
      {stage0_38[483]},
      {stage1_38[262]}
   );
   gpc1_1 gpc3886 (
      {stage0_38[484]},
      {stage1_38[263]}
   );
   gpc1_1 gpc3887 (
      {stage0_38[485]},
      {stage1_38[264]}
   );
   gpc1_1 gpc3888 (
      {stage0_39[447]},
      {stage1_39[174]}
   );
   gpc1_1 gpc3889 (
      {stage0_39[448]},
      {stage1_39[175]}
   );
   gpc1_1 gpc3890 (
      {stage0_39[449]},
      {stage1_39[176]}
   );
   gpc1_1 gpc3891 (
      {stage0_39[450]},
      {stage1_39[177]}
   );
   gpc1_1 gpc3892 (
      {stage0_39[451]},
      {stage1_39[178]}
   );
   gpc1_1 gpc3893 (
      {stage0_39[452]},
      {stage1_39[179]}
   );
   gpc1_1 gpc3894 (
      {stage0_39[453]},
      {stage1_39[180]}
   );
   gpc1_1 gpc3895 (
      {stage0_39[454]},
      {stage1_39[181]}
   );
   gpc1_1 gpc3896 (
      {stage0_39[455]},
      {stage1_39[182]}
   );
   gpc1_1 gpc3897 (
      {stage0_39[456]},
      {stage1_39[183]}
   );
   gpc1_1 gpc3898 (
      {stage0_39[457]},
      {stage1_39[184]}
   );
   gpc1_1 gpc3899 (
      {stage0_39[458]},
      {stage1_39[185]}
   );
   gpc1_1 gpc3900 (
      {stage0_39[459]},
      {stage1_39[186]}
   );
   gpc1_1 gpc3901 (
      {stage0_39[460]},
      {stage1_39[187]}
   );
   gpc1_1 gpc3902 (
      {stage0_39[461]},
      {stage1_39[188]}
   );
   gpc1_1 gpc3903 (
      {stage0_39[462]},
      {stage1_39[189]}
   );
   gpc1_1 gpc3904 (
      {stage0_39[463]},
      {stage1_39[190]}
   );
   gpc1_1 gpc3905 (
      {stage0_39[464]},
      {stage1_39[191]}
   );
   gpc1_1 gpc3906 (
      {stage0_39[465]},
      {stage1_39[192]}
   );
   gpc1_1 gpc3907 (
      {stage0_39[466]},
      {stage1_39[193]}
   );
   gpc1_1 gpc3908 (
      {stage0_39[467]},
      {stage1_39[194]}
   );
   gpc1_1 gpc3909 (
      {stage0_39[468]},
      {stage1_39[195]}
   );
   gpc1_1 gpc3910 (
      {stage0_39[469]},
      {stage1_39[196]}
   );
   gpc1_1 gpc3911 (
      {stage0_39[470]},
      {stage1_39[197]}
   );
   gpc1_1 gpc3912 (
      {stage0_39[471]},
      {stage1_39[198]}
   );
   gpc1_1 gpc3913 (
      {stage0_39[472]},
      {stage1_39[199]}
   );
   gpc1_1 gpc3914 (
      {stage0_39[473]},
      {stage1_39[200]}
   );
   gpc1_1 gpc3915 (
      {stage0_39[474]},
      {stage1_39[201]}
   );
   gpc1_1 gpc3916 (
      {stage0_39[475]},
      {stage1_39[202]}
   );
   gpc1_1 gpc3917 (
      {stage0_39[476]},
      {stage1_39[203]}
   );
   gpc1_1 gpc3918 (
      {stage0_39[477]},
      {stage1_39[204]}
   );
   gpc1_1 gpc3919 (
      {stage0_39[478]},
      {stage1_39[205]}
   );
   gpc1_1 gpc3920 (
      {stage0_39[479]},
      {stage1_39[206]}
   );
   gpc1_1 gpc3921 (
      {stage0_39[480]},
      {stage1_39[207]}
   );
   gpc1_1 gpc3922 (
      {stage0_39[481]},
      {stage1_39[208]}
   );
   gpc1_1 gpc3923 (
      {stage0_39[482]},
      {stage1_39[209]}
   );
   gpc1_1 gpc3924 (
      {stage0_39[483]},
      {stage1_39[210]}
   );
   gpc1_1 gpc3925 (
      {stage0_39[484]},
      {stage1_39[211]}
   );
   gpc1_1 gpc3926 (
      {stage0_39[485]},
      {stage1_39[212]}
   );
   gpc1_1 gpc3927 (
      {stage0_40[380]},
      {stage1_40[198]}
   );
   gpc1_1 gpc3928 (
      {stage0_40[381]},
      {stage1_40[199]}
   );
   gpc1_1 gpc3929 (
      {stage0_40[382]},
      {stage1_40[200]}
   );
   gpc1_1 gpc3930 (
      {stage0_40[383]},
      {stage1_40[201]}
   );
   gpc1_1 gpc3931 (
      {stage0_40[384]},
      {stage1_40[202]}
   );
   gpc1_1 gpc3932 (
      {stage0_40[385]},
      {stage1_40[203]}
   );
   gpc1_1 gpc3933 (
      {stage0_40[386]},
      {stage1_40[204]}
   );
   gpc1_1 gpc3934 (
      {stage0_40[387]},
      {stage1_40[205]}
   );
   gpc1_1 gpc3935 (
      {stage0_40[388]},
      {stage1_40[206]}
   );
   gpc1_1 gpc3936 (
      {stage0_40[389]},
      {stage1_40[207]}
   );
   gpc1_1 gpc3937 (
      {stage0_40[390]},
      {stage1_40[208]}
   );
   gpc1_1 gpc3938 (
      {stage0_40[391]},
      {stage1_40[209]}
   );
   gpc1_1 gpc3939 (
      {stage0_40[392]},
      {stage1_40[210]}
   );
   gpc1_1 gpc3940 (
      {stage0_40[393]},
      {stage1_40[211]}
   );
   gpc1_1 gpc3941 (
      {stage0_40[394]},
      {stage1_40[212]}
   );
   gpc1_1 gpc3942 (
      {stage0_40[395]},
      {stage1_40[213]}
   );
   gpc1_1 gpc3943 (
      {stage0_40[396]},
      {stage1_40[214]}
   );
   gpc1_1 gpc3944 (
      {stage0_40[397]},
      {stage1_40[215]}
   );
   gpc1_1 gpc3945 (
      {stage0_40[398]},
      {stage1_40[216]}
   );
   gpc1_1 gpc3946 (
      {stage0_40[399]},
      {stage1_40[217]}
   );
   gpc1_1 gpc3947 (
      {stage0_40[400]},
      {stage1_40[218]}
   );
   gpc1_1 gpc3948 (
      {stage0_40[401]},
      {stage1_40[219]}
   );
   gpc1_1 gpc3949 (
      {stage0_40[402]},
      {stage1_40[220]}
   );
   gpc1_1 gpc3950 (
      {stage0_40[403]},
      {stage1_40[221]}
   );
   gpc1_1 gpc3951 (
      {stage0_40[404]},
      {stage1_40[222]}
   );
   gpc1_1 gpc3952 (
      {stage0_40[405]},
      {stage1_40[223]}
   );
   gpc1_1 gpc3953 (
      {stage0_40[406]},
      {stage1_40[224]}
   );
   gpc1_1 gpc3954 (
      {stage0_40[407]},
      {stage1_40[225]}
   );
   gpc1_1 gpc3955 (
      {stage0_40[408]},
      {stage1_40[226]}
   );
   gpc1_1 gpc3956 (
      {stage0_40[409]},
      {stage1_40[227]}
   );
   gpc1_1 gpc3957 (
      {stage0_40[410]},
      {stage1_40[228]}
   );
   gpc1_1 gpc3958 (
      {stage0_40[411]},
      {stage1_40[229]}
   );
   gpc1_1 gpc3959 (
      {stage0_40[412]},
      {stage1_40[230]}
   );
   gpc1_1 gpc3960 (
      {stage0_40[413]},
      {stage1_40[231]}
   );
   gpc1_1 gpc3961 (
      {stage0_40[414]},
      {stage1_40[232]}
   );
   gpc1_1 gpc3962 (
      {stage0_40[415]},
      {stage1_40[233]}
   );
   gpc1_1 gpc3963 (
      {stage0_40[416]},
      {stage1_40[234]}
   );
   gpc1_1 gpc3964 (
      {stage0_40[417]},
      {stage1_40[235]}
   );
   gpc1_1 gpc3965 (
      {stage0_40[418]},
      {stage1_40[236]}
   );
   gpc1_1 gpc3966 (
      {stage0_40[419]},
      {stage1_40[237]}
   );
   gpc1_1 gpc3967 (
      {stage0_40[420]},
      {stage1_40[238]}
   );
   gpc1_1 gpc3968 (
      {stage0_40[421]},
      {stage1_40[239]}
   );
   gpc1_1 gpc3969 (
      {stage0_40[422]},
      {stage1_40[240]}
   );
   gpc1_1 gpc3970 (
      {stage0_40[423]},
      {stage1_40[241]}
   );
   gpc1_1 gpc3971 (
      {stage0_40[424]},
      {stage1_40[242]}
   );
   gpc1_1 gpc3972 (
      {stage0_40[425]},
      {stage1_40[243]}
   );
   gpc1_1 gpc3973 (
      {stage0_40[426]},
      {stage1_40[244]}
   );
   gpc1_1 gpc3974 (
      {stage0_40[427]},
      {stage1_40[245]}
   );
   gpc1_1 gpc3975 (
      {stage0_40[428]},
      {stage1_40[246]}
   );
   gpc1_1 gpc3976 (
      {stage0_40[429]},
      {stage1_40[247]}
   );
   gpc1_1 gpc3977 (
      {stage0_40[430]},
      {stage1_40[248]}
   );
   gpc1_1 gpc3978 (
      {stage0_40[431]},
      {stage1_40[249]}
   );
   gpc1_1 gpc3979 (
      {stage0_40[432]},
      {stage1_40[250]}
   );
   gpc1_1 gpc3980 (
      {stage0_40[433]},
      {stage1_40[251]}
   );
   gpc1_1 gpc3981 (
      {stage0_40[434]},
      {stage1_40[252]}
   );
   gpc1_1 gpc3982 (
      {stage0_40[435]},
      {stage1_40[253]}
   );
   gpc1_1 gpc3983 (
      {stage0_40[436]},
      {stage1_40[254]}
   );
   gpc1_1 gpc3984 (
      {stage0_40[437]},
      {stage1_40[255]}
   );
   gpc1_1 gpc3985 (
      {stage0_40[438]},
      {stage1_40[256]}
   );
   gpc1_1 gpc3986 (
      {stage0_40[439]},
      {stage1_40[257]}
   );
   gpc1_1 gpc3987 (
      {stage0_40[440]},
      {stage1_40[258]}
   );
   gpc1_1 gpc3988 (
      {stage0_40[441]},
      {stage1_40[259]}
   );
   gpc1_1 gpc3989 (
      {stage0_40[442]},
      {stage1_40[260]}
   );
   gpc1_1 gpc3990 (
      {stage0_40[443]},
      {stage1_40[261]}
   );
   gpc1_1 gpc3991 (
      {stage0_40[444]},
      {stage1_40[262]}
   );
   gpc1_1 gpc3992 (
      {stage0_40[445]},
      {stage1_40[263]}
   );
   gpc1_1 gpc3993 (
      {stage0_40[446]},
      {stage1_40[264]}
   );
   gpc1_1 gpc3994 (
      {stage0_40[447]},
      {stage1_40[265]}
   );
   gpc1_1 gpc3995 (
      {stage0_40[448]},
      {stage1_40[266]}
   );
   gpc1_1 gpc3996 (
      {stage0_40[449]},
      {stage1_40[267]}
   );
   gpc1_1 gpc3997 (
      {stage0_40[450]},
      {stage1_40[268]}
   );
   gpc1_1 gpc3998 (
      {stage0_40[451]},
      {stage1_40[269]}
   );
   gpc1_1 gpc3999 (
      {stage0_40[452]},
      {stage1_40[270]}
   );
   gpc1_1 gpc4000 (
      {stage0_40[453]},
      {stage1_40[271]}
   );
   gpc1_1 gpc4001 (
      {stage0_40[454]},
      {stage1_40[272]}
   );
   gpc1_1 gpc4002 (
      {stage0_40[455]},
      {stage1_40[273]}
   );
   gpc1_1 gpc4003 (
      {stage0_40[456]},
      {stage1_40[274]}
   );
   gpc1_1 gpc4004 (
      {stage0_40[457]},
      {stage1_40[275]}
   );
   gpc1_1 gpc4005 (
      {stage0_40[458]},
      {stage1_40[276]}
   );
   gpc1_1 gpc4006 (
      {stage0_40[459]},
      {stage1_40[277]}
   );
   gpc1_1 gpc4007 (
      {stage0_40[460]},
      {stage1_40[278]}
   );
   gpc1_1 gpc4008 (
      {stage0_40[461]},
      {stage1_40[279]}
   );
   gpc1_1 gpc4009 (
      {stage0_40[462]},
      {stage1_40[280]}
   );
   gpc1_1 gpc4010 (
      {stage0_40[463]},
      {stage1_40[281]}
   );
   gpc1_1 gpc4011 (
      {stage0_40[464]},
      {stage1_40[282]}
   );
   gpc1_1 gpc4012 (
      {stage0_40[465]},
      {stage1_40[283]}
   );
   gpc1_1 gpc4013 (
      {stage0_40[466]},
      {stage1_40[284]}
   );
   gpc1_1 gpc4014 (
      {stage0_40[467]},
      {stage1_40[285]}
   );
   gpc1_1 gpc4015 (
      {stage0_40[468]},
      {stage1_40[286]}
   );
   gpc1_1 gpc4016 (
      {stage0_40[469]},
      {stage1_40[287]}
   );
   gpc1_1 gpc4017 (
      {stage0_40[470]},
      {stage1_40[288]}
   );
   gpc1_1 gpc4018 (
      {stage0_40[471]},
      {stage1_40[289]}
   );
   gpc1_1 gpc4019 (
      {stage0_40[472]},
      {stage1_40[290]}
   );
   gpc1_1 gpc4020 (
      {stage0_40[473]},
      {stage1_40[291]}
   );
   gpc1_1 gpc4021 (
      {stage0_40[474]},
      {stage1_40[292]}
   );
   gpc1_1 gpc4022 (
      {stage0_40[475]},
      {stage1_40[293]}
   );
   gpc1_1 gpc4023 (
      {stage0_40[476]},
      {stage1_40[294]}
   );
   gpc1_1 gpc4024 (
      {stage0_40[477]},
      {stage1_40[295]}
   );
   gpc1_1 gpc4025 (
      {stage0_40[478]},
      {stage1_40[296]}
   );
   gpc1_1 gpc4026 (
      {stage0_40[479]},
      {stage1_40[297]}
   );
   gpc1_1 gpc4027 (
      {stage0_40[480]},
      {stage1_40[298]}
   );
   gpc1_1 gpc4028 (
      {stage0_40[481]},
      {stage1_40[299]}
   );
   gpc1_1 gpc4029 (
      {stage0_40[482]},
      {stage1_40[300]}
   );
   gpc1_1 gpc4030 (
      {stage0_40[483]},
      {stage1_40[301]}
   );
   gpc1_1 gpc4031 (
      {stage0_40[484]},
      {stage1_40[302]}
   );
   gpc1_1 gpc4032 (
      {stage0_40[485]},
      {stage1_40[303]}
   );
   gpc1_1 gpc4033 (
      {stage0_41[477]},
      {stage1_41[162]}
   );
   gpc1_1 gpc4034 (
      {stage0_41[478]},
      {stage1_41[163]}
   );
   gpc1_1 gpc4035 (
      {stage0_41[479]},
      {stage1_41[164]}
   );
   gpc1_1 gpc4036 (
      {stage0_41[480]},
      {stage1_41[165]}
   );
   gpc1_1 gpc4037 (
      {stage0_41[481]},
      {stage1_41[166]}
   );
   gpc1_1 gpc4038 (
      {stage0_41[482]},
      {stage1_41[167]}
   );
   gpc1_1 gpc4039 (
      {stage0_41[483]},
      {stage1_41[168]}
   );
   gpc1_1 gpc4040 (
      {stage0_41[484]},
      {stage1_41[169]}
   );
   gpc1_1 gpc4041 (
      {stage0_41[485]},
      {stage1_41[170]}
   );
   gpc1_1 gpc4042 (
      {stage0_42[483]},
      {stage1_42[171]}
   );
   gpc1_1 gpc4043 (
      {stage0_42[484]},
      {stage1_42[172]}
   );
   gpc1_1 gpc4044 (
      {stage0_42[485]},
      {stage1_42[173]}
   );
   gpc1_1 gpc4045 (
      {stage0_43[451]},
      {stage1_43[219]}
   );
   gpc1_1 gpc4046 (
      {stage0_43[452]},
      {stage1_43[220]}
   );
   gpc1_1 gpc4047 (
      {stage0_43[453]},
      {stage1_43[221]}
   );
   gpc1_1 gpc4048 (
      {stage0_43[454]},
      {stage1_43[222]}
   );
   gpc1_1 gpc4049 (
      {stage0_43[455]},
      {stage1_43[223]}
   );
   gpc1_1 gpc4050 (
      {stage0_43[456]},
      {stage1_43[224]}
   );
   gpc1_1 gpc4051 (
      {stage0_43[457]},
      {stage1_43[225]}
   );
   gpc1_1 gpc4052 (
      {stage0_43[458]},
      {stage1_43[226]}
   );
   gpc1_1 gpc4053 (
      {stage0_43[459]},
      {stage1_43[227]}
   );
   gpc1_1 gpc4054 (
      {stage0_43[460]},
      {stage1_43[228]}
   );
   gpc1_1 gpc4055 (
      {stage0_43[461]},
      {stage1_43[229]}
   );
   gpc1_1 gpc4056 (
      {stage0_43[462]},
      {stage1_43[230]}
   );
   gpc1_1 gpc4057 (
      {stage0_43[463]},
      {stage1_43[231]}
   );
   gpc1_1 gpc4058 (
      {stage0_43[464]},
      {stage1_43[232]}
   );
   gpc1_1 gpc4059 (
      {stage0_43[465]},
      {stage1_43[233]}
   );
   gpc1_1 gpc4060 (
      {stage0_43[466]},
      {stage1_43[234]}
   );
   gpc1_1 gpc4061 (
      {stage0_43[467]},
      {stage1_43[235]}
   );
   gpc1_1 gpc4062 (
      {stage0_43[468]},
      {stage1_43[236]}
   );
   gpc1_1 gpc4063 (
      {stage0_43[469]},
      {stage1_43[237]}
   );
   gpc1_1 gpc4064 (
      {stage0_43[470]},
      {stage1_43[238]}
   );
   gpc1_1 gpc4065 (
      {stage0_43[471]},
      {stage1_43[239]}
   );
   gpc1_1 gpc4066 (
      {stage0_43[472]},
      {stage1_43[240]}
   );
   gpc1_1 gpc4067 (
      {stage0_43[473]},
      {stage1_43[241]}
   );
   gpc1_1 gpc4068 (
      {stage0_43[474]},
      {stage1_43[242]}
   );
   gpc1_1 gpc4069 (
      {stage0_43[475]},
      {stage1_43[243]}
   );
   gpc1_1 gpc4070 (
      {stage0_43[476]},
      {stage1_43[244]}
   );
   gpc1_1 gpc4071 (
      {stage0_43[477]},
      {stage1_43[245]}
   );
   gpc1_1 gpc4072 (
      {stage0_43[478]},
      {stage1_43[246]}
   );
   gpc1_1 gpc4073 (
      {stage0_43[479]},
      {stage1_43[247]}
   );
   gpc1_1 gpc4074 (
      {stage0_43[480]},
      {stage1_43[248]}
   );
   gpc1_1 gpc4075 (
      {stage0_43[481]},
      {stage1_43[249]}
   );
   gpc1_1 gpc4076 (
      {stage0_43[482]},
      {stage1_43[250]}
   );
   gpc1_1 gpc4077 (
      {stage0_43[483]},
      {stage1_43[251]}
   );
   gpc1_1 gpc4078 (
      {stage0_43[484]},
      {stage1_43[252]}
   );
   gpc1_1 gpc4079 (
      {stage0_43[485]},
      {stage1_43[253]}
   );
   gpc1_1 gpc4080 (
      {stage0_44[424]},
      {stage1_44[194]}
   );
   gpc1_1 gpc4081 (
      {stage0_44[425]},
      {stage1_44[195]}
   );
   gpc1_1 gpc4082 (
      {stage0_44[426]},
      {stage1_44[196]}
   );
   gpc1_1 gpc4083 (
      {stage0_44[427]},
      {stage1_44[197]}
   );
   gpc1_1 gpc4084 (
      {stage0_44[428]},
      {stage1_44[198]}
   );
   gpc1_1 gpc4085 (
      {stage0_44[429]},
      {stage1_44[199]}
   );
   gpc1_1 gpc4086 (
      {stage0_44[430]},
      {stage1_44[200]}
   );
   gpc1_1 gpc4087 (
      {stage0_44[431]},
      {stage1_44[201]}
   );
   gpc1_1 gpc4088 (
      {stage0_44[432]},
      {stage1_44[202]}
   );
   gpc1_1 gpc4089 (
      {stage0_44[433]},
      {stage1_44[203]}
   );
   gpc1_1 gpc4090 (
      {stage0_44[434]},
      {stage1_44[204]}
   );
   gpc1_1 gpc4091 (
      {stage0_44[435]},
      {stage1_44[205]}
   );
   gpc1_1 gpc4092 (
      {stage0_44[436]},
      {stage1_44[206]}
   );
   gpc1_1 gpc4093 (
      {stage0_44[437]},
      {stage1_44[207]}
   );
   gpc1_1 gpc4094 (
      {stage0_44[438]},
      {stage1_44[208]}
   );
   gpc1_1 gpc4095 (
      {stage0_44[439]},
      {stage1_44[209]}
   );
   gpc1_1 gpc4096 (
      {stage0_44[440]},
      {stage1_44[210]}
   );
   gpc1_1 gpc4097 (
      {stage0_44[441]},
      {stage1_44[211]}
   );
   gpc1_1 gpc4098 (
      {stage0_44[442]},
      {stage1_44[212]}
   );
   gpc1_1 gpc4099 (
      {stage0_44[443]},
      {stage1_44[213]}
   );
   gpc1_1 gpc4100 (
      {stage0_44[444]},
      {stage1_44[214]}
   );
   gpc1_1 gpc4101 (
      {stage0_44[445]},
      {stage1_44[215]}
   );
   gpc1_1 gpc4102 (
      {stage0_44[446]},
      {stage1_44[216]}
   );
   gpc1_1 gpc4103 (
      {stage0_44[447]},
      {stage1_44[217]}
   );
   gpc1_1 gpc4104 (
      {stage0_44[448]},
      {stage1_44[218]}
   );
   gpc1_1 gpc4105 (
      {stage0_44[449]},
      {stage1_44[219]}
   );
   gpc1_1 gpc4106 (
      {stage0_44[450]},
      {stage1_44[220]}
   );
   gpc1_1 gpc4107 (
      {stage0_44[451]},
      {stage1_44[221]}
   );
   gpc1_1 gpc4108 (
      {stage0_44[452]},
      {stage1_44[222]}
   );
   gpc1_1 gpc4109 (
      {stage0_44[453]},
      {stage1_44[223]}
   );
   gpc1_1 gpc4110 (
      {stage0_44[454]},
      {stage1_44[224]}
   );
   gpc1_1 gpc4111 (
      {stage0_44[455]},
      {stage1_44[225]}
   );
   gpc1_1 gpc4112 (
      {stage0_44[456]},
      {stage1_44[226]}
   );
   gpc1_1 gpc4113 (
      {stage0_44[457]},
      {stage1_44[227]}
   );
   gpc1_1 gpc4114 (
      {stage0_44[458]},
      {stage1_44[228]}
   );
   gpc1_1 gpc4115 (
      {stage0_44[459]},
      {stage1_44[229]}
   );
   gpc1_1 gpc4116 (
      {stage0_44[460]},
      {stage1_44[230]}
   );
   gpc1_1 gpc4117 (
      {stage0_44[461]},
      {stage1_44[231]}
   );
   gpc1_1 gpc4118 (
      {stage0_44[462]},
      {stage1_44[232]}
   );
   gpc1_1 gpc4119 (
      {stage0_44[463]},
      {stage1_44[233]}
   );
   gpc1_1 gpc4120 (
      {stage0_44[464]},
      {stage1_44[234]}
   );
   gpc1_1 gpc4121 (
      {stage0_44[465]},
      {stage1_44[235]}
   );
   gpc1_1 gpc4122 (
      {stage0_44[466]},
      {stage1_44[236]}
   );
   gpc1_1 gpc4123 (
      {stage0_44[467]},
      {stage1_44[237]}
   );
   gpc1_1 gpc4124 (
      {stage0_44[468]},
      {stage1_44[238]}
   );
   gpc1_1 gpc4125 (
      {stage0_44[469]},
      {stage1_44[239]}
   );
   gpc1_1 gpc4126 (
      {stage0_44[470]},
      {stage1_44[240]}
   );
   gpc1_1 gpc4127 (
      {stage0_44[471]},
      {stage1_44[241]}
   );
   gpc1_1 gpc4128 (
      {stage0_44[472]},
      {stage1_44[242]}
   );
   gpc1_1 gpc4129 (
      {stage0_44[473]},
      {stage1_44[243]}
   );
   gpc1_1 gpc4130 (
      {stage0_44[474]},
      {stage1_44[244]}
   );
   gpc1_1 gpc4131 (
      {stage0_44[475]},
      {stage1_44[245]}
   );
   gpc1_1 gpc4132 (
      {stage0_44[476]},
      {stage1_44[246]}
   );
   gpc1_1 gpc4133 (
      {stage0_44[477]},
      {stage1_44[247]}
   );
   gpc1_1 gpc4134 (
      {stage0_44[478]},
      {stage1_44[248]}
   );
   gpc1_1 gpc4135 (
      {stage0_44[479]},
      {stage1_44[249]}
   );
   gpc1_1 gpc4136 (
      {stage0_44[480]},
      {stage1_44[250]}
   );
   gpc1_1 gpc4137 (
      {stage0_44[481]},
      {stage1_44[251]}
   );
   gpc1_1 gpc4138 (
      {stage0_44[482]},
      {stage1_44[252]}
   );
   gpc1_1 gpc4139 (
      {stage0_44[483]},
      {stage1_44[253]}
   );
   gpc1_1 gpc4140 (
      {stage0_44[484]},
      {stage1_44[254]}
   );
   gpc1_1 gpc4141 (
      {stage0_44[485]},
      {stage1_44[255]}
   );
   gpc1_1 gpc4142 (
      {stage0_45[433]},
      {stage1_45[159]}
   );
   gpc1_1 gpc4143 (
      {stage0_45[434]},
      {stage1_45[160]}
   );
   gpc1_1 gpc4144 (
      {stage0_45[435]},
      {stage1_45[161]}
   );
   gpc1_1 gpc4145 (
      {stage0_45[436]},
      {stage1_45[162]}
   );
   gpc1_1 gpc4146 (
      {stage0_45[437]},
      {stage1_45[163]}
   );
   gpc1_1 gpc4147 (
      {stage0_45[438]},
      {stage1_45[164]}
   );
   gpc1_1 gpc4148 (
      {stage0_45[439]},
      {stage1_45[165]}
   );
   gpc1_1 gpc4149 (
      {stage0_45[440]},
      {stage1_45[166]}
   );
   gpc1_1 gpc4150 (
      {stage0_45[441]},
      {stage1_45[167]}
   );
   gpc1_1 gpc4151 (
      {stage0_45[442]},
      {stage1_45[168]}
   );
   gpc1_1 gpc4152 (
      {stage0_45[443]},
      {stage1_45[169]}
   );
   gpc1_1 gpc4153 (
      {stage0_45[444]},
      {stage1_45[170]}
   );
   gpc1_1 gpc4154 (
      {stage0_45[445]},
      {stage1_45[171]}
   );
   gpc1_1 gpc4155 (
      {stage0_45[446]},
      {stage1_45[172]}
   );
   gpc1_1 gpc4156 (
      {stage0_45[447]},
      {stage1_45[173]}
   );
   gpc1_1 gpc4157 (
      {stage0_45[448]},
      {stage1_45[174]}
   );
   gpc1_1 gpc4158 (
      {stage0_45[449]},
      {stage1_45[175]}
   );
   gpc1_1 gpc4159 (
      {stage0_45[450]},
      {stage1_45[176]}
   );
   gpc1_1 gpc4160 (
      {stage0_45[451]},
      {stage1_45[177]}
   );
   gpc1_1 gpc4161 (
      {stage0_45[452]},
      {stage1_45[178]}
   );
   gpc1_1 gpc4162 (
      {stage0_45[453]},
      {stage1_45[179]}
   );
   gpc1_1 gpc4163 (
      {stage0_45[454]},
      {stage1_45[180]}
   );
   gpc1_1 gpc4164 (
      {stage0_45[455]},
      {stage1_45[181]}
   );
   gpc1_1 gpc4165 (
      {stage0_45[456]},
      {stage1_45[182]}
   );
   gpc1_1 gpc4166 (
      {stage0_45[457]},
      {stage1_45[183]}
   );
   gpc1_1 gpc4167 (
      {stage0_45[458]},
      {stage1_45[184]}
   );
   gpc1_1 gpc4168 (
      {stage0_45[459]},
      {stage1_45[185]}
   );
   gpc1_1 gpc4169 (
      {stage0_45[460]},
      {stage1_45[186]}
   );
   gpc1_1 gpc4170 (
      {stage0_45[461]},
      {stage1_45[187]}
   );
   gpc1_1 gpc4171 (
      {stage0_45[462]},
      {stage1_45[188]}
   );
   gpc1_1 gpc4172 (
      {stage0_45[463]},
      {stage1_45[189]}
   );
   gpc1_1 gpc4173 (
      {stage0_45[464]},
      {stage1_45[190]}
   );
   gpc1_1 gpc4174 (
      {stage0_45[465]},
      {stage1_45[191]}
   );
   gpc1_1 gpc4175 (
      {stage0_45[466]},
      {stage1_45[192]}
   );
   gpc1_1 gpc4176 (
      {stage0_45[467]},
      {stage1_45[193]}
   );
   gpc1_1 gpc4177 (
      {stage0_45[468]},
      {stage1_45[194]}
   );
   gpc1_1 gpc4178 (
      {stage0_45[469]},
      {stage1_45[195]}
   );
   gpc1_1 gpc4179 (
      {stage0_45[470]},
      {stage1_45[196]}
   );
   gpc1_1 gpc4180 (
      {stage0_45[471]},
      {stage1_45[197]}
   );
   gpc1_1 gpc4181 (
      {stage0_45[472]},
      {stage1_45[198]}
   );
   gpc1_1 gpc4182 (
      {stage0_45[473]},
      {stage1_45[199]}
   );
   gpc1_1 gpc4183 (
      {stage0_45[474]},
      {stage1_45[200]}
   );
   gpc1_1 gpc4184 (
      {stage0_45[475]},
      {stage1_45[201]}
   );
   gpc1_1 gpc4185 (
      {stage0_45[476]},
      {stage1_45[202]}
   );
   gpc1_1 gpc4186 (
      {stage0_45[477]},
      {stage1_45[203]}
   );
   gpc1_1 gpc4187 (
      {stage0_45[478]},
      {stage1_45[204]}
   );
   gpc1_1 gpc4188 (
      {stage0_45[479]},
      {stage1_45[205]}
   );
   gpc1_1 gpc4189 (
      {stage0_45[480]},
      {stage1_45[206]}
   );
   gpc1_1 gpc4190 (
      {stage0_45[481]},
      {stage1_45[207]}
   );
   gpc1_1 gpc4191 (
      {stage0_45[482]},
      {stage1_45[208]}
   );
   gpc1_1 gpc4192 (
      {stage0_45[483]},
      {stage1_45[209]}
   );
   gpc1_1 gpc4193 (
      {stage0_45[484]},
      {stage1_45[210]}
   );
   gpc1_1 gpc4194 (
      {stage0_45[485]},
      {stage1_45[211]}
   );
   gpc1_1 gpc4195 (
      {stage0_46[356]},
      {stage1_46[168]}
   );
   gpc1_1 gpc4196 (
      {stage0_46[357]},
      {stage1_46[169]}
   );
   gpc1_1 gpc4197 (
      {stage0_46[358]},
      {stage1_46[170]}
   );
   gpc1_1 gpc4198 (
      {stage0_46[359]},
      {stage1_46[171]}
   );
   gpc1_1 gpc4199 (
      {stage0_46[360]},
      {stage1_46[172]}
   );
   gpc1_1 gpc4200 (
      {stage0_46[361]},
      {stage1_46[173]}
   );
   gpc1_1 gpc4201 (
      {stage0_46[362]},
      {stage1_46[174]}
   );
   gpc1_1 gpc4202 (
      {stage0_46[363]},
      {stage1_46[175]}
   );
   gpc1_1 gpc4203 (
      {stage0_46[364]},
      {stage1_46[176]}
   );
   gpc1_1 gpc4204 (
      {stage0_46[365]},
      {stage1_46[177]}
   );
   gpc1_1 gpc4205 (
      {stage0_46[366]},
      {stage1_46[178]}
   );
   gpc1_1 gpc4206 (
      {stage0_46[367]},
      {stage1_46[179]}
   );
   gpc1_1 gpc4207 (
      {stage0_46[368]},
      {stage1_46[180]}
   );
   gpc1_1 gpc4208 (
      {stage0_46[369]},
      {stage1_46[181]}
   );
   gpc1_1 gpc4209 (
      {stage0_46[370]},
      {stage1_46[182]}
   );
   gpc1_1 gpc4210 (
      {stage0_46[371]},
      {stage1_46[183]}
   );
   gpc1_1 gpc4211 (
      {stage0_46[372]},
      {stage1_46[184]}
   );
   gpc1_1 gpc4212 (
      {stage0_46[373]},
      {stage1_46[185]}
   );
   gpc1_1 gpc4213 (
      {stage0_46[374]},
      {stage1_46[186]}
   );
   gpc1_1 gpc4214 (
      {stage0_46[375]},
      {stage1_46[187]}
   );
   gpc1_1 gpc4215 (
      {stage0_46[376]},
      {stage1_46[188]}
   );
   gpc1_1 gpc4216 (
      {stage0_46[377]},
      {stage1_46[189]}
   );
   gpc1_1 gpc4217 (
      {stage0_46[378]},
      {stage1_46[190]}
   );
   gpc1_1 gpc4218 (
      {stage0_46[379]},
      {stage1_46[191]}
   );
   gpc1_1 gpc4219 (
      {stage0_46[380]},
      {stage1_46[192]}
   );
   gpc1_1 gpc4220 (
      {stage0_46[381]},
      {stage1_46[193]}
   );
   gpc1_1 gpc4221 (
      {stage0_46[382]},
      {stage1_46[194]}
   );
   gpc1_1 gpc4222 (
      {stage0_46[383]},
      {stage1_46[195]}
   );
   gpc1_1 gpc4223 (
      {stage0_46[384]},
      {stage1_46[196]}
   );
   gpc1_1 gpc4224 (
      {stage0_46[385]},
      {stage1_46[197]}
   );
   gpc1_1 gpc4225 (
      {stage0_46[386]},
      {stage1_46[198]}
   );
   gpc1_1 gpc4226 (
      {stage0_46[387]},
      {stage1_46[199]}
   );
   gpc1_1 gpc4227 (
      {stage0_46[388]},
      {stage1_46[200]}
   );
   gpc1_1 gpc4228 (
      {stage0_46[389]},
      {stage1_46[201]}
   );
   gpc1_1 gpc4229 (
      {stage0_46[390]},
      {stage1_46[202]}
   );
   gpc1_1 gpc4230 (
      {stage0_46[391]},
      {stage1_46[203]}
   );
   gpc1_1 gpc4231 (
      {stage0_46[392]},
      {stage1_46[204]}
   );
   gpc1_1 gpc4232 (
      {stage0_46[393]},
      {stage1_46[205]}
   );
   gpc1_1 gpc4233 (
      {stage0_46[394]},
      {stage1_46[206]}
   );
   gpc1_1 gpc4234 (
      {stage0_46[395]},
      {stage1_46[207]}
   );
   gpc1_1 gpc4235 (
      {stage0_46[396]},
      {stage1_46[208]}
   );
   gpc1_1 gpc4236 (
      {stage0_46[397]},
      {stage1_46[209]}
   );
   gpc1_1 gpc4237 (
      {stage0_46[398]},
      {stage1_46[210]}
   );
   gpc1_1 gpc4238 (
      {stage0_46[399]},
      {stage1_46[211]}
   );
   gpc1_1 gpc4239 (
      {stage0_46[400]},
      {stage1_46[212]}
   );
   gpc1_1 gpc4240 (
      {stage0_46[401]},
      {stage1_46[213]}
   );
   gpc1_1 gpc4241 (
      {stage0_46[402]},
      {stage1_46[214]}
   );
   gpc1_1 gpc4242 (
      {stage0_46[403]},
      {stage1_46[215]}
   );
   gpc1_1 gpc4243 (
      {stage0_46[404]},
      {stage1_46[216]}
   );
   gpc1_1 gpc4244 (
      {stage0_46[405]},
      {stage1_46[217]}
   );
   gpc1_1 gpc4245 (
      {stage0_46[406]},
      {stage1_46[218]}
   );
   gpc1_1 gpc4246 (
      {stage0_46[407]},
      {stage1_46[219]}
   );
   gpc1_1 gpc4247 (
      {stage0_46[408]},
      {stage1_46[220]}
   );
   gpc1_1 gpc4248 (
      {stage0_46[409]},
      {stage1_46[221]}
   );
   gpc1_1 gpc4249 (
      {stage0_46[410]},
      {stage1_46[222]}
   );
   gpc1_1 gpc4250 (
      {stage0_46[411]},
      {stage1_46[223]}
   );
   gpc1_1 gpc4251 (
      {stage0_46[412]},
      {stage1_46[224]}
   );
   gpc1_1 gpc4252 (
      {stage0_46[413]},
      {stage1_46[225]}
   );
   gpc1_1 gpc4253 (
      {stage0_46[414]},
      {stage1_46[226]}
   );
   gpc1_1 gpc4254 (
      {stage0_46[415]},
      {stage1_46[227]}
   );
   gpc1_1 gpc4255 (
      {stage0_46[416]},
      {stage1_46[228]}
   );
   gpc1_1 gpc4256 (
      {stage0_46[417]},
      {stage1_46[229]}
   );
   gpc1_1 gpc4257 (
      {stage0_46[418]},
      {stage1_46[230]}
   );
   gpc1_1 gpc4258 (
      {stage0_46[419]},
      {stage1_46[231]}
   );
   gpc1_1 gpc4259 (
      {stage0_46[420]},
      {stage1_46[232]}
   );
   gpc1_1 gpc4260 (
      {stage0_46[421]},
      {stage1_46[233]}
   );
   gpc1_1 gpc4261 (
      {stage0_46[422]},
      {stage1_46[234]}
   );
   gpc1_1 gpc4262 (
      {stage0_46[423]},
      {stage1_46[235]}
   );
   gpc1_1 gpc4263 (
      {stage0_46[424]},
      {stage1_46[236]}
   );
   gpc1_1 gpc4264 (
      {stage0_46[425]},
      {stage1_46[237]}
   );
   gpc1_1 gpc4265 (
      {stage0_46[426]},
      {stage1_46[238]}
   );
   gpc1_1 gpc4266 (
      {stage0_46[427]},
      {stage1_46[239]}
   );
   gpc1_1 gpc4267 (
      {stage0_46[428]},
      {stage1_46[240]}
   );
   gpc1_1 gpc4268 (
      {stage0_46[429]},
      {stage1_46[241]}
   );
   gpc1_1 gpc4269 (
      {stage0_46[430]},
      {stage1_46[242]}
   );
   gpc1_1 gpc4270 (
      {stage0_46[431]},
      {stage1_46[243]}
   );
   gpc1_1 gpc4271 (
      {stage0_46[432]},
      {stage1_46[244]}
   );
   gpc1_1 gpc4272 (
      {stage0_46[433]},
      {stage1_46[245]}
   );
   gpc1_1 gpc4273 (
      {stage0_46[434]},
      {stage1_46[246]}
   );
   gpc1_1 gpc4274 (
      {stage0_46[435]},
      {stage1_46[247]}
   );
   gpc1_1 gpc4275 (
      {stage0_46[436]},
      {stage1_46[248]}
   );
   gpc1_1 gpc4276 (
      {stage0_46[437]},
      {stage1_46[249]}
   );
   gpc1_1 gpc4277 (
      {stage0_46[438]},
      {stage1_46[250]}
   );
   gpc1_1 gpc4278 (
      {stage0_46[439]},
      {stage1_46[251]}
   );
   gpc1_1 gpc4279 (
      {stage0_46[440]},
      {stage1_46[252]}
   );
   gpc1_1 gpc4280 (
      {stage0_46[441]},
      {stage1_46[253]}
   );
   gpc1_1 gpc4281 (
      {stage0_46[442]},
      {stage1_46[254]}
   );
   gpc1_1 gpc4282 (
      {stage0_46[443]},
      {stage1_46[255]}
   );
   gpc1_1 gpc4283 (
      {stage0_46[444]},
      {stage1_46[256]}
   );
   gpc1_1 gpc4284 (
      {stage0_46[445]},
      {stage1_46[257]}
   );
   gpc1_1 gpc4285 (
      {stage0_46[446]},
      {stage1_46[258]}
   );
   gpc1_1 gpc4286 (
      {stage0_46[447]},
      {stage1_46[259]}
   );
   gpc1_1 gpc4287 (
      {stage0_46[448]},
      {stage1_46[260]}
   );
   gpc1_1 gpc4288 (
      {stage0_46[449]},
      {stage1_46[261]}
   );
   gpc1_1 gpc4289 (
      {stage0_46[450]},
      {stage1_46[262]}
   );
   gpc1_1 gpc4290 (
      {stage0_46[451]},
      {stage1_46[263]}
   );
   gpc1_1 gpc4291 (
      {stage0_46[452]},
      {stage1_46[264]}
   );
   gpc1_1 gpc4292 (
      {stage0_46[453]},
      {stage1_46[265]}
   );
   gpc1_1 gpc4293 (
      {stage0_46[454]},
      {stage1_46[266]}
   );
   gpc1_1 gpc4294 (
      {stage0_46[455]},
      {stage1_46[267]}
   );
   gpc1_1 gpc4295 (
      {stage0_46[456]},
      {stage1_46[268]}
   );
   gpc1_1 gpc4296 (
      {stage0_46[457]},
      {stage1_46[269]}
   );
   gpc1_1 gpc4297 (
      {stage0_46[458]},
      {stage1_46[270]}
   );
   gpc1_1 gpc4298 (
      {stage0_46[459]},
      {stage1_46[271]}
   );
   gpc1_1 gpc4299 (
      {stage0_46[460]},
      {stage1_46[272]}
   );
   gpc1_1 gpc4300 (
      {stage0_46[461]},
      {stage1_46[273]}
   );
   gpc1_1 gpc4301 (
      {stage0_46[462]},
      {stage1_46[274]}
   );
   gpc1_1 gpc4302 (
      {stage0_46[463]},
      {stage1_46[275]}
   );
   gpc1_1 gpc4303 (
      {stage0_46[464]},
      {stage1_46[276]}
   );
   gpc1_1 gpc4304 (
      {stage0_46[465]},
      {stage1_46[277]}
   );
   gpc1_1 gpc4305 (
      {stage0_46[466]},
      {stage1_46[278]}
   );
   gpc1_1 gpc4306 (
      {stage0_46[467]},
      {stage1_46[279]}
   );
   gpc1_1 gpc4307 (
      {stage0_46[468]},
      {stage1_46[280]}
   );
   gpc1_1 gpc4308 (
      {stage0_46[469]},
      {stage1_46[281]}
   );
   gpc1_1 gpc4309 (
      {stage0_46[470]},
      {stage1_46[282]}
   );
   gpc1_1 gpc4310 (
      {stage0_46[471]},
      {stage1_46[283]}
   );
   gpc1_1 gpc4311 (
      {stage0_46[472]},
      {stage1_46[284]}
   );
   gpc1_1 gpc4312 (
      {stage0_46[473]},
      {stage1_46[285]}
   );
   gpc1_1 gpc4313 (
      {stage0_46[474]},
      {stage1_46[286]}
   );
   gpc1_1 gpc4314 (
      {stage0_46[475]},
      {stage1_46[287]}
   );
   gpc1_1 gpc4315 (
      {stage0_46[476]},
      {stage1_46[288]}
   );
   gpc1_1 gpc4316 (
      {stage0_46[477]},
      {stage1_46[289]}
   );
   gpc1_1 gpc4317 (
      {stage0_46[478]},
      {stage1_46[290]}
   );
   gpc1_1 gpc4318 (
      {stage0_46[479]},
      {stage1_46[291]}
   );
   gpc1_1 gpc4319 (
      {stage0_46[480]},
      {stage1_46[292]}
   );
   gpc1_1 gpc4320 (
      {stage0_46[481]},
      {stage1_46[293]}
   );
   gpc1_1 gpc4321 (
      {stage0_46[482]},
      {stage1_46[294]}
   );
   gpc1_1 gpc4322 (
      {stage0_46[483]},
      {stage1_46[295]}
   );
   gpc1_1 gpc4323 (
      {stage0_46[484]},
      {stage1_46[296]}
   );
   gpc1_1 gpc4324 (
      {stage0_46[485]},
      {stage1_46[297]}
   );
   gpc1_1 gpc4325 (
      {stage0_47[443]},
      {stage1_47[193]}
   );
   gpc1_1 gpc4326 (
      {stage0_47[444]},
      {stage1_47[194]}
   );
   gpc1_1 gpc4327 (
      {stage0_47[445]},
      {stage1_47[195]}
   );
   gpc1_1 gpc4328 (
      {stage0_47[446]},
      {stage1_47[196]}
   );
   gpc1_1 gpc4329 (
      {stage0_47[447]},
      {stage1_47[197]}
   );
   gpc1_1 gpc4330 (
      {stage0_47[448]},
      {stage1_47[198]}
   );
   gpc1_1 gpc4331 (
      {stage0_47[449]},
      {stage1_47[199]}
   );
   gpc1_1 gpc4332 (
      {stage0_47[450]},
      {stage1_47[200]}
   );
   gpc1_1 gpc4333 (
      {stage0_47[451]},
      {stage1_47[201]}
   );
   gpc1_1 gpc4334 (
      {stage0_47[452]},
      {stage1_47[202]}
   );
   gpc1_1 gpc4335 (
      {stage0_47[453]},
      {stage1_47[203]}
   );
   gpc1_1 gpc4336 (
      {stage0_47[454]},
      {stage1_47[204]}
   );
   gpc1_1 gpc4337 (
      {stage0_47[455]},
      {stage1_47[205]}
   );
   gpc1_1 gpc4338 (
      {stage0_47[456]},
      {stage1_47[206]}
   );
   gpc1_1 gpc4339 (
      {stage0_47[457]},
      {stage1_47[207]}
   );
   gpc1_1 gpc4340 (
      {stage0_47[458]},
      {stage1_47[208]}
   );
   gpc1_1 gpc4341 (
      {stage0_47[459]},
      {stage1_47[209]}
   );
   gpc1_1 gpc4342 (
      {stage0_47[460]},
      {stage1_47[210]}
   );
   gpc1_1 gpc4343 (
      {stage0_47[461]},
      {stage1_47[211]}
   );
   gpc1_1 gpc4344 (
      {stage0_47[462]},
      {stage1_47[212]}
   );
   gpc1_1 gpc4345 (
      {stage0_47[463]},
      {stage1_47[213]}
   );
   gpc1_1 gpc4346 (
      {stage0_47[464]},
      {stage1_47[214]}
   );
   gpc1_1 gpc4347 (
      {stage0_47[465]},
      {stage1_47[215]}
   );
   gpc1_1 gpc4348 (
      {stage0_47[466]},
      {stage1_47[216]}
   );
   gpc1_1 gpc4349 (
      {stage0_47[467]},
      {stage1_47[217]}
   );
   gpc1_1 gpc4350 (
      {stage0_47[468]},
      {stage1_47[218]}
   );
   gpc1_1 gpc4351 (
      {stage0_47[469]},
      {stage1_47[219]}
   );
   gpc1_1 gpc4352 (
      {stage0_47[470]},
      {stage1_47[220]}
   );
   gpc1_1 gpc4353 (
      {stage0_47[471]},
      {stage1_47[221]}
   );
   gpc1_1 gpc4354 (
      {stage0_47[472]},
      {stage1_47[222]}
   );
   gpc1_1 gpc4355 (
      {stage0_47[473]},
      {stage1_47[223]}
   );
   gpc1_1 gpc4356 (
      {stage0_47[474]},
      {stage1_47[224]}
   );
   gpc1_1 gpc4357 (
      {stage0_47[475]},
      {stage1_47[225]}
   );
   gpc1_1 gpc4358 (
      {stage0_47[476]},
      {stage1_47[226]}
   );
   gpc1_1 gpc4359 (
      {stage0_47[477]},
      {stage1_47[227]}
   );
   gpc1_1 gpc4360 (
      {stage0_47[478]},
      {stage1_47[228]}
   );
   gpc1_1 gpc4361 (
      {stage0_47[479]},
      {stage1_47[229]}
   );
   gpc1_1 gpc4362 (
      {stage0_47[480]},
      {stage1_47[230]}
   );
   gpc1_1 gpc4363 (
      {stage0_47[481]},
      {stage1_47[231]}
   );
   gpc1_1 gpc4364 (
      {stage0_47[482]},
      {stage1_47[232]}
   );
   gpc1_1 gpc4365 (
      {stage0_47[483]},
      {stage1_47[233]}
   );
   gpc1_1 gpc4366 (
      {stage0_47[484]},
      {stage1_47[234]}
   );
   gpc1_1 gpc4367 (
      {stage0_47[485]},
      {stage1_47[235]}
   );
   gpc1_1 gpc4368 (
      {stage0_48[478]},
      {stage1_48[190]}
   );
   gpc1_1 gpc4369 (
      {stage0_48[479]},
      {stage1_48[191]}
   );
   gpc1_1 gpc4370 (
      {stage0_48[480]},
      {stage1_48[192]}
   );
   gpc1_1 gpc4371 (
      {stage0_48[481]},
      {stage1_48[193]}
   );
   gpc1_1 gpc4372 (
      {stage0_48[482]},
      {stage1_48[194]}
   );
   gpc1_1 gpc4373 (
      {stage0_48[483]},
      {stage1_48[195]}
   );
   gpc1_1 gpc4374 (
      {stage0_48[484]},
      {stage1_48[196]}
   );
   gpc1_1 gpc4375 (
      {stage0_48[485]},
      {stage1_48[197]}
   );
   gpc1_1 gpc4376 (
      {stage0_50[481]},
      {stage1_50[185]}
   );
   gpc1_1 gpc4377 (
      {stage0_50[482]},
      {stage1_50[186]}
   );
   gpc1_1 gpc4378 (
      {stage0_50[483]},
      {stage1_50[187]}
   );
   gpc1_1 gpc4379 (
      {stage0_50[484]},
      {stage1_50[188]}
   );
   gpc1_1 gpc4380 (
      {stage0_50[485]},
      {stage1_50[189]}
   );
   gpc1_1 gpc4381 (
      {stage0_51[435]},
      {stage1_51[224]}
   );
   gpc1_1 gpc4382 (
      {stage0_51[436]},
      {stage1_51[225]}
   );
   gpc1_1 gpc4383 (
      {stage0_51[437]},
      {stage1_51[226]}
   );
   gpc1_1 gpc4384 (
      {stage0_51[438]},
      {stage1_51[227]}
   );
   gpc1_1 gpc4385 (
      {stage0_51[439]},
      {stage1_51[228]}
   );
   gpc1_1 gpc4386 (
      {stage0_51[440]},
      {stage1_51[229]}
   );
   gpc1_1 gpc4387 (
      {stage0_51[441]},
      {stage1_51[230]}
   );
   gpc1_1 gpc4388 (
      {stage0_51[442]},
      {stage1_51[231]}
   );
   gpc1_1 gpc4389 (
      {stage0_51[443]},
      {stage1_51[232]}
   );
   gpc1_1 gpc4390 (
      {stage0_51[444]},
      {stage1_51[233]}
   );
   gpc1_1 gpc4391 (
      {stage0_51[445]},
      {stage1_51[234]}
   );
   gpc1_1 gpc4392 (
      {stage0_51[446]},
      {stage1_51[235]}
   );
   gpc1_1 gpc4393 (
      {stage0_51[447]},
      {stage1_51[236]}
   );
   gpc1_1 gpc4394 (
      {stage0_51[448]},
      {stage1_51[237]}
   );
   gpc1_1 gpc4395 (
      {stage0_51[449]},
      {stage1_51[238]}
   );
   gpc1_1 gpc4396 (
      {stage0_51[450]},
      {stage1_51[239]}
   );
   gpc1_1 gpc4397 (
      {stage0_51[451]},
      {stage1_51[240]}
   );
   gpc1_1 gpc4398 (
      {stage0_51[452]},
      {stage1_51[241]}
   );
   gpc1_1 gpc4399 (
      {stage0_51[453]},
      {stage1_51[242]}
   );
   gpc1_1 gpc4400 (
      {stage0_51[454]},
      {stage1_51[243]}
   );
   gpc1_1 gpc4401 (
      {stage0_51[455]},
      {stage1_51[244]}
   );
   gpc1_1 gpc4402 (
      {stage0_51[456]},
      {stage1_51[245]}
   );
   gpc1_1 gpc4403 (
      {stage0_51[457]},
      {stage1_51[246]}
   );
   gpc1_1 gpc4404 (
      {stage0_51[458]},
      {stage1_51[247]}
   );
   gpc1_1 gpc4405 (
      {stage0_51[459]},
      {stage1_51[248]}
   );
   gpc1_1 gpc4406 (
      {stage0_51[460]},
      {stage1_51[249]}
   );
   gpc1_1 gpc4407 (
      {stage0_51[461]},
      {stage1_51[250]}
   );
   gpc1_1 gpc4408 (
      {stage0_51[462]},
      {stage1_51[251]}
   );
   gpc1_1 gpc4409 (
      {stage0_51[463]},
      {stage1_51[252]}
   );
   gpc1_1 gpc4410 (
      {stage0_51[464]},
      {stage1_51[253]}
   );
   gpc1_1 gpc4411 (
      {stage0_51[465]},
      {stage1_51[254]}
   );
   gpc1_1 gpc4412 (
      {stage0_51[466]},
      {stage1_51[255]}
   );
   gpc1_1 gpc4413 (
      {stage0_51[467]},
      {stage1_51[256]}
   );
   gpc1_1 gpc4414 (
      {stage0_51[468]},
      {stage1_51[257]}
   );
   gpc1_1 gpc4415 (
      {stage0_51[469]},
      {stage1_51[258]}
   );
   gpc1_1 gpc4416 (
      {stage0_51[470]},
      {stage1_51[259]}
   );
   gpc1_1 gpc4417 (
      {stage0_51[471]},
      {stage1_51[260]}
   );
   gpc1_1 gpc4418 (
      {stage0_51[472]},
      {stage1_51[261]}
   );
   gpc1_1 gpc4419 (
      {stage0_51[473]},
      {stage1_51[262]}
   );
   gpc1_1 gpc4420 (
      {stage0_51[474]},
      {stage1_51[263]}
   );
   gpc1_1 gpc4421 (
      {stage0_51[475]},
      {stage1_51[264]}
   );
   gpc1_1 gpc4422 (
      {stage0_51[476]},
      {stage1_51[265]}
   );
   gpc1_1 gpc4423 (
      {stage0_51[477]},
      {stage1_51[266]}
   );
   gpc1_1 gpc4424 (
      {stage0_51[478]},
      {stage1_51[267]}
   );
   gpc1_1 gpc4425 (
      {stage0_51[479]},
      {stage1_51[268]}
   );
   gpc1_1 gpc4426 (
      {stage0_51[480]},
      {stage1_51[269]}
   );
   gpc1_1 gpc4427 (
      {stage0_51[481]},
      {stage1_51[270]}
   );
   gpc1_1 gpc4428 (
      {stage0_51[482]},
      {stage1_51[271]}
   );
   gpc1_1 gpc4429 (
      {stage0_51[483]},
      {stage1_51[272]}
   );
   gpc1_1 gpc4430 (
      {stage0_51[484]},
      {stage1_51[273]}
   );
   gpc1_1 gpc4431 (
      {stage0_51[485]},
      {stage1_51[274]}
   );
   gpc1_1 gpc4432 (
      {stage0_54[453]},
      {stage1_54[198]}
   );
   gpc1_1 gpc4433 (
      {stage0_54[454]},
      {stage1_54[199]}
   );
   gpc1_1 gpc4434 (
      {stage0_54[455]},
      {stage1_54[200]}
   );
   gpc1_1 gpc4435 (
      {stage0_54[456]},
      {stage1_54[201]}
   );
   gpc1_1 gpc4436 (
      {stage0_54[457]},
      {stage1_54[202]}
   );
   gpc1_1 gpc4437 (
      {stage0_54[458]},
      {stage1_54[203]}
   );
   gpc1_1 gpc4438 (
      {stage0_54[459]},
      {stage1_54[204]}
   );
   gpc1_1 gpc4439 (
      {stage0_54[460]},
      {stage1_54[205]}
   );
   gpc1_1 gpc4440 (
      {stage0_54[461]},
      {stage1_54[206]}
   );
   gpc1_1 gpc4441 (
      {stage0_54[462]},
      {stage1_54[207]}
   );
   gpc1_1 gpc4442 (
      {stage0_54[463]},
      {stage1_54[208]}
   );
   gpc1_1 gpc4443 (
      {stage0_54[464]},
      {stage1_54[209]}
   );
   gpc1_1 gpc4444 (
      {stage0_54[465]},
      {stage1_54[210]}
   );
   gpc1_1 gpc4445 (
      {stage0_54[466]},
      {stage1_54[211]}
   );
   gpc1_1 gpc4446 (
      {stage0_54[467]},
      {stage1_54[212]}
   );
   gpc1_1 gpc4447 (
      {stage0_54[468]},
      {stage1_54[213]}
   );
   gpc1_1 gpc4448 (
      {stage0_54[469]},
      {stage1_54[214]}
   );
   gpc1_1 gpc4449 (
      {stage0_54[470]},
      {stage1_54[215]}
   );
   gpc1_1 gpc4450 (
      {stage0_54[471]},
      {stage1_54[216]}
   );
   gpc1_1 gpc4451 (
      {stage0_54[472]},
      {stage1_54[217]}
   );
   gpc1_1 gpc4452 (
      {stage0_54[473]},
      {stage1_54[218]}
   );
   gpc1_1 gpc4453 (
      {stage0_54[474]},
      {stage1_54[219]}
   );
   gpc1_1 gpc4454 (
      {stage0_54[475]},
      {stage1_54[220]}
   );
   gpc1_1 gpc4455 (
      {stage0_54[476]},
      {stage1_54[221]}
   );
   gpc1_1 gpc4456 (
      {stage0_54[477]},
      {stage1_54[222]}
   );
   gpc1_1 gpc4457 (
      {stage0_54[478]},
      {stage1_54[223]}
   );
   gpc1_1 gpc4458 (
      {stage0_54[479]},
      {stage1_54[224]}
   );
   gpc1_1 gpc4459 (
      {stage0_54[480]},
      {stage1_54[225]}
   );
   gpc1_1 gpc4460 (
      {stage0_54[481]},
      {stage1_54[226]}
   );
   gpc1_1 gpc4461 (
      {stage0_54[482]},
      {stage1_54[227]}
   );
   gpc1_1 gpc4462 (
      {stage0_54[483]},
      {stage1_54[228]}
   );
   gpc1_1 gpc4463 (
      {stage0_54[484]},
      {stage1_54[229]}
   );
   gpc1_1 gpc4464 (
      {stage0_54[485]},
      {stage1_54[230]}
   );
   gpc1_1 gpc4465 (
      {stage0_55[425]},
      {stage1_55[206]}
   );
   gpc1_1 gpc4466 (
      {stage0_55[426]},
      {stage1_55[207]}
   );
   gpc1_1 gpc4467 (
      {stage0_55[427]},
      {stage1_55[208]}
   );
   gpc1_1 gpc4468 (
      {stage0_55[428]},
      {stage1_55[209]}
   );
   gpc1_1 gpc4469 (
      {stage0_55[429]},
      {stage1_55[210]}
   );
   gpc1_1 gpc4470 (
      {stage0_55[430]},
      {stage1_55[211]}
   );
   gpc1_1 gpc4471 (
      {stage0_55[431]},
      {stage1_55[212]}
   );
   gpc1_1 gpc4472 (
      {stage0_55[432]},
      {stage1_55[213]}
   );
   gpc1_1 gpc4473 (
      {stage0_55[433]},
      {stage1_55[214]}
   );
   gpc1_1 gpc4474 (
      {stage0_55[434]},
      {stage1_55[215]}
   );
   gpc1_1 gpc4475 (
      {stage0_55[435]},
      {stage1_55[216]}
   );
   gpc1_1 gpc4476 (
      {stage0_55[436]},
      {stage1_55[217]}
   );
   gpc1_1 gpc4477 (
      {stage0_55[437]},
      {stage1_55[218]}
   );
   gpc1_1 gpc4478 (
      {stage0_55[438]},
      {stage1_55[219]}
   );
   gpc1_1 gpc4479 (
      {stage0_55[439]},
      {stage1_55[220]}
   );
   gpc1_1 gpc4480 (
      {stage0_55[440]},
      {stage1_55[221]}
   );
   gpc1_1 gpc4481 (
      {stage0_55[441]},
      {stage1_55[222]}
   );
   gpc1_1 gpc4482 (
      {stage0_55[442]},
      {stage1_55[223]}
   );
   gpc1_1 gpc4483 (
      {stage0_55[443]},
      {stage1_55[224]}
   );
   gpc1_1 gpc4484 (
      {stage0_55[444]},
      {stage1_55[225]}
   );
   gpc1_1 gpc4485 (
      {stage0_55[445]},
      {stage1_55[226]}
   );
   gpc1_1 gpc4486 (
      {stage0_55[446]},
      {stage1_55[227]}
   );
   gpc1_1 gpc4487 (
      {stage0_55[447]},
      {stage1_55[228]}
   );
   gpc1_1 gpc4488 (
      {stage0_55[448]},
      {stage1_55[229]}
   );
   gpc1_1 gpc4489 (
      {stage0_55[449]},
      {stage1_55[230]}
   );
   gpc1_1 gpc4490 (
      {stage0_55[450]},
      {stage1_55[231]}
   );
   gpc1_1 gpc4491 (
      {stage0_55[451]},
      {stage1_55[232]}
   );
   gpc1_1 gpc4492 (
      {stage0_55[452]},
      {stage1_55[233]}
   );
   gpc1_1 gpc4493 (
      {stage0_55[453]},
      {stage1_55[234]}
   );
   gpc1_1 gpc4494 (
      {stage0_55[454]},
      {stage1_55[235]}
   );
   gpc1_1 gpc4495 (
      {stage0_55[455]},
      {stage1_55[236]}
   );
   gpc1_1 gpc4496 (
      {stage0_55[456]},
      {stage1_55[237]}
   );
   gpc1_1 gpc4497 (
      {stage0_55[457]},
      {stage1_55[238]}
   );
   gpc1_1 gpc4498 (
      {stage0_55[458]},
      {stage1_55[239]}
   );
   gpc1_1 gpc4499 (
      {stage0_55[459]},
      {stage1_55[240]}
   );
   gpc1_1 gpc4500 (
      {stage0_55[460]},
      {stage1_55[241]}
   );
   gpc1_1 gpc4501 (
      {stage0_55[461]},
      {stage1_55[242]}
   );
   gpc1_1 gpc4502 (
      {stage0_55[462]},
      {stage1_55[243]}
   );
   gpc1_1 gpc4503 (
      {stage0_55[463]},
      {stage1_55[244]}
   );
   gpc1_1 gpc4504 (
      {stage0_55[464]},
      {stage1_55[245]}
   );
   gpc1_1 gpc4505 (
      {stage0_55[465]},
      {stage1_55[246]}
   );
   gpc1_1 gpc4506 (
      {stage0_55[466]},
      {stage1_55[247]}
   );
   gpc1_1 gpc4507 (
      {stage0_55[467]},
      {stage1_55[248]}
   );
   gpc1_1 gpc4508 (
      {stage0_55[468]},
      {stage1_55[249]}
   );
   gpc1_1 gpc4509 (
      {stage0_55[469]},
      {stage1_55[250]}
   );
   gpc1_1 gpc4510 (
      {stage0_55[470]},
      {stage1_55[251]}
   );
   gpc1_1 gpc4511 (
      {stage0_55[471]},
      {stage1_55[252]}
   );
   gpc1_1 gpc4512 (
      {stage0_55[472]},
      {stage1_55[253]}
   );
   gpc1_1 gpc4513 (
      {stage0_55[473]},
      {stage1_55[254]}
   );
   gpc1_1 gpc4514 (
      {stage0_55[474]},
      {stage1_55[255]}
   );
   gpc1_1 gpc4515 (
      {stage0_55[475]},
      {stage1_55[256]}
   );
   gpc1_1 gpc4516 (
      {stage0_55[476]},
      {stage1_55[257]}
   );
   gpc1_1 gpc4517 (
      {stage0_55[477]},
      {stage1_55[258]}
   );
   gpc1_1 gpc4518 (
      {stage0_55[478]},
      {stage1_55[259]}
   );
   gpc1_1 gpc4519 (
      {stage0_55[479]},
      {stage1_55[260]}
   );
   gpc1_1 gpc4520 (
      {stage0_55[480]},
      {stage1_55[261]}
   );
   gpc1_1 gpc4521 (
      {stage0_55[481]},
      {stage1_55[262]}
   );
   gpc1_1 gpc4522 (
      {stage0_55[482]},
      {stage1_55[263]}
   );
   gpc1_1 gpc4523 (
      {stage0_55[483]},
      {stage1_55[264]}
   );
   gpc1_1 gpc4524 (
      {stage0_55[484]},
      {stage1_55[265]}
   );
   gpc1_1 gpc4525 (
      {stage0_55[485]},
      {stage1_55[266]}
   );
   gpc1_1 gpc4526 (
      {stage0_58[460]},
      {stage1_58[194]}
   );
   gpc1_1 gpc4527 (
      {stage0_58[461]},
      {stage1_58[195]}
   );
   gpc1_1 gpc4528 (
      {stage0_58[462]},
      {stage1_58[196]}
   );
   gpc1_1 gpc4529 (
      {stage0_58[463]},
      {stage1_58[197]}
   );
   gpc1_1 gpc4530 (
      {stage0_58[464]},
      {stage1_58[198]}
   );
   gpc1_1 gpc4531 (
      {stage0_58[465]},
      {stage1_58[199]}
   );
   gpc1_1 gpc4532 (
      {stage0_58[466]},
      {stage1_58[200]}
   );
   gpc1_1 gpc4533 (
      {stage0_58[467]},
      {stage1_58[201]}
   );
   gpc1_1 gpc4534 (
      {stage0_58[468]},
      {stage1_58[202]}
   );
   gpc1_1 gpc4535 (
      {stage0_58[469]},
      {stage1_58[203]}
   );
   gpc1_1 gpc4536 (
      {stage0_58[470]},
      {stage1_58[204]}
   );
   gpc1_1 gpc4537 (
      {stage0_58[471]},
      {stage1_58[205]}
   );
   gpc1_1 gpc4538 (
      {stage0_58[472]},
      {stage1_58[206]}
   );
   gpc1_1 gpc4539 (
      {stage0_58[473]},
      {stage1_58[207]}
   );
   gpc1_1 gpc4540 (
      {stage0_58[474]},
      {stage1_58[208]}
   );
   gpc1_1 gpc4541 (
      {stage0_58[475]},
      {stage1_58[209]}
   );
   gpc1_1 gpc4542 (
      {stage0_58[476]},
      {stage1_58[210]}
   );
   gpc1_1 gpc4543 (
      {stage0_58[477]},
      {stage1_58[211]}
   );
   gpc1_1 gpc4544 (
      {stage0_58[478]},
      {stage1_58[212]}
   );
   gpc1_1 gpc4545 (
      {stage0_58[479]},
      {stage1_58[213]}
   );
   gpc1_1 gpc4546 (
      {stage0_58[480]},
      {stage1_58[214]}
   );
   gpc1_1 gpc4547 (
      {stage0_58[481]},
      {stage1_58[215]}
   );
   gpc1_1 gpc4548 (
      {stage0_58[482]},
      {stage1_58[216]}
   );
   gpc1_1 gpc4549 (
      {stage0_58[483]},
      {stage1_58[217]}
   );
   gpc1_1 gpc4550 (
      {stage0_58[484]},
      {stage1_58[218]}
   );
   gpc1_1 gpc4551 (
      {stage0_58[485]},
      {stage1_58[219]}
   );
   gpc1_1 gpc4552 (
      {stage0_59[469]},
      {stage1_59[189]}
   );
   gpc1_1 gpc4553 (
      {stage0_59[470]},
      {stage1_59[190]}
   );
   gpc1_1 gpc4554 (
      {stage0_59[471]},
      {stage1_59[191]}
   );
   gpc1_1 gpc4555 (
      {stage0_59[472]},
      {stage1_59[192]}
   );
   gpc1_1 gpc4556 (
      {stage0_59[473]},
      {stage1_59[193]}
   );
   gpc1_1 gpc4557 (
      {stage0_59[474]},
      {stage1_59[194]}
   );
   gpc1_1 gpc4558 (
      {stage0_59[475]},
      {stage1_59[195]}
   );
   gpc1_1 gpc4559 (
      {stage0_59[476]},
      {stage1_59[196]}
   );
   gpc1_1 gpc4560 (
      {stage0_59[477]},
      {stage1_59[197]}
   );
   gpc1_1 gpc4561 (
      {stage0_59[478]},
      {stage1_59[198]}
   );
   gpc1_1 gpc4562 (
      {stage0_59[479]},
      {stage1_59[199]}
   );
   gpc1_1 gpc4563 (
      {stage0_59[480]},
      {stage1_59[200]}
   );
   gpc1_1 gpc4564 (
      {stage0_59[481]},
      {stage1_59[201]}
   );
   gpc1_1 gpc4565 (
      {stage0_59[482]},
      {stage1_59[202]}
   );
   gpc1_1 gpc4566 (
      {stage0_59[483]},
      {stage1_59[203]}
   );
   gpc1_1 gpc4567 (
      {stage0_59[484]},
      {stage1_59[204]}
   );
   gpc1_1 gpc4568 (
      {stage0_59[485]},
      {stage1_59[205]}
   );
   gpc1_1 gpc4569 (
      {stage0_62[474]},
      {stage1_62[181]}
   );
   gpc1_1 gpc4570 (
      {stage0_62[475]},
      {stage1_62[182]}
   );
   gpc1_1 gpc4571 (
      {stage0_62[476]},
      {stage1_62[183]}
   );
   gpc1_1 gpc4572 (
      {stage0_62[477]},
      {stage1_62[184]}
   );
   gpc1_1 gpc4573 (
      {stage0_62[478]},
      {stage1_62[185]}
   );
   gpc1_1 gpc4574 (
      {stage0_62[479]},
      {stage1_62[186]}
   );
   gpc1_1 gpc4575 (
      {stage0_62[480]},
      {stage1_62[187]}
   );
   gpc1_1 gpc4576 (
      {stage0_62[481]},
      {stage1_62[188]}
   );
   gpc1_1 gpc4577 (
      {stage0_62[482]},
      {stage1_62[189]}
   );
   gpc1_1 gpc4578 (
      {stage0_62[483]},
      {stage1_62[190]}
   );
   gpc1_1 gpc4579 (
      {stage0_62[484]},
      {stage1_62[191]}
   );
   gpc1_1 gpc4580 (
      {stage0_62[485]},
      {stage1_62[192]}
   );
   gpc1_1 gpc4581 (
      {stage0_63[324]},
      {stage1_63[146]}
   );
   gpc1_1 gpc4582 (
      {stage0_63[325]},
      {stage1_63[147]}
   );
   gpc1_1 gpc4583 (
      {stage0_63[326]},
      {stage1_63[148]}
   );
   gpc1_1 gpc4584 (
      {stage0_63[327]},
      {stage1_63[149]}
   );
   gpc1_1 gpc4585 (
      {stage0_63[328]},
      {stage1_63[150]}
   );
   gpc1_1 gpc4586 (
      {stage0_63[329]},
      {stage1_63[151]}
   );
   gpc1_1 gpc4587 (
      {stage0_63[330]},
      {stage1_63[152]}
   );
   gpc1_1 gpc4588 (
      {stage0_63[331]},
      {stage1_63[153]}
   );
   gpc1_1 gpc4589 (
      {stage0_63[332]},
      {stage1_63[154]}
   );
   gpc1_1 gpc4590 (
      {stage0_63[333]},
      {stage1_63[155]}
   );
   gpc1_1 gpc4591 (
      {stage0_63[334]},
      {stage1_63[156]}
   );
   gpc1_1 gpc4592 (
      {stage0_63[335]},
      {stage1_63[157]}
   );
   gpc1_1 gpc4593 (
      {stage0_63[336]},
      {stage1_63[158]}
   );
   gpc1_1 gpc4594 (
      {stage0_63[337]},
      {stage1_63[159]}
   );
   gpc1_1 gpc4595 (
      {stage0_63[338]},
      {stage1_63[160]}
   );
   gpc1_1 gpc4596 (
      {stage0_63[339]},
      {stage1_63[161]}
   );
   gpc1_1 gpc4597 (
      {stage0_63[340]},
      {stage1_63[162]}
   );
   gpc1_1 gpc4598 (
      {stage0_63[341]},
      {stage1_63[163]}
   );
   gpc1_1 gpc4599 (
      {stage0_63[342]},
      {stage1_63[164]}
   );
   gpc1_1 gpc4600 (
      {stage0_63[343]},
      {stage1_63[165]}
   );
   gpc1_1 gpc4601 (
      {stage0_63[344]},
      {stage1_63[166]}
   );
   gpc1_1 gpc4602 (
      {stage0_63[345]},
      {stage1_63[167]}
   );
   gpc1_1 gpc4603 (
      {stage0_63[346]},
      {stage1_63[168]}
   );
   gpc1_1 gpc4604 (
      {stage0_63[347]},
      {stage1_63[169]}
   );
   gpc1_1 gpc4605 (
      {stage0_63[348]},
      {stage1_63[170]}
   );
   gpc1_1 gpc4606 (
      {stage0_63[349]},
      {stage1_63[171]}
   );
   gpc1_1 gpc4607 (
      {stage0_63[350]},
      {stage1_63[172]}
   );
   gpc1_1 gpc4608 (
      {stage0_63[351]},
      {stage1_63[173]}
   );
   gpc1_1 gpc4609 (
      {stage0_63[352]},
      {stage1_63[174]}
   );
   gpc1_1 gpc4610 (
      {stage0_63[353]},
      {stage1_63[175]}
   );
   gpc1_1 gpc4611 (
      {stage0_63[354]},
      {stage1_63[176]}
   );
   gpc1_1 gpc4612 (
      {stage0_63[355]},
      {stage1_63[177]}
   );
   gpc1_1 gpc4613 (
      {stage0_63[356]},
      {stage1_63[178]}
   );
   gpc1_1 gpc4614 (
      {stage0_63[357]},
      {stage1_63[179]}
   );
   gpc1_1 gpc4615 (
      {stage0_63[358]},
      {stage1_63[180]}
   );
   gpc1_1 gpc4616 (
      {stage0_63[359]},
      {stage1_63[181]}
   );
   gpc1_1 gpc4617 (
      {stage0_63[360]},
      {stage1_63[182]}
   );
   gpc1_1 gpc4618 (
      {stage0_63[361]},
      {stage1_63[183]}
   );
   gpc1_1 gpc4619 (
      {stage0_63[362]},
      {stage1_63[184]}
   );
   gpc1_1 gpc4620 (
      {stage0_63[363]},
      {stage1_63[185]}
   );
   gpc1_1 gpc4621 (
      {stage0_63[364]},
      {stage1_63[186]}
   );
   gpc1_1 gpc4622 (
      {stage0_63[365]},
      {stage1_63[187]}
   );
   gpc1_1 gpc4623 (
      {stage0_63[366]},
      {stage1_63[188]}
   );
   gpc1_1 gpc4624 (
      {stage0_63[367]},
      {stage1_63[189]}
   );
   gpc1_1 gpc4625 (
      {stage0_63[368]},
      {stage1_63[190]}
   );
   gpc1_1 gpc4626 (
      {stage0_63[369]},
      {stage1_63[191]}
   );
   gpc1_1 gpc4627 (
      {stage0_63[370]},
      {stage1_63[192]}
   );
   gpc1_1 gpc4628 (
      {stage0_63[371]},
      {stage1_63[193]}
   );
   gpc1_1 gpc4629 (
      {stage0_63[372]},
      {stage1_63[194]}
   );
   gpc1_1 gpc4630 (
      {stage0_63[373]},
      {stage1_63[195]}
   );
   gpc1_1 gpc4631 (
      {stage0_63[374]},
      {stage1_63[196]}
   );
   gpc1_1 gpc4632 (
      {stage0_63[375]},
      {stage1_63[197]}
   );
   gpc1_1 gpc4633 (
      {stage0_63[376]},
      {stage1_63[198]}
   );
   gpc1_1 gpc4634 (
      {stage0_63[377]},
      {stage1_63[199]}
   );
   gpc1_1 gpc4635 (
      {stage0_63[378]},
      {stage1_63[200]}
   );
   gpc1_1 gpc4636 (
      {stage0_63[379]},
      {stage1_63[201]}
   );
   gpc1_1 gpc4637 (
      {stage0_63[380]},
      {stage1_63[202]}
   );
   gpc1_1 gpc4638 (
      {stage0_63[381]},
      {stage1_63[203]}
   );
   gpc1_1 gpc4639 (
      {stage0_63[382]},
      {stage1_63[204]}
   );
   gpc1_1 gpc4640 (
      {stage0_63[383]},
      {stage1_63[205]}
   );
   gpc1_1 gpc4641 (
      {stage0_63[384]},
      {stage1_63[206]}
   );
   gpc1_1 gpc4642 (
      {stage0_63[385]},
      {stage1_63[207]}
   );
   gpc1_1 gpc4643 (
      {stage0_63[386]},
      {stage1_63[208]}
   );
   gpc1_1 gpc4644 (
      {stage0_63[387]},
      {stage1_63[209]}
   );
   gpc1_1 gpc4645 (
      {stage0_63[388]},
      {stage1_63[210]}
   );
   gpc1_1 gpc4646 (
      {stage0_63[389]},
      {stage1_63[211]}
   );
   gpc1_1 gpc4647 (
      {stage0_63[390]},
      {stage1_63[212]}
   );
   gpc1_1 gpc4648 (
      {stage0_63[391]},
      {stage1_63[213]}
   );
   gpc1_1 gpc4649 (
      {stage0_63[392]},
      {stage1_63[214]}
   );
   gpc1_1 gpc4650 (
      {stage0_63[393]},
      {stage1_63[215]}
   );
   gpc1_1 gpc4651 (
      {stage0_63[394]},
      {stage1_63[216]}
   );
   gpc1_1 gpc4652 (
      {stage0_63[395]},
      {stage1_63[217]}
   );
   gpc1_1 gpc4653 (
      {stage0_63[396]},
      {stage1_63[218]}
   );
   gpc1_1 gpc4654 (
      {stage0_63[397]},
      {stage1_63[219]}
   );
   gpc1_1 gpc4655 (
      {stage0_63[398]},
      {stage1_63[220]}
   );
   gpc1_1 gpc4656 (
      {stage0_63[399]},
      {stage1_63[221]}
   );
   gpc1_1 gpc4657 (
      {stage0_63[400]},
      {stage1_63[222]}
   );
   gpc1_1 gpc4658 (
      {stage0_63[401]},
      {stage1_63[223]}
   );
   gpc1_1 gpc4659 (
      {stage0_63[402]},
      {stage1_63[224]}
   );
   gpc1_1 gpc4660 (
      {stage0_63[403]},
      {stage1_63[225]}
   );
   gpc1_1 gpc4661 (
      {stage0_63[404]},
      {stage1_63[226]}
   );
   gpc1_1 gpc4662 (
      {stage0_63[405]},
      {stage1_63[227]}
   );
   gpc1_1 gpc4663 (
      {stage0_63[406]},
      {stage1_63[228]}
   );
   gpc1_1 gpc4664 (
      {stage0_63[407]},
      {stage1_63[229]}
   );
   gpc1_1 gpc4665 (
      {stage0_63[408]},
      {stage1_63[230]}
   );
   gpc1_1 gpc4666 (
      {stage0_63[409]},
      {stage1_63[231]}
   );
   gpc1_1 gpc4667 (
      {stage0_63[410]},
      {stage1_63[232]}
   );
   gpc1_1 gpc4668 (
      {stage0_63[411]},
      {stage1_63[233]}
   );
   gpc1_1 gpc4669 (
      {stage0_63[412]},
      {stage1_63[234]}
   );
   gpc1_1 gpc4670 (
      {stage0_63[413]},
      {stage1_63[235]}
   );
   gpc1_1 gpc4671 (
      {stage0_63[414]},
      {stage1_63[236]}
   );
   gpc1_1 gpc4672 (
      {stage0_63[415]},
      {stage1_63[237]}
   );
   gpc1_1 gpc4673 (
      {stage0_63[416]},
      {stage1_63[238]}
   );
   gpc1_1 gpc4674 (
      {stage0_63[417]},
      {stage1_63[239]}
   );
   gpc1_1 gpc4675 (
      {stage0_63[418]},
      {stage1_63[240]}
   );
   gpc1_1 gpc4676 (
      {stage0_63[419]},
      {stage1_63[241]}
   );
   gpc1_1 gpc4677 (
      {stage0_63[420]},
      {stage1_63[242]}
   );
   gpc1_1 gpc4678 (
      {stage0_63[421]},
      {stage1_63[243]}
   );
   gpc1_1 gpc4679 (
      {stage0_63[422]},
      {stage1_63[244]}
   );
   gpc1_1 gpc4680 (
      {stage0_63[423]},
      {stage1_63[245]}
   );
   gpc1_1 gpc4681 (
      {stage0_63[424]},
      {stage1_63[246]}
   );
   gpc1_1 gpc4682 (
      {stage0_63[425]},
      {stage1_63[247]}
   );
   gpc1_1 gpc4683 (
      {stage0_63[426]},
      {stage1_63[248]}
   );
   gpc1_1 gpc4684 (
      {stage0_63[427]},
      {stage1_63[249]}
   );
   gpc1_1 gpc4685 (
      {stage0_63[428]},
      {stage1_63[250]}
   );
   gpc1_1 gpc4686 (
      {stage0_63[429]},
      {stage1_63[251]}
   );
   gpc1_1 gpc4687 (
      {stage0_63[430]},
      {stage1_63[252]}
   );
   gpc1_1 gpc4688 (
      {stage0_63[431]},
      {stage1_63[253]}
   );
   gpc1_1 gpc4689 (
      {stage0_63[432]},
      {stage1_63[254]}
   );
   gpc1_1 gpc4690 (
      {stage0_63[433]},
      {stage1_63[255]}
   );
   gpc1_1 gpc4691 (
      {stage0_63[434]},
      {stage1_63[256]}
   );
   gpc1_1 gpc4692 (
      {stage0_63[435]},
      {stage1_63[257]}
   );
   gpc1_1 gpc4693 (
      {stage0_63[436]},
      {stage1_63[258]}
   );
   gpc1_1 gpc4694 (
      {stage0_63[437]},
      {stage1_63[259]}
   );
   gpc1_1 gpc4695 (
      {stage0_63[438]},
      {stage1_63[260]}
   );
   gpc1_1 gpc4696 (
      {stage0_63[439]},
      {stage1_63[261]}
   );
   gpc1_1 gpc4697 (
      {stage0_63[440]},
      {stage1_63[262]}
   );
   gpc1_1 gpc4698 (
      {stage0_63[441]},
      {stage1_63[263]}
   );
   gpc1_1 gpc4699 (
      {stage0_63[442]},
      {stage1_63[264]}
   );
   gpc1_1 gpc4700 (
      {stage0_63[443]},
      {stage1_63[265]}
   );
   gpc1_1 gpc4701 (
      {stage0_63[444]},
      {stage1_63[266]}
   );
   gpc1_1 gpc4702 (
      {stage0_63[445]},
      {stage1_63[267]}
   );
   gpc1_1 gpc4703 (
      {stage0_63[446]},
      {stage1_63[268]}
   );
   gpc1_1 gpc4704 (
      {stage0_63[447]},
      {stage1_63[269]}
   );
   gpc1_1 gpc4705 (
      {stage0_63[448]},
      {stage1_63[270]}
   );
   gpc1_1 gpc4706 (
      {stage0_63[449]},
      {stage1_63[271]}
   );
   gpc1_1 gpc4707 (
      {stage0_63[450]},
      {stage1_63[272]}
   );
   gpc1_1 gpc4708 (
      {stage0_63[451]},
      {stage1_63[273]}
   );
   gpc1_1 gpc4709 (
      {stage0_63[452]},
      {stage1_63[274]}
   );
   gpc1_1 gpc4710 (
      {stage0_63[453]},
      {stage1_63[275]}
   );
   gpc1_1 gpc4711 (
      {stage0_63[454]},
      {stage1_63[276]}
   );
   gpc1_1 gpc4712 (
      {stage0_63[455]},
      {stage1_63[277]}
   );
   gpc1_1 gpc4713 (
      {stage0_63[456]},
      {stage1_63[278]}
   );
   gpc1_1 gpc4714 (
      {stage0_63[457]},
      {stage1_63[279]}
   );
   gpc1_1 gpc4715 (
      {stage0_63[458]},
      {stage1_63[280]}
   );
   gpc1_1 gpc4716 (
      {stage0_63[459]},
      {stage1_63[281]}
   );
   gpc1_1 gpc4717 (
      {stage0_63[460]},
      {stage1_63[282]}
   );
   gpc1_1 gpc4718 (
      {stage0_63[461]},
      {stage1_63[283]}
   );
   gpc1_1 gpc4719 (
      {stage0_63[462]},
      {stage1_63[284]}
   );
   gpc1_1 gpc4720 (
      {stage0_63[463]},
      {stage1_63[285]}
   );
   gpc1_1 gpc4721 (
      {stage0_63[464]},
      {stage1_63[286]}
   );
   gpc1_1 gpc4722 (
      {stage0_63[465]},
      {stage1_63[287]}
   );
   gpc1_1 gpc4723 (
      {stage0_63[466]},
      {stage1_63[288]}
   );
   gpc1_1 gpc4724 (
      {stage0_63[467]},
      {stage1_63[289]}
   );
   gpc1_1 gpc4725 (
      {stage0_63[468]},
      {stage1_63[290]}
   );
   gpc1_1 gpc4726 (
      {stage0_63[469]},
      {stage1_63[291]}
   );
   gpc1_1 gpc4727 (
      {stage0_63[470]},
      {stage1_63[292]}
   );
   gpc1_1 gpc4728 (
      {stage0_63[471]},
      {stage1_63[293]}
   );
   gpc1_1 gpc4729 (
      {stage0_63[472]},
      {stage1_63[294]}
   );
   gpc1_1 gpc4730 (
      {stage0_63[473]},
      {stage1_63[295]}
   );
   gpc1_1 gpc4731 (
      {stage0_63[474]},
      {stage1_63[296]}
   );
   gpc1_1 gpc4732 (
      {stage0_63[475]},
      {stage1_63[297]}
   );
   gpc1_1 gpc4733 (
      {stage0_63[476]},
      {stage1_63[298]}
   );
   gpc1_1 gpc4734 (
      {stage0_63[477]},
      {stage1_63[299]}
   );
   gpc1_1 gpc4735 (
      {stage0_63[478]},
      {stage1_63[300]}
   );
   gpc1_1 gpc4736 (
      {stage0_63[479]},
      {stage1_63[301]}
   );
   gpc1_1 gpc4737 (
      {stage0_63[480]},
      {stage1_63[302]}
   );
   gpc1_1 gpc4738 (
      {stage0_63[481]},
      {stage1_63[303]}
   );
   gpc1_1 gpc4739 (
      {stage0_63[482]},
      {stage1_63[304]}
   );
   gpc1_1 gpc4740 (
      {stage0_63[483]},
      {stage1_63[305]}
   );
   gpc1_1 gpc4741 (
      {stage0_63[484]},
      {stage1_63[306]}
   );
   gpc1_1 gpc4742 (
      {stage0_63[485]},
      {stage1_63[307]}
   );
   gpc606_5 gpc4743 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc4744 (
      {stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc606_5 gpc4745 (
      {stage1_0[12], stage1_0[13], stage1_0[14], stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc615_5 gpc4746 (
      {stage1_0[18], stage1_0[19], stage1_0[20], stage1_0[21], stage1_0[22]},
      {stage1_1[0]},
      {stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc615_5 gpc4747 (
      {stage1_0[23], stage1_0[24], stage1_0[25], stage1_0[26], stage1_0[27]},
      {stage1_1[1]},
      {stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27], stage1_2[28], stage1_2[29]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc615_5 gpc4748 (
      {stage1_0[28], stage1_0[29], stage1_0[30], stage1_0[31], stage1_0[32]},
      {stage1_1[2]},
      {stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33], stage1_2[34], stage1_2[35]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc615_5 gpc4749 (
      {stage1_0[33], stage1_0[34], stage1_0[35], stage1_0[36], stage1_0[37]},
      {stage1_1[3]},
      {stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39], stage1_2[40], stage1_2[41]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc615_5 gpc4750 (
      {stage1_0[38], stage1_0[39], stage1_0[40], stage1_0[41], stage1_0[42]},
      {stage1_1[4]},
      {stage1_2[42], stage1_2[43], stage1_2[44], stage1_2[45], stage1_2[46], stage1_2[47]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc615_5 gpc4751 (
      {stage1_0[43], stage1_0[44], stage1_0[45], stage1_0[46], stage1_0[47]},
      {stage1_1[5]},
      {stage1_2[48], stage1_2[49], stage1_2[50], stage1_2[51], stage1_2[52], stage1_2[53]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc615_5 gpc4752 (
      {stage1_0[48], stage1_0[49], stage1_0[50], stage1_0[51], stage1_0[52]},
      {stage1_1[6]},
      {stage1_2[54], stage1_2[55], stage1_2[56], stage1_2[57], stage1_2[58], stage1_2[59]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc615_5 gpc4753 (
      {stage1_0[53], stage1_0[54], stage1_0[55], stage1_0[56], stage1_0[57]},
      {stage1_1[7]},
      {stage1_2[60], stage1_2[61], stage1_2[62], stage1_2[63], stage1_2[64], stage1_2[65]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc615_5 gpc4754 (
      {stage1_0[58], stage1_0[59], stage1_0[60], stage1_0[61], stage1_0[62]},
      {stage1_1[8]},
      {stage1_2[66], stage1_2[67], stage1_2[68], stage1_2[69], stage1_2[70], stage1_2[71]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc615_5 gpc4755 (
      {stage1_0[63], stage1_0[64], stage1_0[65], stage1_0[66], stage1_0[67]},
      {stage1_1[9]},
      {stage1_2[72], stage1_2[73], stage1_2[74], stage1_2[75], stage1_2[76], stage1_2[77]},
      {stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12],stage2_0[12]}
   );
   gpc615_5 gpc4756 (
      {stage1_0[68], stage1_0[69], stage1_0[70], stage1_0[71], stage1_0[72]},
      {stage1_1[10]},
      {stage1_2[78], stage1_2[79], stage1_2[80], stage1_2[81], stage1_2[82], stage1_2[83]},
      {stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13],stage2_0[13]}
   );
   gpc615_5 gpc4757 (
      {stage1_0[73], stage1_0[74], stage1_0[75], stage1_0[76], stage1_0[77]},
      {stage1_1[11]},
      {stage1_2[84], stage1_2[85], stage1_2[86], stage1_2[87], stage1_2[88], stage1_2[89]},
      {stage2_4[14],stage2_3[14],stage2_2[14],stage2_1[14],stage2_0[14]}
   );
   gpc615_5 gpc4758 (
      {stage1_0[78], stage1_0[79], stage1_0[80], stage1_0[81], stage1_0[82]},
      {stage1_1[12]},
      {stage1_2[90], stage1_2[91], stage1_2[92], stage1_2[93], stage1_2[94], stage1_2[95]},
      {stage2_4[15],stage2_3[15],stage2_2[15],stage2_1[15],stage2_0[15]}
   );
   gpc615_5 gpc4759 (
      {stage1_0[83], stage1_0[84], stage1_0[85], stage1_0[86], stage1_0[87]},
      {stage1_1[13]},
      {stage1_2[96], stage1_2[97], stage1_2[98], stage1_2[99], stage1_2[100], stage1_2[101]},
      {stage2_4[16],stage2_3[16],stage2_2[16],stage2_1[16],stage2_0[16]}
   );
   gpc615_5 gpc4760 (
      {stage1_0[88], stage1_0[89], stage1_0[90], stage1_0[91], stage1_0[92]},
      {stage1_1[14]},
      {stage1_2[102], stage1_2[103], stage1_2[104], stage1_2[105], stage1_2[106], stage1_2[107]},
      {stage2_4[17],stage2_3[17],stage2_2[17],stage2_1[17],stage2_0[17]}
   );
   gpc615_5 gpc4761 (
      {stage1_0[93], stage1_0[94], stage1_0[95], stage1_0[96], stage1_0[97]},
      {stage1_1[15]},
      {stage1_2[108], stage1_2[109], stage1_2[110], stage1_2[111], stage1_2[112], stage1_2[113]},
      {stage2_4[18],stage2_3[18],stage2_2[18],stage2_1[18],stage2_0[18]}
   );
   gpc615_5 gpc4762 (
      {stage1_0[98], stage1_0[99], stage1_0[100], stage1_0[101], stage1_0[102]},
      {stage1_1[16]},
      {stage1_2[114], stage1_2[115], stage1_2[116], stage1_2[117], stage1_2[118], stage1_2[119]},
      {stage2_4[19],stage2_3[19],stage2_2[19],stage2_1[19],stage2_0[19]}
   );
   gpc615_5 gpc4763 (
      {stage1_0[103], stage1_0[104], stage1_0[105], stage1_0[106], stage1_0[107]},
      {stage1_1[17]},
      {stage1_2[120], stage1_2[121], stage1_2[122], stage1_2[123], stage1_2[124], stage1_2[125]},
      {stage2_4[20],stage2_3[20],stage2_2[20],stage2_1[20],stage2_0[20]}
   );
   gpc606_5 gpc4764 (
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage2_5[0],stage2_4[21],stage2_3[21],stage2_2[21],stage2_1[21]}
   );
   gpc606_5 gpc4765 (
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage2_5[1],stage2_4[22],stage2_3[22],stage2_2[22],stage2_1[22]}
   );
   gpc606_5 gpc4766 (
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage2_5[2],stage2_4[23],stage2_3[23],stage2_2[23],stage2_1[23]}
   );
   gpc606_5 gpc4767 (
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23]},
      {stage2_5[3],stage2_4[24],stage2_3[24],stage2_2[24],stage2_1[24]}
   );
   gpc606_5 gpc4768 (
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27], stage1_3[28], stage1_3[29]},
      {stage2_5[4],stage2_4[25],stage2_3[25],stage2_2[25],stage2_1[25]}
   );
   gpc606_5 gpc4769 (
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_3[30], stage1_3[31], stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35]},
      {stage2_5[5],stage2_4[26],stage2_3[26],stage2_2[26],stage2_1[26]}
   );
   gpc606_5 gpc4770 (
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59]},
      {stage1_3[36], stage1_3[37], stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41]},
      {stage2_5[6],stage2_4[27],stage2_3[27],stage2_2[27],stage2_1[27]}
   );
   gpc606_5 gpc4771 (
      {stage1_1[60], stage1_1[61], stage1_1[62], stage1_1[63], stage1_1[64], stage1_1[65]},
      {stage1_3[42], stage1_3[43], stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47]},
      {stage2_5[7],stage2_4[28],stage2_3[28],stage2_2[28],stage2_1[28]}
   );
   gpc606_5 gpc4772 (
      {stage1_1[66], stage1_1[67], stage1_1[68], stage1_1[69], stage1_1[70], stage1_1[71]},
      {stage1_3[48], stage1_3[49], stage1_3[50], stage1_3[51], stage1_3[52], stage1_3[53]},
      {stage2_5[8],stage2_4[29],stage2_3[29],stage2_2[29],stage2_1[29]}
   );
   gpc606_5 gpc4773 (
      {stage1_1[72], stage1_1[73], stage1_1[74], stage1_1[75], stage1_1[76], stage1_1[77]},
      {stage1_3[54], stage1_3[55], stage1_3[56], stage1_3[57], stage1_3[58], stage1_3[59]},
      {stage2_5[9],stage2_4[30],stage2_3[30],stage2_2[30],stage2_1[30]}
   );
   gpc606_5 gpc4774 (
      {stage1_1[78], stage1_1[79], stage1_1[80], stage1_1[81], stage1_1[82], stage1_1[83]},
      {stage1_3[60], stage1_3[61], stage1_3[62], stage1_3[63], stage1_3[64], stage1_3[65]},
      {stage2_5[10],stage2_4[31],stage2_3[31],stage2_2[31],stage2_1[31]}
   );
   gpc606_5 gpc4775 (
      {stage1_1[84], stage1_1[85], stage1_1[86], stage1_1[87], stage1_1[88], stage1_1[89]},
      {stage1_3[66], stage1_3[67], stage1_3[68], stage1_3[69], stage1_3[70], stage1_3[71]},
      {stage2_5[11],stage2_4[32],stage2_3[32],stage2_2[32],stage2_1[32]}
   );
   gpc606_5 gpc4776 (
      {stage1_1[90], stage1_1[91], stage1_1[92], stage1_1[93], stage1_1[94], stage1_1[95]},
      {stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75], stage1_3[76], stage1_3[77]},
      {stage2_5[12],stage2_4[33],stage2_3[33],stage2_2[33],stage2_1[33]}
   );
   gpc606_5 gpc4777 (
      {stage1_1[96], stage1_1[97], stage1_1[98], stage1_1[99], stage1_1[100], stage1_1[101]},
      {stage1_3[78], stage1_3[79], stage1_3[80], stage1_3[81], stage1_3[82], stage1_3[83]},
      {stage2_5[13],stage2_4[34],stage2_3[34],stage2_2[34],stage2_1[34]}
   );
   gpc606_5 gpc4778 (
      {stage1_1[102], stage1_1[103], stage1_1[104], stage1_1[105], stage1_1[106], stage1_1[107]},
      {stage1_3[84], stage1_3[85], stage1_3[86], stage1_3[87], stage1_3[88], stage1_3[89]},
      {stage2_5[14],stage2_4[35],stage2_3[35],stage2_2[35],stage2_1[35]}
   );
   gpc606_5 gpc4779 (
      {stage1_1[108], stage1_1[109], stage1_1[110], stage1_1[111], stage1_1[112], stage1_1[113]},
      {stage1_3[90], stage1_3[91], stage1_3[92], stage1_3[93], stage1_3[94], stage1_3[95]},
      {stage2_5[15],stage2_4[36],stage2_3[36],stage2_2[36],stage2_1[36]}
   );
   gpc606_5 gpc4780 (
      {stage1_1[114], stage1_1[115], stage1_1[116], stage1_1[117], stage1_1[118], stage1_1[119]},
      {stage1_3[96], stage1_3[97], stage1_3[98], stage1_3[99], stage1_3[100], stage1_3[101]},
      {stage2_5[16],stage2_4[37],stage2_3[37],stage2_2[37],stage2_1[37]}
   );
   gpc606_5 gpc4781 (
      {stage1_1[120], stage1_1[121], stage1_1[122], stage1_1[123], stage1_1[124], stage1_1[125]},
      {stage1_3[102], stage1_3[103], stage1_3[104], stage1_3[105], stage1_3[106], stage1_3[107]},
      {stage2_5[17],stage2_4[38],stage2_3[38],stage2_2[38],stage2_1[38]}
   );
   gpc606_5 gpc4782 (
      {stage1_1[126], stage1_1[127], stage1_1[128], stage1_1[129], stage1_1[130], stage1_1[131]},
      {stage1_3[108], stage1_3[109], stage1_3[110], stage1_3[111], stage1_3[112], stage1_3[113]},
      {stage2_5[18],stage2_4[39],stage2_3[39],stage2_2[39],stage2_1[39]}
   );
   gpc606_5 gpc4783 (
      {stage1_1[132], stage1_1[133], stage1_1[134], stage1_1[135], stage1_1[136], stage1_1[137]},
      {stage1_3[114], stage1_3[115], stage1_3[116], stage1_3[117], stage1_3[118], stage1_3[119]},
      {stage2_5[19],stage2_4[40],stage2_3[40],stage2_2[40],stage2_1[40]}
   );
   gpc606_5 gpc4784 (
      {stage1_1[138], stage1_1[139], stage1_1[140], stage1_1[141], stage1_1[142], stage1_1[143]},
      {stage1_3[120], stage1_3[121], stage1_3[122], stage1_3[123], stage1_3[124], stage1_3[125]},
      {stage2_5[20],stage2_4[41],stage2_3[41],stage2_2[41],stage2_1[41]}
   );
   gpc606_5 gpc4785 (
      {stage1_1[144], stage1_1[145], stage1_1[146], stage1_1[147], stage1_1[148], stage1_1[149]},
      {stage1_3[126], stage1_3[127], stage1_3[128], stage1_3[129], stage1_3[130], stage1_3[131]},
      {stage2_5[21],stage2_4[42],stage2_3[42],stage2_2[42],stage2_1[42]}
   );
   gpc606_5 gpc4786 (
      {stage1_1[150], stage1_1[151], stage1_1[152], stage1_1[153], stage1_1[154], stage1_1[155]},
      {stage1_3[132], stage1_3[133], stage1_3[134], stage1_3[135], stage1_3[136], stage1_3[137]},
      {stage2_5[22],stage2_4[43],stage2_3[43],stage2_2[43],stage2_1[43]}
   );
   gpc606_5 gpc4787 (
      {stage1_1[156], stage1_1[157], stage1_1[158], stage1_1[159], stage1_1[160], stage1_1[161]},
      {stage1_3[138], stage1_3[139], stage1_3[140], stage1_3[141], stage1_3[142], stage1_3[143]},
      {stage2_5[23],stage2_4[44],stage2_3[44],stage2_2[44],stage2_1[44]}
   );
   gpc606_5 gpc4788 (
      {stage1_1[162], stage1_1[163], stage1_1[164], stage1_1[165], stage1_1[166], stage1_1[167]},
      {stage1_3[144], stage1_3[145], stage1_3[146], stage1_3[147], stage1_3[148], stage1_3[149]},
      {stage2_5[24],stage2_4[45],stage2_3[45],stage2_2[45],stage2_1[45]}
   );
   gpc606_5 gpc4789 (
      {stage1_2[126], stage1_2[127], stage1_2[128], stage1_2[129], stage1_2[130], stage1_2[131]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[25],stage2_4[46],stage2_3[46],stage2_2[46]}
   );
   gpc606_5 gpc4790 (
      {stage1_2[132], stage1_2[133], stage1_2[134], stage1_2[135], stage1_2[136], stage1_2[137]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[26],stage2_4[47],stage2_3[47],stage2_2[47]}
   );
   gpc606_5 gpc4791 (
      {stage1_2[138], stage1_2[139], stage1_2[140], stage1_2[141], stage1_2[142], stage1_2[143]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[27],stage2_4[48],stage2_3[48],stage2_2[48]}
   );
   gpc1343_5 gpc4792 (
      {stage1_4[18], stage1_4[19], stage1_4[20]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3]},
      {stage1_6[0], stage1_6[1], stage1_6[2]},
      {stage1_7[0]},
      {stage2_8[0],stage2_7[0],stage2_6[3],stage2_5[28],stage2_4[49]}
   );
   gpc1406_5 gpc4793 (
      {stage1_4[21], stage1_4[22], stage1_4[23], stage1_4[24], stage1_4[25], stage1_4[26]},
      {stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6]},
      {stage1_7[1]},
      {stage2_8[1],stage2_7[1],stage2_6[4],stage2_5[29],stage2_4[50]}
   );
   gpc606_5 gpc4794 (
      {stage1_4[27], stage1_4[28], stage1_4[29], stage1_4[30], stage1_4[31], stage1_4[32]},
      {stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12]},
      {stage2_8[2],stage2_7[2],stage2_6[5],stage2_5[30],stage2_4[51]}
   );
   gpc606_5 gpc4795 (
      {stage1_4[33], stage1_4[34], stage1_4[35], stage1_4[36], stage1_4[37], stage1_4[38]},
      {stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17], stage1_6[18]},
      {stage2_8[3],stage2_7[3],stage2_6[6],stage2_5[31],stage2_4[52]}
   );
   gpc606_5 gpc4796 (
      {stage1_4[39], stage1_4[40], stage1_4[41], stage1_4[42], stage1_4[43], stage1_4[44]},
      {stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23], stage1_6[24]},
      {stage2_8[4],stage2_7[4],stage2_6[7],stage2_5[32],stage2_4[53]}
   );
   gpc606_5 gpc4797 (
      {stage1_4[45], stage1_4[46], stage1_4[47], stage1_4[48], stage1_4[49], stage1_4[50]},
      {stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29], stage1_6[30]},
      {stage2_8[5],stage2_7[5],stage2_6[8],stage2_5[33],stage2_4[54]}
   );
   gpc606_5 gpc4798 (
      {stage1_4[51], stage1_4[52], stage1_4[53], stage1_4[54], stage1_4[55], stage1_4[56]},
      {stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35], stage1_6[36]},
      {stage2_8[6],stage2_7[6],stage2_6[9],stage2_5[34],stage2_4[55]}
   );
   gpc606_5 gpc4799 (
      {stage1_4[57], stage1_4[58], stage1_4[59], stage1_4[60], stage1_4[61], stage1_4[62]},
      {stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41], stage1_6[42]},
      {stage2_8[7],stage2_7[7],stage2_6[10],stage2_5[35],stage2_4[56]}
   );
   gpc606_5 gpc4800 (
      {stage1_4[63], stage1_4[64], stage1_4[65], stage1_4[66], stage1_4[67], stage1_4[68]},
      {stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47], stage1_6[48]},
      {stage2_8[8],stage2_7[8],stage2_6[11],stage2_5[36],stage2_4[57]}
   );
   gpc606_5 gpc4801 (
      {stage1_4[69], stage1_4[70], stage1_4[71], stage1_4[72], stage1_4[73], stage1_4[74]},
      {stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53], stage1_6[54]},
      {stage2_8[9],stage2_7[9],stage2_6[12],stage2_5[37],stage2_4[58]}
   );
   gpc606_5 gpc4802 (
      {stage1_4[75], stage1_4[76], stage1_4[77], stage1_4[78], stage1_4[79], stage1_4[80]},
      {stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59], stage1_6[60]},
      {stage2_8[10],stage2_7[10],stage2_6[13],stage2_5[38],stage2_4[59]}
   );
   gpc606_5 gpc4803 (
      {stage1_4[81], stage1_4[82], stage1_4[83], stage1_4[84], stage1_4[85], stage1_4[86]},
      {stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65], stage1_6[66]},
      {stage2_8[11],stage2_7[11],stage2_6[14],stage2_5[39],stage2_4[60]}
   );
   gpc606_5 gpc4804 (
      {stage1_4[87], stage1_4[88], stage1_4[89], stage1_4[90], stage1_4[91], stage1_4[92]},
      {stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71], stage1_6[72]},
      {stage2_8[12],stage2_7[12],stage2_6[15],stage2_5[40],stage2_4[61]}
   );
   gpc606_5 gpc4805 (
      {stage1_4[93], stage1_4[94], stage1_4[95], stage1_4[96], stage1_4[97], stage1_4[98]},
      {stage1_6[73], stage1_6[74], stage1_6[75], stage1_6[76], stage1_6[77], stage1_6[78]},
      {stage2_8[13],stage2_7[13],stage2_6[16],stage2_5[41],stage2_4[62]}
   );
   gpc606_5 gpc4806 (
      {stage1_4[99], stage1_4[100], stage1_4[101], stage1_4[102], stage1_4[103], stage1_4[104]},
      {stage1_6[79], stage1_6[80], stage1_6[81], stage1_6[82], stage1_6[83], stage1_6[84]},
      {stage2_8[14],stage2_7[14],stage2_6[17],stage2_5[42],stage2_4[63]}
   );
   gpc606_5 gpc4807 (
      {stage1_4[105], stage1_4[106], stage1_4[107], stage1_4[108], stage1_4[109], stage1_4[110]},
      {stage1_6[85], stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89], stage1_6[90]},
      {stage2_8[15],stage2_7[15],stage2_6[18],stage2_5[43],stage2_4[64]}
   );
   gpc606_5 gpc4808 (
      {stage1_4[111], stage1_4[112], stage1_4[113], stage1_4[114], stage1_4[115], stage1_4[116]},
      {stage1_6[91], stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95], stage1_6[96]},
      {stage2_8[16],stage2_7[16],stage2_6[19],stage2_5[44],stage2_4[65]}
   );
   gpc606_5 gpc4809 (
      {stage1_4[117], stage1_4[118], stage1_4[119], stage1_4[120], stage1_4[121], stage1_4[122]},
      {stage1_6[97], stage1_6[98], stage1_6[99], stage1_6[100], stage1_6[101], stage1_6[102]},
      {stage2_8[17],stage2_7[17],stage2_6[20],stage2_5[45],stage2_4[66]}
   );
   gpc606_5 gpc4810 (
      {stage1_4[123], stage1_4[124], stage1_4[125], stage1_4[126], stage1_4[127], stage1_4[128]},
      {stage1_6[103], stage1_6[104], stage1_6[105], stage1_6[106], stage1_6[107], stage1_6[108]},
      {stage2_8[18],stage2_7[18],stage2_6[21],stage2_5[46],stage2_4[67]}
   );
   gpc606_5 gpc4811 (
      {stage1_4[129], stage1_4[130], stage1_4[131], stage1_4[132], stage1_4[133], stage1_4[134]},
      {stage1_6[109], stage1_6[110], stage1_6[111], stage1_6[112], stage1_6[113], stage1_6[114]},
      {stage2_8[19],stage2_7[19],stage2_6[22],stage2_5[47],stage2_4[68]}
   );
   gpc606_5 gpc4812 (
      {stage1_4[135], stage1_4[136], stage1_4[137], stage1_4[138], stage1_4[139], stage1_4[140]},
      {stage1_6[115], stage1_6[116], stage1_6[117], stage1_6[118], stage1_6[119], stage1_6[120]},
      {stage2_8[20],stage2_7[20],stage2_6[23],stage2_5[48],stage2_4[69]}
   );
   gpc606_5 gpc4813 (
      {stage1_4[141], stage1_4[142], stage1_4[143], stage1_4[144], stage1_4[145], stage1_4[146]},
      {stage1_6[121], stage1_6[122], stage1_6[123], stage1_6[124], stage1_6[125], stage1_6[126]},
      {stage2_8[21],stage2_7[21],stage2_6[24],stage2_5[49],stage2_4[70]}
   );
   gpc606_5 gpc4814 (
      {stage1_4[147], stage1_4[148], stage1_4[149], stage1_4[150], stage1_4[151], stage1_4[152]},
      {stage1_6[127], stage1_6[128], stage1_6[129], stage1_6[130], stage1_6[131], stage1_6[132]},
      {stage2_8[22],stage2_7[22],stage2_6[25],stage2_5[50],stage2_4[71]}
   );
   gpc606_5 gpc4815 (
      {stage1_4[153], stage1_4[154], stage1_4[155], stage1_4[156], stage1_4[157], stage1_4[158]},
      {stage1_6[133], stage1_6[134], stage1_6[135], stage1_6[136], stage1_6[137], stage1_6[138]},
      {stage2_8[23],stage2_7[23],stage2_6[26],stage2_5[51],stage2_4[72]}
   );
   gpc606_5 gpc4816 (
      {stage1_4[159], stage1_4[160], stage1_4[161], stage1_4[162], stage1_4[163], stage1_4[164]},
      {stage1_6[139], stage1_6[140], stage1_6[141], stage1_6[142], stage1_6[143], stage1_6[144]},
      {stage2_8[24],stage2_7[24],stage2_6[27],stage2_5[52],stage2_4[73]}
   );
   gpc606_5 gpc4817 (
      {stage1_4[165], stage1_4[166], stage1_4[167], stage1_4[168], stage1_4[169], stage1_4[170]},
      {stage1_6[145], stage1_6[146], stage1_6[147], stage1_6[148], stage1_6[149], stage1_6[150]},
      {stage2_8[25],stage2_7[25],stage2_6[28],stage2_5[53],stage2_4[74]}
   );
   gpc606_5 gpc4818 (
      {stage1_4[171], stage1_4[172], stage1_4[173], stage1_4[174], stage1_4[175], stage1_4[176]},
      {stage1_6[151], stage1_6[152], stage1_6[153], stage1_6[154], stage1_6[155], stage1_6[156]},
      {stage2_8[26],stage2_7[26],stage2_6[29],stage2_5[54],stage2_4[75]}
   );
   gpc606_5 gpc4819 (
      {stage1_4[177], stage1_4[178], stage1_4[179], stage1_4[180], stage1_4[181], stage1_4[182]},
      {stage1_6[157], stage1_6[158], stage1_6[159], stage1_6[160], stage1_6[161], stage1_6[162]},
      {stage2_8[27],stage2_7[27],stage2_6[30],stage2_5[55],stage2_4[76]}
   );
   gpc606_5 gpc4820 (
      {stage1_4[183], stage1_4[184], stage1_4[185], stage1_4[186], stage1_4[187], stage1_4[188]},
      {stage1_6[163], stage1_6[164], stage1_6[165], stage1_6[166], stage1_6[167], stage1_6[168]},
      {stage2_8[28],stage2_7[28],stage2_6[31],stage2_5[56],stage2_4[77]}
   );
   gpc606_5 gpc4821 (
      {stage1_4[189], stage1_4[190], stage1_4[191], stage1_4[192], stage1_4[193], stage1_4[194]},
      {stage1_6[169], stage1_6[170], stage1_6[171], stage1_6[172], stage1_6[173], stage1_6[174]},
      {stage2_8[29],stage2_7[29],stage2_6[32],stage2_5[57],stage2_4[78]}
   );
   gpc606_5 gpc4822 (
      {stage1_5[4], stage1_5[5], stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9]},
      {stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5], stage1_7[6], stage1_7[7]},
      {stage2_9[0],stage2_8[30],stage2_7[30],stage2_6[33],stage2_5[58]}
   );
   gpc606_5 gpc4823 (
      {stage1_5[10], stage1_5[11], stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15]},
      {stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12], stage1_7[13]},
      {stage2_9[1],stage2_8[31],stage2_7[31],stage2_6[34],stage2_5[59]}
   );
   gpc606_5 gpc4824 (
      {stage1_5[16], stage1_5[17], stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21]},
      {stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17], stage1_7[18], stage1_7[19]},
      {stage2_9[2],stage2_8[32],stage2_7[32],stage2_6[35],stage2_5[60]}
   );
   gpc606_5 gpc4825 (
      {stage1_5[22], stage1_5[23], stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27]},
      {stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23], stage1_7[24], stage1_7[25]},
      {stage2_9[3],stage2_8[33],stage2_7[33],stage2_6[36],stage2_5[61]}
   );
   gpc606_5 gpc4826 (
      {stage1_5[28], stage1_5[29], stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33]},
      {stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29], stage1_7[30], stage1_7[31]},
      {stage2_9[4],stage2_8[34],stage2_7[34],stage2_6[37],stage2_5[62]}
   );
   gpc606_5 gpc4827 (
      {stage1_5[34], stage1_5[35], stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39]},
      {stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35], stage1_7[36], stage1_7[37]},
      {stage2_9[5],stage2_8[35],stage2_7[35],stage2_6[38],stage2_5[63]}
   );
   gpc606_5 gpc4828 (
      {stage1_5[40], stage1_5[41], stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45]},
      {stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41], stage1_7[42], stage1_7[43]},
      {stage2_9[6],stage2_8[36],stage2_7[36],stage2_6[39],stage2_5[64]}
   );
   gpc606_5 gpc4829 (
      {stage1_5[46], stage1_5[47], stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51]},
      {stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47], stage1_7[48], stage1_7[49]},
      {stage2_9[7],stage2_8[37],stage2_7[37],stage2_6[40],stage2_5[65]}
   );
   gpc606_5 gpc4830 (
      {stage1_5[52], stage1_5[53], stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57]},
      {stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53], stage1_7[54], stage1_7[55]},
      {stage2_9[8],stage2_8[38],stage2_7[38],stage2_6[41],stage2_5[66]}
   );
   gpc606_5 gpc4831 (
      {stage1_5[58], stage1_5[59], stage1_5[60], stage1_5[61], stage1_5[62], stage1_5[63]},
      {stage1_7[56], stage1_7[57], stage1_7[58], stage1_7[59], stage1_7[60], stage1_7[61]},
      {stage2_9[9],stage2_8[39],stage2_7[39],stage2_6[42],stage2_5[67]}
   );
   gpc606_5 gpc4832 (
      {stage1_5[64], stage1_5[65], stage1_5[66], stage1_5[67], stage1_5[68], stage1_5[69]},
      {stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65], stage1_7[66], stage1_7[67]},
      {stage2_9[10],stage2_8[40],stage2_7[40],stage2_6[43],stage2_5[68]}
   );
   gpc606_5 gpc4833 (
      {stage1_5[70], stage1_5[71], stage1_5[72], stage1_5[73], stage1_5[74], stage1_5[75]},
      {stage1_7[68], stage1_7[69], stage1_7[70], stage1_7[71], stage1_7[72], stage1_7[73]},
      {stage2_9[11],stage2_8[41],stage2_7[41],stage2_6[44],stage2_5[69]}
   );
   gpc606_5 gpc4834 (
      {stage1_5[76], stage1_5[77], stage1_5[78], stage1_5[79], stage1_5[80], stage1_5[81]},
      {stage1_7[74], stage1_7[75], stage1_7[76], stage1_7[77], stage1_7[78], stage1_7[79]},
      {stage2_9[12],stage2_8[42],stage2_7[42],stage2_6[45],stage2_5[70]}
   );
   gpc606_5 gpc4835 (
      {stage1_5[82], stage1_5[83], stage1_5[84], stage1_5[85], stage1_5[86], stage1_5[87]},
      {stage1_7[80], stage1_7[81], stage1_7[82], stage1_7[83], stage1_7[84], stage1_7[85]},
      {stage2_9[13],stage2_8[43],stage2_7[43],stage2_6[46],stage2_5[71]}
   );
   gpc606_5 gpc4836 (
      {stage1_5[88], stage1_5[89], stage1_5[90], stage1_5[91], stage1_5[92], stage1_5[93]},
      {stage1_7[86], stage1_7[87], stage1_7[88], stage1_7[89], stage1_7[90], stage1_7[91]},
      {stage2_9[14],stage2_8[44],stage2_7[44],stage2_6[47],stage2_5[72]}
   );
   gpc606_5 gpc4837 (
      {stage1_5[94], stage1_5[95], stage1_5[96], stage1_5[97], stage1_5[98], stage1_5[99]},
      {stage1_7[92], stage1_7[93], stage1_7[94], stage1_7[95], stage1_7[96], stage1_7[97]},
      {stage2_9[15],stage2_8[45],stage2_7[45],stage2_6[48],stage2_5[73]}
   );
   gpc606_5 gpc4838 (
      {stage1_5[100], stage1_5[101], stage1_5[102], stage1_5[103], stage1_5[104], stage1_5[105]},
      {stage1_7[98], stage1_7[99], stage1_7[100], stage1_7[101], stage1_7[102], stage1_7[103]},
      {stage2_9[16],stage2_8[46],stage2_7[46],stage2_6[49],stage2_5[74]}
   );
   gpc606_5 gpc4839 (
      {stage1_5[106], stage1_5[107], stage1_5[108], stage1_5[109], stage1_5[110], stage1_5[111]},
      {stage1_7[104], stage1_7[105], stage1_7[106], stage1_7[107], stage1_7[108], stage1_7[109]},
      {stage2_9[17],stage2_8[47],stage2_7[47],stage2_6[50],stage2_5[75]}
   );
   gpc606_5 gpc4840 (
      {stage1_5[112], stage1_5[113], stage1_5[114], stage1_5[115], stage1_5[116], stage1_5[117]},
      {stage1_7[110], stage1_7[111], stage1_7[112], stage1_7[113], stage1_7[114], stage1_7[115]},
      {stage2_9[18],stage2_8[48],stage2_7[48],stage2_6[51],stage2_5[76]}
   );
   gpc606_5 gpc4841 (
      {stage1_5[118], stage1_5[119], stage1_5[120], stage1_5[121], stage1_5[122], stage1_5[123]},
      {stage1_7[116], stage1_7[117], stage1_7[118], stage1_7[119], stage1_7[120], stage1_7[121]},
      {stage2_9[19],stage2_8[49],stage2_7[49],stage2_6[52],stage2_5[77]}
   );
   gpc615_5 gpc4842 (
      {stage1_7[122], stage1_7[123], stage1_7[124], stage1_7[125], stage1_7[126]},
      {stage1_8[0]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[0],stage2_9[20],stage2_8[50],stage2_7[50]}
   );
   gpc615_5 gpc4843 (
      {stage1_7[127], stage1_7[128], stage1_7[129], stage1_7[130], stage1_7[131]},
      {stage1_8[1]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[1],stage2_9[21],stage2_8[51],stage2_7[51]}
   );
   gpc615_5 gpc4844 (
      {stage1_7[132], stage1_7[133], stage1_7[134], stage1_7[135], stage1_7[136]},
      {stage1_8[2]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[2],stage2_9[22],stage2_8[52],stage2_7[52]}
   );
   gpc615_5 gpc4845 (
      {stage1_7[137], stage1_7[138], stage1_7[139], stage1_7[140], stage1_7[141]},
      {stage1_8[3]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[3],stage2_9[23],stage2_8[53],stage2_7[53]}
   );
   gpc615_5 gpc4846 (
      {stage1_7[142], stage1_7[143], stage1_7[144], stage1_7[145], stage1_7[146]},
      {stage1_8[4]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[4],stage2_9[24],stage2_8[54],stage2_7[54]}
   );
   gpc615_5 gpc4847 (
      {stage1_7[147], stage1_7[148], stage1_7[149], stage1_7[150], stage1_7[151]},
      {stage1_8[5]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[5],stage2_9[25],stage2_8[55],stage2_7[55]}
   );
   gpc615_5 gpc4848 (
      {stage1_7[152], stage1_7[153], stage1_7[154], stage1_7[155], stage1_7[156]},
      {stage1_8[6]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[6],stage2_9[26],stage2_8[56],stage2_7[56]}
   );
   gpc615_5 gpc4849 (
      {stage1_7[157], stage1_7[158], stage1_7[159], stage1_7[160], stage1_7[161]},
      {stage1_8[7]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[7],stage2_9[27],stage2_8[57],stage2_7[57]}
   );
   gpc615_5 gpc4850 (
      {stage1_7[162], stage1_7[163], stage1_7[164], stage1_7[165], stage1_7[166]},
      {stage1_8[8]},
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage2_11[8],stage2_10[8],stage2_9[28],stage2_8[58],stage2_7[58]}
   );
   gpc615_5 gpc4851 (
      {stage1_7[167], stage1_7[168], stage1_7[169], stage1_7[170], stage1_7[171]},
      {stage1_8[9]},
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage2_11[9],stage2_10[9],stage2_9[29],stage2_8[59],stage2_7[59]}
   );
   gpc615_5 gpc4852 (
      {stage1_7[172], stage1_7[173], stage1_7[174], stage1_7[175], stage1_7[176]},
      {stage1_8[10]},
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage2_11[10],stage2_10[10],stage2_9[30],stage2_8[60],stage2_7[60]}
   );
   gpc615_5 gpc4853 (
      {stage1_7[177], stage1_7[178], stage1_7[179], stage1_7[180], stage1_7[181]},
      {stage1_8[11]},
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage2_11[11],stage2_10[11],stage2_9[31],stage2_8[61],stage2_7[61]}
   );
   gpc615_5 gpc4854 (
      {stage1_7[182], stage1_7[183], stage1_7[184], stage1_7[185], stage1_7[186]},
      {stage1_8[12]},
      {stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77]},
      {stage2_11[12],stage2_10[12],stage2_9[32],stage2_8[62],stage2_7[62]}
   );
   gpc615_5 gpc4855 (
      {stage1_7[187], stage1_7[188], stage1_7[189], stage1_7[190], stage1_7[191]},
      {stage1_8[13]},
      {stage1_9[78], stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83]},
      {stage2_11[13],stage2_10[13],stage2_9[33],stage2_8[63],stage2_7[63]}
   );
   gpc615_5 gpc4856 (
      {stage1_7[192], stage1_7[193], stage1_7[194], stage1_7[195], stage1_7[196]},
      {stage1_8[14]},
      {stage1_9[84], stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89]},
      {stage2_11[14],stage2_10[14],stage2_9[34],stage2_8[64],stage2_7[64]}
   );
   gpc615_5 gpc4857 (
      {stage1_7[197], stage1_7[198], stage1_7[199], stage1_7[200], stage1_7[201]},
      {stage1_8[15]},
      {stage1_9[90], stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95]},
      {stage2_11[15],stage2_10[15],stage2_9[35],stage2_8[65],stage2_7[65]}
   );
   gpc615_5 gpc4858 (
      {stage1_7[202], stage1_7[203], stage1_7[204], stage1_7[205], stage1_7[206]},
      {stage1_8[16]},
      {stage1_9[96], stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100], stage1_9[101]},
      {stage2_11[16],stage2_10[16],stage2_9[36],stage2_8[66],stage2_7[66]}
   );
   gpc615_5 gpc4859 (
      {stage1_7[207], stage1_7[208], stage1_7[209], stage1_7[210], stage1_7[211]},
      {stage1_8[17]},
      {stage1_9[102], stage1_9[103], stage1_9[104], stage1_9[105], stage1_9[106], stage1_9[107]},
      {stage2_11[17],stage2_10[17],stage2_9[37],stage2_8[67],stage2_7[67]}
   );
   gpc615_5 gpc4860 (
      {stage1_7[212], stage1_7[213], stage1_7[214], stage1_7[215], stage1_7[216]},
      {stage1_8[18]},
      {stage1_9[108], stage1_9[109], stage1_9[110], stage1_9[111], stage1_9[112], stage1_9[113]},
      {stage2_11[18],stage2_10[18],stage2_9[38],stage2_8[68],stage2_7[68]}
   );
   gpc207_4 gpc4861 (
      {stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23], stage1_8[24], stage1_8[25]},
      {stage1_10[0], stage1_10[1]},
      {stage2_11[19],stage2_10[19],stage2_9[39],stage2_8[69]}
   );
   gpc606_5 gpc4862 (
      {stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29], stage1_8[30], stage1_8[31]},
      {stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5], stage1_10[6], stage1_10[7]},
      {stage2_12[0],stage2_11[20],stage2_10[20],stage2_9[40],stage2_8[70]}
   );
   gpc606_5 gpc4863 (
      {stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35], stage1_8[36], stage1_8[37]},
      {stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11], stage1_10[12], stage1_10[13]},
      {stage2_12[1],stage2_11[21],stage2_10[21],stage2_9[41],stage2_8[71]}
   );
   gpc606_5 gpc4864 (
      {stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41], stage1_8[42], stage1_8[43]},
      {stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17], stage1_10[18], stage1_10[19]},
      {stage2_12[2],stage2_11[22],stage2_10[22],stage2_9[42],stage2_8[72]}
   );
   gpc606_5 gpc4865 (
      {stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47], stage1_8[48], stage1_8[49]},
      {stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23], stage1_10[24], stage1_10[25]},
      {stage2_12[3],stage2_11[23],stage2_10[23],stage2_9[43],stage2_8[73]}
   );
   gpc606_5 gpc4866 (
      {stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53], stage1_8[54], stage1_8[55]},
      {stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29], stage1_10[30], stage1_10[31]},
      {stage2_12[4],stage2_11[24],stage2_10[24],stage2_9[44],stage2_8[74]}
   );
   gpc606_5 gpc4867 (
      {stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59], stage1_8[60], stage1_8[61]},
      {stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35], stage1_10[36], stage1_10[37]},
      {stage2_12[5],stage2_11[25],stage2_10[25],stage2_9[45],stage2_8[75]}
   );
   gpc606_5 gpc4868 (
      {stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65], stage1_8[66], stage1_8[67]},
      {stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41], stage1_10[42], stage1_10[43]},
      {stage2_12[6],stage2_11[26],stage2_10[26],stage2_9[46],stage2_8[76]}
   );
   gpc606_5 gpc4869 (
      {stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71], stage1_8[72], stage1_8[73]},
      {stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47], stage1_10[48], stage1_10[49]},
      {stage2_12[7],stage2_11[27],stage2_10[27],stage2_9[47],stage2_8[77]}
   );
   gpc606_5 gpc4870 (
      {stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77], stage1_8[78], stage1_8[79]},
      {stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53], stage1_10[54], stage1_10[55]},
      {stage2_12[8],stage2_11[28],stage2_10[28],stage2_9[48],stage2_8[78]}
   );
   gpc606_5 gpc4871 (
      {stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83], stage1_8[84], stage1_8[85]},
      {stage1_10[56], stage1_10[57], stage1_10[58], stage1_10[59], stage1_10[60], stage1_10[61]},
      {stage2_12[9],stage2_11[29],stage2_10[29],stage2_9[49],stage2_8[79]}
   );
   gpc606_5 gpc4872 (
      {stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89], stage1_8[90], stage1_8[91]},
      {stage1_10[62], stage1_10[63], stage1_10[64], stage1_10[65], stage1_10[66], stage1_10[67]},
      {stage2_12[10],stage2_11[30],stage2_10[30],stage2_9[50],stage2_8[80]}
   );
   gpc606_5 gpc4873 (
      {stage1_8[92], stage1_8[93], stage1_8[94], stage1_8[95], stage1_8[96], stage1_8[97]},
      {stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71], stage1_10[72], stage1_10[73]},
      {stage2_12[11],stage2_11[31],stage2_10[31],stage2_9[51],stage2_8[81]}
   );
   gpc606_5 gpc4874 (
      {stage1_8[98], stage1_8[99], stage1_8[100], stage1_8[101], stage1_8[102], stage1_8[103]},
      {stage1_10[74], stage1_10[75], stage1_10[76], stage1_10[77], stage1_10[78], stage1_10[79]},
      {stage2_12[12],stage2_11[32],stage2_10[32],stage2_9[52],stage2_8[82]}
   );
   gpc606_5 gpc4875 (
      {stage1_8[104], stage1_8[105], stage1_8[106], stage1_8[107], stage1_8[108], stage1_8[109]},
      {stage1_10[80], stage1_10[81], stage1_10[82], stage1_10[83], stage1_10[84], stage1_10[85]},
      {stage2_12[13],stage2_11[33],stage2_10[33],stage2_9[53],stage2_8[83]}
   );
   gpc606_5 gpc4876 (
      {stage1_8[110], stage1_8[111], stage1_8[112], stage1_8[113], stage1_8[114], stage1_8[115]},
      {stage1_10[86], stage1_10[87], stage1_10[88], stage1_10[89], stage1_10[90], stage1_10[91]},
      {stage2_12[14],stage2_11[34],stage2_10[34],stage2_9[54],stage2_8[84]}
   );
   gpc606_5 gpc4877 (
      {stage1_8[116], stage1_8[117], stage1_8[118], stage1_8[119], stage1_8[120], stage1_8[121]},
      {stage1_10[92], stage1_10[93], stage1_10[94], stage1_10[95], stage1_10[96], stage1_10[97]},
      {stage2_12[15],stage2_11[35],stage2_10[35],stage2_9[55],stage2_8[85]}
   );
   gpc606_5 gpc4878 (
      {stage1_8[122], stage1_8[123], stage1_8[124], stage1_8[125], stage1_8[126], stage1_8[127]},
      {stage1_10[98], stage1_10[99], stage1_10[100], stage1_10[101], stage1_10[102], stage1_10[103]},
      {stage2_12[16],stage2_11[36],stage2_10[36],stage2_9[56],stage2_8[86]}
   );
   gpc606_5 gpc4879 (
      {stage1_8[128], stage1_8[129], stage1_8[130], stage1_8[131], stage1_8[132], stage1_8[133]},
      {stage1_10[104], stage1_10[105], stage1_10[106], stage1_10[107], stage1_10[108], stage1_10[109]},
      {stage2_12[17],stage2_11[37],stage2_10[37],stage2_9[57],stage2_8[87]}
   );
   gpc606_5 gpc4880 (
      {stage1_9[114], stage1_9[115], stage1_9[116], stage1_9[117], stage1_9[118], stage1_9[119]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[18],stage2_11[38],stage2_10[38],stage2_9[58]}
   );
   gpc606_5 gpc4881 (
      {stage1_9[120], stage1_9[121], stage1_9[122], stage1_9[123], stage1_9[124], stage1_9[125]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[19],stage2_11[39],stage2_10[39],stage2_9[59]}
   );
   gpc606_5 gpc4882 (
      {stage1_9[126], stage1_9[127], stage1_9[128], stage1_9[129], stage1_9[130], stage1_9[131]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[20],stage2_11[40],stage2_10[40],stage2_9[60]}
   );
   gpc615_5 gpc4883 (
      {stage1_10[110], stage1_10[111], stage1_10[112], stage1_10[113], stage1_10[114]},
      {stage1_11[18]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[3],stage2_12[21],stage2_11[41],stage2_10[41]}
   );
   gpc615_5 gpc4884 (
      {stage1_10[115], stage1_10[116], stage1_10[117], stage1_10[118], stage1_10[119]},
      {stage1_11[19]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[4],stage2_12[22],stage2_11[42],stage2_10[42]}
   );
   gpc615_5 gpc4885 (
      {stage1_10[120], stage1_10[121], stage1_10[122], stage1_10[123], stage1_10[124]},
      {stage1_11[20]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[5],stage2_12[23],stage2_11[43],stage2_10[43]}
   );
   gpc615_5 gpc4886 (
      {stage1_10[125], stage1_10[126], stage1_10[127], stage1_10[128], stage1_10[129]},
      {stage1_11[21]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[6],stage2_12[24],stage2_11[44],stage2_10[44]}
   );
   gpc615_5 gpc4887 (
      {stage1_10[130], stage1_10[131], stage1_10[132], stage1_10[133], stage1_10[134]},
      {stage1_11[22]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[7],stage2_12[25],stage2_11[45],stage2_10[45]}
   );
   gpc615_5 gpc4888 (
      {stage1_10[135], stage1_10[136], stage1_10[137], stage1_10[138], stage1_10[139]},
      {stage1_11[23]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[8],stage2_12[26],stage2_11[46],stage2_10[46]}
   );
   gpc615_5 gpc4889 (
      {stage1_10[140], stage1_10[141], stage1_10[142], stage1_10[143], stage1_10[144]},
      {stage1_11[24]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[9],stage2_12[27],stage2_11[47],stage2_10[47]}
   );
   gpc615_5 gpc4890 (
      {stage1_10[145], stage1_10[146], stage1_10[147], stage1_10[148], stage1_10[149]},
      {stage1_11[25]},
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage2_14[7],stage2_13[10],stage2_12[28],stage2_11[48],stage2_10[48]}
   );
   gpc615_5 gpc4891 (
      {stage1_10[150], stage1_10[151], stage1_10[152], stage1_10[153], stage1_10[154]},
      {stage1_11[26]},
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage2_14[8],stage2_13[11],stage2_12[29],stage2_11[49],stage2_10[49]}
   );
   gpc615_5 gpc4892 (
      {stage1_10[155], stage1_10[156], stage1_10[157], stage1_10[158], stage1_10[159]},
      {stage1_11[27]},
      {stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage2_14[9],stage2_13[12],stage2_12[30],stage2_11[50],stage2_10[50]}
   );
   gpc615_5 gpc4893 (
      {stage1_10[160], stage1_10[161], stage1_10[162], stage1_10[163], stage1_10[164]},
      {stage1_11[28]},
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64], stage1_12[65]},
      {stage2_14[10],stage2_13[13],stage2_12[31],stage2_11[51],stage2_10[51]}
   );
   gpc615_5 gpc4894 (
      {stage1_10[165], stage1_10[166], stage1_10[167], stage1_10[168], stage1_10[169]},
      {stage1_11[29]},
      {stage1_12[66], stage1_12[67], stage1_12[68], stage1_12[69], stage1_12[70], stage1_12[71]},
      {stage2_14[11],stage2_13[14],stage2_12[32],stage2_11[52],stage2_10[52]}
   );
   gpc615_5 gpc4895 (
      {stage1_10[170], stage1_10[171], stage1_10[172], stage1_10[173], stage1_10[174]},
      {stage1_11[30]},
      {stage1_12[72], stage1_12[73], stage1_12[74], stage1_12[75], stage1_12[76], stage1_12[77]},
      {stage2_14[12],stage2_13[15],stage2_12[33],stage2_11[53],stage2_10[53]}
   );
   gpc606_5 gpc4896 (
      {stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35], stage1_11[36]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[13],stage2_13[16],stage2_12[34],stage2_11[54]}
   );
   gpc606_5 gpc4897 (
      {stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41], stage1_11[42]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[14],stage2_13[17],stage2_12[35],stage2_11[55]}
   );
   gpc606_5 gpc4898 (
      {stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47], stage1_11[48]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[15],stage2_13[18],stage2_12[36],stage2_11[56]}
   );
   gpc606_5 gpc4899 (
      {stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53], stage1_11[54]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[16],stage2_13[19],stage2_12[37],stage2_11[57]}
   );
   gpc606_5 gpc4900 (
      {stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58], stage1_11[59], stage1_11[60]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[17],stage2_13[20],stage2_12[38],stage2_11[58]}
   );
   gpc606_5 gpc4901 (
      {stage1_11[61], stage1_11[62], stage1_11[63], stage1_11[64], stage1_11[65], stage1_11[66]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[18],stage2_13[21],stage2_12[39],stage2_11[59]}
   );
   gpc606_5 gpc4902 (
      {stage1_11[67], stage1_11[68], stage1_11[69], stage1_11[70], stage1_11[71], stage1_11[72]},
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage2_15[6],stage2_14[19],stage2_13[22],stage2_12[40],stage2_11[60]}
   );
   gpc606_5 gpc4903 (
      {stage1_11[73], stage1_11[74], stage1_11[75], stage1_11[76], stage1_11[77], stage1_11[78]},
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage2_15[7],stage2_14[20],stage2_13[23],stage2_12[41],stage2_11[61]}
   );
   gpc606_5 gpc4904 (
      {stage1_11[79], stage1_11[80], stage1_11[81], stage1_11[82], stage1_11[83], stage1_11[84]},
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage2_15[8],stage2_14[21],stage2_13[24],stage2_12[42],stage2_11[62]}
   );
   gpc606_5 gpc4905 (
      {stage1_11[85], stage1_11[86], stage1_11[87], stage1_11[88], stage1_11[89], stage1_11[90]},
      {stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59]},
      {stage2_15[9],stage2_14[22],stage2_13[25],stage2_12[43],stage2_11[63]}
   );
   gpc606_5 gpc4906 (
      {stage1_11[91], stage1_11[92], stage1_11[93], stage1_11[94], stage1_11[95], stage1_11[96]},
      {stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage2_15[10],stage2_14[23],stage2_13[26],stage2_12[44],stage2_11[64]}
   );
   gpc606_5 gpc4907 (
      {stage1_11[97], stage1_11[98], stage1_11[99], stage1_11[100], stage1_11[101], stage1_11[102]},
      {stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69], stage1_13[70], stage1_13[71]},
      {stage2_15[11],stage2_14[24],stage2_13[27],stage2_12[45],stage2_11[65]}
   );
   gpc606_5 gpc4908 (
      {stage1_11[103], stage1_11[104], stage1_11[105], stage1_11[106], stage1_11[107], stage1_11[108]},
      {stage1_13[72], stage1_13[73], stage1_13[74], stage1_13[75], stage1_13[76], stage1_13[77]},
      {stage2_15[12],stage2_14[25],stage2_13[28],stage2_12[46],stage2_11[66]}
   );
   gpc606_5 gpc4909 (
      {stage1_11[109], stage1_11[110], stage1_11[111], stage1_11[112], stage1_11[113], stage1_11[114]},
      {stage1_13[78], stage1_13[79], stage1_13[80], stage1_13[81], stage1_13[82], stage1_13[83]},
      {stage2_15[13],stage2_14[26],stage2_13[29],stage2_12[47],stage2_11[67]}
   );
   gpc606_5 gpc4910 (
      {stage1_11[115], stage1_11[116], stage1_11[117], stage1_11[118], stage1_11[119], stage1_11[120]},
      {stage1_13[84], stage1_13[85], stage1_13[86], stage1_13[87], stage1_13[88], stage1_13[89]},
      {stage2_15[14],stage2_14[27],stage2_13[30],stage2_12[48],stage2_11[68]}
   );
   gpc606_5 gpc4911 (
      {stage1_11[121], stage1_11[122], stage1_11[123], stage1_11[124], stage1_11[125], stage1_11[126]},
      {stage1_13[90], stage1_13[91], stage1_13[92], stage1_13[93], stage1_13[94], stage1_13[95]},
      {stage2_15[15],stage2_14[28],stage2_13[31],stage2_12[49],stage2_11[69]}
   );
   gpc606_5 gpc4912 (
      {stage1_11[127], stage1_11[128], stage1_11[129], stage1_11[130], stage1_11[131], stage1_11[132]},
      {stage1_13[96], stage1_13[97], stage1_13[98], stage1_13[99], stage1_13[100], stage1_13[101]},
      {stage2_15[16],stage2_14[29],stage2_13[32],stage2_12[50],stage2_11[70]}
   );
   gpc615_5 gpc4913 (
      {stage1_11[133], stage1_11[134], stage1_11[135], stage1_11[136], stage1_11[137]},
      {stage1_12[78]},
      {stage1_13[102], stage1_13[103], stage1_13[104], stage1_13[105], stage1_13[106], stage1_13[107]},
      {stage2_15[17],stage2_14[30],stage2_13[33],stage2_12[51],stage2_11[71]}
   );
   gpc615_5 gpc4914 (
      {stage1_11[138], stage1_11[139], stage1_11[140], stage1_11[141], stage1_11[142]},
      {stage1_12[79]},
      {stage1_13[108], stage1_13[109], stage1_13[110], stage1_13[111], stage1_13[112], stage1_13[113]},
      {stage2_15[18],stage2_14[31],stage2_13[34],stage2_12[52],stage2_11[72]}
   );
   gpc615_5 gpc4915 (
      {stage1_11[143], stage1_11[144], stage1_11[145], stage1_11[146], stage1_11[147]},
      {stage1_12[80]},
      {stage1_13[114], stage1_13[115], stage1_13[116], stage1_13[117], stage1_13[118], stage1_13[119]},
      {stage2_15[19],stage2_14[32],stage2_13[35],stage2_12[53],stage2_11[73]}
   );
   gpc615_5 gpc4916 (
      {stage1_11[148], stage1_11[149], stage1_11[150], stage1_11[151], stage1_11[152]},
      {stage1_12[81]},
      {stage1_13[120], stage1_13[121], stage1_13[122], stage1_13[123], stage1_13[124], stage1_13[125]},
      {stage2_15[20],stage2_14[33],stage2_13[36],stage2_12[54],stage2_11[74]}
   );
   gpc615_5 gpc4917 (
      {stage1_11[153], stage1_11[154], stage1_11[155], stage1_11[156], stage1_11[157]},
      {stage1_12[82]},
      {stage1_13[126], stage1_13[127], stage1_13[128], stage1_13[129], stage1_13[130], stage1_13[131]},
      {stage2_15[21],stage2_14[34],stage2_13[37],stage2_12[55],stage2_11[75]}
   );
   gpc615_5 gpc4918 (
      {stage1_11[158], stage1_11[159], stage1_11[160], stage1_11[161], stage1_11[162]},
      {stage1_12[83]},
      {stage1_13[132], stage1_13[133], stage1_13[134], stage1_13[135], stage1_13[136], stage1_13[137]},
      {stage2_15[22],stage2_14[35],stage2_13[38],stage2_12[56],stage2_11[76]}
   );
   gpc615_5 gpc4919 (
      {stage1_11[163], stage1_11[164], stage1_11[165], stage1_11[166], stage1_11[167]},
      {stage1_12[84]},
      {stage1_13[138], stage1_13[139], stage1_13[140], stage1_13[141], stage1_13[142], stage1_13[143]},
      {stage2_15[23],stage2_14[36],stage2_13[39],stage2_12[57],stage2_11[77]}
   );
   gpc615_5 gpc4920 (
      {stage1_11[168], stage1_11[169], stage1_11[170], stage1_11[171], stage1_11[172]},
      {stage1_12[85]},
      {stage1_13[144], stage1_13[145], stage1_13[146], stage1_13[147], stage1_13[148], stage1_13[149]},
      {stage2_15[24],stage2_14[37],stage2_13[40],stage2_12[58],stage2_11[78]}
   );
   gpc615_5 gpc4921 (
      {stage1_11[173], stage1_11[174], stage1_11[175], stage1_11[176], stage1_11[177]},
      {stage1_12[86]},
      {stage1_13[150], stage1_13[151], stage1_13[152], stage1_13[153], stage1_13[154], stage1_13[155]},
      {stage2_15[25],stage2_14[38],stage2_13[41],stage2_12[59],stage2_11[79]}
   );
   gpc615_5 gpc4922 (
      {stage1_11[178], stage1_11[179], stage1_11[180], stage1_11[181], stage1_11[182]},
      {stage1_12[87]},
      {stage1_13[156], stage1_13[157], stage1_13[158], stage1_13[159], stage1_13[160], stage1_13[161]},
      {stage2_15[26],stage2_14[39],stage2_13[42],stage2_12[60],stage2_11[80]}
   );
   gpc615_5 gpc4923 (
      {stage1_11[183], stage1_11[184], stage1_11[185], stage1_11[186], stage1_11[187]},
      {stage1_12[88]},
      {stage1_13[162], stage1_13[163], stage1_13[164], stage1_13[165], stage1_13[166], stage1_13[167]},
      {stage2_15[27],stage2_14[40],stage2_13[43],stage2_12[61],stage2_11[81]}
   );
   gpc615_5 gpc4924 (
      {stage1_11[188], stage1_11[189], stage1_11[190], stage1_11[191], stage1_11[192]},
      {stage1_12[89]},
      {stage1_13[168], stage1_13[169], stage1_13[170], stage1_13[171], stage1_13[172], stage1_13[173]},
      {stage2_15[28],stage2_14[41],stage2_13[44],stage2_12[62],stage2_11[82]}
   );
   gpc615_5 gpc4925 (
      {stage1_11[193], stage1_11[194], stage1_11[195], stage1_11[196], stage1_11[197]},
      {stage1_12[90]},
      {stage1_13[174], stage1_13[175], stage1_13[176], stage1_13[177], stage1_13[178], stage1_13[179]},
      {stage2_15[29],stage2_14[42],stage2_13[45],stage2_12[63],stage2_11[83]}
   );
   gpc615_5 gpc4926 (
      {stage1_11[198], stage1_11[199], stage1_11[200], stage1_11[201], stage1_11[202]},
      {stage1_12[91]},
      {stage1_13[180], stage1_13[181], stage1_13[182], stage1_13[183], stage1_13[184], stage1_13[185]},
      {stage2_15[30],stage2_14[43],stage2_13[46],stage2_12[64],stage2_11[84]}
   );
   gpc615_5 gpc4927 (
      {stage1_11[203], stage1_11[204], stage1_11[205], stage1_11[206], stage1_11[207]},
      {stage1_12[92]},
      {stage1_13[186], stage1_13[187], stage1_13[188], stage1_13[189], stage1_13[190], stage1_13[191]},
      {stage2_15[31],stage2_14[44],stage2_13[47],stage2_12[65],stage2_11[85]}
   );
   gpc615_5 gpc4928 (
      {stage1_11[208], stage1_11[209], stage1_11[210], stage1_11[211], stage1_11[212]},
      {stage1_12[93]},
      {stage1_13[192], stage1_13[193], stage1_13[194], stage1_13[195], stage1_13[196], stage1_13[197]},
      {stage2_15[32],stage2_14[45],stage2_13[48],stage2_12[66],stage2_11[86]}
   );
   gpc615_5 gpc4929 (
      {stage1_11[213], stage1_11[214], stage1_11[215], stage1_11[216], stage1_11[217]},
      {stage1_12[94]},
      {stage1_13[198], stage1_13[199], stage1_13[200], stage1_13[201], stage1_13[202], stage1_13[203]},
      {stage2_15[33],stage2_14[46],stage2_13[49],stage2_12[67],stage2_11[87]}
   );
   gpc615_5 gpc4930 (
      {stage1_11[218], stage1_11[219], stage1_11[220], stage1_11[221], stage1_11[222]},
      {stage1_12[95]},
      {stage1_13[204], stage1_13[205], stage1_13[206], stage1_13[207], stage1_13[208], stage1_13[209]},
      {stage2_15[34],stage2_14[47],stage2_13[50],stage2_12[68],stage2_11[88]}
   );
   gpc1325_5 gpc4931 (
      {stage1_11[223], stage1_11[224], stage1_11[225], stage1_11[226], stage1_11[227]},
      {stage1_12[96], stage1_12[97]},
      {stage1_13[210], stage1_13[211], stage1_13[212]},
      {stage1_14[0]},
      {stage2_15[35],stage2_14[48],stage2_13[51],stage2_12[69],stage2_11[89]}
   );
   gpc2135_5 gpc4932 (
      {stage1_12[98], stage1_12[99], stage1_12[100], stage1_12[101], stage1_12[102]},
      {stage1_13[213], stage1_13[214], stage1_13[215]},
      {stage1_14[1]},
      {stage1_15[0], stage1_15[1]},
      {stage2_16[0],stage2_15[36],stage2_14[49],stage2_13[52],stage2_12[70]}
   );
   gpc606_5 gpc4933 (
      {stage1_12[103], stage1_12[104], stage1_12[105], stage1_12[106], stage1_12[107], stage1_12[108]},
      {stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5], stage1_14[6], stage1_14[7]},
      {stage2_16[1],stage2_15[37],stage2_14[50],stage2_13[53],stage2_12[71]}
   );
   gpc606_5 gpc4934 (
      {stage1_12[109], stage1_12[110], stage1_12[111], stage1_12[112], stage1_12[113], stage1_12[114]},
      {stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11], stage1_14[12], stage1_14[13]},
      {stage2_16[2],stage2_15[38],stage2_14[51],stage2_13[54],stage2_12[72]}
   );
   gpc606_5 gpc4935 (
      {stage1_12[115], stage1_12[116], stage1_12[117], stage1_12[118], stage1_12[119], stage1_12[120]},
      {stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17], stage1_14[18], stage1_14[19]},
      {stage2_16[3],stage2_15[39],stage2_14[52],stage2_13[55],stage2_12[73]}
   );
   gpc606_5 gpc4936 (
      {stage1_12[121], stage1_12[122], stage1_12[123], stage1_12[124], stage1_12[125], stage1_12[126]},
      {stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23], stage1_14[24], stage1_14[25]},
      {stage2_16[4],stage2_15[40],stage2_14[53],stage2_13[56],stage2_12[74]}
   );
   gpc606_5 gpc4937 (
      {stage1_12[127], stage1_12[128], stage1_12[129], stage1_12[130], stage1_12[131], stage1_12[132]},
      {stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29], stage1_14[30], stage1_14[31]},
      {stage2_16[5],stage2_15[41],stage2_14[54],stage2_13[57],stage2_12[75]}
   );
   gpc606_5 gpc4938 (
      {stage1_12[133], stage1_12[134], stage1_12[135], stage1_12[136], stage1_12[137], stage1_12[138]},
      {stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35], stage1_14[36], stage1_14[37]},
      {stage2_16[6],stage2_15[42],stage2_14[55],stage2_13[58],stage2_12[76]}
   );
   gpc606_5 gpc4939 (
      {stage1_12[139], stage1_12[140], stage1_12[141], stage1_12[142], stage1_12[143], stage1_12[144]},
      {stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41], stage1_14[42], stage1_14[43]},
      {stage2_16[7],stage2_15[43],stage2_14[56],stage2_13[59],stage2_12[77]}
   );
   gpc606_5 gpc4940 (
      {stage1_12[145], stage1_12[146], stage1_12[147], stage1_12[148], stage1_12[149], stage1_12[150]},
      {stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47], stage1_14[48], stage1_14[49]},
      {stage2_16[8],stage2_15[44],stage2_14[57],stage2_13[60],stage2_12[78]}
   );
   gpc606_5 gpc4941 (
      {stage1_12[151], stage1_12[152], stage1_12[153], stage1_12[154], stage1_12[155], stage1_12[156]},
      {stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53], stage1_14[54], stage1_14[55]},
      {stage2_16[9],stage2_15[45],stage2_14[58],stage2_13[61],stage2_12[79]}
   );
   gpc606_5 gpc4942 (
      {stage1_12[157], stage1_12[158], stage1_12[159], stage1_12[160], stage1_12[161], stage1_12[162]},
      {stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59], stage1_14[60], stage1_14[61]},
      {stage2_16[10],stage2_15[46],stage2_14[59],stage2_13[62],stage2_12[80]}
   );
   gpc606_5 gpc4943 (
      {stage1_13[216], stage1_13[217], stage1_13[218], stage1_13[219], stage1_13[220], stage1_13[221]},
      {stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5], stage1_15[6], stage1_15[7]},
      {stage2_17[0],stage2_16[11],stage2_15[47],stage2_14[60],stage2_13[63]}
   );
   gpc606_5 gpc4944 (
      {stage1_13[222], stage1_13[223], stage1_13[224], stage1_13[225], stage1_13[226], stage1_13[227]},
      {stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11], stage1_15[12], stage1_15[13]},
      {stage2_17[1],stage2_16[12],stage2_15[48],stage2_14[61],stage2_13[64]}
   );
   gpc606_5 gpc4945 (
      {stage1_13[228], stage1_13[229], stage1_13[230], stage1_13[231], stage1_13[232], stage1_13[233]},
      {stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17], stage1_15[18], stage1_15[19]},
      {stage2_17[2],stage2_16[13],stage2_15[49],stage2_14[62],stage2_13[65]}
   );
   gpc606_5 gpc4946 (
      {stage1_13[234], stage1_13[235], stage1_13[236], stage1_13[237], stage1_13[238], stage1_13[239]},
      {stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23], stage1_15[24], stage1_15[25]},
      {stage2_17[3],stage2_16[14],stage2_15[50],stage2_14[63],stage2_13[66]}
   );
   gpc606_5 gpc4947 (
      {stage1_13[240], stage1_13[241], stage1_13[242], stage1_13[243], stage1_13[244], stage1_13[245]},
      {stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29], stage1_15[30], stage1_15[31]},
      {stage2_17[4],stage2_16[15],stage2_15[51],stage2_14[64],stage2_13[67]}
   );
   gpc606_5 gpc4948 (
      {stage1_13[246], stage1_13[247], stage1_13[248], stage1_13[249], stage1_13[250], stage1_13[251]},
      {stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35], stage1_15[36], stage1_15[37]},
      {stage2_17[5],stage2_16[16],stage2_15[52],stage2_14[65],stage2_13[68]}
   );
   gpc606_5 gpc4949 (
      {stage1_13[252], stage1_13[253], stage1_13[254], stage1_13[255], stage1_13[256], stage1_13[257]},
      {stage1_15[38], stage1_15[39], stage1_15[40], stage1_15[41], stage1_15[42], stage1_15[43]},
      {stage2_17[6],stage2_16[17],stage2_15[53],stage2_14[66],stage2_13[69]}
   );
   gpc606_5 gpc4950 (
      {stage1_13[258], stage1_13[259], stage1_13[260], stage1_13[261], stage1_13[262], stage1_13[263]},
      {stage1_15[44], stage1_15[45], stage1_15[46], stage1_15[47], stage1_15[48], stage1_15[49]},
      {stage2_17[7],stage2_16[18],stage2_15[54],stage2_14[67],stage2_13[70]}
   );
   gpc606_5 gpc4951 (
      {stage1_13[264], stage1_13[265], stage1_13[266], stage1_13[267], stage1_13[268], stage1_13[269]},
      {stage1_15[50], stage1_15[51], stage1_15[52], stage1_15[53], stage1_15[54], stage1_15[55]},
      {stage2_17[8],stage2_16[19],stage2_15[55],stage2_14[68],stage2_13[71]}
   );
   gpc606_5 gpc4952 (
      {stage1_13[270], stage1_13[271], stage1_13[272], stage1_13[273], stage1_13[274], stage1_13[275]},
      {stage1_15[56], stage1_15[57], stage1_15[58], stage1_15[59], stage1_15[60], stage1_15[61]},
      {stage2_17[9],stage2_16[20],stage2_15[56],stage2_14[69],stage2_13[72]}
   );
   gpc606_5 gpc4953 (
      {stage1_13[276], stage1_13[277], stage1_13[278], stage1_13[279], stage1_13[280], stage1_13[281]},
      {stage1_15[62], stage1_15[63], stage1_15[64], stage1_15[65], stage1_15[66], stage1_15[67]},
      {stage2_17[10],stage2_16[21],stage2_15[57],stage2_14[70],stage2_13[73]}
   );
   gpc606_5 gpc4954 (
      {stage1_13[282], stage1_13[283], stage1_13[284], stage1_13[285], stage1_13[286], stage1_13[287]},
      {stage1_15[68], stage1_15[69], stage1_15[70], stage1_15[71], stage1_15[72], stage1_15[73]},
      {stage2_17[11],stage2_16[22],stage2_15[58],stage2_14[71],stage2_13[74]}
   );
   gpc606_5 gpc4955 (
      {stage1_13[288], stage1_13[289], stage1_13[290], stage1_13[291], stage1_13[292], stage1_13[293]},
      {stage1_15[74], stage1_15[75], stage1_15[76], stage1_15[77], stage1_15[78], stage1_15[79]},
      {stage2_17[12],stage2_16[23],stage2_15[59],stage2_14[72],stage2_13[75]}
   );
   gpc606_5 gpc4956 (
      {stage1_13[294], stage1_13[295], stage1_13[296], stage1_13[297], stage1_13[298], stage1_13[299]},
      {stage1_15[80], stage1_15[81], stage1_15[82], stage1_15[83], stage1_15[84], stage1_15[85]},
      {stage2_17[13],stage2_16[24],stage2_15[60],stage2_14[73],stage2_13[76]}
   );
   gpc606_5 gpc4957 (
      {stage1_13[300], stage1_13[301], stage1_13[302], stage1_13[303], stage1_13[304], 1'b0},
      {stage1_15[86], stage1_15[87], stage1_15[88], stage1_15[89], stage1_15[90], stage1_15[91]},
      {stage2_17[14],stage2_16[25],stage2_15[61],stage2_14[74],stage2_13[77]}
   );
   gpc615_5 gpc4958 (
      {stage1_14[62], stage1_14[63], stage1_14[64], stage1_14[65], stage1_14[66]},
      {stage1_15[92]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[15],stage2_16[26],stage2_15[62],stage2_14[75]}
   );
   gpc615_5 gpc4959 (
      {stage1_14[67], stage1_14[68], stage1_14[69], stage1_14[70], stage1_14[71]},
      {stage1_15[93]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[16],stage2_16[27],stage2_15[63],stage2_14[76]}
   );
   gpc615_5 gpc4960 (
      {stage1_14[72], stage1_14[73], stage1_14[74], stage1_14[75], stage1_14[76]},
      {stage1_15[94]},
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage2_18[2],stage2_17[17],stage2_16[28],stage2_15[64],stage2_14[77]}
   );
   gpc615_5 gpc4961 (
      {stage1_14[77], stage1_14[78], stage1_14[79], stage1_14[80], stage1_14[81]},
      {stage1_15[95]},
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage2_18[3],stage2_17[18],stage2_16[29],stage2_15[65],stage2_14[78]}
   );
   gpc615_5 gpc4962 (
      {stage1_14[82], stage1_14[83], stage1_14[84], stage1_14[85], stage1_14[86]},
      {stage1_15[96]},
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage2_18[4],stage2_17[19],stage2_16[30],stage2_15[66],stage2_14[79]}
   );
   gpc615_5 gpc4963 (
      {stage1_14[87], stage1_14[88], stage1_14[89], stage1_14[90], stage1_14[91]},
      {stage1_15[97]},
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage2_18[5],stage2_17[20],stage2_16[31],stage2_15[67],stage2_14[80]}
   );
   gpc615_5 gpc4964 (
      {stage1_14[92], stage1_14[93], stage1_14[94], stage1_14[95], stage1_14[96]},
      {stage1_15[98]},
      {stage1_16[36], stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41]},
      {stage2_18[6],stage2_17[21],stage2_16[32],stage2_15[68],stage2_14[81]}
   );
   gpc615_5 gpc4965 (
      {stage1_14[97], stage1_14[98], stage1_14[99], stage1_14[100], stage1_14[101]},
      {stage1_15[99]},
      {stage1_16[42], stage1_16[43], stage1_16[44], stage1_16[45], stage1_16[46], stage1_16[47]},
      {stage2_18[7],stage2_17[22],stage2_16[33],stage2_15[69],stage2_14[82]}
   );
   gpc615_5 gpc4966 (
      {stage1_14[102], stage1_14[103], stage1_14[104], stage1_14[105], stage1_14[106]},
      {stage1_15[100]},
      {stage1_16[48], stage1_16[49], stage1_16[50], stage1_16[51], stage1_16[52], stage1_16[53]},
      {stage2_18[8],stage2_17[23],stage2_16[34],stage2_15[70],stage2_14[83]}
   );
   gpc615_5 gpc4967 (
      {stage1_14[107], stage1_14[108], stage1_14[109], stage1_14[110], stage1_14[111]},
      {stage1_15[101]},
      {stage1_16[54], stage1_16[55], stage1_16[56], stage1_16[57], stage1_16[58], stage1_16[59]},
      {stage2_18[9],stage2_17[24],stage2_16[35],stage2_15[71],stage2_14[84]}
   );
   gpc615_5 gpc4968 (
      {stage1_14[112], stage1_14[113], stage1_14[114], stage1_14[115], stage1_14[116]},
      {stage1_15[102]},
      {stage1_16[60], stage1_16[61], stage1_16[62], stage1_16[63], stage1_16[64], stage1_16[65]},
      {stage2_18[10],stage2_17[25],stage2_16[36],stage2_15[72],stage2_14[85]}
   );
   gpc615_5 gpc4969 (
      {stage1_14[117], stage1_14[118], stage1_14[119], stage1_14[120], stage1_14[121]},
      {stage1_15[103]},
      {stage1_16[66], stage1_16[67], stage1_16[68], stage1_16[69], stage1_16[70], stage1_16[71]},
      {stage2_18[11],stage2_17[26],stage2_16[37],stage2_15[73],stage2_14[86]}
   );
   gpc615_5 gpc4970 (
      {stage1_14[122], stage1_14[123], stage1_14[124], stage1_14[125], stage1_14[126]},
      {stage1_15[104]},
      {stage1_16[72], stage1_16[73], stage1_16[74], stage1_16[75], stage1_16[76], stage1_16[77]},
      {stage2_18[12],stage2_17[27],stage2_16[38],stage2_15[74],stage2_14[87]}
   );
   gpc615_5 gpc4971 (
      {stage1_14[127], stage1_14[128], stage1_14[129], stage1_14[130], stage1_14[131]},
      {stage1_15[105]},
      {stage1_16[78], stage1_16[79], stage1_16[80], stage1_16[81], stage1_16[82], stage1_16[83]},
      {stage2_18[13],stage2_17[28],stage2_16[39],stage2_15[75],stage2_14[88]}
   );
   gpc615_5 gpc4972 (
      {stage1_14[132], stage1_14[133], stage1_14[134], stage1_14[135], stage1_14[136]},
      {stage1_15[106]},
      {stage1_16[84], stage1_16[85], stage1_16[86], stage1_16[87], stage1_16[88], stage1_16[89]},
      {stage2_18[14],stage2_17[29],stage2_16[40],stage2_15[76],stage2_14[89]}
   );
   gpc615_5 gpc4973 (
      {stage1_14[137], stage1_14[138], stage1_14[139], stage1_14[140], stage1_14[141]},
      {stage1_15[107]},
      {stage1_16[90], stage1_16[91], stage1_16[92], stage1_16[93], stage1_16[94], stage1_16[95]},
      {stage2_18[15],stage2_17[30],stage2_16[41],stage2_15[77],stage2_14[90]}
   );
   gpc615_5 gpc4974 (
      {stage1_14[142], stage1_14[143], stage1_14[144], stage1_14[145], stage1_14[146]},
      {stage1_15[108]},
      {stage1_16[96], stage1_16[97], stage1_16[98], stage1_16[99], stage1_16[100], stage1_16[101]},
      {stage2_18[16],stage2_17[31],stage2_16[42],stage2_15[78],stage2_14[91]}
   );
   gpc615_5 gpc4975 (
      {stage1_14[147], stage1_14[148], stage1_14[149], stage1_14[150], stage1_14[151]},
      {stage1_15[109]},
      {stage1_16[102], stage1_16[103], stage1_16[104], stage1_16[105], stage1_16[106], stage1_16[107]},
      {stage2_18[17],stage2_17[32],stage2_16[43],stage2_15[79],stage2_14[92]}
   );
   gpc615_5 gpc4976 (
      {stage1_14[152], stage1_14[153], stage1_14[154], stage1_14[155], stage1_14[156]},
      {stage1_15[110]},
      {stage1_16[108], stage1_16[109], stage1_16[110], stage1_16[111], stage1_16[112], stage1_16[113]},
      {stage2_18[18],stage2_17[33],stage2_16[44],stage2_15[80],stage2_14[93]}
   );
   gpc615_5 gpc4977 (
      {stage1_14[157], stage1_14[158], stage1_14[159], stage1_14[160], stage1_14[161]},
      {stage1_15[111]},
      {stage1_16[114], stage1_16[115], stage1_16[116], stage1_16[117], stage1_16[118], stage1_16[119]},
      {stage2_18[19],stage2_17[34],stage2_16[45],stage2_15[81],stage2_14[94]}
   );
   gpc615_5 gpc4978 (
      {stage1_14[162], stage1_14[163], stage1_14[164], stage1_14[165], stage1_14[166]},
      {stage1_15[112]},
      {stage1_16[120], stage1_16[121], stage1_16[122], stage1_16[123], stage1_16[124], stage1_16[125]},
      {stage2_18[20],stage2_17[35],stage2_16[46],stage2_15[82],stage2_14[95]}
   );
   gpc615_5 gpc4979 (
      {stage1_14[167], stage1_14[168], stage1_14[169], stage1_14[170], stage1_14[171]},
      {stage1_15[113]},
      {stage1_16[126], stage1_16[127], stage1_16[128], stage1_16[129], stage1_16[130], stage1_16[131]},
      {stage2_18[21],stage2_17[36],stage2_16[47],stage2_15[83],stage2_14[96]}
   );
   gpc615_5 gpc4980 (
      {stage1_14[172], stage1_14[173], stage1_14[174], stage1_14[175], stage1_14[176]},
      {stage1_15[114]},
      {stage1_16[132], stage1_16[133], stage1_16[134], stage1_16[135], stage1_16[136], stage1_16[137]},
      {stage2_18[22],stage2_17[37],stage2_16[48],stage2_15[84],stage2_14[97]}
   );
   gpc615_5 gpc4981 (
      {stage1_14[177], stage1_14[178], stage1_14[179], stage1_14[180], stage1_14[181]},
      {stage1_15[115]},
      {stage1_16[138], stage1_16[139], stage1_16[140], stage1_16[141], stage1_16[142], stage1_16[143]},
      {stage2_18[23],stage2_17[38],stage2_16[49],stage2_15[85],stage2_14[98]}
   );
   gpc615_5 gpc4982 (
      {stage1_14[182], stage1_14[183], stage1_14[184], stage1_14[185], stage1_14[186]},
      {stage1_15[116]},
      {stage1_16[144], stage1_16[145], stage1_16[146], stage1_16[147], stage1_16[148], stage1_16[149]},
      {stage2_18[24],stage2_17[39],stage2_16[50],stage2_15[86],stage2_14[99]}
   );
   gpc615_5 gpc4983 (
      {stage1_14[187], stage1_14[188], stage1_14[189], stage1_14[190], stage1_14[191]},
      {stage1_15[117]},
      {stage1_16[150], stage1_16[151], stage1_16[152], stage1_16[153], stage1_16[154], stage1_16[155]},
      {stage2_18[25],stage2_17[40],stage2_16[51],stage2_15[87],stage2_14[100]}
   );
   gpc615_5 gpc4984 (
      {stage1_14[192], stage1_14[193], stage1_14[194], stage1_14[195], stage1_14[196]},
      {stage1_15[118]},
      {stage1_16[156], stage1_16[157], stage1_16[158], stage1_16[159], stage1_16[160], stage1_16[161]},
      {stage2_18[26],stage2_17[41],stage2_16[52],stage2_15[88],stage2_14[101]}
   );
   gpc615_5 gpc4985 (
      {stage1_14[197], stage1_14[198], stage1_14[199], stage1_14[200], stage1_14[201]},
      {stage1_15[119]},
      {stage1_16[162], stage1_16[163], stage1_16[164], stage1_16[165], stage1_16[166], stage1_16[167]},
      {stage2_18[27],stage2_17[42],stage2_16[53],stage2_15[89],stage2_14[102]}
   );
   gpc615_5 gpc4986 (
      {stage1_14[202], stage1_14[203], stage1_14[204], stage1_14[205], stage1_14[206]},
      {stage1_15[120]},
      {stage1_16[168], stage1_16[169], stage1_16[170], stage1_16[171], stage1_16[172], stage1_16[173]},
      {stage2_18[28],stage2_17[43],stage2_16[54],stage2_15[90],stage2_14[103]}
   );
   gpc615_5 gpc4987 (
      {stage1_14[207], stage1_14[208], stage1_14[209], stage1_14[210], stage1_14[211]},
      {stage1_15[121]},
      {stage1_16[174], stage1_16[175], stage1_16[176], stage1_16[177], stage1_16[178], stage1_16[179]},
      {stage2_18[29],stage2_17[44],stage2_16[55],stage2_15[91],stage2_14[104]}
   );
   gpc615_5 gpc4988 (
      {stage1_14[212], stage1_14[213], stage1_14[214], stage1_14[215], stage1_14[216]},
      {stage1_15[122]},
      {stage1_16[180], stage1_16[181], stage1_16[182], stage1_16[183], stage1_16[184], stage1_16[185]},
      {stage2_18[30],stage2_17[45],stage2_16[56],stage2_15[92],stage2_14[105]}
   );
   gpc606_5 gpc4989 (
      {stage1_16[186], stage1_16[187], stage1_16[188], stage1_16[189], stage1_16[190], stage1_16[191]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[0],stage2_18[31],stage2_17[46],stage2_16[57]}
   );
   gpc606_5 gpc4990 (
      {stage1_16[192], stage1_16[193], stage1_16[194], stage1_16[195], stage1_16[196], stage1_16[197]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[1],stage2_18[32],stage2_17[47],stage2_16[58]}
   );
   gpc606_5 gpc4991 (
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[2],stage2_19[2],stage2_18[33],stage2_17[48]}
   );
   gpc606_5 gpc4992 (
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[3],stage2_19[3],stage2_18[34],stage2_17[49]}
   );
   gpc606_5 gpc4993 (
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17]},
      {stage2_21[2],stage2_20[4],stage2_19[4],stage2_18[35],stage2_17[50]}
   );
   gpc606_5 gpc4994 (
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage1_19[18], stage1_19[19], stage1_19[20], stage1_19[21], stage1_19[22], stage1_19[23]},
      {stage2_21[3],stage2_20[5],stage2_19[5],stage2_18[36],stage2_17[51]}
   );
   gpc606_5 gpc4995 (
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage1_19[24], stage1_19[25], stage1_19[26], stage1_19[27], stage1_19[28], stage1_19[29]},
      {stage2_21[4],stage2_20[6],stage2_19[6],stage2_18[37],stage2_17[52]}
   );
   gpc606_5 gpc4996 (
      {stage1_17[30], stage1_17[31], stage1_17[32], stage1_17[33], stage1_17[34], stage1_17[35]},
      {stage1_19[30], stage1_19[31], stage1_19[32], stage1_19[33], stage1_19[34], stage1_19[35]},
      {stage2_21[5],stage2_20[7],stage2_19[7],stage2_18[38],stage2_17[53]}
   );
   gpc606_5 gpc4997 (
      {stage1_17[36], stage1_17[37], stage1_17[38], stage1_17[39], stage1_17[40], stage1_17[41]},
      {stage1_19[36], stage1_19[37], stage1_19[38], stage1_19[39], stage1_19[40], stage1_19[41]},
      {stage2_21[6],stage2_20[8],stage2_19[8],stage2_18[39],stage2_17[54]}
   );
   gpc606_5 gpc4998 (
      {stage1_17[42], stage1_17[43], stage1_17[44], stage1_17[45], stage1_17[46], stage1_17[47]},
      {stage1_19[42], stage1_19[43], stage1_19[44], stage1_19[45], stage1_19[46], stage1_19[47]},
      {stage2_21[7],stage2_20[9],stage2_19[9],stage2_18[40],stage2_17[55]}
   );
   gpc606_5 gpc4999 (
      {stage1_17[48], stage1_17[49], stage1_17[50], stage1_17[51], stage1_17[52], stage1_17[53]},
      {stage1_19[48], stage1_19[49], stage1_19[50], stage1_19[51], stage1_19[52], stage1_19[53]},
      {stage2_21[8],stage2_20[10],stage2_19[10],stage2_18[41],stage2_17[56]}
   );
   gpc606_5 gpc5000 (
      {stage1_17[54], stage1_17[55], stage1_17[56], stage1_17[57], stage1_17[58], stage1_17[59]},
      {stage1_19[54], stage1_19[55], stage1_19[56], stage1_19[57], stage1_19[58], stage1_19[59]},
      {stage2_21[9],stage2_20[11],stage2_19[11],stage2_18[42],stage2_17[57]}
   );
   gpc606_5 gpc5001 (
      {stage1_17[60], stage1_17[61], stage1_17[62], stage1_17[63], stage1_17[64], stage1_17[65]},
      {stage1_19[60], stage1_19[61], stage1_19[62], stage1_19[63], stage1_19[64], stage1_19[65]},
      {stage2_21[10],stage2_20[12],stage2_19[12],stage2_18[43],stage2_17[58]}
   );
   gpc606_5 gpc5002 (
      {stage1_17[66], stage1_17[67], stage1_17[68], stage1_17[69], stage1_17[70], stage1_17[71]},
      {stage1_19[66], stage1_19[67], stage1_19[68], stage1_19[69], stage1_19[70], stage1_19[71]},
      {stage2_21[11],stage2_20[13],stage2_19[13],stage2_18[44],stage2_17[59]}
   );
   gpc606_5 gpc5003 (
      {stage1_17[72], stage1_17[73], stage1_17[74], stage1_17[75], stage1_17[76], stage1_17[77]},
      {stage1_19[72], stage1_19[73], stage1_19[74], stage1_19[75], stage1_19[76], stage1_19[77]},
      {stage2_21[12],stage2_20[14],stage2_19[14],stage2_18[45],stage2_17[60]}
   );
   gpc606_5 gpc5004 (
      {stage1_17[78], stage1_17[79], stage1_17[80], stage1_17[81], stage1_17[82], stage1_17[83]},
      {stage1_19[78], stage1_19[79], stage1_19[80], stage1_19[81], stage1_19[82], stage1_19[83]},
      {stage2_21[13],stage2_20[15],stage2_19[15],stage2_18[46],stage2_17[61]}
   );
   gpc606_5 gpc5005 (
      {stage1_17[84], stage1_17[85], stage1_17[86], stage1_17[87], stage1_17[88], stage1_17[89]},
      {stage1_19[84], stage1_19[85], stage1_19[86], stage1_19[87], stage1_19[88], stage1_19[89]},
      {stage2_21[14],stage2_20[16],stage2_19[16],stage2_18[47],stage2_17[62]}
   );
   gpc606_5 gpc5006 (
      {stage1_17[90], stage1_17[91], stage1_17[92], stage1_17[93], stage1_17[94], stage1_17[95]},
      {stage1_19[90], stage1_19[91], stage1_19[92], stage1_19[93], stage1_19[94], stage1_19[95]},
      {stage2_21[15],stage2_20[17],stage2_19[17],stage2_18[48],stage2_17[63]}
   );
   gpc606_5 gpc5007 (
      {stage1_17[96], stage1_17[97], stage1_17[98], stage1_17[99], stage1_17[100], stage1_17[101]},
      {stage1_19[96], stage1_19[97], stage1_19[98], stage1_19[99], stage1_19[100], stage1_19[101]},
      {stage2_21[16],stage2_20[18],stage2_19[18],stage2_18[49],stage2_17[64]}
   );
   gpc606_5 gpc5008 (
      {stage1_17[102], stage1_17[103], stage1_17[104], stage1_17[105], stage1_17[106], stage1_17[107]},
      {stage1_19[102], stage1_19[103], stage1_19[104], stage1_19[105], stage1_19[106], stage1_19[107]},
      {stage2_21[17],stage2_20[19],stage2_19[19],stage2_18[50],stage2_17[65]}
   );
   gpc606_5 gpc5009 (
      {stage1_17[108], stage1_17[109], stage1_17[110], stage1_17[111], stage1_17[112], stage1_17[113]},
      {stage1_19[108], stage1_19[109], stage1_19[110], stage1_19[111], stage1_19[112], stage1_19[113]},
      {stage2_21[18],stage2_20[20],stage2_19[20],stage2_18[51],stage2_17[66]}
   );
   gpc606_5 gpc5010 (
      {stage1_17[114], stage1_17[115], stage1_17[116], stage1_17[117], stage1_17[118], stage1_17[119]},
      {stage1_19[114], stage1_19[115], stage1_19[116], stage1_19[117], stage1_19[118], stage1_19[119]},
      {stage2_21[19],stage2_20[21],stage2_19[21],stage2_18[52],stage2_17[67]}
   );
   gpc606_5 gpc5011 (
      {stage1_17[120], stage1_17[121], stage1_17[122], stage1_17[123], stage1_17[124], stage1_17[125]},
      {stage1_19[120], stage1_19[121], stage1_19[122], stage1_19[123], stage1_19[124], stage1_19[125]},
      {stage2_21[20],stage2_20[22],stage2_19[22],stage2_18[53],stage2_17[68]}
   );
   gpc606_5 gpc5012 (
      {stage1_17[126], stage1_17[127], stage1_17[128], stage1_17[129], stage1_17[130], stage1_17[131]},
      {stage1_19[126], stage1_19[127], stage1_19[128], stage1_19[129], stage1_19[130], stage1_19[131]},
      {stage2_21[21],stage2_20[23],stage2_19[23],stage2_18[54],stage2_17[69]}
   );
   gpc606_5 gpc5013 (
      {stage1_17[132], stage1_17[133], stage1_17[134], stage1_17[135], stage1_17[136], stage1_17[137]},
      {stage1_19[132], stage1_19[133], stage1_19[134], stage1_19[135], stage1_19[136], stage1_19[137]},
      {stage2_21[22],stage2_20[24],stage2_19[24],stage2_18[55],stage2_17[70]}
   );
   gpc606_5 gpc5014 (
      {stage1_17[138], stage1_17[139], stage1_17[140], stage1_17[141], stage1_17[142], stage1_17[143]},
      {stage1_19[138], stage1_19[139], stage1_19[140], stage1_19[141], stage1_19[142], stage1_19[143]},
      {stage2_21[23],stage2_20[25],stage2_19[25],stage2_18[56],stage2_17[71]}
   );
   gpc606_5 gpc5015 (
      {stage1_17[144], stage1_17[145], stage1_17[146], stage1_17[147], stage1_17[148], stage1_17[149]},
      {stage1_19[144], stage1_19[145], stage1_19[146], stage1_19[147], stage1_19[148], stage1_19[149]},
      {stage2_21[24],stage2_20[26],stage2_19[26],stage2_18[57],stage2_17[72]}
   );
   gpc606_5 gpc5016 (
      {stage1_17[150], stage1_17[151], stage1_17[152], stage1_17[153], stage1_17[154], stage1_17[155]},
      {stage1_19[150], stage1_19[151], stage1_19[152], stage1_19[153], stage1_19[154], stage1_19[155]},
      {stage2_21[25],stage2_20[27],stage2_19[27],stage2_18[58],stage2_17[73]}
   );
   gpc606_5 gpc5017 (
      {stage1_17[156], stage1_17[157], stage1_17[158], stage1_17[159], stage1_17[160], stage1_17[161]},
      {stage1_19[156], stage1_19[157], stage1_19[158], stage1_19[159], stage1_19[160], stage1_19[161]},
      {stage2_21[26],stage2_20[28],stage2_19[28],stage2_18[59],stage2_17[74]}
   );
   gpc606_5 gpc5018 (
      {stage1_17[162], stage1_17[163], stage1_17[164], stage1_17[165], stage1_17[166], stage1_17[167]},
      {stage1_19[162], stage1_19[163], stage1_19[164], stage1_19[165], stage1_19[166], stage1_19[167]},
      {stage2_21[27],stage2_20[29],stage2_19[29],stage2_18[60],stage2_17[75]}
   );
   gpc606_5 gpc5019 (
      {stage1_17[168], stage1_17[169], stage1_17[170], stage1_17[171], stage1_17[172], stage1_17[173]},
      {stage1_19[168], stage1_19[169], stage1_19[170], stage1_19[171], stage1_19[172], stage1_19[173]},
      {stage2_21[28],stage2_20[30],stage2_19[30],stage2_18[61],stage2_17[76]}
   );
   gpc606_5 gpc5020 (
      {stage1_17[174], stage1_17[175], stage1_17[176], stage1_17[177], stage1_17[178], stage1_17[179]},
      {stage1_19[174], stage1_19[175], stage1_19[176], stage1_19[177], stage1_19[178], stage1_19[179]},
      {stage2_21[29],stage2_20[31],stage2_19[31],stage2_18[62],stage2_17[77]}
   );
   gpc606_5 gpc5021 (
      {stage1_17[180], stage1_17[181], stage1_17[182], stage1_17[183], stage1_17[184], stage1_17[185]},
      {stage1_19[180], stage1_19[181], stage1_19[182], stage1_19[183], stage1_19[184], stage1_19[185]},
      {stage2_21[30],stage2_20[32],stage2_19[32],stage2_18[63],stage2_17[78]}
   );
   gpc606_5 gpc5022 (
      {stage1_17[186], stage1_17[187], stage1_17[188], stage1_17[189], stage1_17[190], stage1_17[191]},
      {stage1_19[186], stage1_19[187], stage1_19[188], stage1_19[189], stage1_19[190], stage1_19[191]},
      {stage2_21[31],stage2_20[33],stage2_19[33],stage2_18[64],stage2_17[79]}
   );
   gpc606_5 gpc5023 (
      {stage1_17[192], stage1_17[193], stage1_17[194], stage1_17[195], stage1_17[196], stage1_17[197]},
      {stage1_19[192], stage1_19[193], stage1_19[194], stage1_19[195], stage1_19[196], stage1_19[197]},
      {stage2_21[32],stage2_20[34],stage2_19[34],stage2_18[65],stage2_17[80]}
   );
   gpc606_5 gpc5024 (
      {stage1_17[198], stage1_17[199], stage1_17[200], stage1_17[201], stage1_17[202], stage1_17[203]},
      {stage1_19[198], stage1_19[199], stage1_19[200], stage1_19[201], stage1_19[202], stage1_19[203]},
      {stage2_21[33],stage2_20[35],stage2_19[35],stage2_18[66],stage2_17[81]}
   );
   gpc606_5 gpc5025 (
      {stage1_17[204], stage1_17[205], stage1_17[206], stage1_17[207], stage1_17[208], stage1_17[209]},
      {stage1_19[204], stage1_19[205], stage1_19[206], stage1_19[207], stage1_19[208], stage1_19[209]},
      {stage2_21[34],stage2_20[36],stage2_19[36],stage2_18[67],stage2_17[82]}
   );
   gpc606_5 gpc5026 (
      {stage1_17[210], stage1_17[211], stage1_17[212], stage1_17[213], stage1_17[214], stage1_17[215]},
      {stage1_19[210], stage1_19[211], stage1_19[212], stage1_19[213], stage1_19[214], stage1_19[215]},
      {stage2_21[35],stage2_20[37],stage2_19[37],stage2_18[68],stage2_17[83]}
   );
   gpc606_5 gpc5027 (
      {stage1_17[216], stage1_17[217], stage1_17[218], stage1_17[219], stage1_17[220], stage1_17[221]},
      {stage1_19[216], stage1_19[217], stage1_19[218], stage1_19[219], stage1_19[220], stage1_19[221]},
      {stage2_21[36],stage2_20[38],stage2_19[38],stage2_18[69],stage2_17[84]}
   );
   gpc606_5 gpc5028 (
      {stage1_17[222], stage1_17[223], stage1_17[224], stage1_17[225], stage1_17[226], stage1_17[227]},
      {stage1_19[222], stage1_19[223], stage1_19[224], stage1_19[225], stage1_19[226], stage1_19[227]},
      {stage2_21[37],stage2_20[39],stage2_19[39],stage2_18[70],stage2_17[85]}
   );
   gpc606_5 gpc5029 (
      {stage1_18[12], stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[38],stage2_20[40],stage2_19[40],stage2_18[71]}
   );
   gpc606_5 gpc5030 (
      {stage1_18[18], stage1_18[19], stage1_18[20], stage1_18[21], stage1_18[22], stage1_18[23]},
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage2_22[1],stage2_21[39],stage2_20[41],stage2_19[41],stage2_18[72]}
   );
   gpc606_5 gpc5031 (
      {stage1_18[24], stage1_18[25], stage1_18[26], stage1_18[27], stage1_18[28], stage1_18[29]},
      {stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15], stage1_20[16], stage1_20[17]},
      {stage2_22[2],stage2_21[40],stage2_20[42],stage2_19[42],stage2_18[73]}
   );
   gpc606_5 gpc5032 (
      {stage1_18[30], stage1_18[31], stage1_18[32], stage1_18[33], stage1_18[34], stage1_18[35]},
      {stage1_20[18], stage1_20[19], stage1_20[20], stage1_20[21], stage1_20[22], stage1_20[23]},
      {stage2_22[3],stage2_21[41],stage2_20[43],stage2_19[43],stage2_18[74]}
   );
   gpc606_5 gpc5033 (
      {stage1_18[36], stage1_18[37], stage1_18[38], stage1_18[39], stage1_18[40], stage1_18[41]},
      {stage1_20[24], stage1_20[25], stage1_20[26], stage1_20[27], stage1_20[28], stage1_20[29]},
      {stage2_22[4],stage2_21[42],stage2_20[44],stage2_19[44],stage2_18[75]}
   );
   gpc606_5 gpc5034 (
      {stage1_18[42], stage1_18[43], stage1_18[44], stage1_18[45], stage1_18[46], stage1_18[47]},
      {stage1_20[30], stage1_20[31], stage1_20[32], stage1_20[33], stage1_20[34], stage1_20[35]},
      {stage2_22[5],stage2_21[43],stage2_20[45],stage2_19[45],stage2_18[76]}
   );
   gpc606_5 gpc5035 (
      {stage1_18[48], stage1_18[49], stage1_18[50], stage1_18[51], stage1_18[52], stage1_18[53]},
      {stage1_20[36], stage1_20[37], stage1_20[38], stage1_20[39], stage1_20[40], stage1_20[41]},
      {stage2_22[6],stage2_21[44],stage2_20[46],stage2_19[46],stage2_18[77]}
   );
   gpc606_5 gpc5036 (
      {stage1_18[54], stage1_18[55], stage1_18[56], stage1_18[57], stage1_18[58], stage1_18[59]},
      {stage1_20[42], stage1_20[43], stage1_20[44], stage1_20[45], stage1_20[46], stage1_20[47]},
      {stage2_22[7],stage2_21[45],stage2_20[47],stage2_19[47],stage2_18[78]}
   );
   gpc606_5 gpc5037 (
      {stage1_18[60], stage1_18[61], stage1_18[62], stage1_18[63], stage1_18[64], stage1_18[65]},
      {stage1_20[48], stage1_20[49], stage1_20[50], stage1_20[51], stage1_20[52], stage1_20[53]},
      {stage2_22[8],stage2_21[46],stage2_20[48],stage2_19[48],stage2_18[79]}
   );
   gpc606_5 gpc5038 (
      {stage1_18[66], stage1_18[67], stage1_18[68], stage1_18[69], stage1_18[70], stage1_18[71]},
      {stage1_20[54], stage1_20[55], stage1_20[56], stage1_20[57], stage1_20[58], stage1_20[59]},
      {stage2_22[9],stage2_21[47],stage2_20[49],stage2_19[49],stage2_18[80]}
   );
   gpc606_5 gpc5039 (
      {stage1_18[72], stage1_18[73], stage1_18[74], stage1_18[75], stage1_18[76], stage1_18[77]},
      {stage1_20[60], stage1_20[61], stage1_20[62], stage1_20[63], stage1_20[64], stage1_20[65]},
      {stage2_22[10],stage2_21[48],stage2_20[50],stage2_19[50],stage2_18[81]}
   );
   gpc606_5 gpc5040 (
      {stage1_18[78], stage1_18[79], stage1_18[80], stage1_18[81], stage1_18[82], stage1_18[83]},
      {stage1_20[66], stage1_20[67], stage1_20[68], stage1_20[69], stage1_20[70], stage1_20[71]},
      {stage2_22[11],stage2_21[49],stage2_20[51],stage2_19[51],stage2_18[82]}
   );
   gpc606_5 gpc5041 (
      {stage1_18[84], stage1_18[85], stage1_18[86], stage1_18[87], stage1_18[88], stage1_18[89]},
      {stage1_20[72], stage1_20[73], stage1_20[74], stage1_20[75], stage1_20[76], stage1_20[77]},
      {stage2_22[12],stage2_21[50],stage2_20[52],stage2_19[52],stage2_18[83]}
   );
   gpc606_5 gpc5042 (
      {stage1_18[90], stage1_18[91], stage1_18[92], stage1_18[93], stage1_18[94], stage1_18[95]},
      {stage1_20[78], stage1_20[79], stage1_20[80], stage1_20[81], stage1_20[82], stage1_20[83]},
      {stage2_22[13],stage2_21[51],stage2_20[53],stage2_19[53],stage2_18[84]}
   );
   gpc606_5 gpc5043 (
      {stage1_18[96], stage1_18[97], stage1_18[98], stage1_18[99], stage1_18[100], stage1_18[101]},
      {stage1_20[84], stage1_20[85], stage1_20[86], stage1_20[87], stage1_20[88], stage1_20[89]},
      {stage2_22[14],stage2_21[52],stage2_20[54],stage2_19[54],stage2_18[85]}
   );
   gpc606_5 gpc5044 (
      {stage1_18[102], stage1_18[103], stage1_18[104], stage1_18[105], stage1_18[106], stage1_18[107]},
      {stage1_20[90], stage1_20[91], stage1_20[92], stage1_20[93], stage1_20[94], stage1_20[95]},
      {stage2_22[15],stage2_21[53],stage2_20[55],stage2_19[55],stage2_18[86]}
   );
   gpc606_5 gpc5045 (
      {stage1_18[108], stage1_18[109], stage1_18[110], stage1_18[111], stage1_18[112], stage1_18[113]},
      {stage1_20[96], stage1_20[97], stage1_20[98], stage1_20[99], stage1_20[100], stage1_20[101]},
      {stage2_22[16],stage2_21[54],stage2_20[56],stage2_19[56],stage2_18[87]}
   );
   gpc606_5 gpc5046 (
      {stage1_18[114], stage1_18[115], stage1_18[116], stage1_18[117], stage1_18[118], stage1_18[119]},
      {stage1_20[102], stage1_20[103], stage1_20[104], stage1_20[105], stage1_20[106], stage1_20[107]},
      {stage2_22[17],stage2_21[55],stage2_20[57],stage2_19[57],stage2_18[88]}
   );
   gpc606_5 gpc5047 (
      {stage1_18[120], stage1_18[121], stage1_18[122], stage1_18[123], stage1_18[124], stage1_18[125]},
      {stage1_20[108], stage1_20[109], stage1_20[110], stage1_20[111], stage1_20[112], stage1_20[113]},
      {stage2_22[18],stage2_21[56],stage2_20[58],stage2_19[58],stage2_18[89]}
   );
   gpc606_5 gpc5048 (
      {stage1_18[126], stage1_18[127], stage1_18[128], stage1_18[129], stage1_18[130], stage1_18[131]},
      {stage1_20[114], stage1_20[115], stage1_20[116], stage1_20[117], stage1_20[118], stage1_20[119]},
      {stage2_22[19],stage2_21[57],stage2_20[59],stage2_19[59],stage2_18[90]}
   );
   gpc606_5 gpc5049 (
      {stage1_18[132], stage1_18[133], stage1_18[134], stage1_18[135], stage1_18[136], stage1_18[137]},
      {stage1_20[120], stage1_20[121], stage1_20[122], stage1_20[123], stage1_20[124], stage1_20[125]},
      {stage2_22[20],stage2_21[58],stage2_20[60],stage2_19[60],stage2_18[91]}
   );
   gpc606_5 gpc5050 (
      {stage1_18[138], stage1_18[139], stage1_18[140], stage1_18[141], stage1_18[142], stage1_18[143]},
      {stage1_20[126], stage1_20[127], stage1_20[128], stage1_20[129], stage1_20[130], stage1_20[131]},
      {stage2_22[21],stage2_21[59],stage2_20[61],stage2_19[61],stage2_18[92]}
   );
   gpc606_5 gpc5051 (
      {stage1_18[144], stage1_18[145], stage1_18[146], stage1_18[147], stage1_18[148], stage1_18[149]},
      {stage1_20[132], stage1_20[133], stage1_20[134], stage1_20[135], stage1_20[136], stage1_20[137]},
      {stage2_22[22],stage2_21[60],stage2_20[62],stage2_19[62],stage2_18[93]}
   );
   gpc606_5 gpc5052 (
      {stage1_18[150], stage1_18[151], stage1_18[152], stage1_18[153], stage1_18[154], stage1_18[155]},
      {stage1_20[138], stage1_20[139], stage1_20[140], stage1_20[141], stage1_20[142], stage1_20[143]},
      {stage2_22[23],stage2_21[61],stage2_20[63],stage2_19[63],stage2_18[94]}
   );
   gpc606_5 gpc5053 (
      {stage1_18[156], stage1_18[157], stage1_18[158], stage1_18[159], stage1_18[160], stage1_18[161]},
      {stage1_20[144], stage1_20[145], stage1_20[146], stage1_20[147], stage1_20[148], stage1_20[149]},
      {stage2_22[24],stage2_21[62],stage2_20[64],stage2_19[64],stage2_18[95]}
   );
   gpc606_5 gpc5054 (
      {stage1_18[162], stage1_18[163], stage1_18[164], stage1_18[165], stage1_18[166], stage1_18[167]},
      {stage1_20[150], stage1_20[151], stage1_20[152], stage1_20[153], stage1_20[154], stage1_20[155]},
      {stage2_22[25],stage2_21[63],stage2_20[65],stage2_19[65],stage2_18[96]}
   );
   gpc606_5 gpc5055 (
      {stage1_18[168], stage1_18[169], stage1_18[170], stage1_18[171], stage1_18[172], stage1_18[173]},
      {stage1_20[156], stage1_20[157], stage1_20[158], stage1_20[159], stage1_20[160], stage1_20[161]},
      {stage2_22[26],stage2_21[64],stage2_20[66],stage2_19[66],stage2_18[97]}
   );
   gpc606_5 gpc5056 (
      {stage1_18[174], stage1_18[175], stage1_18[176], stage1_18[177], stage1_18[178], stage1_18[179]},
      {stage1_20[162], stage1_20[163], stage1_20[164], stage1_20[165], stage1_20[166], stage1_20[167]},
      {stage2_22[27],stage2_21[65],stage2_20[67],stage2_19[67],stage2_18[98]}
   );
   gpc606_5 gpc5057 (
      {stage1_18[180], stage1_18[181], stage1_18[182], stage1_18[183], stage1_18[184], stage1_18[185]},
      {stage1_20[168], stage1_20[169], stage1_20[170], stage1_20[171], stage1_20[172], stage1_20[173]},
      {stage2_22[28],stage2_21[66],stage2_20[68],stage2_19[68],stage2_18[99]}
   );
   gpc615_5 gpc5058 (
      {stage1_18[186], stage1_18[187], stage1_18[188], stage1_18[189], stage1_18[190]},
      {stage1_19[228]},
      {stage1_20[174], stage1_20[175], stage1_20[176], stage1_20[177], stage1_20[178], stage1_20[179]},
      {stage2_22[29],stage2_21[67],stage2_20[69],stage2_19[69],stage2_18[100]}
   );
   gpc615_5 gpc5059 (
      {stage1_19[229], stage1_19[230], stage1_19[231], stage1_19[232], stage1_19[233]},
      {stage1_20[180]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[30],stage2_21[68],stage2_20[70],stage2_19[70]}
   );
   gpc606_5 gpc5060 (
      {stage1_20[181], stage1_20[182], stage1_20[183], stage1_20[184], stage1_20[185], stage1_20[186]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[1],stage2_22[31],stage2_21[69],stage2_20[71]}
   );
   gpc615_5 gpc5061 (
      {stage1_20[187], stage1_20[188], stage1_20[189], stage1_20[190], stage1_20[191]},
      {stage1_21[6]},
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage2_24[1],stage2_23[2],stage2_22[32],stage2_21[70],stage2_20[72]}
   );
   gpc615_5 gpc5062 (
      {stage1_20[192], stage1_20[193], stage1_20[194], stage1_20[195], stage1_20[196]},
      {stage1_21[7]},
      {stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage2_24[2],stage2_23[3],stage2_22[33],stage2_21[71],stage2_20[73]}
   );
   gpc615_5 gpc5063 (
      {stage1_20[197], stage1_20[198], stage1_20[199], stage1_20[200], stage1_20[201]},
      {stage1_21[8]},
      {stage1_22[18], stage1_22[19], stage1_22[20], stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage2_24[3],stage2_23[4],stage2_22[34],stage2_21[72],stage2_20[74]}
   );
   gpc615_5 gpc5064 (
      {stage1_20[202], stage1_20[203], stage1_20[204], stage1_20[205], stage1_20[206]},
      {stage1_21[9]},
      {stage1_22[24], stage1_22[25], stage1_22[26], stage1_22[27], stage1_22[28], stage1_22[29]},
      {stage2_24[4],stage2_23[5],stage2_22[35],stage2_21[73],stage2_20[75]}
   );
   gpc615_5 gpc5065 (
      {stage1_20[207], stage1_20[208], stage1_20[209], stage1_20[210], stage1_20[211]},
      {stage1_21[10]},
      {stage1_22[30], stage1_22[31], stage1_22[32], stage1_22[33], stage1_22[34], stage1_22[35]},
      {stage2_24[5],stage2_23[6],stage2_22[36],stage2_21[74],stage2_20[76]}
   );
   gpc615_5 gpc5066 (
      {stage1_20[212], stage1_20[213], stage1_20[214], stage1_20[215], stage1_20[216]},
      {stage1_21[11]},
      {stage1_22[36], stage1_22[37], stage1_22[38], stage1_22[39], stage1_22[40], stage1_22[41]},
      {stage2_24[6],stage2_23[7],stage2_22[37],stage2_21[75],stage2_20[77]}
   );
   gpc615_5 gpc5067 (
      {stage1_20[217], stage1_20[218], stage1_20[219], stage1_20[220], stage1_20[221]},
      {stage1_21[12]},
      {stage1_22[42], stage1_22[43], stage1_22[44], stage1_22[45], stage1_22[46], stage1_22[47]},
      {stage2_24[7],stage2_23[8],stage2_22[38],stage2_21[76],stage2_20[78]}
   );
   gpc615_5 gpc5068 (
      {stage1_20[222], stage1_20[223], stage1_20[224], stage1_20[225], stage1_20[226]},
      {stage1_21[13]},
      {stage1_22[48], stage1_22[49], stage1_22[50], stage1_22[51], stage1_22[52], stage1_22[53]},
      {stage2_24[8],stage2_23[9],stage2_22[39],stage2_21[77],stage2_20[79]}
   );
   gpc615_5 gpc5069 (
      {stage1_20[227], stage1_20[228], stage1_20[229], stage1_20[230], stage1_20[231]},
      {stage1_21[14]},
      {stage1_22[54], stage1_22[55], stage1_22[56], stage1_22[57], stage1_22[58], stage1_22[59]},
      {stage2_24[9],stage2_23[10],stage2_22[40],stage2_21[78],stage2_20[80]}
   );
   gpc615_5 gpc5070 (
      {stage1_20[232], stage1_20[233], stage1_20[234], stage1_20[235], stage1_20[236]},
      {stage1_21[15]},
      {stage1_22[60], stage1_22[61], stage1_22[62], stage1_22[63], stage1_22[64], stage1_22[65]},
      {stage2_24[10],stage2_23[11],stage2_22[41],stage2_21[79],stage2_20[81]}
   );
   gpc615_5 gpc5071 (
      {stage1_20[237], stage1_20[238], stage1_20[239], stage1_20[240], stage1_20[241]},
      {stage1_21[16]},
      {stage1_22[66], stage1_22[67], stage1_22[68], stage1_22[69], stage1_22[70], stage1_22[71]},
      {stage2_24[11],stage2_23[12],stage2_22[42],stage2_21[80],stage2_20[82]}
   );
   gpc615_5 gpc5072 (
      {stage1_20[242], stage1_20[243], stage1_20[244], stage1_20[245], stage1_20[246]},
      {stage1_21[17]},
      {stage1_22[72], stage1_22[73], stage1_22[74], stage1_22[75], stage1_22[76], stage1_22[77]},
      {stage2_24[12],stage2_23[13],stage2_22[43],stage2_21[81],stage2_20[83]}
   );
   gpc615_5 gpc5073 (
      {stage1_20[247], stage1_20[248], stage1_20[249], stage1_20[250], stage1_20[251]},
      {stage1_21[18]},
      {stage1_22[78], stage1_22[79], stage1_22[80], stage1_22[81], stage1_22[82], stage1_22[83]},
      {stage2_24[13],stage2_23[14],stage2_22[44],stage2_21[82],stage2_20[84]}
   );
   gpc615_5 gpc5074 (
      {stage1_20[252], stage1_20[253], stage1_20[254], stage1_20[255], stage1_20[256]},
      {stage1_21[19]},
      {stage1_22[84], stage1_22[85], stage1_22[86], stage1_22[87], stage1_22[88], stage1_22[89]},
      {stage2_24[14],stage2_23[15],stage2_22[45],stage2_21[83],stage2_20[85]}
   );
   gpc615_5 gpc5075 (
      {stage1_20[257], stage1_20[258], stage1_20[259], stage1_20[260], stage1_20[261]},
      {stage1_21[20]},
      {stage1_22[90], stage1_22[91], stage1_22[92], stage1_22[93], stage1_22[94], stage1_22[95]},
      {stage2_24[15],stage2_23[16],stage2_22[46],stage2_21[84],stage2_20[86]}
   );
   gpc606_5 gpc5076 (
      {stage1_21[21], stage1_21[22], stage1_21[23], stage1_21[24], stage1_21[25], stage1_21[26]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[16],stage2_23[17],stage2_22[47],stage2_21[85]}
   );
   gpc606_5 gpc5077 (
      {stage1_21[27], stage1_21[28], stage1_21[29], stage1_21[30], stage1_21[31], stage1_21[32]},
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage2_25[1],stage2_24[17],stage2_23[18],stage2_22[48],stage2_21[86]}
   );
   gpc606_5 gpc5078 (
      {stage1_21[33], stage1_21[34], stage1_21[35], stage1_21[36], stage1_21[37], stage1_21[38]},
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage2_25[2],stage2_24[18],stage2_23[19],stage2_22[49],stage2_21[87]}
   );
   gpc606_5 gpc5079 (
      {stage1_21[39], stage1_21[40], stage1_21[41], stage1_21[42], stage1_21[43], stage1_21[44]},
      {stage1_23[18], stage1_23[19], stage1_23[20], stage1_23[21], stage1_23[22], stage1_23[23]},
      {stage2_25[3],stage2_24[19],stage2_23[20],stage2_22[50],stage2_21[88]}
   );
   gpc606_5 gpc5080 (
      {stage1_21[45], stage1_21[46], stage1_21[47], stage1_21[48], stage1_21[49], stage1_21[50]},
      {stage1_23[24], stage1_23[25], stage1_23[26], stage1_23[27], stage1_23[28], stage1_23[29]},
      {stage2_25[4],stage2_24[20],stage2_23[21],stage2_22[51],stage2_21[89]}
   );
   gpc606_5 gpc5081 (
      {stage1_21[51], stage1_21[52], stage1_21[53], stage1_21[54], stage1_21[55], stage1_21[56]},
      {stage1_23[30], stage1_23[31], stage1_23[32], stage1_23[33], stage1_23[34], stage1_23[35]},
      {stage2_25[5],stage2_24[21],stage2_23[22],stage2_22[52],stage2_21[90]}
   );
   gpc606_5 gpc5082 (
      {stage1_21[57], stage1_21[58], stage1_21[59], stage1_21[60], stage1_21[61], stage1_21[62]},
      {stage1_23[36], stage1_23[37], stage1_23[38], stage1_23[39], stage1_23[40], stage1_23[41]},
      {stage2_25[6],stage2_24[22],stage2_23[23],stage2_22[53],stage2_21[91]}
   );
   gpc606_5 gpc5083 (
      {stage1_21[63], stage1_21[64], stage1_21[65], stage1_21[66], stage1_21[67], stage1_21[68]},
      {stage1_23[42], stage1_23[43], stage1_23[44], stage1_23[45], stage1_23[46], stage1_23[47]},
      {stage2_25[7],stage2_24[23],stage2_23[24],stage2_22[54],stage2_21[92]}
   );
   gpc606_5 gpc5084 (
      {stage1_21[69], stage1_21[70], stage1_21[71], stage1_21[72], stage1_21[73], stage1_21[74]},
      {stage1_23[48], stage1_23[49], stage1_23[50], stage1_23[51], stage1_23[52], stage1_23[53]},
      {stage2_25[8],stage2_24[24],stage2_23[25],stage2_22[55],stage2_21[93]}
   );
   gpc606_5 gpc5085 (
      {stage1_21[75], stage1_21[76], stage1_21[77], stage1_21[78], stage1_21[79], stage1_21[80]},
      {stage1_23[54], stage1_23[55], stage1_23[56], stage1_23[57], stage1_23[58], stage1_23[59]},
      {stage2_25[9],stage2_24[25],stage2_23[26],stage2_22[56],stage2_21[94]}
   );
   gpc606_5 gpc5086 (
      {stage1_21[81], stage1_21[82], stage1_21[83], stage1_21[84], stage1_21[85], stage1_21[86]},
      {stage1_23[60], stage1_23[61], stage1_23[62], stage1_23[63], stage1_23[64], stage1_23[65]},
      {stage2_25[10],stage2_24[26],stage2_23[27],stage2_22[57],stage2_21[95]}
   );
   gpc606_5 gpc5087 (
      {stage1_21[87], stage1_21[88], stage1_21[89], stage1_21[90], stage1_21[91], stage1_21[92]},
      {stage1_23[66], stage1_23[67], stage1_23[68], stage1_23[69], stage1_23[70], stage1_23[71]},
      {stage2_25[11],stage2_24[27],stage2_23[28],stage2_22[58],stage2_21[96]}
   );
   gpc606_5 gpc5088 (
      {stage1_21[93], stage1_21[94], stage1_21[95], stage1_21[96], stage1_21[97], stage1_21[98]},
      {stage1_23[72], stage1_23[73], stage1_23[74], stage1_23[75], stage1_23[76], stage1_23[77]},
      {stage2_25[12],stage2_24[28],stage2_23[29],stage2_22[59],stage2_21[97]}
   );
   gpc606_5 gpc5089 (
      {stage1_21[99], stage1_21[100], stage1_21[101], stage1_21[102], stage1_21[103], stage1_21[104]},
      {stage1_23[78], stage1_23[79], stage1_23[80], stage1_23[81], stage1_23[82], stage1_23[83]},
      {stage2_25[13],stage2_24[29],stage2_23[30],stage2_22[60],stage2_21[98]}
   );
   gpc606_5 gpc5090 (
      {stage1_21[105], stage1_21[106], stage1_21[107], stage1_21[108], stage1_21[109], stage1_21[110]},
      {stage1_23[84], stage1_23[85], stage1_23[86], stage1_23[87], stage1_23[88], stage1_23[89]},
      {stage2_25[14],stage2_24[30],stage2_23[31],stage2_22[61],stage2_21[99]}
   );
   gpc606_5 gpc5091 (
      {stage1_21[111], stage1_21[112], stage1_21[113], stage1_21[114], stage1_21[115], stage1_21[116]},
      {stage1_23[90], stage1_23[91], stage1_23[92], stage1_23[93], stage1_23[94], stage1_23[95]},
      {stage2_25[15],stage2_24[31],stage2_23[32],stage2_22[62],stage2_21[100]}
   );
   gpc606_5 gpc5092 (
      {stage1_21[117], stage1_21[118], stage1_21[119], stage1_21[120], stage1_21[121], stage1_21[122]},
      {stage1_23[96], stage1_23[97], stage1_23[98], stage1_23[99], stage1_23[100], stage1_23[101]},
      {stage2_25[16],stage2_24[32],stage2_23[33],stage2_22[63],stage2_21[101]}
   );
   gpc606_5 gpc5093 (
      {stage1_21[123], stage1_21[124], stage1_21[125], stage1_21[126], stage1_21[127], stage1_21[128]},
      {stage1_23[102], stage1_23[103], stage1_23[104], stage1_23[105], stage1_23[106], stage1_23[107]},
      {stage2_25[17],stage2_24[33],stage2_23[34],stage2_22[64],stage2_21[102]}
   );
   gpc615_5 gpc5094 (
      {stage1_21[129], stage1_21[130], stage1_21[131], stage1_21[132], stage1_21[133]},
      {stage1_22[96]},
      {stage1_23[108], stage1_23[109], stage1_23[110], stage1_23[111], stage1_23[112], stage1_23[113]},
      {stage2_25[18],stage2_24[34],stage2_23[35],stage2_22[65],stage2_21[103]}
   );
   gpc615_5 gpc5095 (
      {stage1_21[134], stage1_21[135], stage1_21[136], stage1_21[137], stage1_21[138]},
      {stage1_22[97]},
      {stage1_23[114], stage1_23[115], stage1_23[116], stage1_23[117], stage1_23[118], stage1_23[119]},
      {stage2_25[19],stage2_24[35],stage2_23[36],stage2_22[66],stage2_21[104]}
   );
   gpc615_5 gpc5096 (
      {stage1_21[139], stage1_21[140], stage1_21[141], stage1_21[142], stage1_21[143]},
      {stage1_22[98]},
      {stage1_23[120], stage1_23[121], stage1_23[122], stage1_23[123], stage1_23[124], stage1_23[125]},
      {stage2_25[20],stage2_24[36],stage2_23[37],stage2_22[67],stage2_21[105]}
   );
   gpc615_5 gpc5097 (
      {stage1_21[144], stage1_21[145], stage1_21[146], stage1_21[147], stage1_21[148]},
      {stage1_22[99]},
      {stage1_23[126], stage1_23[127], stage1_23[128], stage1_23[129], stage1_23[130], stage1_23[131]},
      {stage2_25[21],stage2_24[37],stage2_23[38],stage2_22[68],stage2_21[106]}
   );
   gpc615_5 gpc5098 (
      {stage1_21[149], stage1_21[150], stage1_21[151], stage1_21[152], stage1_21[153]},
      {stage1_22[100]},
      {stage1_23[132], stage1_23[133], stage1_23[134], stage1_23[135], stage1_23[136], stage1_23[137]},
      {stage2_25[22],stage2_24[38],stage2_23[39],stage2_22[69],stage2_21[107]}
   );
   gpc615_5 gpc5099 (
      {stage1_21[154], stage1_21[155], stage1_21[156], stage1_21[157], stage1_21[158]},
      {stage1_22[101]},
      {stage1_23[138], stage1_23[139], stage1_23[140], stage1_23[141], stage1_23[142], stage1_23[143]},
      {stage2_25[23],stage2_24[39],stage2_23[40],stage2_22[70],stage2_21[108]}
   );
   gpc615_5 gpc5100 (
      {stage1_21[159], stage1_21[160], stage1_21[161], stage1_21[162], stage1_21[163]},
      {stage1_22[102]},
      {stage1_23[144], stage1_23[145], stage1_23[146], stage1_23[147], stage1_23[148], stage1_23[149]},
      {stage2_25[24],stage2_24[40],stage2_23[41],stage2_22[71],stage2_21[109]}
   );
   gpc615_5 gpc5101 (
      {stage1_21[164], stage1_21[165], stage1_21[166], stage1_21[167], stage1_21[168]},
      {stage1_22[103]},
      {stage1_23[150], stage1_23[151], stage1_23[152], stage1_23[153], stage1_23[154], stage1_23[155]},
      {stage2_25[25],stage2_24[41],stage2_23[42],stage2_22[72],stage2_21[110]}
   );
   gpc615_5 gpc5102 (
      {stage1_21[169], stage1_21[170], stage1_21[171], stage1_21[172], stage1_21[173]},
      {stage1_22[104]},
      {stage1_23[156], stage1_23[157], stage1_23[158], stage1_23[159], stage1_23[160], stage1_23[161]},
      {stage2_25[26],stage2_24[42],stage2_23[43],stage2_22[73],stage2_21[111]}
   );
   gpc615_5 gpc5103 (
      {stage1_22[105], stage1_22[106], stage1_22[107], stage1_22[108], stage1_22[109]},
      {stage1_23[162]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5]},
      {stage2_26[0],stage2_25[27],stage2_24[43],stage2_23[44],stage2_22[74]}
   );
   gpc615_5 gpc5104 (
      {stage1_22[110], stage1_22[111], stage1_22[112], stage1_22[113], stage1_22[114]},
      {stage1_23[163]},
      {stage1_24[6], stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11]},
      {stage2_26[1],stage2_25[28],stage2_24[44],stage2_23[45],stage2_22[75]}
   );
   gpc615_5 gpc5105 (
      {stage1_22[115], stage1_22[116], stage1_22[117], stage1_22[118], stage1_22[119]},
      {stage1_23[164]},
      {stage1_24[12], stage1_24[13], stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17]},
      {stage2_26[2],stage2_25[29],stage2_24[45],stage2_23[46],stage2_22[76]}
   );
   gpc615_5 gpc5106 (
      {stage1_22[120], stage1_22[121], stage1_22[122], stage1_22[123], stage1_22[124]},
      {stage1_23[165]},
      {stage1_24[18], stage1_24[19], stage1_24[20], stage1_24[21], stage1_24[22], stage1_24[23]},
      {stage2_26[3],stage2_25[30],stage2_24[46],stage2_23[47],stage2_22[77]}
   );
   gpc615_5 gpc5107 (
      {stage1_22[125], stage1_22[126], stage1_22[127], stage1_22[128], stage1_22[129]},
      {stage1_23[166]},
      {stage1_24[24], stage1_24[25], stage1_24[26], stage1_24[27], stage1_24[28], stage1_24[29]},
      {stage2_26[4],stage2_25[31],stage2_24[47],stage2_23[48],stage2_22[78]}
   );
   gpc615_5 gpc5108 (
      {stage1_22[130], stage1_22[131], stage1_22[132], stage1_22[133], stage1_22[134]},
      {stage1_23[167]},
      {stage1_24[30], stage1_24[31], stage1_24[32], stage1_24[33], stage1_24[34], stage1_24[35]},
      {stage2_26[5],stage2_25[32],stage2_24[48],stage2_23[49],stage2_22[79]}
   );
   gpc615_5 gpc5109 (
      {stage1_22[135], stage1_22[136], stage1_22[137], stage1_22[138], stage1_22[139]},
      {stage1_23[168]},
      {stage1_24[36], stage1_24[37], stage1_24[38], stage1_24[39], stage1_24[40], stage1_24[41]},
      {stage2_26[6],stage2_25[33],stage2_24[49],stage2_23[50],stage2_22[80]}
   );
   gpc615_5 gpc5110 (
      {stage1_22[140], stage1_22[141], stage1_22[142], stage1_22[143], stage1_22[144]},
      {stage1_23[169]},
      {stage1_24[42], stage1_24[43], stage1_24[44], stage1_24[45], stage1_24[46], stage1_24[47]},
      {stage2_26[7],stage2_25[34],stage2_24[50],stage2_23[51],stage2_22[81]}
   );
   gpc615_5 gpc5111 (
      {stage1_23[170], stage1_23[171], stage1_23[172], stage1_23[173], stage1_23[174]},
      {stage1_24[48]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[8],stage2_25[35],stage2_24[51],stage2_23[52]}
   );
   gpc615_5 gpc5112 (
      {stage1_23[175], stage1_23[176], stage1_23[177], stage1_23[178], stage1_23[179]},
      {stage1_24[49]},
      {stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11]},
      {stage2_27[1],stage2_26[9],stage2_25[36],stage2_24[52],stage2_23[53]}
   );
   gpc615_5 gpc5113 (
      {stage1_23[180], stage1_23[181], stage1_23[182], stage1_23[183], stage1_23[184]},
      {stage1_24[50]},
      {stage1_25[12], stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {stage2_27[2],stage2_26[10],stage2_25[37],stage2_24[53],stage2_23[54]}
   );
   gpc615_5 gpc5114 (
      {stage1_23[185], stage1_23[186], stage1_23[187], stage1_23[188], stage1_23[189]},
      {stage1_24[51]},
      {stage1_25[18], stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23]},
      {stage2_27[3],stage2_26[11],stage2_25[38],stage2_24[54],stage2_23[55]}
   );
   gpc615_5 gpc5115 (
      {stage1_23[190], stage1_23[191], stage1_23[192], stage1_23[193], stage1_23[194]},
      {stage1_24[52]},
      {stage1_25[24], stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29]},
      {stage2_27[4],stage2_26[12],stage2_25[39],stage2_24[55],stage2_23[56]}
   );
   gpc615_5 gpc5116 (
      {stage1_23[195], stage1_23[196], stage1_23[197], stage1_23[198], stage1_23[199]},
      {stage1_24[53]},
      {stage1_25[30], stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35]},
      {stage2_27[5],stage2_26[13],stage2_25[40],stage2_24[56],stage2_23[57]}
   );
   gpc615_5 gpc5117 (
      {stage1_23[200], stage1_23[201], stage1_23[202], stage1_23[203], stage1_23[204]},
      {stage1_24[54]},
      {stage1_25[36], stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41]},
      {stage2_27[6],stage2_26[14],stage2_25[41],stage2_24[57],stage2_23[58]}
   );
   gpc615_5 gpc5118 (
      {stage1_23[205], stage1_23[206], stage1_23[207], stage1_23[208], stage1_23[209]},
      {stage1_24[55]},
      {stage1_25[42], stage1_25[43], stage1_25[44], stage1_25[45], stage1_25[46], stage1_25[47]},
      {stage2_27[7],stage2_26[15],stage2_25[42],stage2_24[58],stage2_23[59]}
   );
   gpc615_5 gpc5119 (
      {stage1_23[210], stage1_23[211], stage1_23[212], stage1_23[213], stage1_23[214]},
      {stage1_24[56]},
      {stage1_25[48], stage1_25[49], stage1_25[50], stage1_25[51], stage1_25[52], stage1_25[53]},
      {stage2_27[8],stage2_26[16],stage2_25[43],stage2_24[59],stage2_23[60]}
   );
   gpc615_5 gpc5120 (
      {stage1_23[215], stage1_23[216], stage1_23[217], stage1_23[218], stage1_23[219]},
      {stage1_24[57]},
      {stage1_25[54], stage1_25[55], stage1_25[56], stage1_25[57], stage1_25[58], stage1_25[59]},
      {stage2_27[9],stage2_26[17],stage2_25[44],stage2_24[60],stage2_23[61]}
   );
   gpc615_5 gpc5121 (
      {stage1_23[220], stage1_23[221], stage1_23[222], stage1_23[223], stage1_23[224]},
      {stage1_24[58]},
      {stage1_25[60], stage1_25[61], stage1_25[62], stage1_25[63], stage1_25[64], stage1_25[65]},
      {stage2_27[10],stage2_26[18],stage2_25[45],stage2_24[61],stage2_23[62]}
   );
   gpc615_5 gpc5122 (
      {stage1_23[225], stage1_23[226], stage1_23[227], stage1_23[228], stage1_23[229]},
      {stage1_24[59]},
      {stage1_25[66], stage1_25[67], stage1_25[68], stage1_25[69], stage1_25[70], stage1_25[71]},
      {stage2_27[11],stage2_26[19],stage2_25[46],stage2_24[62],stage2_23[63]}
   );
   gpc615_5 gpc5123 (
      {stage1_23[230], stage1_23[231], stage1_23[232], stage1_23[233], stage1_23[234]},
      {stage1_24[60]},
      {stage1_25[72], stage1_25[73], stage1_25[74], stage1_25[75], stage1_25[76], stage1_25[77]},
      {stage2_27[12],stage2_26[20],stage2_25[47],stage2_24[63],stage2_23[64]}
   );
   gpc615_5 gpc5124 (
      {stage1_23[235], stage1_23[236], stage1_23[237], stage1_23[238], stage1_23[239]},
      {stage1_24[61]},
      {stage1_25[78], stage1_25[79], stage1_25[80], stage1_25[81], stage1_25[82], stage1_25[83]},
      {stage2_27[13],stage2_26[21],stage2_25[48],stage2_24[64],stage2_23[65]}
   );
   gpc615_5 gpc5125 (
      {stage1_23[240], stage1_23[241], stage1_23[242], stage1_23[243], stage1_23[244]},
      {stage1_24[62]},
      {stage1_25[84], stage1_25[85], stage1_25[86], stage1_25[87], stage1_25[88], stage1_25[89]},
      {stage2_27[14],stage2_26[22],stage2_25[49],stage2_24[65],stage2_23[66]}
   );
   gpc615_5 gpc5126 (
      {stage1_23[245], stage1_23[246], stage1_23[247], stage1_23[248], stage1_23[249]},
      {stage1_24[63]},
      {stage1_25[90], stage1_25[91], stage1_25[92], stage1_25[93], stage1_25[94], stage1_25[95]},
      {stage2_27[15],stage2_26[23],stage2_25[50],stage2_24[66],stage2_23[67]}
   );
   gpc615_5 gpc5127 (
      {stage1_23[250], stage1_23[251], stage1_23[252], stage1_23[253], stage1_23[254]},
      {stage1_24[64]},
      {stage1_25[96], stage1_25[97], stage1_25[98], stage1_25[99], stage1_25[100], stage1_25[101]},
      {stage2_27[16],stage2_26[24],stage2_25[51],stage2_24[67],stage2_23[68]}
   );
   gpc615_5 gpc5128 (
      {stage1_23[255], stage1_23[256], stage1_23[257], stage1_23[258], stage1_23[259]},
      {stage1_24[65]},
      {stage1_25[102], stage1_25[103], stage1_25[104], stage1_25[105], stage1_25[106], stage1_25[107]},
      {stage2_27[17],stage2_26[25],stage2_25[52],stage2_24[68],stage2_23[69]}
   );
   gpc615_5 gpc5129 (
      {stage1_23[260], stage1_23[261], stage1_23[262], stage1_23[263], stage1_23[264]},
      {stage1_24[66]},
      {stage1_25[108], stage1_25[109], stage1_25[110], stage1_25[111], stage1_25[112], stage1_25[113]},
      {stage2_27[18],stage2_26[26],stage2_25[53],stage2_24[69],stage2_23[70]}
   );
   gpc615_5 gpc5130 (
      {stage1_23[265], stage1_23[266], stage1_23[267], stage1_23[268], stage1_23[269]},
      {stage1_24[67]},
      {stage1_25[114], stage1_25[115], stage1_25[116], stage1_25[117], stage1_25[118], stage1_25[119]},
      {stage2_27[19],stage2_26[27],stage2_25[54],stage2_24[70],stage2_23[71]}
   );
   gpc615_5 gpc5131 (
      {stage1_23[270], stage1_23[271], stage1_23[272], stage1_23[273], stage1_23[274]},
      {stage1_24[68]},
      {stage1_25[120], stage1_25[121], stage1_25[122], stage1_25[123], stage1_25[124], stage1_25[125]},
      {stage2_27[20],stage2_26[28],stage2_25[55],stage2_24[71],stage2_23[72]}
   );
   gpc615_5 gpc5132 (
      {stage1_23[275], stage1_23[276], stage1_23[277], stage1_23[278], stage1_23[279]},
      {stage1_24[69]},
      {stage1_25[126], stage1_25[127], stage1_25[128], stage1_25[129], stage1_25[130], stage1_25[131]},
      {stage2_27[21],stage2_26[29],stage2_25[56],stage2_24[72],stage2_23[73]}
   );
   gpc615_5 gpc5133 (
      {stage1_23[280], stage1_23[281], stage1_23[282], stage1_23[283], stage1_23[284]},
      {stage1_24[70]},
      {stage1_25[132], stage1_25[133], stage1_25[134], stage1_25[135], stage1_25[136], stage1_25[137]},
      {stage2_27[22],stage2_26[30],stage2_25[57],stage2_24[73],stage2_23[74]}
   );
   gpc615_5 gpc5134 (
      {stage1_23[285], stage1_23[286], 1'b0, 1'b0, 1'b0},
      {stage1_24[71]},
      {stage1_25[138], stage1_25[139], stage1_25[140], stage1_25[141], stage1_25[142], stage1_25[143]},
      {stage2_27[23],stage2_26[31],stage2_25[58],stage2_24[74],stage2_23[75]}
   );
   gpc606_5 gpc5135 (
      {stage1_24[72], stage1_24[73], stage1_24[74], stage1_24[75], stage1_24[76], stage1_24[77]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[24],stage2_26[32],stage2_25[59],stage2_24[75]}
   );
   gpc606_5 gpc5136 (
      {stage1_24[78], stage1_24[79], stage1_24[80], stage1_24[81], stage1_24[82], stage1_24[83]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[25],stage2_26[33],stage2_25[60],stage2_24[76]}
   );
   gpc606_5 gpc5137 (
      {stage1_24[84], stage1_24[85], stage1_24[86], stage1_24[87], stage1_24[88], stage1_24[89]},
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17]},
      {stage2_28[2],stage2_27[26],stage2_26[34],stage2_25[61],stage2_24[77]}
   );
   gpc606_5 gpc5138 (
      {stage1_24[90], stage1_24[91], stage1_24[92], stage1_24[93], stage1_24[94], stage1_24[95]},
      {stage1_26[18], stage1_26[19], stage1_26[20], stage1_26[21], stage1_26[22], stage1_26[23]},
      {stage2_28[3],stage2_27[27],stage2_26[35],stage2_25[62],stage2_24[78]}
   );
   gpc606_5 gpc5139 (
      {stage1_24[96], stage1_24[97], stage1_24[98], stage1_24[99], stage1_24[100], stage1_24[101]},
      {stage1_26[24], stage1_26[25], stage1_26[26], stage1_26[27], stage1_26[28], stage1_26[29]},
      {stage2_28[4],stage2_27[28],stage2_26[36],stage2_25[63],stage2_24[79]}
   );
   gpc606_5 gpc5140 (
      {stage1_24[102], stage1_24[103], stage1_24[104], stage1_24[105], stage1_24[106], stage1_24[107]},
      {stage1_26[30], stage1_26[31], stage1_26[32], stage1_26[33], stage1_26[34], stage1_26[35]},
      {stage2_28[5],stage2_27[29],stage2_26[37],stage2_25[64],stage2_24[80]}
   );
   gpc606_5 gpc5141 (
      {stage1_24[108], stage1_24[109], stage1_24[110], stage1_24[111], stage1_24[112], stage1_24[113]},
      {stage1_26[36], stage1_26[37], stage1_26[38], stage1_26[39], stage1_26[40], stage1_26[41]},
      {stage2_28[6],stage2_27[30],stage2_26[38],stage2_25[65],stage2_24[81]}
   );
   gpc606_5 gpc5142 (
      {stage1_24[114], stage1_24[115], stage1_24[116], stage1_24[117], stage1_24[118], stage1_24[119]},
      {stage1_26[42], stage1_26[43], stage1_26[44], stage1_26[45], stage1_26[46], stage1_26[47]},
      {stage2_28[7],stage2_27[31],stage2_26[39],stage2_25[66],stage2_24[82]}
   );
   gpc606_5 gpc5143 (
      {stage1_24[120], stage1_24[121], stage1_24[122], stage1_24[123], stage1_24[124], stage1_24[125]},
      {stage1_26[48], stage1_26[49], stage1_26[50], stage1_26[51], stage1_26[52], stage1_26[53]},
      {stage2_28[8],stage2_27[32],stage2_26[40],stage2_25[67],stage2_24[83]}
   );
   gpc606_5 gpc5144 (
      {stage1_24[126], stage1_24[127], stage1_24[128], stage1_24[129], stage1_24[130], stage1_24[131]},
      {stage1_26[54], stage1_26[55], stage1_26[56], stage1_26[57], stage1_26[58], stage1_26[59]},
      {stage2_28[9],stage2_27[33],stage2_26[41],stage2_25[68],stage2_24[84]}
   );
   gpc606_5 gpc5145 (
      {stage1_24[132], stage1_24[133], stage1_24[134], stage1_24[135], stage1_24[136], stage1_24[137]},
      {stage1_26[60], stage1_26[61], stage1_26[62], stage1_26[63], stage1_26[64], stage1_26[65]},
      {stage2_28[10],stage2_27[34],stage2_26[42],stage2_25[69],stage2_24[85]}
   );
   gpc606_5 gpc5146 (
      {stage1_24[138], stage1_24[139], stage1_24[140], stage1_24[141], stage1_24[142], stage1_24[143]},
      {stage1_26[66], stage1_26[67], stage1_26[68], stage1_26[69], stage1_26[70], stage1_26[71]},
      {stage2_28[11],stage2_27[35],stage2_26[43],stage2_25[70],stage2_24[86]}
   );
   gpc606_5 gpc5147 (
      {stage1_24[144], stage1_24[145], stage1_24[146], stage1_24[147], stage1_24[148], stage1_24[149]},
      {stage1_26[72], stage1_26[73], stage1_26[74], stage1_26[75], stage1_26[76], stage1_26[77]},
      {stage2_28[12],stage2_27[36],stage2_26[44],stage2_25[71],stage2_24[87]}
   );
   gpc606_5 gpc5148 (
      {stage1_24[150], stage1_24[151], stage1_24[152], stage1_24[153], stage1_24[154], stage1_24[155]},
      {stage1_26[78], stage1_26[79], stage1_26[80], stage1_26[81], stage1_26[82], stage1_26[83]},
      {stage2_28[13],stage2_27[37],stage2_26[45],stage2_25[72],stage2_24[88]}
   );
   gpc606_5 gpc5149 (
      {stage1_24[156], stage1_24[157], stage1_24[158], stage1_24[159], stage1_24[160], stage1_24[161]},
      {stage1_26[84], stage1_26[85], stage1_26[86], stage1_26[87], stage1_26[88], stage1_26[89]},
      {stage2_28[14],stage2_27[38],stage2_26[46],stage2_25[73],stage2_24[89]}
   );
   gpc606_5 gpc5150 (
      {stage1_24[162], stage1_24[163], stage1_24[164], stage1_24[165], stage1_24[166], stage1_24[167]},
      {stage1_26[90], stage1_26[91], stage1_26[92], stage1_26[93], stage1_26[94], stage1_26[95]},
      {stage2_28[15],stage2_27[39],stage2_26[47],stage2_25[74],stage2_24[90]}
   );
   gpc606_5 gpc5151 (
      {stage1_24[168], stage1_24[169], stage1_24[170], stage1_24[171], stage1_24[172], stage1_24[173]},
      {stage1_26[96], stage1_26[97], stage1_26[98], stage1_26[99], stage1_26[100], stage1_26[101]},
      {stage2_28[16],stage2_27[40],stage2_26[48],stage2_25[75],stage2_24[91]}
   );
   gpc606_5 gpc5152 (
      {stage1_24[174], stage1_24[175], stage1_24[176], stage1_24[177], stage1_24[178], stage1_24[179]},
      {stage1_26[102], stage1_26[103], stage1_26[104], stage1_26[105], stage1_26[106], stage1_26[107]},
      {stage2_28[17],stage2_27[41],stage2_26[49],stage2_25[76],stage2_24[92]}
   );
   gpc606_5 gpc5153 (
      {stage1_24[180], stage1_24[181], stage1_24[182], stage1_24[183], stage1_24[184], stage1_24[185]},
      {stage1_26[108], stage1_26[109], stage1_26[110], stage1_26[111], stage1_26[112], stage1_26[113]},
      {stage2_28[18],stage2_27[42],stage2_26[50],stage2_25[77],stage2_24[93]}
   );
   gpc606_5 gpc5154 (
      {stage1_24[186], stage1_24[187], stage1_24[188], stage1_24[189], stage1_24[190], stage1_24[191]},
      {stage1_26[114], stage1_26[115], stage1_26[116], stage1_26[117], stage1_26[118], stage1_26[119]},
      {stage2_28[19],stage2_27[43],stage2_26[51],stage2_25[78],stage2_24[94]}
   );
   gpc606_5 gpc5155 (
      {stage1_24[192], stage1_24[193], stage1_24[194], stage1_24[195], stage1_24[196], stage1_24[197]},
      {stage1_26[120], stage1_26[121], stage1_26[122], stage1_26[123], stage1_26[124], stage1_26[125]},
      {stage2_28[20],stage2_27[44],stage2_26[52],stage2_25[79],stage2_24[95]}
   );
   gpc606_5 gpc5156 (
      {stage1_24[198], stage1_24[199], stage1_24[200], stage1_24[201], stage1_24[202], stage1_24[203]},
      {stage1_26[126], stage1_26[127], stage1_26[128], stage1_26[129], stage1_26[130], stage1_26[131]},
      {stage2_28[21],stage2_27[45],stage2_26[53],stage2_25[80],stage2_24[96]}
   );
   gpc606_5 gpc5157 (
      {stage1_24[204], stage1_24[205], stage1_24[206], stage1_24[207], stage1_24[208], stage1_24[209]},
      {stage1_26[132], stage1_26[133], stage1_26[134], stage1_26[135], stage1_26[136], stage1_26[137]},
      {stage2_28[22],stage2_27[46],stage2_26[54],stage2_25[81],stage2_24[97]}
   );
   gpc207_4 gpc5158 (
      {stage1_25[144], stage1_25[145], stage1_25[146], stage1_25[147], stage1_25[148], stage1_25[149], stage1_25[150]},
      {stage1_27[0], stage1_27[1]},
      {stage2_28[23],stage2_27[47],stage2_26[55],stage2_25[82]}
   );
   gpc606_5 gpc5159 (
      {stage1_25[151], stage1_25[152], stage1_25[153], stage1_25[154], stage1_25[155], stage1_25[156]},
      {stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5], stage1_27[6], stage1_27[7]},
      {stage2_29[0],stage2_28[24],stage2_27[48],stage2_26[56],stage2_25[83]}
   );
   gpc606_5 gpc5160 (
      {stage1_25[157], stage1_25[158], stage1_25[159], stage1_25[160], stage1_25[161], stage1_25[162]},
      {stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11], stage1_27[12], stage1_27[13]},
      {stage2_29[1],stage2_28[25],stage2_27[49],stage2_26[57],stage2_25[84]}
   );
   gpc606_5 gpc5161 (
      {stage1_25[163], stage1_25[164], stage1_25[165], stage1_25[166], stage1_25[167], stage1_25[168]},
      {stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17], stage1_27[18], stage1_27[19]},
      {stage2_29[2],stage2_28[26],stage2_27[50],stage2_26[58],stage2_25[85]}
   );
   gpc606_5 gpc5162 (
      {stage1_25[169], stage1_25[170], stage1_25[171], stage1_25[172], stage1_25[173], stage1_25[174]},
      {stage1_27[20], stage1_27[21], stage1_27[22], stage1_27[23], stage1_27[24], stage1_27[25]},
      {stage2_29[3],stage2_28[27],stage2_27[51],stage2_26[59],stage2_25[86]}
   );
   gpc615_5 gpc5163 (
      {stage1_26[138], stage1_26[139], stage1_26[140], stage1_26[141], stage1_26[142]},
      {stage1_27[26]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[4],stage2_28[28],stage2_27[52],stage2_26[60]}
   );
   gpc615_5 gpc5164 (
      {stage1_26[143], stage1_26[144], stage1_26[145], stage1_26[146], stage1_26[147]},
      {stage1_27[27]},
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11]},
      {stage2_30[1],stage2_29[5],stage2_28[29],stage2_27[53],stage2_26[61]}
   );
   gpc615_5 gpc5165 (
      {stage1_26[148], stage1_26[149], stage1_26[150], stage1_26[151], stage1_26[152]},
      {stage1_27[28]},
      {stage1_28[12], stage1_28[13], stage1_28[14], stage1_28[15], stage1_28[16], stage1_28[17]},
      {stage2_30[2],stage2_29[6],stage2_28[30],stage2_27[54],stage2_26[62]}
   );
   gpc615_5 gpc5166 (
      {stage1_26[153], stage1_26[154], stage1_26[155], stage1_26[156], stage1_26[157]},
      {stage1_27[29]},
      {stage1_28[18], stage1_28[19], stage1_28[20], stage1_28[21], stage1_28[22], stage1_28[23]},
      {stage2_30[3],stage2_29[7],stage2_28[31],stage2_27[55],stage2_26[63]}
   );
   gpc615_5 gpc5167 (
      {stage1_26[158], stage1_26[159], stage1_26[160], stage1_26[161], stage1_26[162]},
      {stage1_27[30]},
      {stage1_28[24], stage1_28[25], stage1_28[26], stage1_28[27], stage1_28[28], stage1_28[29]},
      {stage2_30[4],stage2_29[8],stage2_28[32],stage2_27[56],stage2_26[64]}
   );
   gpc615_5 gpc5168 (
      {stage1_26[163], stage1_26[164], stage1_26[165], stage1_26[166], stage1_26[167]},
      {stage1_27[31]},
      {stage1_28[30], stage1_28[31], stage1_28[32], stage1_28[33], stage1_28[34], stage1_28[35]},
      {stage2_30[5],stage2_29[9],stage2_28[33],stage2_27[57],stage2_26[65]}
   );
   gpc615_5 gpc5169 (
      {stage1_26[168], stage1_26[169], stage1_26[170], stage1_26[171], stage1_26[172]},
      {stage1_27[32]},
      {stage1_28[36], stage1_28[37], stage1_28[38], stage1_28[39], stage1_28[40], stage1_28[41]},
      {stage2_30[6],stage2_29[10],stage2_28[34],stage2_27[58],stage2_26[66]}
   );
   gpc615_5 gpc5170 (
      {stage1_26[173], stage1_26[174], stage1_26[175], stage1_26[176], stage1_26[177]},
      {stage1_27[33]},
      {stage1_28[42], stage1_28[43], stage1_28[44], stage1_28[45], stage1_28[46], stage1_28[47]},
      {stage2_30[7],stage2_29[11],stage2_28[35],stage2_27[59],stage2_26[67]}
   );
   gpc615_5 gpc5171 (
      {stage1_26[178], stage1_26[179], stage1_26[180], stage1_26[181], stage1_26[182]},
      {stage1_27[34]},
      {stage1_28[48], stage1_28[49], stage1_28[50], stage1_28[51], stage1_28[52], stage1_28[53]},
      {stage2_30[8],stage2_29[12],stage2_28[36],stage2_27[60],stage2_26[68]}
   );
   gpc615_5 gpc5172 (
      {stage1_26[183], stage1_26[184], stage1_26[185], stage1_26[186], stage1_26[187]},
      {stage1_27[35]},
      {stage1_28[54], stage1_28[55], stage1_28[56], stage1_28[57], stage1_28[58], stage1_28[59]},
      {stage2_30[9],stage2_29[13],stage2_28[37],stage2_27[61],stage2_26[69]}
   );
   gpc615_5 gpc5173 (
      {stage1_26[188], stage1_26[189], stage1_26[190], stage1_26[191], stage1_26[192]},
      {stage1_27[36]},
      {stage1_28[60], stage1_28[61], stage1_28[62], stage1_28[63], stage1_28[64], stage1_28[65]},
      {stage2_30[10],stage2_29[14],stage2_28[38],stage2_27[62],stage2_26[70]}
   );
   gpc615_5 gpc5174 (
      {stage1_26[193], stage1_26[194], stage1_26[195], stage1_26[196], stage1_26[197]},
      {stage1_27[37]},
      {stage1_28[66], stage1_28[67], stage1_28[68], stage1_28[69], stage1_28[70], stage1_28[71]},
      {stage2_30[11],stage2_29[15],stage2_28[39],stage2_27[63],stage2_26[71]}
   );
   gpc615_5 gpc5175 (
      {stage1_26[198], stage1_26[199], stage1_26[200], stage1_26[201], stage1_26[202]},
      {stage1_27[38]},
      {stage1_28[72], stage1_28[73], stage1_28[74], stage1_28[75], stage1_28[76], stage1_28[77]},
      {stage2_30[12],stage2_29[16],stage2_28[40],stage2_27[64],stage2_26[72]}
   );
   gpc615_5 gpc5176 (
      {stage1_26[203], stage1_26[204], stage1_26[205], stage1_26[206], stage1_26[207]},
      {stage1_27[39]},
      {stage1_28[78], stage1_28[79], stage1_28[80], stage1_28[81], stage1_28[82], stage1_28[83]},
      {stage2_30[13],stage2_29[17],stage2_28[41],stage2_27[65],stage2_26[73]}
   );
   gpc615_5 gpc5177 (
      {stage1_26[208], stage1_26[209], stage1_26[210], stage1_26[211], stage1_26[212]},
      {stage1_27[40]},
      {stage1_28[84], stage1_28[85], stage1_28[86], stage1_28[87], stage1_28[88], stage1_28[89]},
      {stage2_30[14],stage2_29[18],stage2_28[42],stage2_27[66],stage2_26[74]}
   );
   gpc615_5 gpc5178 (
      {stage1_26[213], stage1_26[214], stage1_26[215], stage1_26[216], stage1_26[217]},
      {stage1_27[41]},
      {stage1_28[90], stage1_28[91], stage1_28[92], stage1_28[93], stage1_28[94], stage1_28[95]},
      {stage2_30[15],stage2_29[19],stage2_28[43],stage2_27[67],stage2_26[75]}
   );
   gpc615_5 gpc5179 (
      {stage1_26[218], stage1_26[219], stage1_26[220], stage1_26[221], stage1_26[222]},
      {stage1_27[42]},
      {stage1_28[96], stage1_28[97], stage1_28[98], stage1_28[99], stage1_28[100], stage1_28[101]},
      {stage2_30[16],stage2_29[20],stage2_28[44],stage2_27[68],stage2_26[76]}
   );
   gpc615_5 gpc5180 (
      {stage1_26[223], stage1_26[224], stage1_26[225], stage1_26[226], stage1_26[227]},
      {stage1_27[43]},
      {stage1_28[102], stage1_28[103], stage1_28[104], stage1_28[105], stage1_28[106], stage1_28[107]},
      {stage2_30[17],stage2_29[21],stage2_28[45],stage2_27[69],stage2_26[77]}
   );
   gpc615_5 gpc5181 (
      {stage1_26[228], stage1_26[229], stage1_26[230], stage1_26[231], stage1_26[232]},
      {stage1_27[44]},
      {stage1_28[108], stage1_28[109], stage1_28[110], stage1_28[111], stage1_28[112], stage1_28[113]},
      {stage2_30[18],stage2_29[22],stage2_28[46],stage2_27[70],stage2_26[78]}
   );
   gpc615_5 gpc5182 (
      {stage1_26[233], stage1_26[234], stage1_26[235], stage1_26[236], stage1_26[237]},
      {stage1_27[45]},
      {stage1_28[114], stage1_28[115], stage1_28[116], stage1_28[117], stage1_28[118], stage1_28[119]},
      {stage2_30[19],stage2_29[23],stage2_28[47],stage2_27[71],stage2_26[79]}
   );
   gpc615_5 gpc5183 (
      {stage1_26[238], stage1_26[239], stage1_26[240], stage1_26[241], stage1_26[242]},
      {stage1_27[46]},
      {stage1_28[120], stage1_28[121], stage1_28[122], stage1_28[123], stage1_28[124], stage1_28[125]},
      {stage2_30[20],stage2_29[24],stage2_28[48],stage2_27[72],stage2_26[80]}
   );
   gpc615_5 gpc5184 (
      {stage1_26[243], stage1_26[244], stage1_26[245], stage1_26[246], stage1_26[247]},
      {stage1_27[47]},
      {stage1_28[126], stage1_28[127], stage1_28[128], stage1_28[129], stage1_28[130], stage1_28[131]},
      {stage2_30[21],stage2_29[25],stage2_28[49],stage2_27[73],stage2_26[81]}
   );
   gpc615_5 gpc5185 (
      {stage1_27[48], stage1_27[49], stage1_27[50], stage1_27[51], stage1_27[52]},
      {stage1_28[132]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[22],stage2_29[26],stage2_28[50],stage2_27[74]}
   );
   gpc615_5 gpc5186 (
      {stage1_27[53], stage1_27[54], stage1_27[55], stage1_27[56], stage1_27[57]},
      {stage1_28[133]},
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage2_31[1],stage2_30[23],stage2_29[27],stage2_28[51],stage2_27[75]}
   );
   gpc615_5 gpc5187 (
      {stage1_27[58], stage1_27[59], stage1_27[60], stage1_27[61], stage1_27[62]},
      {stage1_28[134]},
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17]},
      {stage2_31[2],stage2_30[24],stage2_29[28],stage2_28[52],stage2_27[76]}
   );
   gpc615_5 gpc5188 (
      {stage1_27[63], stage1_27[64], stage1_27[65], stage1_27[66], stage1_27[67]},
      {stage1_28[135]},
      {stage1_29[18], stage1_29[19], stage1_29[20], stage1_29[21], stage1_29[22], stage1_29[23]},
      {stage2_31[3],stage2_30[25],stage2_29[29],stage2_28[53],stage2_27[77]}
   );
   gpc615_5 gpc5189 (
      {stage1_27[68], stage1_27[69], stage1_27[70], stage1_27[71], stage1_27[72]},
      {stage1_28[136]},
      {stage1_29[24], stage1_29[25], stage1_29[26], stage1_29[27], stage1_29[28], stage1_29[29]},
      {stage2_31[4],stage2_30[26],stage2_29[30],stage2_28[54],stage2_27[78]}
   );
   gpc615_5 gpc5190 (
      {stage1_27[73], stage1_27[74], stage1_27[75], stage1_27[76], stage1_27[77]},
      {stage1_28[137]},
      {stage1_29[30], stage1_29[31], stage1_29[32], stage1_29[33], stage1_29[34], stage1_29[35]},
      {stage2_31[5],stage2_30[27],stage2_29[31],stage2_28[55],stage2_27[79]}
   );
   gpc615_5 gpc5191 (
      {stage1_27[78], stage1_27[79], stage1_27[80], stage1_27[81], stage1_27[82]},
      {stage1_28[138]},
      {stage1_29[36], stage1_29[37], stage1_29[38], stage1_29[39], stage1_29[40], stage1_29[41]},
      {stage2_31[6],stage2_30[28],stage2_29[32],stage2_28[56],stage2_27[80]}
   );
   gpc615_5 gpc5192 (
      {stage1_27[83], stage1_27[84], stage1_27[85], stage1_27[86], stage1_27[87]},
      {stage1_28[139]},
      {stage1_29[42], stage1_29[43], stage1_29[44], stage1_29[45], stage1_29[46], stage1_29[47]},
      {stage2_31[7],stage2_30[29],stage2_29[33],stage2_28[57],stage2_27[81]}
   );
   gpc615_5 gpc5193 (
      {stage1_27[88], stage1_27[89], stage1_27[90], stage1_27[91], stage1_27[92]},
      {stage1_28[140]},
      {stage1_29[48], stage1_29[49], stage1_29[50], stage1_29[51], stage1_29[52], stage1_29[53]},
      {stage2_31[8],stage2_30[30],stage2_29[34],stage2_28[58],stage2_27[82]}
   );
   gpc615_5 gpc5194 (
      {stage1_27[93], stage1_27[94], stage1_27[95], stage1_27[96], stage1_27[97]},
      {stage1_28[141]},
      {stage1_29[54], stage1_29[55], stage1_29[56], stage1_29[57], stage1_29[58], stage1_29[59]},
      {stage2_31[9],stage2_30[31],stage2_29[35],stage2_28[59],stage2_27[83]}
   );
   gpc615_5 gpc5195 (
      {stage1_27[98], stage1_27[99], stage1_27[100], stage1_27[101], stage1_27[102]},
      {stage1_28[142]},
      {stage1_29[60], stage1_29[61], stage1_29[62], stage1_29[63], stage1_29[64], stage1_29[65]},
      {stage2_31[10],stage2_30[32],stage2_29[36],stage2_28[60],stage2_27[84]}
   );
   gpc615_5 gpc5196 (
      {stage1_27[103], stage1_27[104], stage1_27[105], stage1_27[106], stage1_27[107]},
      {stage1_28[143]},
      {stage1_29[66], stage1_29[67], stage1_29[68], stage1_29[69], stage1_29[70], stage1_29[71]},
      {stage2_31[11],stage2_30[33],stage2_29[37],stage2_28[61],stage2_27[85]}
   );
   gpc615_5 gpc5197 (
      {stage1_27[108], stage1_27[109], stage1_27[110], stage1_27[111], stage1_27[112]},
      {stage1_28[144]},
      {stage1_29[72], stage1_29[73], stage1_29[74], stage1_29[75], stage1_29[76], stage1_29[77]},
      {stage2_31[12],stage2_30[34],stage2_29[38],stage2_28[62],stage2_27[86]}
   );
   gpc615_5 gpc5198 (
      {stage1_27[113], stage1_27[114], stage1_27[115], stage1_27[116], stage1_27[117]},
      {stage1_28[145]},
      {stage1_29[78], stage1_29[79], stage1_29[80], stage1_29[81], stage1_29[82], stage1_29[83]},
      {stage2_31[13],stage2_30[35],stage2_29[39],stage2_28[63],stage2_27[87]}
   );
   gpc615_5 gpc5199 (
      {stage1_27[118], stage1_27[119], stage1_27[120], stage1_27[121], stage1_27[122]},
      {stage1_28[146]},
      {stage1_29[84], stage1_29[85], stage1_29[86], stage1_29[87], stage1_29[88], stage1_29[89]},
      {stage2_31[14],stage2_30[36],stage2_29[40],stage2_28[64],stage2_27[88]}
   );
   gpc615_5 gpc5200 (
      {stage1_27[123], stage1_27[124], stage1_27[125], stage1_27[126], stage1_27[127]},
      {stage1_28[147]},
      {stage1_29[90], stage1_29[91], stage1_29[92], stage1_29[93], stage1_29[94], stage1_29[95]},
      {stage2_31[15],stage2_30[37],stage2_29[41],stage2_28[65],stage2_27[89]}
   );
   gpc615_5 gpc5201 (
      {stage1_27[128], stage1_27[129], stage1_27[130], stage1_27[131], stage1_27[132]},
      {stage1_28[148]},
      {stage1_29[96], stage1_29[97], stage1_29[98], stage1_29[99], stage1_29[100], stage1_29[101]},
      {stage2_31[16],stage2_30[38],stage2_29[42],stage2_28[66],stage2_27[90]}
   );
   gpc615_5 gpc5202 (
      {stage1_27[133], stage1_27[134], stage1_27[135], stage1_27[136], stage1_27[137]},
      {stage1_28[149]},
      {stage1_29[102], stage1_29[103], stage1_29[104], stage1_29[105], stage1_29[106], stage1_29[107]},
      {stage2_31[17],stage2_30[39],stage2_29[43],stage2_28[67],stage2_27[91]}
   );
   gpc615_5 gpc5203 (
      {stage1_27[138], stage1_27[139], stage1_27[140], stage1_27[141], stage1_27[142]},
      {stage1_28[150]},
      {stage1_29[108], stage1_29[109], stage1_29[110], stage1_29[111], stage1_29[112], stage1_29[113]},
      {stage2_31[18],stage2_30[40],stage2_29[44],stage2_28[68],stage2_27[92]}
   );
   gpc615_5 gpc5204 (
      {stage1_27[143], stage1_27[144], stage1_27[145], stage1_27[146], stage1_27[147]},
      {stage1_28[151]},
      {stage1_29[114], stage1_29[115], stage1_29[116], stage1_29[117], stage1_29[118], stage1_29[119]},
      {stage2_31[19],stage2_30[41],stage2_29[45],stage2_28[69],stage2_27[93]}
   );
   gpc615_5 gpc5205 (
      {stage1_27[148], stage1_27[149], stage1_27[150], stage1_27[151], stage1_27[152]},
      {stage1_28[152]},
      {stage1_29[120], stage1_29[121], stage1_29[122], stage1_29[123], stage1_29[124], stage1_29[125]},
      {stage2_31[20],stage2_30[42],stage2_29[46],stage2_28[70],stage2_27[94]}
   );
   gpc615_5 gpc5206 (
      {stage1_27[153], stage1_27[154], stage1_27[155], stage1_27[156], stage1_27[157]},
      {stage1_28[153]},
      {stage1_29[126], stage1_29[127], stage1_29[128], stage1_29[129], stage1_29[130], stage1_29[131]},
      {stage2_31[21],stage2_30[43],stage2_29[47],stage2_28[71],stage2_27[95]}
   );
   gpc615_5 gpc5207 (
      {stage1_27[158], stage1_27[159], stage1_27[160], stage1_27[161], stage1_27[162]},
      {stage1_28[154]},
      {stage1_29[132], stage1_29[133], stage1_29[134], stage1_29[135], stage1_29[136], stage1_29[137]},
      {stage2_31[22],stage2_30[44],stage2_29[48],stage2_28[72],stage2_27[96]}
   );
   gpc615_5 gpc5208 (
      {stage1_27[163], stage1_27[164], stage1_27[165], stage1_27[166], stage1_27[167]},
      {stage1_28[155]},
      {stage1_29[138], stage1_29[139], stage1_29[140], stage1_29[141], stage1_29[142], stage1_29[143]},
      {stage2_31[23],stage2_30[45],stage2_29[49],stage2_28[73],stage2_27[97]}
   );
   gpc615_5 gpc5209 (
      {stage1_27[168], stage1_27[169], stage1_27[170], stage1_27[171], stage1_27[172]},
      {stage1_28[156]},
      {stage1_29[144], stage1_29[145], stage1_29[146], stage1_29[147], stage1_29[148], stage1_29[149]},
      {stage2_31[24],stage2_30[46],stage2_29[50],stage2_28[74],stage2_27[98]}
   );
   gpc615_5 gpc5210 (
      {stage1_27[173], stage1_27[174], stage1_27[175], stage1_27[176], stage1_27[177]},
      {stage1_28[157]},
      {stage1_29[150], stage1_29[151], stage1_29[152], stage1_29[153], stage1_29[154], stage1_29[155]},
      {stage2_31[25],stage2_30[47],stage2_29[51],stage2_28[75],stage2_27[99]}
   );
   gpc615_5 gpc5211 (
      {stage1_27[178], stage1_27[179], stage1_27[180], stage1_27[181], stage1_27[182]},
      {stage1_28[158]},
      {stage1_29[156], stage1_29[157], stage1_29[158], stage1_29[159], stage1_29[160], stage1_29[161]},
      {stage2_31[26],stage2_30[48],stage2_29[52],stage2_28[76],stage2_27[100]}
   );
   gpc615_5 gpc5212 (
      {stage1_27[183], stage1_27[184], stage1_27[185], stage1_27[186], stage1_27[187]},
      {stage1_28[159]},
      {stage1_29[162], stage1_29[163], stage1_29[164], stage1_29[165], stage1_29[166], stage1_29[167]},
      {stage2_31[27],stage2_30[49],stage2_29[53],stage2_28[77],stage2_27[101]}
   );
   gpc615_5 gpc5213 (
      {stage1_27[188], stage1_27[189], stage1_27[190], stage1_27[191], stage1_27[192]},
      {stage1_28[160]},
      {stage1_29[168], stage1_29[169], stage1_29[170], stage1_29[171], stage1_29[172], stage1_29[173]},
      {stage2_31[28],stage2_30[50],stage2_29[54],stage2_28[78],stage2_27[102]}
   );
   gpc615_5 gpc5214 (
      {stage1_27[193], stage1_27[194], stage1_27[195], stage1_27[196], stage1_27[197]},
      {stage1_28[161]},
      {stage1_29[174], stage1_29[175], stage1_29[176], stage1_29[177], stage1_29[178], stage1_29[179]},
      {stage2_31[29],stage2_30[51],stage2_29[55],stage2_28[79],stage2_27[103]}
   );
   gpc615_5 gpc5215 (
      {stage1_27[198], stage1_27[199], stage1_27[200], stage1_27[201], stage1_27[202]},
      {stage1_28[162]},
      {stage1_29[180], stage1_29[181], stage1_29[182], stage1_29[183], stage1_29[184], stage1_29[185]},
      {stage2_31[30],stage2_30[52],stage2_29[56],stage2_28[80],stage2_27[104]}
   );
   gpc615_5 gpc5216 (
      {stage1_27[203], stage1_27[204], stage1_27[205], 1'b0, 1'b0},
      {stage1_28[163]},
      {stage1_29[186], stage1_29[187], stage1_29[188], stage1_29[189], stage1_29[190], stage1_29[191]},
      {stage2_31[31],stage2_30[53],stage2_29[57],stage2_28[81],stage2_27[105]}
   );
   gpc606_5 gpc5217 (
      {stage1_28[164], stage1_28[165], stage1_28[166], stage1_28[167], stage1_28[168], stage1_28[169]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[32],stage2_30[54],stage2_29[58],stage2_28[82]}
   );
   gpc606_5 gpc5218 (
      {stage1_28[170], stage1_28[171], stage1_28[172], stage1_28[173], stage1_28[174], stage1_28[175]},
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage2_32[1],stage2_31[33],stage2_30[55],stage2_29[59],stage2_28[83]}
   );
   gpc606_5 gpc5219 (
      {stage1_28[176], stage1_28[177], stage1_28[178], stage1_28[179], stage1_28[180], stage1_28[181]},
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage2_32[2],stage2_31[34],stage2_30[56],stage2_29[60],stage2_28[84]}
   );
   gpc606_5 gpc5220 (
      {stage1_28[182], stage1_28[183], stage1_28[184], stage1_28[185], stage1_28[186], stage1_28[187]},
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22], stage1_30[23]},
      {stage2_32[3],stage2_31[35],stage2_30[57],stage2_29[61],stage2_28[85]}
   );
   gpc606_5 gpc5221 (
      {stage1_28[188], stage1_28[189], stage1_28[190], stage1_28[191], stage1_28[192], stage1_28[193]},
      {stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27], stage1_30[28], stage1_30[29]},
      {stage2_32[4],stage2_31[36],stage2_30[58],stage2_29[62],stage2_28[86]}
   );
   gpc606_5 gpc5222 (
      {stage1_28[194], stage1_28[195], stage1_28[196], stage1_28[197], stage1_28[198], stage1_28[199]},
      {stage1_30[30], stage1_30[31], stage1_30[32], stage1_30[33], stage1_30[34], stage1_30[35]},
      {stage2_32[5],stage2_31[37],stage2_30[59],stage2_29[63],stage2_28[87]}
   );
   gpc606_5 gpc5223 (
      {stage1_28[200], stage1_28[201], stage1_28[202], stage1_28[203], stage1_28[204], stage1_28[205]},
      {stage1_30[36], stage1_30[37], stage1_30[38], stage1_30[39], stage1_30[40], stage1_30[41]},
      {stage2_32[6],stage2_31[38],stage2_30[60],stage2_29[64],stage2_28[88]}
   );
   gpc606_5 gpc5224 (
      {stage1_28[206], stage1_28[207], stage1_28[208], stage1_28[209], stage1_28[210], stage1_28[211]},
      {stage1_30[42], stage1_30[43], stage1_30[44], stage1_30[45], stage1_30[46], stage1_30[47]},
      {stage2_32[7],stage2_31[39],stage2_30[61],stage2_29[65],stage2_28[89]}
   );
   gpc606_5 gpc5225 (
      {stage1_28[212], stage1_28[213], stage1_28[214], stage1_28[215], stage1_28[216], stage1_28[217]},
      {stage1_30[48], stage1_30[49], stage1_30[50], stage1_30[51], stage1_30[52], stage1_30[53]},
      {stage2_32[8],stage2_31[40],stage2_30[62],stage2_29[66],stage2_28[90]}
   );
   gpc606_5 gpc5226 (
      {stage1_28[218], stage1_28[219], stage1_28[220], stage1_28[221], stage1_28[222], stage1_28[223]},
      {stage1_30[54], stage1_30[55], stage1_30[56], stage1_30[57], stage1_30[58], stage1_30[59]},
      {stage2_32[9],stage2_31[41],stage2_30[63],stage2_29[67],stage2_28[91]}
   );
   gpc1163_5 gpc5227 (
      {stage1_29[192], stage1_29[193], stage1_29[194]},
      {stage1_30[60], stage1_30[61], stage1_30[62], stage1_30[63], stage1_30[64], stage1_30[65]},
      {stage1_31[0]},
      {stage1_32[0]},
      {stage2_33[0],stage2_32[10],stage2_31[42],stage2_30[64],stage2_29[68]}
   );
   gpc1163_5 gpc5228 (
      {stage1_29[195], stage1_29[196], stage1_29[197]},
      {stage1_30[66], stage1_30[67], stage1_30[68], stage1_30[69], stage1_30[70], stage1_30[71]},
      {stage1_31[1]},
      {stage1_32[1]},
      {stage2_33[1],stage2_32[11],stage2_31[43],stage2_30[65],stage2_29[69]}
   );
   gpc1163_5 gpc5229 (
      {stage1_29[198], stage1_29[199], stage1_29[200]},
      {stage1_30[72], stage1_30[73], stage1_30[74], stage1_30[75], stage1_30[76], stage1_30[77]},
      {stage1_31[2]},
      {stage1_32[2]},
      {stage2_33[2],stage2_32[12],stage2_31[44],stage2_30[66],stage2_29[70]}
   );
   gpc1163_5 gpc5230 (
      {stage1_29[201], stage1_29[202], stage1_29[203]},
      {stage1_30[78], stage1_30[79], stage1_30[80], stage1_30[81], stage1_30[82], stage1_30[83]},
      {stage1_31[3]},
      {stage1_32[3]},
      {stage2_33[3],stage2_32[13],stage2_31[45],stage2_30[67],stage2_29[71]}
   );
   gpc606_5 gpc5231 (
      {stage1_29[204], stage1_29[205], stage1_29[206], stage1_29[207], stage1_29[208], stage1_29[209]},
      {stage1_31[4], stage1_31[5], stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9]},
      {stage2_33[4],stage2_32[14],stage2_31[46],stage2_30[68],stage2_29[72]}
   );
   gpc606_5 gpc5232 (
      {stage1_29[210], stage1_29[211], stage1_29[212], stage1_29[213], stage1_29[214], stage1_29[215]},
      {stage1_31[10], stage1_31[11], stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15]},
      {stage2_33[5],stage2_32[15],stage2_31[47],stage2_30[69],stage2_29[73]}
   );
   gpc606_5 gpc5233 (
      {stage1_30[84], stage1_30[85], stage1_30[86], stage1_30[87], stage1_30[88], stage1_30[89]},
      {stage1_32[4], stage1_32[5], stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9]},
      {stage2_34[0],stage2_33[6],stage2_32[16],stage2_31[48],stage2_30[70]}
   );
   gpc615_5 gpc5234 (
      {stage1_30[90], stage1_30[91], stage1_30[92], stage1_30[93], stage1_30[94]},
      {stage1_31[16]},
      {stage1_32[10], stage1_32[11], stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15]},
      {stage2_34[1],stage2_33[7],stage2_32[17],stage2_31[49],stage2_30[71]}
   );
   gpc615_5 gpc5235 (
      {stage1_30[95], stage1_30[96], stage1_30[97], stage1_30[98], stage1_30[99]},
      {stage1_31[17]},
      {stage1_32[16], stage1_32[17], stage1_32[18], stage1_32[19], stage1_32[20], stage1_32[21]},
      {stage2_34[2],stage2_33[8],stage2_32[18],stage2_31[50],stage2_30[72]}
   );
   gpc615_5 gpc5236 (
      {stage1_30[100], stage1_30[101], stage1_30[102], stage1_30[103], stage1_30[104]},
      {stage1_31[18]},
      {stage1_32[22], stage1_32[23], stage1_32[24], stage1_32[25], stage1_32[26], stage1_32[27]},
      {stage2_34[3],stage2_33[9],stage2_32[19],stage2_31[51],stage2_30[73]}
   );
   gpc615_5 gpc5237 (
      {stage1_30[105], stage1_30[106], stage1_30[107], stage1_30[108], stage1_30[109]},
      {stage1_31[19]},
      {stage1_32[28], stage1_32[29], stage1_32[30], stage1_32[31], stage1_32[32], stage1_32[33]},
      {stage2_34[4],stage2_33[10],stage2_32[20],stage2_31[52],stage2_30[74]}
   );
   gpc615_5 gpc5238 (
      {stage1_30[110], stage1_30[111], stage1_30[112], stage1_30[113], stage1_30[114]},
      {stage1_31[20]},
      {stage1_32[34], stage1_32[35], stage1_32[36], stage1_32[37], stage1_32[38], stage1_32[39]},
      {stage2_34[5],stage2_33[11],stage2_32[21],stage2_31[53],stage2_30[75]}
   );
   gpc615_5 gpc5239 (
      {stage1_30[115], stage1_30[116], stage1_30[117], stage1_30[118], stage1_30[119]},
      {stage1_31[21]},
      {stage1_32[40], stage1_32[41], stage1_32[42], stage1_32[43], stage1_32[44], stage1_32[45]},
      {stage2_34[6],stage2_33[12],stage2_32[22],stage2_31[54],stage2_30[76]}
   );
   gpc615_5 gpc5240 (
      {stage1_30[120], stage1_30[121], stage1_30[122], stage1_30[123], stage1_30[124]},
      {stage1_31[22]},
      {stage1_32[46], stage1_32[47], stage1_32[48], stage1_32[49], stage1_32[50], stage1_32[51]},
      {stage2_34[7],stage2_33[13],stage2_32[23],stage2_31[55],stage2_30[77]}
   );
   gpc615_5 gpc5241 (
      {stage1_30[125], stage1_30[126], stage1_30[127], stage1_30[128], stage1_30[129]},
      {stage1_31[23]},
      {stage1_32[52], stage1_32[53], stage1_32[54], stage1_32[55], stage1_32[56], stage1_32[57]},
      {stage2_34[8],stage2_33[14],stage2_32[24],stage2_31[56],stage2_30[78]}
   );
   gpc615_5 gpc5242 (
      {stage1_30[130], stage1_30[131], stage1_30[132], stage1_30[133], stage1_30[134]},
      {stage1_31[24]},
      {stage1_32[58], stage1_32[59], stage1_32[60], stage1_32[61], stage1_32[62], stage1_32[63]},
      {stage2_34[9],stage2_33[15],stage2_32[25],stage2_31[57],stage2_30[79]}
   );
   gpc615_5 gpc5243 (
      {stage1_30[135], stage1_30[136], stage1_30[137], stage1_30[138], stage1_30[139]},
      {stage1_31[25]},
      {stage1_32[64], stage1_32[65], stage1_32[66], stage1_32[67], stage1_32[68], stage1_32[69]},
      {stage2_34[10],stage2_33[16],stage2_32[26],stage2_31[58],stage2_30[80]}
   );
   gpc615_5 gpc5244 (
      {stage1_30[140], stage1_30[141], stage1_30[142], stage1_30[143], stage1_30[144]},
      {stage1_31[26]},
      {stage1_32[70], stage1_32[71], stage1_32[72], stage1_32[73], stage1_32[74], stage1_32[75]},
      {stage2_34[11],stage2_33[17],stage2_32[27],stage2_31[59],stage2_30[81]}
   );
   gpc615_5 gpc5245 (
      {stage1_30[145], stage1_30[146], stage1_30[147], stage1_30[148], stage1_30[149]},
      {stage1_31[27]},
      {stage1_32[76], stage1_32[77], stage1_32[78], stage1_32[79], stage1_32[80], stage1_32[81]},
      {stage2_34[12],stage2_33[18],stage2_32[28],stage2_31[60],stage2_30[82]}
   );
   gpc615_5 gpc5246 (
      {stage1_30[150], stage1_30[151], stage1_30[152], stage1_30[153], stage1_30[154]},
      {stage1_31[28]},
      {stage1_32[82], stage1_32[83], stage1_32[84], stage1_32[85], stage1_32[86], stage1_32[87]},
      {stage2_34[13],stage2_33[19],stage2_32[29],stage2_31[61],stage2_30[83]}
   );
   gpc615_5 gpc5247 (
      {stage1_30[155], stage1_30[156], stage1_30[157], stage1_30[158], stage1_30[159]},
      {stage1_31[29]},
      {stage1_32[88], stage1_32[89], stage1_32[90], stage1_32[91], stage1_32[92], stage1_32[93]},
      {stage2_34[14],stage2_33[20],stage2_32[30],stage2_31[62],stage2_30[84]}
   );
   gpc1163_5 gpc5248 (
      {stage1_31[30], stage1_31[31], stage1_31[32]},
      {stage1_32[94], stage1_32[95], stage1_32[96], stage1_32[97], stage1_32[98], stage1_32[99]},
      {stage1_33[0]},
      {stage1_34[0]},
      {stage2_35[0],stage2_34[15],stage2_33[21],stage2_32[31],stage2_31[63]}
   );
   gpc606_5 gpc5249 (
      {stage1_31[33], stage1_31[34], stage1_31[35], stage1_31[36], stage1_31[37], stage1_31[38]},
      {stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5], stage1_33[6]},
      {stage2_35[1],stage2_34[16],stage2_33[22],stage2_32[32],stage2_31[64]}
   );
   gpc606_5 gpc5250 (
      {stage1_31[39], stage1_31[40], stage1_31[41], stage1_31[42], stage1_31[43], stage1_31[44]},
      {stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11], stage1_33[12]},
      {stage2_35[2],stage2_34[17],stage2_33[23],stage2_32[33],stage2_31[65]}
   );
   gpc606_5 gpc5251 (
      {stage1_31[45], stage1_31[46], stage1_31[47], stage1_31[48], stage1_31[49], stage1_31[50]},
      {stage1_33[13], stage1_33[14], stage1_33[15], stage1_33[16], stage1_33[17], stage1_33[18]},
      {stage2_35[3],stage2_34[18],stage2_33[24],stage2_32[34],stage2_31[66]}
   );
   gpc606_5 gpc5252 (
      {stage1_31[51], stage1_31[52], stage1_31[53], stage1_31[54], stage1_31[55], stage1_31[56]},
      {stage1_33[19], stage1_33[20], stage1_33[21], stage1_33[22], stage1_33[23], stage1_33[24]},
      {stage2_35[4],stage2_34[19],stage2_33[25],stage2_32[35],stage2_31[67]}
   );
   gpc606_5 gpc5253 (
      {stage1_31[57], stage1_31[58], stage1_31[59], stage1_31[60], stage1_31[61], stage1_31[62]},
      {stage1_33[25], stage1_33[26], stage1_33[27], stage1_33[28], stage1_33[29], stage1_33[30]},
      {stage2_35[5],stage2_34[20],stage2_33[26],stage2_32[36],stage2_31[68]}
   );
   gpc606_5 gpc5254 (
      {stage1_31[63], stage1_31[64], stage1_31[65], stage1_31[66], stage1_31[67], stage1_31[68]},
      {stage1_33[31], stage1_33[32], stage1_33[33], stage1_33[34], stage1_33[35], stage1_33[36]},
      {stage2_35[6],stage2_34[21],stage2_33[27],stage2_32[37],stage2_31[69]}
   );
   gpc606_5 gpc5255 (
      {stage1_31[69], stage1_31[70], stage1_31[71], stage1_31[72], stage1_31[73], stage1_31[74]},
      {stage1_33[37], stage1_33[38], stage1_33[39], stage1_33[40], stage1_33[41], stage1_33[42]},
      {stage2_35[7],stage2_34[22],stage2_33[28],stage2_32[38],stage2_31[70]}
   );
   gpc606_5 gpc5256 (
      {stage1_31[75], stage1_31[76], stage1_31[77], stage1_31[78], stage1_31[79], stage1_31[80]},
      {stage1_33[43], stage1_33[44], stage1_33[45], stage1_33[46], stage1_33[47], stage1_33[48]},
      {stage2_35[8],stage2_34[23],stage2_33[29],stage2_32[39],stage2_31[71]}
   );
   gpc606_5 gpc5257 (
      {stage1_31[81], stage1_31[82], stage1_31[83], stage1_31[84], stage1_31[85], stage1_31[86]},
      {stage1_33[49], stage1_33[50], stage1_33[51], stage1_33[52], stage1_33[53], stage1_33[54]},
      {stage2_35[9],stage2_34[24],stage2_33[30],stage2_32[40],stage2_31[72]}
   );
   gpc606_5 gpc5258 (
      {stage1_31[87], stage1_31[88], stage1_31[89], stage1_31[90], stage1_31[91], stage1_31[92]},
      {stage1_33[55], stage1_33[56], stage1_33[57], stage1_33[58], stage1_33[59], stage1_33[60]},
      {stage2_35[10],stage2_34[25],stage2_33[31],stage2_32[41],stage2_31[73]}
   );
   gpc606_5 gpc5259 (
      {stage1_31[93], stage1_31[94], stage1_31[95], stage1_31[96], stage1_31[97], stage1_31[98]},
      {stage1_33[61], stage1_33[62], stage1_33[63], stage1_33[64], stage1_33[65], stage1_33[66]},
      {stage2_35[11],stage2_34[26],stage2_33[32],stage2_32[42],stage2_31[74]}
   );
   gpc606_5 gpc5260 (
      {stage1_31[99], stage1_31[100], stage1_31[101], stage1_31[102], stage1_31[103], stage1_31[104]},
      {stage1_33[67], stage1_33[68], stage1_33[69], stage1_33[70], stage1_33[71], stage1_33[72]},
      {stage2_35[12],stage2_34[27],stage2_33[33],stage2_32[43],stage2_31[75]}
   );
   gpc615_5 gpc5261 (
      {stage1_31[105], stage1_31[106], stage1_31[107], stage1_31[108], stage1_31[109]},
      {stage1_32[100]},
      {stage1_33[73], stage1_33[74], stage1_33[75], stage1_33[76], stage1_33[77], stage1_33[78]},
      {stage2_35[13],stage2_34[28],stage2_33[34],stage2_32[44],stage2_31[76]}
   );
   gpc615_5 gpc5262 (
      {stage1_31[110], stage1_31[111], stage1_31[112], stage1_31[113], stage1_31[114]},
      {stage1_32[101]},
      {stage1_33[79], stage1_33[80], stage1_33[81], stage1_33[82], stage1_33[83], stage1_33[84]},
      {stage2_35[14],stage2_34[29],stage2_33[35],stage2_32[45],stage2_31[77]}
   );
   gpc615_5 gpc5263 (
      {stage1_31[115], stage1_31[116], stage1_31[117], stage1_31[118], stage1_31[119]},
      {stage1_32[102]},
      {stage1_33[85], stage1_33[86], stage1_33[87], stage1_33[88], stage1_33[89], stage1_33[90]},
      {stage2_35[15],stage2_34[30],stage2_33[36],stage2_32[46],stage2_31[78]}
   );
   gpc615_5 gpc5264 (
      {stage1_31[120], stage1_31[121], stage1_31[122], stage1_31[123], stage1_31[124]},
      {stage1_32[103]},
      {stage1_33[91], stage1_33[92], stage1_33[93], stage1_33[94], stage1_33[95], stage1_33[96]},
      {stage2_35[16],stage2_34[31],stage2_33[37],stage2_32[47],stage2_31[79]}
   );
   gpc615_5 gpc5265 (
      {stage1_31[125], stage1_31[126], stage1_31[127], stage1_31[128], stage1_31[129]},
      {stage1_32[104]},
      {stage1_33[97], stage1_33[98], stage1_33[99], stage1_33[100], stage1_33[101], stage1_33[102]},
      {stage2_35[17],stage2_34[32],stage2_33[38],stage2_32[48],stage2_31[80]}
   );
   gpc615_5 gpc5266 (
      {stage1_31[130], stage1_31[131], stage1_31[132], stage1_31[133], stage1_31[134]},
      {stage1_32[105]},
      {stage1_33[103], stage1_33[104], stage1_33[105], stage1_33[106], stage1_33[107], stage1_33[108]},
      {stage2_35[18],stage2_34[33],stage2_33[39],stage2_32[49],stage2_31[81]}
   );
   gpc615_5 gpc5267 (
      {stage1_31[135], stage1_31[136], stage1_31[137], stage1_31[138], stage1_31[139]},
      {stage1_32[106]},
      {stage1_33[109], stage1_33[110], stage1_33[111], stage1_33[112], stage1_33[113], stage1_33[114]},
      {stage2_35[19],stage2_34[34],stage2_33[40],stage2_32[50],stage2_31[82]}
   );
   gpc615_5 gpc5268 (
      {stage1_31[140], stage1_31[141], stage1_31[142], stage1_31[143], stage1_31[144]},
      {stage1_32[107]},
      {stage1_33[115], stage1_33[116], stage1_33[117], stage1_33[118], stage1_33[119], stage1_33[120]},
      {stage2_35[20],stage2_34[35],stage2_33[41],stage2_32[51],stage2_31[83]}
   );
   gpc615_5 gpc5269 (
      {stage1_31[145], stage1_31[146], stage1_31[147], stage1_31[148], stage1_31[149]},
      {stage1_32[108]},
      {stage1_33[121], stage1_33[122], stage1_33[123], stage1_33[124], stage1_33[125], stage1_33[126]},
      {stage2_35[21],stage2_34[36],stage2_33[42],stage2_32[52],stage2_31[84]}
   );
   gpc615_5 gpc5270 (
      {stage1_31[150], stage1_31[151], stage1_31[152], stage1_31[153], stage1_31[154]},
      {stage1_32[109]},
      {stage1_33[127], stage1_33[128], stage1_33[129], stage1_33[130], stage1_33[131], stage1_33[132]},
      {stage2_35[22],stage2_34[37],stage2_33[43],stage2_32[53],stage2_31[85]}
   );
   gpc615_5 gpc5271 (
      {stage1_31[155], stage1_31[156], stage1_31[157], stage1_31[158], stage1_31[159]},
      {stage1_32[110]},
      {stage1_33[133], stage1_33[134], stage1_33[135], stage1_33[136], stage1_33[137], stage1_33[138]},
      {stage2_35[23],stage2_34[38],stage2_33[44],stage2_32[54],stage2_31[86]}
   );
   gpc615_5 gpc5272 (
      {stage1_31[160], stage1_31[161], stage1_31[162], stage1_31[163], stage1_31[164]},
      {stage1_32[111]},
      {stage1_33[139], stage1_33[140], stage1_33[141], stage1_33[142], stage1_33[143], stage1_33[144]},
      {stage2_35[24],stage2_34[39],stage2_33[45],stage2_32[55],stage2_31[87]}
   );
   gpc615_5 gpc5273 (
      {stage1_31[165], stage1_31[166], stage1_31[167], stage1_31[168], stage1_31[169]},
      {stage1_32[112]},
      {stage1_33[145], stage1_33[146], stage1_33[147], stage1_33[148], stage1_33[149], stage1_33[150]},
      {stage2_35[25],stage2_34[40],stage2_33[46],stage2_32[56],stage2_31[88]}
   );
   gpc615_5 gpc5274 (
      {stage1_31[170], stage1_31[171], stage1_31[172], stage1_31[173], stage1_31[174]},
      {stage1_32[113]},
      {stage1_33[151], stage1_33[152], stage1_33[153], stage1_33[154], stage1_33[155], stage1_33[156]},
      {stage2_35[26],stage2_34[41],stage2_33[47],stage2_32[57],stage2_31[89]}
   );
   gpc615_5 gpc5275 (
      {stage1_31[175], stage1_31[176], stage1_31[177], stage1_31[178], stage1_31[179]},
      {stage1_32[114]},
      {stage1_33[157], stage1_33[158], stage1_33[159], stage1_33[160], stage1_33[161], stage1_33[162]},
      {stage2_35[27],stage2_34[42],stage2_33[48],stage2_32[58],stage2_31[90]}
   );
   gpc615_5 gpc5276 (
      {stage1_31[180], stage1_31[181], stage1_31[182], stage1_31[183], stage1_31[184]},
      {stage1_32[115]},
      {stage1_33[163], stage1_33[164], stage1_33[165], stage1_33[166], stage1_33[167], stage1_33[168]},
      {stage2_35[28],stage2_34[43],stage2_33[49],stage2_32[59],stage2_31[91]}
   );
   gpc615_5 gpc5277 (
      {stage1_31[185], stage1_31[186], stage1_31[187], stage1_31[188], stage1_31[189]},
      {stage1_32[116]},
      {stage1_33[169], stage1_33[170], stage1_33[171], stage1_33[172], stage1_33[173], stage1_33[174]},
      {stage2_35[29],stage2_34[44],stage2_33[50],stage2_32[60],stage2_31[92]}
   );
   gpc615_5 gpc5278 (
      {stage1_31[190], stage1_31[191], stage1_31[192], stage1_31[193], stage1_31[194]},
      {stage1_32[117]},
      {stage1_33[175], stage1_33[176], stage1_33[177], stage1_33[178], stage1_33[179], stage1_33[180]},
      {stage2_35[30],stage2_34[45],stage2_33[51],stage2_32[61],stage2_31[93]}
   );
   gpc615_5 gpc5279 (
      {stage1_31[195], stage1_31[196], stage1_31[197], stage1_31[198], stage1_31[199]},
      {stage1_32[118]},
      {stage1_33[181], stage1_33[182], stage1_33[183], stage1_33[184], stage1_33[185], stage1_33[186]},
      {stage2_35[31],stage2_34[46],stage2_33[52],stage2_32[62],stage2_31[94]}
   );
   gpc615_5 gpc5280 (
      {stage1_31[200], stage1_31[201], stage1_31[202], stage1_31[203], stage1_31[204]},
      {stage1_32[119]},
      {stage1_33[187], stage1_33[188], stage1_33[189], stage1_33[190], stage1_33[191], stage1_33[192]},
      {stage2_35[32],stage2_34[47],stage2_33[53],stage2_32[63],stage2_31[95]}
   );
   gpc615_5 gpc5281 (
      {stage1_31[205], stage1_31[206], stage1_31[207], stage1_31[208], stage1_31[209]},
      {stage1_32[120]},
      {stage1_33[193], stage1_33[194], stage1_33[195], stage1_33[196], stage1_33[197], stage1_33[198]},
      {stage2_35[33],stage2_34[48],stage2_33[54],stage2_32[64],stage2_31[96]}
   );
   gpc615_5 gpc5282 (
      {stage1_31[210], stage1_31[211], stage1_31[212], stage1_31[213], stage1_31[214]},
      {stage1_32[121]},
      {stage1_33[199], stage1_33[200], stage1_33[201], stage1_33[202], stage1_33[203], stage1_33[204]},
      {stage2_35[34],stage2_34[49],stage2_33[55],stage2_32[65],stage2_31[97]}
   );
   gpc615_5 gpc5283 (
      {stage1_31[215], stage1_31[216], stage1_31[217], 1'b0, 1'b0},
      {stage1_32[122]},
      {stage1_33[205], stage1_33[206], stage1_33[207], stage1_33[208], stage1_33[209], stage1_33[210]},
      {stage2_35[35],stage2_34[50],stage2_33[56],stage2_32[66],stage2_31[98]}
   );
   gpc606_5 gpc5284 (
      {stage1_32[123], stage1_32[124], stage1_32[125], stage1_32[126], stage1_32[127], stage1_32[128]},
      {stage1_34[1], stage1_34[2], stage1_34[3], stage1_34[4], stage1_34[5], stage1_34[6]},
      {stage2_36[0],stage2_35[36],stage2_34[51],stage2_33[57],stage2_32[67]}
   );
   gpc606_5 gpc5285 (
      {stage1_32[129], stage1_32[130], stage1_32[131], stage1_32[132], stage1_32[133], stage1_32[134]},
      {stage1_34[7], stage1_34[8], stage1_34[9], stage1_34[10], stage1_34[11], stage1_34[12]},
      {stage2_36[1],stage2_35[37],stage2_34[52],stage2_33[58],stage2_32[68]}
   );
   gpc606_5 gpc5286 (
      {stage1_32[135], stage1_32[136], stage1_32[137], stage1_32[138], stage1_32[139], stage1_32[140]},
      {stage1_34[13], stage1_34[14], stage1_34[15], stage1_34[16], stage1_34[17], stage1_34[18]},
      {stage2_36[2],stage2_35[38],stage2_34[53],stage2_33[59],stage2_32[69]}
   );
   gpc606_5 gpc5287 (
      {stage1_32[141], stage1_32[142], stage1_32[143], stage1_32[144], stage1_32[145], stage1_32[146]},
      {stage1_34[19], stage1_34[20], stage1_34[21], stage1_34[22], stage1_34[23], stage1_34[24]},
      {stage2_36[3],stage2_35[39],stage2_34[54],stage2_33[60],stage2_32[70]}
   );
   gpc606_5 gpc5288 (
      {stage1_32[147], stage1_32[148], stage1_32[149], stage1_32[150], stage1_32[151], stage1_32[152]},
      {stage1_34[25], stage1_34[26], stage1_34[27], stage1_34[28], stage1_34[29], stage1_34[30]},
      {stage2_36[4],stage2_35[40],stage2_34[55],stage2_33[61],stage2_32[71]}
   );
   gpc606_5 gpc5289 (
      {stage1_32[153], stage1_32[154], stage1_32[155], stage1_32[156], stage1_32[157], stage1_32[158]},
      {stage1_34[31], stage1_34[32], stage1_34[33], stage1_34[34], stage1_34[35], stage1_34[36]},
      {stage2_36[5],stage2_35[41],stage2_34[56],stage2_33[62],stage2_32[72]}
   );
   gpc606_5 gpc5290 (
      {stage1_32[159], stage1_32[160], stage1_32[161], stage1_32[162], stage1_32[163], stage1_32[164]},
      {stage1_34[37], stage1_34[38], stage1_34[39], stage1_34[40], stage1_34[41], stage1_34[42]},
      {stage2_36[6],stage2_35[42],stage2_34[57],stage2_33[63],stage2_32[73]}
   );
   gpc606_5 gpc5291 (
      {stage1_32[165], stage1_32[166], stage1_32[167], stage1_32[168], stage1_32[169], stage1_32[170]},
      {stage1_34[43], stage1_34[44], stage1_34[45], stage1_34[46], stage1_34[47], stage1_34[48]},
      {stage2_36[7],stage2_35[43],stage2_34[58],stage2_33[64],stage2_32[74]}
   );
   gpc606_5 gpc5292 (
      {stage1_32[171], stage1_32[172], stage1_32[173], stage1_32[174], stage1_32[175], stage1_32[176]},
      {stage1_34[49], stage1_34[50], stage1_34[51], stage1_34[52], stage1_34[53], stage1_34[54]},
      {stage2_36[8],stage2_35[44],stage2_34[59],stage2_33[65],stage2_32[75]}
   );
   gpc606_5 gpc5293 (
      {stage1_32[177], stage1_32[178], stage1_32[179], stage1_32[180], stage1_32[181], stage1_32[182]},
      {stage1_34[55], stage1_34[56], stage1_34[57], stage1_34[58], stage1_34[59], stage1_34[60]},
      {stage2_36[9],stage2_35[45],stage2_34[60],stage2_33[66],stage2_32[76]}
   );
   gpc606_5 gpc5294 (
      {stage1_32[183], stage1_32[184], stage1_32[185], stage1_32[186], stage1_32[187], stage1_32[188]},
      {stage1_34[61], stage1_34[62], stage1_34[63], stage1_34[64], stage1_34[65], stage1_34[66]},
      {stage2_36[10],stage2_35[46],stage2_34[61],stage2_33[67],stage2_32[77]}
   );
   gpc2116_5 gpc5295 (
      {stage1_33[211], stage1_33[212], stage1_33[213], stage1_33[214], stage1_33[215], stage1_33[216]},
      {stage1_34[67]},
      {stage1_35[0]},
      {stage1_36[0], stage1_36[1]},
      {stage2_37[0],stage2_36[11],stage2_35[47],stage2_34[62],stage2_33[68]}
   );
   gpc606_5 gpc5296 (
      {stage1_33[217], stage1_33[218], stage1_33[219], stage1_33[220], stage1_33[221], stage1_33[222]},
      {stage1_35[1], stage1_35[2], stage1_35[3], stage1_35[4], stage1_35[5], stage1_35[6]},
      {stage2_37[1],stage2_36[12],stage2_35[48],stage2_34[63],stage2_33[69]}
   );
   gpc606_5 gpc5297 (
      {stage1_33[223], stage1_33[224], stage1_33[225], stage1_33[226], stage1_33[227], stage1_33[228]},
      {stage1_35[7], stage1_35[8], stage1_35[9], stage1_35[10], stage1_35[11], stage1_35[12]},
      {stage2_37[2],stage2_36[13],stage2_35[49],stage2_34[64],stage2_33[70]}
   );
   gpc606_5 gpc5298 (
      {stage1_33[229], stage1_33[230], stage1_33[231], stage1_33[232], stage1_33[233], stage1_33[234]},
      {stage1_35[13], stage1_35[14], stage1_35[15], stage1_35[16], stage1_35[17], stage1_35[18]},
      {stage2_37[3],stage2_36[14],stage2_35[50],stage2_34[65],stage2_33[71]}
   );
   gpc606_5 gpc5299 (
      {stage1_33[235], stage1_33[236], stage1_33[237], stage1_33[238], stage1_33[239], stage1_33[240]},
      {stage1_35[19], stage1_35[20], stage1_35[21], stage1_35[22], stage1_35[23], stage1_35[24]},
      {stage2_37[4],stage2_36[15],stage2_35[51],stage2_34[66],stage2_33[72]}
   );
   gpc606_5 gpc5300 (
      {stage1_33[241], stage1_33[242], stage1_33[243], stage1_33[244], stage1_33[245], stage1_33[246]},
      {stage1_35[25], stage1_35[26], stage1_35[27], stage1_35[28], stage1_35[29], stage1_35[30]},
      {stage2_37[5],stage2_36[16],stage2_35[52],stage2_34[67],stage2_33[73]}
   );
   gpc606_5 gpc5301 (
      {stage1_33[247], stage1_33[248], stage1_33[249], stage1_33[250], stage1_33[251], stage1_33[252]},
      {stage1_35[31], stage1_35[32], stage1_35[33], stage1_35[34], stage1_35[35], stage1_35[36]},
      {stage2_37[6],stage2_36[17],stage2_35[53],stage2_34[68],stage2_33[74]}
   );
   gpc606_5 gpc5302 (
      {stage1_33[253], stage1_33[254], stage1_33[255], stage1_33[256], stage1_33[257], stage1_33[258]},
      {stage1_35[37], stage1_35[38], stage1_35[39], stage1_35[40], stage1_35[41], stage1_35[42]},
      {stage2_37[7],stage2_36[18],stage2_35[54],stage2_34[69],stage2_33[75]}
   );
   gpc606_5 gpc5303 (
      {stage1_34[68], stage1_34[69], stage1_34[70], stage1_34[71], stage1_34[72], stage1_34[73]},
      {stage1_36[2], stage1_36[3], stage1_36[4], stage1_36[5], stage1_36[6], stage1_36[7]},
      {stage2_38[0],stage2_37[8],stage2_36[19],stage2_35[55],stage2_34[70]}
   );
   gpc606_5 gpc5304 (
      {stage1_34[74], stage1_34[75], stage1_34[76], stage1_34[77], stage1_34[78], stage1_34[79]},
      {stage1_36[8], stage1_36[9], stage1_36[10], stage1_36[11], stage1_36[12], stage1_36[13]},
      {stage2_38[1],stage2_37[9],stage2_36[20],stage2_35[56],stage2_34[71]}
   );
   gpc606_5 gpc5305 (
      {stage1_34[80], stage1_34[81], stage1_34[82], stage1_34[83], stage1_34[84], stage1_34[85]},
      {stage1_36[14], stage1_36[15], stage1_36[16], stage1_36[17], stage1_36[18], stage1_36[19]},
      {stage2_38[2],stage2_37[10],stage2_36[21],stage2_35[57],stage2_34[72]}
   );
   gpc606_5 gpc5306 (
      {stage1_34[86], stage1_34[87], stage1_34[88], stage1_34[89], stage1_34[90], stage1_34[91]},
      {stage1_36[20], stage1_36[21], stage1_36[22], stage1_36[23], stage1_36[24], stage1_36[25]},
      {stage2_38[3],stage2_37[11],stage2_36[22],stage2_35[58],stage2_34[73]}
   );
   gpc606_5 gpc5307 (
      {stage1_34[92], stage1_34[93], stage1_34[94], stage1_34[95], stage1_34[96], stage1_34[97]},
      {stage1_36[26], stage1_36[27], stage1_36[28], stage1_36[29], stage1_36[30], stage1_36[31]},
      {stage2_38[4],stage2_37[12],stage2_36[23],stage2_35[59],stage2_34[74]}
   );
   gpc606_5 gpc5308 (
      {stage1_34[98], stage1_34[99], stage1_34[100], stage1_34[101], stage1_34[102], stage1_34[103]},
      {stage1_36[32], stage1_36[33], stage1_36[34], stage1_36[35], stage1_36[36], stage1_36[37]},
      {stage2_38[5],stage2_37[13],stage2_36[24],stage2_35[60],stage2_34[75]}
   );
   gpc606_5 gpc5309 (
      {stage1_34[104], stage1_34[105], stage1_34[106], stage1_34[107], stage1_34[108], stage1_34[109]},
      {stage1_36[38], stage1_36[39], stage1_36[40], stage1_36[41], stage1_36[42], stage1_36[43]},
      {stage2_38[6],stage2_37[14],stage2_36[25],stage2_35[61],stage2_34[76]}
   );
   gpc606_5 gpc5310 (
      {stage1_34[110], stage1_34[111], stage1_34[112], stage1_34[113], stage1_34[114], stage1_34[115]},
      {stage1_36[44], stage1_36[45], stage1_36[46], stage1_36[47], stage1_36[48], stage1_36[49]},
      {stage2_38[7],stage2_37[15],stage2_36[26],stage2_35[62],stage2_34[77]}
   );
   gpc606_5 gpc5311 (
      {stage1_34[116], stage1_34[117], stage1_34[118], stage1_34[119], stage1_34[120], stage1_34[121]},
      {stage1_36[50], stage1_36[51], stage1_36[52], stage1_36[53], stage1_36[54], stage1_36[55]},
      {stage2_38[8],stage2_37[16],stage2_36[27],stage2_35[63],stage2_34[78]}
   );
   gpc606_5 gpc5312 (
      {stage1_34[122], stage1_34[123], stage1_34[124], stage1_34[125], stage1_34[126], stage1_34[127]},
      {stage1_36[56], stage1_36[57], stage1_36[58], stage1_36[59], stage1_36[60], stage1_36[61]},
      {stage2_38[9],stage2_37[17],stage2_36[28],stage2_35[64],stage2_34[79]}
   );
   gpc606_5 gpc5313 (
      {stage1_34[128], stage1_34[129], stage1_34[130], stage1_34[131], stage1_34[132], stage1_34[133]},
      {stage1_36[62], stage1_36[63], stage1_36[64], stage1_36[65], stage1_36[66], stage1_36[67]},
      {stage2_38[10],stage2_37[18],stage2_36[29],stage2_35[65],stage2_34[80]}
   );
   gpc606_5 gpc5314 (
      {stage1_34[134], stage1_34[135], stage1_34[136], stage1_34[137], stage1_34[138], stage1_34[139]},
      {stage1_36[68], stage1_36[69], stage1_36[70], stage1_36[71], stage1_36[72], stage1_36[73]},
      {stage2_38[11],stage2_37[19],stage2_36[30],stage2_35[66],stage2_34[81]}
   );
   gpc615_5 gpc5315 (
      {stage1_35[43], stage1_35[44], stage1_35[45], stage1_35[46], stage1_35[47]},
      {stage1_36[74]},
      {stage1_37[0], stage1_37[1], stage1_37[2], stage1_37[3], stage1_37[4], stage1_37[5]},
      {stage2_39[0],stage2_38[12],stage2_37[20],stage2_36[31],stage2_35[67]}
   );
   gpc615_5 gpc5316 (
      {stage1_35[48], stage1_35[49], stage1_35[50], stage1_35[51], stage1_35[52]},
      {stage1_36[75]},
      {stage1_37[6], stage1_37[7], stage1_37[8], stage1_37[9], stage1_37[10], stage1_37[11]},
      {stage2_39[1],stage2_38[13],stage2_37[21],stage2_36[32],stage2_35[68]}
   );
   gpc615_5 gpc5317 (
      {stage1_35[53], stage1_35[54], stage1_35[55], stage1_35[56], stage1_35[57]},
      {stage1_36[76]},
      {stage1_37[12], stage1_37[13], stage1_37[14], stage1_37[15], stage1_37[16], stage1_37[17]},
      {stage2_39[2],stage2_38[14],stage2_37[22],stage2_36[33],stage2_35[69]}
   );
   gpc615_5 gpc5318 (
      {stage1_35[58], stage1_35[59], stage1_35[60], stage1_35[61], stage1_35[62]},
      {stage1_36[77]},
      {stage1_37[18], stage1_37[19], stage1_37[20], stage1_37[21], stage1_37[22], stage1_37[23]},
      {stage2_39[3],stage2_38[15],stage2_37[23],stage2_36[34],stage2_35[70]}
   );
   gpc615_5 gpc5319 (
      {stage1_35[63], stage1_35[64], stage1_35[65], stage1_35[66], stage1_35[67]},
      {stage1_36[78]},
      {stage1_37[24], stage1_37[25], stage1_37[26], stage1_37[27], stage1_37[28], stage1_37[29]},
      {stage2_39[4],stage2_38[16],stage2_37[24],stage2_36[35],stage2_35[71]}
   );
   gpc615_5 gpc5320 (
      {stage1_35[68], stage1_35[69], stage1_35[70], stage1_35[71], stage1_35[72]},
      {stage1_36[79]},
      {stage1_37[30], stage1_37[31], stage1_37[32], stage1_37[33], stage1_37[34], stage1_37[35]},
      {stage2_39[5],stage2_38[17],stage2_37[25],stage2_36[36],stage2_35[72]}
   );
   gpc615_5 gpc5321 (
      {stage1_35[73], stage1_35[74], stage1_35[75], stage1_35[76], stage1_35[77]},
      {stage1_36[80]},
      {stage1_37[36], stage1_37[37], stage1_37[38], stage1_37[39], stage1_37[40], stage1_37[41]},
      {stage2_39[6],stage2_38[18],stage2_37[26],stage2_36[37],stage2_35[73]}
   );
   gpc615_5 gpc5322 (
      {stage1_35[78], stage1_35[79], stage1_35[80], stage1_35[81], stage1_35[82]},
      {stage1_36[81]},
      {stage1_37[42], stage1_37[43], stage1_37[44], stage1_37[45], stage1_37[46], stage1_37[47]},
      {stage2_39[7],stage2_38[19],stage2_37[27],stage2_36[38],stage2_35[74]}
   );
   gpc615_5 gpc5323 (
      {stage1_35[83], stage1_35[84], stage1_35[85], stage1_35[86], stage1_35[87]},
      {stage1_36[82]},
      {stage1_37[48], stage1_37[49], stage1_37[50], stage1_37[51], stage1_37[52], stage1_37[53]},
      {stage2_39[8],stage2_38[20],stage2_37[28],stage2_36[39],stage2_35[75]}
   );
   gpc615_5 gpc5324 (
      {stage1_35[88], stage1_35[89], stage1_35[90], stage1_35[91], stage1_35[92]},
      {stage1_36[83]},
      {stage1_37[54], stage1_37[55], stage1_37[56], stage1_37[57], stage1_37[58], stage1_37[59]},
      {stage2_39[9],stage2_38[21],stage2_37[29],stage2_36[40],stage2_35[76]}
   );
   gpc615_5 gpc5325 (
      {stage1_35[93], stage1_35[94], stage1_35[95], stage1_35[96], stage1_35[97]},
      {stage1_36[84]},
      {stage1_37[60], stage1_37[61], stage1_37[62], stage1_37[63], stage1_37[64], stage1_37[65]},
      {stage2_39[10],stage2_38[22],stage2_37[30],stage2_36[41],stage2_35[77]}
   );
   gpc615_5 gpc5326 (
      {stage1_35[98], stage1_35[99], stage1_35[100], stage1_35[101], stage1_35[102]},
      {stage1_36[85]},
      {stage1_37[66], stage1_37[67], stage1_37[68], stage1_37[69], stage1_37[70], stage1_37[71]},
      {stage2_39[11],stage2_38[23],stage2_37[31],stage2_36[42],stage2_35[78]}
   );
   gpc615_5 gpc5327 (
      {stage1_35[103], stage1_35[104], stage1_35[105], stage1_35[106], stage1_35[107]},
      {stage1_36[86]},
      {stage1_37[72], stage1_37[73], stage1_37[74], stage1_37[75], stage1_37[76], stage1_37[77]},
      {stage2_39[12],stage2_38[24],stage2_37[32],stage2_36[43],stage2_35[79]}
   );
   gpc615_5 gpc5328 (
      {stage1_35[108], stage1_35[109], stage1_35[110], stage1_35[111], stage1_35[112]},
      {stage1_36[87]},
      {stage1_37[78], stage1_37[79], stage1_37[80], stage1_37[81], stage1_37[82], stage1_37[83]},
      {stage2_39[13],stage2_38[25],stage2_37[33],stage2_36[44],stage2_35[80]}
   );
   gpc615_5 gpc5329 (
      {stage1_35[113], stage1_35[114], stage1_35[115], stage1_35[116], stage1_35[117]},
      {stage1_36[88]},
      {stage1_37[84], stage1_37[85], stage1_37[86], stage1_37[87], stage1_37[88], stage1_37[89]},
      {stage2_39[14],stage2_38[26],stage2_37[34],stage2_36[45],stage2_35[81]}
   );
   gpc615_5 gpc5330 (
      {stage1_35[118], stage1_35[119], stage1_35[120], stage1_35[121], stage1_35[122]},
      {stage1_36[89]},
      {stage1_37[90], stage1_37[91], stage1_37[92], stage1_37[93], stage1_37[94], stage1_37[95]},
      {stage2_39[15],stage2_38[27],stage2_37[35],stage2_36[46],stage2_35[82]}
   );
   gpc615_5 gpc5331 (
      {stage1_35[123], stage1_35[124], stage1_35[125], stage1_35[126], stage1_35[127]},
      {stage1_36[90]},
      {stage1_37[96], stage1_37[97], stage1_37[98], stage1_37[99], stage1_37[100], stage1_37[101]},
      {stage2_39[16],stage2_38[28],stage2_37[36],stage2_36[47],stage2_35[83]}
   );
   gpc615_5 gpc5332 (
      {stage1_35[128], stage1_35[129], stage1_35[130], stage1_35[131], stage1_35[132]},
      {stage1_36[91]},
      {stage1_37[102], stage1_37[103], stage1_37[104], stage1_37[105], stage1_37[106], stage1_37[107]},
      {stage2_39[17],stage2_38[29],stage2_37[37],stage2_36[48],stage2_35[84]}
   );
   gpc615_5 gpc5333 (
      {stage1_35[133], stage1_35[134], stage1_35[135], stage1_35[136], stage1_35[137]},
      {stage1_36[92]},
      {stage1_37[108], stage1_37[109], stage1_37[110], stage1_37[111], stage1_37[112], stage1_37[113]},
      {stage2_39[18],stage2_38[30],stage2_37[38],stage2_36[49],stage2_35[85]}
   );
   gpc615_5 gpc5334 (
      {stage1_35[138], stage1_35[139], stage1_35[140], stage1_35[141], stage1_35[142]},
      {stage1_36[93]},
      {stage1_37[114], stage1_37[115], stage1_37[116], stage1_37[117], stage1_37[118], stage1_37[119]},
      {stage2_39[19],stage2_38[31],stage2_37[39],stage2_36[50],stage2_35[86]}
   );
   gpc615_5 gpc5335 (
      {stage1_35[143], stage1_35[144], stage1_35[145], stage1_35[146], stage1_35[147]},
      {stage1_36[94]},
      {stage1_37[120], stage1_37[121], stage1_37[122], stage1_37[123], stage1_37[124], stage1_37[125]},
      {stage2_39[20],stage2_38[32],stage2_37[40],stage2_36[51],stage2_35[87]}
   );
   gpc615_5 gpc5336 (
      {stage1_35[148], stage1_35[149], stage1_35[150], stage1_35[151], stage1_35[152]},
      {stage1_36[95]},
      {stage1_37[126], stage1_37[127], stage1_37[128], stage1_37[129], stage1_37[130], stage1_37[131]},
      {stage2_39[21],stage2_38[33],stage2_37[41],stage2_36[52],stage2_35[88]}
   );
   gpc615_5 gpc5337 (
      {stage1_35[153], stage1_35[154], stage1_35[155], stage1_35[156], stage1_35[157]},
      {stage1_36[96]},
      {stage1_37[132], stage1_37[133], stage1_37[134], stage1_37[135], stage1_37[136], stage1_37[137]},
      {stage2_39[22],stage2_38[34],stage2_37[42],stage2_36[53],stage2_35[89]}
   );
   gpc615_5 gpc5338 (
      {stage1_35[158], stage1_35[159], stage1_35[160], stage1_35[161], stage1_35[162]},
      {stage1_36[97]},
      {stage1_37[138], stage1_37[139], stage1_37[140], stage1_37[141], stage1_37[142], stage1_37[143]},
      {stage2_39[23],stage2_38[35],stage2_37[43],stage2_36[54],stage2_35[90]}
   );
   gpc615_5 gpc5339 (
      {stage1_35[163], stage1_35[164], stage1_35[165], stage1_35[166], stage1_35[167]},
      {stage1_36[98]},
      {stage1_37[144], stage1_37[145], stage1_37[146], stage1_37[147], stage1_37[148], stage1_37[149]},
      {stage2_39[24],stage2_38[36],stage2_37[44],stage2_36[55],stage2_35[91]}
   );
   gpc615_5 gpc5340 (
      {stage1_35[168], stage1_35[169], stage1_35[170], stage1_35[171], stage1_35[172]},
      {stage1_36[99]},
      {stage1_37[150], stage1_37[151], stage1_37[152], stage1_37[153], stage1_37[154], stage1_37[155]},
      {stage2_39[25],stage2_38[37],stage2_37[45],stage2_36[56],stage2_35[92]}
   );
   gpc615_5 gpc5341 (
      {stage1_35[173], stage1_35[174], stage1_35[175], stage1_35[176], stage1_35[177]},
      {stage1_36[100]},
      {stage1_37[156], stage1_37[157], stage1_37[158], stage1_37[159], stage1_37[160], stage1_37[161]},
      {stage2_39[26],stage2_38[38],stage2_37[46],stage2_36[57],stage2_35[93]}
   );
   gpc1406_5 gpc5342 (
      {stage1_36[101], stage1_36[102], stage1_36[103], stage1_36[104], stage1_36[105], stage1_36[106]},
      {stage1_38[0], stage1_38[1], stage1_38[2], stage1_38[3]},
      {stage1_39[0]},
      {stage2_40[0],stage2_39[27],stage2_38[39],stage2_37[47],stage2_36[58]}
   );
   gpc606_5 gpc5343 (
      {stage1_36[107], stage1_36[108], stage1_36[109], stage1_36[110], stage1_36[111], stage1_36[112]},
      {stage1_38[4], stage1_38[5], stage1_38[6], stage1_38[7], stage1_38[8], stage1_38[9]},
      {stage2_40[1],stage2_39[28],stage2_38[40],stage2_37[48],stage2_36[59]}
   );
   gpc606_5 gpc5344 (
      {stage1_36[113], stage1_36[114], stage1_36[115], stage1_36[116], stage1_36[117], stage1_36[118]},
      {stage1_38[10], stage1_38[11], stage1_38[12], stage1_38[13], stage1_38[14], stage1_38[15]},
      {stage2_40[2],stage2_39[29],stage2_38[41],stage2_37[49],stage2_36[60]}
   );
   gpc606_5 gpc5345 (
      {stage1_36[119], stage1_36[120], stage1_36[121], stage1_36[122], stage1_36[123], stage1_36[124]},
      {stage1_38[16], stage1_38[17], stage1_38[18], stage1_38[19], stage1_38[20], stage1_38[21]},
      {stage2_40[3],stage2_39[30],stage2_38[42],stage2_37[50],stage2_36[61]}
   );
   gpc606_5 gpc5346 (
      {stage1_36[125], stage1_36[126], stage1_36[127], stage1_36[128], stage1_36[129], stage1_36[130]},
      {stage1_38[22], stage1_38[23], stage1_38[24], stage1_38[25], stage1_38[26], stage1_38[27]},
      {stage2_40[4],stage2_39[31],stage2_38[43],stage2_37[51],stage2_36[62]}
   );
   gpc606_5 gpc5347 (
      {stage1_36[131], stage1_36[132], stage1_36[133], stage1_36[134], stage1_36[135], stage1_36[136]},
      {stage1_38[28], stage1_38[29], stage1_38[30], stage1_38[31], stage1_38[32], stage1_38[33]},
      {stage2_40[5],stage2_39[32],stage2_38[44],stage2_37[52],stage2_36[63]}
   );
   gpc606_5 gpc5348 (
      {stage1_36[137], stage1_36[138], stage1_36[139], stage1_36[140], stage1_36[141], stage1_36[142]},
      {stage1_38[34], stage1_38[35], stage1_38[36], stage1_38[37], stage1_38[38], stage1_38[39]},
      {stage2_40[6],stage2_39[33],stage2_38[45],stage2_37[53],stage2_36[64]}
   );
   gpc606_5 gpc5349 (
      {stage1_36[143], stage1_36[144], stage1_36[145], stage1_36[146], stage1_36[147], stage1_36[148]},
      {stage1_38[40], stage1_38[41], stage1_38[42], stage1_38[43], stage1_38[44], stage1_38[45]},
      {stage2_40[7],stage2_39[34],stage2_38[46],stage2_37[54],stage2_36[65]}
   );
   gpc606_5 gpc5350 (
      {stage1_36[149], stage1_36[150], stage1_36[151], stage1_36[152], stage1_36[153], stage1_36[154]},
      {stage1_38[46], stage1_38[47], stage1_38[48], stage1_38[49], stage1_38[50], stage1_38[51]},
      {stage2_40[8],stage2_39[35],stage2_38[47],stage2_37[55],stage2_36[66]}
   );
   gpc606_5 gpc5351 (
      {stage1_36[155], stage1_36[156], stage1_36[157], stage1_36[158], stage1_36[159], stage1_36[160]},
      {stage1_38[52], stage1_38[53], stage1_38[54], stage1_38[55], stage1_38[56], stage1_38[57]},
      {stage2_40[9],stage2_39[36],stage2_38[48],stage2_37[56],stage2_36[67]}
   );
   gpc606_5 gpc5352 (
      {stage1_36[161], stage1_36[162], stage1_36[163], stage1_36[164], stage1_36[165], stage1_36[166]},
      {stage1_38[58], stage1_38[59], stage1_38[60], stage1_38[61], stage1_38[62], stage1_38[63]},
      {stage2_40[10],stage2_39[37],stage2_38[49],stage2_37[57],stage2_36[68]}
   );
   gpc606_5 gpc5353 (
      {stage1_36[167], stage1_36[168], stage1_36[169], stage1_36[170], stage1_36[171], stage1_36[172]},
      {stage1_38[64], stage1_38[65], stage1_38[66], stage1_38[67], stage1_38[68], stage1_38[69]},
      {stage2_40[11],stage2_39[38],stage2_38[50],stage2_37[58],stage2_36[69]}
   );
   gpc606_5 gpc5354 (
      {stage1_36[173], stage1_36[174], stage1_36[175], stage1_36[176], stage1_36[177], stage1_36[178]},
      {stage1_38[70], stage1_38[71], stage1_38[72], stage1_38[73], stage1_38[74], stage1_38[75]},
      {stage2_40[12],stage2_39[39],stage2_38[51],stage2_37[59],stage2_36[70]}
   );
   gpc606_5 gpc5355 (
      {stage1_36[179], stage1_36[180], stage1_36[181], stage1_36[182], stage1_36[183], stage1_36[184]},
      {stage1_38[76], stage1_38[77], stage1_38[78], stage1_38[79], stage1_38[80], stage1_38[81]},
      {stage2_40[13],stage2_39[40],stage2_38[52],stage2_37[60],stage2_36[71]}
   );
   gpc606_5 gpc5356 (
      {stage1_36[185], stage1_36[186], stage1_36[187], stage1_36[188], stage1_36[189], stage1_36[190]},
      {stage1_38[82], stage1_38[83], stage1_38[84], stage1_38[85], stage1_38[86], stage1_38[87]},
      {stage2_40[14],stage2_39[41],stage2_38[53],stage2_37[61],stage2_36[72]}
   );
   gpc606_5 gpc5357 (
      {stage1_36[191], stage1_36[192], stage1_36[193], stage1_36[194], stage1_36[195], stage1_36[196]},
      {stage1_38[88], stage1_38[89], stage1_38[90], stage1_38[91], stage1_38[92], stage1_38[93]},
      {stage2_40[15],stage2_39[42],stage2_38[54],stage2_37[62],stage2_36[73]}
   );
   gpc606_5 gpc5358 (
      {stage1_36[197], stage1_36[198], stage1_36[199], stage1_36[200], stage1_36[201], 1'b0},
      {stage1_38[94], stage1_38[95], stage1_38[96], stage1_38[97], stage1_38[98], stage1_38[99]},
      {stage2_40[16],stage2_39[43],stage2_38[55],stage2_37[63],stage2_36[74]}
   );
   gpc606_5 gpc5359 (
      {stage1_37[162], stage1_37[163], stage1_37[164], stage1_37[165], stage1_37[166], stage1_37[167]},
      {stage1_39[1], stage1_39[2], stage1_39[3], stage1_39[4], stage1_39[5], stage1_39[6]},
      {stage2_41[0],stage2_40[17],stage2_39[44],stage2_38[56],stage2_37[64]}
   );
   gpc606_5 gpc5360 (
      {stage1_37[168], stage1_37[169], stage1_37[170], stage1_37[171], stage1_37[172], stage1_37[173]},
      {stage1_39[7], stage1_39[8], stage1_39[9], stage1_39[10], stage1_39[11], stage1_39[12]},
      {stage2_41[1],stage2_40[18],stage2_39[45],stage2_38[57],stage2_37[65]}
   );
   gpc606_5 gpc5361 (
      {stage1_37[174], stage1_37[175], stage1_37[176], stage1_37[177], stage1_37[178], stage1_37[179]},
      {stage1_39[13], stage1_39[14], stage1_39[15], stage1_39[16], stage1_39[17], stage1_39[18]},
      {stage2_41[2],stage2_40[19],stage2_39[46],stage2_38[58],stage2_37[66]}
   );
   gpc606_5 gpc5362 (
      {stage1_37[180], stage1_37[181], stage1_37[182], stage1_37[183], stage1_37[184], stage1_37[185]},
      {stage1_39[19], stage1_39[20], stage1_39[21], stage1_39[22], stage1_39[23], stage1_39[24]},
      {stage2_41[3],stage2_40[20],stage2_39[47],stage2_38[59],stage2_37[67]}
   );
   gpc606_5 gpc5363 (
      {stage1_37[186], stage1_37[187], stage1_37[188], stage1_37[189], stage1_37[190], stage1_37[191]},
      {stage1_39[25], stage1_39[26], stage1_39[27], stage1_39[28], stage1_39[29], stage1_39[30]},
      {stage2_41[4],stage2_40[21],stage2_39[48],stage2_38[60],stage2_37[68]}
   );
   gpc606_5 gpc5364 (
      {stage1_37[192], stage1_37[193], stage1_37[194], stage1_37[195], stage1_37[196], stage1_37[197]},
      {stage1_39[31], stage1_39[32], stage1_39[33], stage1_39[34], stage1_39[35], stage1_39[36]},
      {stage2_41[5],stage2_40[22],stage2_39[49],stage2_38[61],stage2_37[69]}
   );
   gpc606_5 gpc5365 (
      {stage1_37[198], stage1_37[199], stage1_37[200], stage1_37[201], stage1_37[202], stage1_37[203]},
      {stage1_39[37], stage1_39[38], stage1_39[39], stage1_39[40], stage1_39[41], stage1_39[42]},
      {stage2_41[6],stage2_40[23],stage2_39[50],stage2_38[62],stage2_37[70]}
   );
   gpc606_5 gpc5366 (
      {stage1_37[204], stage1_37[205], stage1_37[206], stage1_37[207], stage1_37[208], stage1_37[209]},
      {stage1_39[43], stage1_39[44], stage1_39[45], stage1_39[46], stage1_39[47], stage1_39[48]},
      {stage2_41[7],stage2_40[24],stage2_39[51],stage2_38[63],stage2_37[71]}
   );
   gpc606_5 gpc5367 (
      {stage1_37[210], stage1_37[211], stage1_37[212], stage1_37[213], stage1_37[214], stage1_37[215]},
      {stage1_39[49], stage1_39[50], stage1_39[51], stage1_39[52], stage1_39[53], stage1_39[54]},
      {stage2_41[8],stage2_40[25],stage2_39[52],stage2_38[64],stage2_37[72]}
   );
   gpc606_5 gpc5368 (
      {stage1_37[216], stage1_37[217], stage1_37[218], stage1_37[219], stage1_37[220], stage1_37[221]},
      {stage1_39[55], stage1_39[56], stage1_39[57], stage1_39[58], stage1_39[59], stage1_39[60]},
      {stage2_41[9],stage2_40[26],stage2_39[53],stage2_38[65],stage2_37[73]}
   );
   gpc606_5 gpc5369 (
      {stage1_37[222], stage1_37[223], stage1_37[224], stage1_37[225], stage1_37[226], stage1_37[227]},
      {stage1_39[61], stage1_39[62], stage1_39[63], stage1_39[64], stage1_39[65], stage1_39[66]},
      {stage2_41[10],stage2_40[27],stage2_39[54],stage2_38[66],stage2_37[74]}
   );
   gpc606_5 gpc5370 (
      {stage1_37[228], stage1_37[229], stage1_37[230], stage1_37[231], stage1_37[232], stage1_37[233]},
      {stage1_39[67], stage1_39[68], stage1_39[69], stage1_39[70], stage1_39[71], stage1_39[72]},
      {stage2_41[11],stage2_40[28],stage2_39[55],stage2_38[67],stage2_37[75]}
   );
   gpc606_5 gpc5371 (
      {stage1_37[234], stage1_37[235], stage1_37[236], stage1_37[237], stage1_37[238], stage1_37[239]},
      {stage1_39[73], stage1_39[74], stage1_39[75], stage1_39[76], stage1_39[77], stage1_39[78]},
      {stage2_41[12],stage2_40[29],stage2_39[56],stage2_38[68],stage2_37[76]}
   );
   gpc606_5 gpc5372 (
      {stage1_37[240], stage1_37[241], stage1_37[242], stage1_37[243], stage1_37[244], stage1_37[245]},
      {stage1_39[79], stage1_39[80], stage1_39[81], stage1_39[82], stage1_39[83], stage1_39[84]},
      {stage2_41[13],stage2_40[30],stage2_39[57],stage2_38[69],stage2_37[77]}
   );
   gpc606_5 gpc5373 (
      {stage1_37[246], stage1_37[247], stage1_37[248], stage1_37[249], stage1_37[250], stage1_37[251]},
      {stage1_39[85], stage1_39[86], stage1_39[87], stage1_39[88], stage1_39[89], stage1_39[90]},
      {stage2_41[14],stage2_40[31],stage2_39[58],stage2_38[70],stage2_37[78]}
   );
   gpc606_5 gpc5374 (
      {stage1_37[252], stage1_37[253], stage1_37[254], stage1_37[255], stage1_37[256], stage1_37[257]},
      {stage1_39[91], stage1_39[92], stage1_39[93], stage1_39[94], stage1_39[95], stage1_39[96]},
      {stage2_41[15],stage2_40[32],stage2_39[59],stage2_38[71],stage2_37[79]}
   );
   gpc606_5 gpc5375 (
      {stage1_37[258], stage1_37[259], stage1_37[260], stage1_37[261], stage1_37[262], stage1_37[263]},
      {stage1_39[97], stage1_39[98], stage1_39[99], stage1_39[100], stage1_39[101], stage1_39[102]},
      {stage2_41[16],stage2_40[33],stage2_39[60],stage2_38[72],stage2_37[80]}
   );
   gpc606_5 gpc5376 (
      {stage1_37[264], stage1_37[265], stage1_37[266], stage1_37[267], stage1_37[268], stage1_37[269]},
      {stage1_39[103], stage1_39[104], stage1_39[105], stage1_39[106], stage1_39[107], stage1_39[108]},
      {stage2_41[17],stage2_40[34],stage2_39[61],stage2_38[73],stage2_37[81]}
   );
   gpc606_5 gpc5377 (
      {stage1_37[270], stage1_37[271], stage1_37[272], stage1_37[273], stage1_37[274], stage1_37[275]},
      {stage1_39[109], stage1_39[110], stage1_39[111], stage1_39[112], stage1_39[113], stage1_39[114]},
      {stage2_41[18],stage2_40[35],stage2_39[62],stage2_38[74],stage2_37[82]}
   );
   gpc606_5 gpc5378 (
      {stage1_37[276], stage1_37[277], stage1_37[278], stage1_37[279], stage1_37[280], stage1_37[281]},
      {stage1_39[115], stage1_39[116], stage1_39[117], stage1_39[118], stage1_39[119], stage1_39[120]},
      {stage2_41[19],stage2_40[36],stage2_39[63],stage2_38[75],stage2_37[83]}
   );
   gpc606_5 gpc5379 (
      {stage1_37[282], stage1_37[283], stage1_37[284], stage1_37[285], stage1_37[286], stage1_37[287]},
      {stage1_39[121], stage1_39[122], stage1_39[123], stage1_39[124], stage1_39[125], stage1_39[126]},
      {stage2_41[20],stage2_40[37],stage2_39[64],stage2_38[76],stage2_37[84]}
   );
   gpc606_5 gpc5380 (
      {stage1_37[288], stage1_37[289], stage1_37[290], stage1_37[291], stage1_37[292], stage1_37[293]},
      {stage1_39[127], stage1_39[128], stage1_39[129], stage1_39[130], stage1_39[131], stage1_39[132]},
      {stage2_41[21],stage2_40[38],stage2_39[65],stage2_38[77],stage2_37[85]}
   );
   gpc606_5 gpc5381 (
      {stage1_37[294], stage1_37[295], stage1_37[296], stage1_37[297], stage1_37[298], stage1_37[299]},
      {stage1_39[133], stage1_39[134], stage1_39[135], stage1_39[136], stage1_39[137], stage1_39[138]},
      {stage2_41[22],stage2_40[39],stage2_39[66],stage2_38[78],stage2_37[86]}
   );
   gpc606_5 gpc5382 (
      {stage1_37[300], stage1_37[301], stage1_37[302], stage1_37[303], stage1_37[304], stage1_37[305]},
      {stage1_39[139], stage1_39[140], stage1_39[141], stage1_39[142], stage1_39[143], stage1_39[144]},
      {stage2_41[23],stage2_40[40],stage2_39[67],stage2_38[79],stage2_37[87]}
   );
   gpc606_5 gpc5383 (
      {stage1_38[100], stage1_38[101], stage1_38[102], stage1_38[103], stage1_38[104], stage1_38[105]},
      {stage1_40[0], stage1_40[1], stage1_40[2], stage1_40[3], stage1_40[4], stage1_40[5]},
      {stage2_42[0],stage2_41[24],stage2_40[41],stage2_39[68],stage2_38[80]}
   );
   gpc615_5 gpc5384 (
      {stage1_38[106], stage1_38[107], stage1_38[108], stage1_38[109], stage1_38[110]},
      {stage1_39[145]},
      {stage1_40[6], stage1_40[7], stage1_40[8], stage1_40[9], stage1_40[10], stage1_40[11]},
      {stage2_42[1],stage2_41[25],stage2_40[42],stage2_39[69],stage2_38[81]}
   );
   gpc615_5 gpc5385 (
      {stage1_38[111], stage1_38[112], stage1_38[113], stage1_38[114], stage1_38[115]},
      {stage1_39[146]},
      {stage1_40[12], stage1_40[13], stage1_40[14], stage1_40[15], stage1_40[16], stage1_40[17]},
      {stage2_42[2],stage2_41[26],stage2_40[43],stage2_39[70],stage2_38[82]}
   );
   gpc615_5 gpc5386 (
      {stage1_38[116], stage1_38[117], stage1_38[118], stage1_38[119], stage1_38[120]},
      {stage1_39[147]},
      {stage1_40[18], stage1_40[19], stage1_40[20], stage1_40[21], stage1_40[22], stage1_40[23]},
      {stage2_42[3],stage2_41[27],stage2_40[44],stage2_39[71],stage2_38[83]}
   );
   gpc615_5 gpc5387 (
      {stage1_38[121], stage1_38[122], stage1_38[123], stage1_38[124], stage1_38[125]},
      {stage1_39[148]},
      {stage1_40[24], stage1_40[25], stage1_40[26], stage1_40[27], stage1_40[28], stage1_40[29]},
      {stage2_42[4],stage2_41[28],stage2_40[45],stage2_39[72],stage2_38[84]}
   );
   gpc615_5 gpc5388 (
      {stage1_38[126], stage1_38[127], stage1_38[128], stage1_38[129], stage1_38[130]},
      {stage1_39[149]},
      {stage1_40[30], stage1_40[31], stage1_40[32], stage1_40[33], stage1_40[34], stage1_40[35]},
      {stage2_42[5],stage2_41[29],stage2_40[46],stage2_39[73],stage2_38[85]}
   );
   gpc615_5 gpc5389 (
      {stage1_38[131], stage1_38[132], stage1_38[133], stage1_38[134], stage1_38[135]},
      {stage1_39[150]},
      {stage1_40[36], stage1_40[37], stage1_40[38], stage1_40[39], stage1_40[40], stage1_40[41]},
      {stage2_42[6],stage2_41[30],stage2_40[47],stage2_39[74],stage2_38[86]}
   );
   gpc615_5 gpc5390 (
      {stage1_38[136], stage1_38[137], stage1_38[138], stage1_38[139], stage1_38[140]},
      {stage1_39[151]},
      {stage1_40[42], stage1_40[43], stage1_40[44], stage1_40[45], stage1_40[46], stage1_40[47]},
      {stage2_42[7],stage2_41[31],stage2_40[48],stage2_39[75],stage2_38[87]}
   );
   gpc615_5 gpc5391 (
      {stage1_38[141], stage1_38[142], stage1_38[143], stage1_38[144], stage1_38[145]},
      {stage1_39[152]},
      {stage1_40[48], stage1_40[49], stage1_40[50], stage1_40[51], stage1_40[52], stage1_40[53]},
      {stage2_42[8],stage2_41[32],stage2_40[49],stage2_39[76],stage2_38[88]}
   );
   gpc615_5 gpc5392 (
      {stage1_38[146], stage1_38[147], stage1_38[148], stage1_38[149], stage1_38[150]},
      {stage1_39[153]},
      {stage1_40[54], stage1_40[55], stage1_40[56], stage1_40[57], stage1_40[58], stage1_40[59]},
      {stage2_42[9],stage2_41[33],stage2_40[50],stage2_39[77],stage2_38[89]}
   );
   gpc615_5 gpc5393 (
      {stage1_38[151], stage1_38[152], stage1_38[153], stage1_38[154], stage1_38[155]},
      {stage1_39[154]},
      {stage1_40[60], stage1_40[61], stage1_40[62], stage1_40[63], stage1_40[64], stage1_40[65]},
      {stage2_42[10],stage2_41[34],stage2_40[51],stage2_39[78],stage2_38[90]}
   );
   gpc615_5 gpc5394 (
      {stage1_38[156], stage1_38[157], stage1_38[158], stage1_38[159], stage1_38[160]},
      {stage1_39[155]},
      {stage1_40[66], stage1_40[67], stage1_40[68], stage1_40[69], stage1_40[70], stage1_40[71]},
      {stage2_42[11],stage2_41[35],stage2_40[52],stage2_39[79],stage2_38[91]}
   );
   gpc615_5 gpc5395 (
      {stage1_38[161], stage1_38[162], stage1_38[163], stage1_38[164], stage1_38[165]},
      {stage1_39[156]},
      {stage1_40[72], stage1_40[73], stage1_40[74], stage1_40[75], stage1_40[76], stage1_40[77]},
      {stage2_42[12],stage2_41[36],stage2_40[53],stage2_39[80],stage2_38[92]}
   );
   gpc615_5 gpc5396 (
      {stage1_38[166], stage1_38[167], stage1_38[168], stage1_38[169], stage1_38[170]},
      {stage1_39[157]},
      {stage1_40[78], stage1_40[79], stage1_40[80], stage1_40[81], stage1_40[82], stage1_40[83]},
      {stage2_42[13],stage2_41[37],stage2_40[54],stage2_39[81],stage2_38[93]}
   );
   gpc615_5 gpc5397 (
      {stage1_38[171], stage1_38[172], stage1_38[173], stage1_38[174], stage1_38[175]},
      {stage1_39[158]},
      {stage1_40[84], stage1_40[85], stage1_40[86], stage1_40[87], stage1_40[88], stage1_40[89]},
      {stage2_42[14],stage2_41[38],stage2_40[55],stage2_39[82],stage2_38[94]}
   );
   gpc615_5 gpc5398 (
      {stage1_38[176], stage1_38[177], stage1_38[178], stage1_38[179], stage1_38[180]},
      {stage1_39[159]},
      {stage1_40[90], stage1_40[91], stage1_40[92], stage1_40[93], stage1_40[94], stage1_40[95]},
      {stage2_42[15],stage2_41[39],stage2_40[56],stage2_39[83],stage2_38[95]}
   );
   gpc615_5 gpc5399 (
      {stage1_38[181], stage1_38[182], stage1_38[183], stage1_38[184], stage1_38[185]},
      {stage1_39[160]},
      {stage1_40[96], stage1_40[97], stage1_40[98], stage1_40[99], stage1_40[100], stage1_40[101]},
      {stage2_42[16],stage2_41[40],stage2_40[57],stage2_39[84],stage2_38[96]}
   );
   gpc615_5 gpc5400 (
      {stage1_38[186], stage1_38[187], stage1_38[188], stage1_38[189], stage1_38[190]},
      {stage1_39[161]},
      {stage1_40[102], stage1_40[103], stage1_40[104], stage1_40[105], stage1_40[106], stage1_40[107]},
      {stage2_42[17],stage2_41[41],stage2_40[58],stage2_39[85],stage2_38[97]}
   );
   gpc615_5 gpc5401 (
      {stage1_38[191], stage1_38[192], stage1_38[193], stage1_38[194], stage1_38[195]},
      {stage1_39[162]},
      {stage1_40[108], stage1_40[109], stage1_40[110], stage1_40[111], stage1_40[112], stage1_40[113]},
      {stage2_42[18],stage2_41[42],stage2_40[59],stage2_39[86],stage2_38[98]}
   );
   gpc615_5 gpc5402 (
      {stage1_38[196], stage1_38[197], stage1_38[198], stage1_38[199], stage1_38[200]},
      {stage1_39[163]},
      {stage1_40[114], stage1_40[115], stage1_40[116], stage1_40[117], stage1_40[118], stage1_40[119]},
      {stage2_42[19],stage2_41[43],stage2_40[60],stage2_39[87],stage2_38[99]}
   );
   gpc615_5 gpc5403 (
      {stage1_38[201], stage1_38[202], stage1_38[203], stage1_38[204], stage1_38[205]},
      {stage1_39[164]},
      {stage1_40[120], stage1_40[121], stage1_40[122], stage1_40[123], stage1_40[124], stage1_40[125]},
      {stage2_42[20],stage2_41[44],stage2_40[61],stage2_39[88],stage2_38[100]}
   );
   gpc615_5 gpc5404 (
      {stage1_38[206], stage1_38[207], stage1_38[208], stage1_38[209], stage1_38[210]},
      {stage1_39[165]},
      {stage1_40[126], stage1_40[127], stage1_40[128], stage1_40[129], stage1_40[130], stage1_40[131]},
      {stage2_42[21],stage2_41[45],stage2_40[62],stage2_39[89],stage2_38[101]}
   );
   gpc615_5 gpc5405 (
      {stage1_38[211], stage1_38[212], stage1_38[213], stage1_38[214], stage1_38[215]},
      {stage1_39[166]},
      {stage1_40[132], stage1_40[133], stage1_40[134], stage1_40[135], stage1_40[136], stage1_40[137]},
      {stage2_42[22],stage2_41[46],stage2_40[63],stage2_39[90],stage2_38[102]}
   );
   gpc615_5 gpc5406 (
      {stage1_38[216], stage1_38[217], stage1_38[218], stage1_38[219], stage1_38[220]},
      {stage1_39[167]},
      {stage1_40[138], stage1_40[139], stage1_40[140], stage1_40[141], stage1_40[142], stage1_40[143]},
      {stage2_42[23],stage2_41[47],stage2_40[64],stage2_39[91],stage2_38[103]}
   );
   gpc615_5 gpc5407 (
      {stage1_38[221], stage1_38[222], stage1_38[223], stage1_38[224], stage1_38[225]},
      {stage1_39[168]},
      {stage1_40[144], stage1_40[145], stage1_40[146], stage1_40[147], stage1_40[148], stage1_40[149]},
      {stage2_42[24],stage2_41[48],stage2_40[65],stage2_39[92],stage2_38[104]}
   );
   gpc615_5 gpc5408 (
      {stage1_38[226], stage1_38[227], stage1_38[228], stage1_38[229], stage1_38[230]},
      {stage1_39[169]},
      {stage1_40[150], stage1_40[151], stage1_40[152], stage1_40[153], stage1_40[154], stage1_40[155]},
      {stage2_42[25],stage2_41[49],stage2_40[66],stage2_39[93],stage2_38[105]}
   );
   gpc606_5 gpc5409 (
      {stage1_40[156], stage1_40[157], stage1_40[158], stage1_40[159], stage1_40[160], stage1_40[161]},
      {stage1_42[0], stage1_42[1], stage1_42[2], stage1_42[3], stage1_42[4], stage1_42[5]},
      {stage2_44[0],stage2_43[0],stage2_42[26],stage2_41[50],stage2_40[67]}
   );
   gpc606_5 gpc5410 (
      {stage1_40[162], stage1_40[163], stage1_40[164], stage1_40[165], stage1_40[166], stage1_40[167]},
      {stage1_42[6], stage1_42[7], stage1_42[8], stage1_42[9], stage1_42[10], stage1_42[11]},
      {stage2_44[1],stage2_43[1],stage2_42[27],stage2_41[51],stage2_40[68]}
   );
   gpc606_5 gpc5411 (
      {stage1_40[168], stage1_40[169], stage1_40[170], stage1_40[171], stage1_40[172], stage1_40[173]},
      {stage1_42[12], stage1_42[13], stage1_42[14], stage1_42[15], stage1_42[16], stage1_42[17]},
      {stage2_44[2],stage2_43[2],stage2_42[28],stage2_41[52],stage2_40[69]}
   );
   gpc606_5 gpc5412 (
      {stage1_40[174], stage1_40[175], stage1_40[176], stage1_40[177], stage1_40[178], stage1_40[179]},
      {stage1_42[18], stage1_42[19], stage1_42[20], stage1_42[21], stage1_42[22], stage1_42[23]},
      {stage2_44[3],stage2_43[3],stage2_42[29],stage2_41[53],stage2_40[70]}
   );
   gpc606_5 gpc5413 (
      {stage1_40[180], stage1_40[181], stage1_40[182], stage1_40[183], stage1_40[184], stage1_40[185]},
      {stage1_42[24], stage1_42[25], stage1_42[26], stage1_42[27], stage1_42[28], stage1_42[29]},
      {stage2_44[4],stage2_43[4],stage2_42[30],stage2_41[54],stage2_40[71]}
   );
   gpc606_5 gpc5414 (
      {stage1_40[186], stage1_40[187], stage1_40[188], stage1_40[189], stage1_40[190], stage1_40[191]},
      {stage1_42[30], stage1_42[31], stage1_42[32], stage1_42[33], stage1_42[34], stage1_42[35]},
      {stage2_44[5],stage2_43[5],stage2_42[31],stage2_41[55],stage2_40[72]}
   );
   gpc606_5 gpc5415 (
      {stage1_40[192], stage1_40[193], stage1_40[194], stage1_40[195], stage1_40[196], stage1_40[197]},
      {stage1_42[36], stage1_42[37], stage1_42[38], stage1_42[39], stage1_42[40], stage1_42[41]},
      {stage2_44[6],stage2_43[6],stage2_42[32],stage2_41[56],stage2_40[73]}
   );
   gpc606_5 gpc5416 (
      {stage1_40[198], stage1_40[199], stage1_40[200], stage1_40[201], stage1_40[202], stage1_40[203]},
      {stage1_42[42], stage1_42[43], stage1_42[44], stage1_42[45], stage1_42[46], stage1_42[47]},
      {stage2_44[7],stage2_43[7],stage2_42[33],stage2_41[57],stage2_40[74]}
   );
   gpc606_5 gpc5417 (
      {stage1_40[204], stage1_40[205], stage1_40[206], stage1_40[207], stage1_40[208], stage1_40[209]},
      {stage1_42[48], stage1_42[49], stage1_42[50], stage1_42[51], stage1_42[52], stage1_42[53]},
      {stage2_44[8],stage2_43[8],stage2_42[34],stage2_41[58],stage2_40[75]}
   );
   gpc606_5 gpc5418 (
      {stage1_40[210], stage1_40[211], stage1_40[212], stage1_40[213], stage1_40[214], stage1_40[215]},
      {stage1_42[54], stage1_42[55], stage1_42[56], stage1_42[57], stage1_42[58], stage1_42[59]},
      {stage2_44[9],stage2_43[9],stage2_42[35],stage2_41[59],stage2_40[76]}
   );
   gpc615_5 gpc5419 (
      {stage1_40[216], stage1_40[217], stage1_40[218], stage1_40[219], stage1_40[220]},
      {stage1_41[0]},
      {stage1_42[60], stage1_42[61], stage1_42[62], stage1_42[63], stage1_42[64], stage1_42[65]},
      {stage2_44[10],stage2_43[10],stage2_42[36],stage2_41[60],stage2_40[77]}
   );
   gpc615_5 gpc5420 (
      {stage1_40[221], stage1_40[222], stage1_40[223], stage1_40[224], stage1_40[225]},
      {stage1_41[1]},
      {stage1_42[66], stage1_42[67], stage1_42[68], stage1_42[69], stage1_42[70], stage1_42[71]},
      {stage2_44[11],stage2_43[11],stage2_42[37],stage2_41[61],stage2_40[78]}
   );
   gpc615_5 gpc5421 (
      {stage1_40[226], stage1_40[227], stage1_40[228], stage1_40[229], stage1_40[230]},
      {stage1_41[2]},
      {stage1_42[72], stage1_42[73], stage1_42[74], stage1_42[75], stage1_42[76], stage1_42[77]},
      {stage2_44[12],stage2_43[12],stage2_42[38],stage2_41[62],stage2_40[79]}
   );
   gpc615_5 gpc5422 (
      {stage1_40[231], stage1_40[232], stage1_40[233], stage1_40[234], stage1_40[235]},
      {stage1_41[3]},
      {stage1_42[78], stage1_42[79], stage1_42[80], stage1_42[81], stage1_42[82], stage1_42[83]},
      {stage2_44[13],stage2_43[13],stage2_42[39],stage2_41[63],stage2_40[80]}
   );
   gpc615_5 gpc5423 (
      {stage1_40[236], stage1_40[237], stage1_40[238], stage1_40[239], stage1_40[240]},
      {stage1_41[4]},
      {stage1_42[84], stage1_42[85], stage1_42[86], stage1_42[87], stage1_42[88], stage1_42[89]},
      {stage2_44[14],stage2_43[14],stage2_42[40],stage2_41[64],stage2_40[81]}
   );
   gpc615_5 gpc5424 (
      {stage1_40[241], stage1_40[242], stage1_40[243], stage1_40[244], stage1_40[245]},
      {stage1_41[5]},
      {stage1_42[90], stage1_42[91], stage1_42[92], stage1_42[93], stage1_42[94], stage1_42[95]},
      {stage2_44[15],stage2_43[15],stage2_42[41],stage2_41[65],stage2_40[82]}
   );
   gpc615_5 gpc5425 (
      {stage1_40[246], stage1_40[247], stage1_40[248], stage1_40[249], stage1_40[250]},
      {stage1_41[6]},
      {stage1_42[96], stage1_42[97], stage1_42[98], stage1_42[99], stage1_42[100], stage1_42[101]},
      {stage2_44[16],stage2_43[16],stage2_42[42],stage2_41[66],stage2_40[83]}
   );
   gpc615_5 gpc5426 (
      {stage1_40[251], stage1_40[252], stage1_40[253], stage1_40[254], stage1_40[255]},
      {stage1_41[7]},
      {stage1_42[102], stage1_42[103], stage1_42[104], stage1_42[105], stage1_42[106], stage1_42[107]},
      {stage2_44[17],stage2_43[17],stage2_42[43],stage2_41[67],stage2_40[84]}
   );
   gpc615_5 gpc5427 (
      {stage1_40[256], stage1_40[257], stage1_40[258], stage1_40[259], stage1_40[260]},
      {stage1_41[8]},
      {stage1_42[108], stage1_42[109], stage1_42[110], stage1_42[111], stage1_42[112], stage1_42[113]},
      {stage2_44[18],stage2_43[18],stage2_42[44],stage2_41[68],stage2_40[85]}
   );
   gpc615_5 gpc5428 (
      {stage1_40[261], stage1_40[262], stage1_40[263], stage1_40[264], stage1_40[265]},
      {stage1_41[9]},
      {stage1_42[114], stage1_42[115], stage1_42[116], stage1_42[117], stage1_42[118], stage1_42[119]},
      {stage2_44[19],stage2_43[19],stage2_42[45],stage2_41[69],stage2_40[86]}
   );
   gpc615_5 gpc5429 (
      {stage1_40[266], stage1_40[267], stage1_40[268], stage1_40[269], stage1_40[270]},
      {stage1_41[10]},
      {stage1_42[120], stage1_42[121], stage1_42[122], stage1_42[123], stage1_42[124], stage1_42[125]},
      {stage2_44[20],stage2_43[20],stage2_42[46],stage2_41[70],stage2_40[87]}
   );
   gpc615_5 gpc5430 (
      {stage1_40[271], stage1_40[272], stage1_40[273], stage1_40[274], stage1_40[275]},
      {stage1_41[11]},
      {stage1_42[126], stage1_42[127], stage1_42[128], stage1_42[129], stage1_42[130], stage1_42[131]},
      {stage2_44[21],stage2_43[21],stage2_42[47],stage2_41[71],stage2_40[88]}
   );
   gpc615_5 gpc5431 (
      {stage1_40[276], stage1_40[277], stage1_40[278], stage1_40[279], stage1_40[280]},
      {stage1_41[12]},
      {stage1_42[132], stage1_42[133], stage1_42[134], stage1_42[135], stage1_42[136], stage1_42[137]},
      {stage2_44[22],stage2_43[22],stage2_42[48],stage2_41[72],stage2_40[89]}
   );
   gpc606_5 gpc5432 (
      {stage1_41[13], stage1_41[14], stage1_41[15], stage1_41[16], stage1_41[17], stage1_41[18]},
      {stage1_43[0], stage1_43[1], stage1_43[2], stage1_43[3], stage1_43[4], stage1_43[5]},
      {stage2_45[0],stage2_44[23],stage2_43[23],stage2_42[49],stage2_41[73]}
   );
   gpc606_5 gpc5433 (
      {stage1_41[19], stage1_41[20], stage1_41[21], stage1_41[22], stage1_41[23], stage1_41[24]},
      {stage1_43[6], stage1_43[7], stage1_43[8], stage1_43[9], stage1_43[10], stage1_43[11]},
      {stage2_45[1],stage2_44[24],stage2_43[24],stage2_42[50],stage2_41[74]}
   );
   gpc606_5 gpc5434 (
      {stage1_41[25], stage1_41[26], stage1_41[27], stage1_41[28], stage1_41[29], stage1_41[30]},
      {stage1_43[12], stage1_43[13], stage1_43[14], stage1_43[15], stage1_43[16], stage1_43[17]},
      {stage2_45[2],stage2_44[25],stage2_43[25],stage2_42[51],stage2_41[75]}
   );
   gpc606_5 gpc5435 (
      {stage1_41[31], stage1_41[32], stage1_41[33], stage1_41[34], stage1_41[35], stage1_41[36]},
      {stage1_43[18], stage1_43[19], stage1_43[20], stage1_43[21], stage1_43[22], stage1_43[23]},
      {stage2_45[3],stage2_44[26],stage2_43[26],stage2_42[52],stage2_41[76]}
   );
   gpc606_5 gpc5436 (
      {stage1_41[37], stage1_41[38], stage1_41[39], stage1_41[40], stage1_41[41], stage1_41[42]},
      {stage1_43[24], stage1_43[25], stage1_43[26], stage1_43[27], stage1_43[28], stage1_43[29]},
      {stage2_45[4],stage2_44[27],stage2_43[27],stage2_42[53],stage2_41[77]}
   );
   gpc615_5 gpc5437 (
      {stage1_41[43], stage1_41[44], stage1_41[45], stage1_41[46], stage1_41[47]},
      {stage1_42[138]},
      {stage1_43[30], stage1_43[31], stage1_43[32], stage1_43[33], stage1_43[34], stage1_43[35]},
      {stage2_45[5],stage2_44[28],stage2_43[28],stage2_42[54],stage2_41[78]}
   );
   gpc615_5 gpc5438 (
      {stage1_41[48], stage1_41[49], stage1_41[50], stage1_41[51], stage1_41[52]},
      {stage1_42[139]},
      {stage1_43[36], stage1_43[37], stage1_43[38], stage1_43[39], stage1_43[40], stage1_43[41]},
      {stage2_45[6],stage2_44[29],stage2_43[29],stage2_42[55],stage2_41[79]}
   );
   gpc615_5 gpc5439 (
      {stage1_41[53], stage1_41[54], stage1_41[55], stage1_41[56], stage1_41[57]},
      {stage1_42[140]},
      {stage1_43[42], stage1_43[43], stage1_43[44], stage1_43[45], stage1_43[46], stage1_43[47]},
      {stage2_45[7],stage2_44[30],stage2_43[30],stage2_42[56],stage2_41[80]}
   );
   gpc615_5 gpc5440 (
      {stage1_41[58], stage1_41[59], stage1_41[60], stage1_41[61], stage1_41[62]},
      {stage1_42[141]},
      {stage1_43[48], stage1_43[49], stage1_43[50], stage1_43[51], stage1_43[52], stage1_43[53]},
      {stage2_45[8],stage2_44[31],stage2_43[31],stage2_42[57],stage2_41[81]}
   );
   gpc615_5 gpc5441 (
      {stage1_41[63], stage1_41[64], stage1_41[65], stage1_41[66], stage1_41[67]},
      {stage1_42[142]},
      {stage1_43[54], stage1_43[55], stage1_43[56], stage1_43[57], stage1_43[58], stage1_43[59]},
      {stage2_45[9],stage2_44[32],stage2_43[32],stage2_42[58],stage2_41[82]}
   );
   gpc615_5 gpc5442 (
      {stage1_41[68], stage1_41[69], stage1_41[70], stage1_41[71], stage1_41[72]},
      {stage1_42[143]},
      {stage1_43[60], stage1_43[61], stage1_43[62], stage1_43[63], stage1_43[64], stage1_43[65]},
      {stage2_45[10],stage2_44[33],stage2_43[33],stage2_42[59],stage2_41[83]}
   );
   gpc615_5 gpc5443 (
      {stage1_41[73], stage1_41[74], stage1_41[75], stage1_41[76], stage1_41[77]},
      {stage1_42[144]},
      {stage1_43[66], stage1_43[67], stage1_43[68], stage1_43[69], stage1_43[70], stage1_43[71]},
      {stage2_45[11],stage2_44[34],stage2_43[34],stage2_42[60],stage2_41[84]}
   );
   gpc615_5 gpc5444 (
      {stage1_41[78], stage1_41[79], stage1_41[80], stage1_41[81], stage1_41[82]},
      {stage1_42[145]},
      {stage1_43[72], stage1_43[73], stage1_43[74], stage1_43[75], stage1_43[76], stage1_43[77]},
      {stage2_45[12],stage2_44[35],stage2_43[35],stage2_42[61],stage2_41[85]}
   );
   gpc615_5 gpc5445 (
      {stage1_41[83], stage1_41[84], stage1_41[85], stage1_41[86], stage1_41[87]},
      {stage1_42[146]},
      {stage1_43[78], stage1_43[79], stage1_43[80], stage1_43[81], stage1_43[82], stage1_43[83]},
      {stage2_45[13],stage2_44[36],stage2_43[36],stage2_42[62],stage2_41[86]}
   );
   gpc615_5 gpc5446 (
      {stage1_41[88], stage1_41[89], stage1_41[90], stage1_41[91], stage1_41[92]},
      {stage1_42[147]},
      {stage1_43[84], stage1_43[85], stage1_43[86], stage1_43[87], stage1_43[88], stage1_43[89]},
      {stage2_45[14],stage2_44[37],stage2_43[37],stage2_42[63],stage2_41[87]}
   );
   gpc615_5 gpc5447 (
      {stage1_41[93], stage1_41[94], stage1_41[95], stage1_41[96], stage1_41[97]},
      {stage1_42[148]},
      {stage1_43[90], stage1_43[91], stage1_43[92], stage1_43[93], stage1_43[94], stage1_43[95]},
      {stage2_45[15],stage2_44[38],stage2_43[38],stage2_42[64],stage2_41[88]}
   );
   gpc615_5 gpc5448 (
      {stage1_41[98], stage1_41[99], stage1_41[100], stage1_41[101], stage1_41[102]},
      {stage1_42[149]},
      {stage1_43[96], stage1_43[97], stage1_43[98], stage1_43[99], stage1_43[100], stage1_43[101]},
      {stage2_45[16],stage2_44[39],stage2_43[39],stage2_42[65],stage2_41[89]}
   );
   gpc615_5 gpc5449 (
      {stage1_41[103], stage1_41[104], stage1_41[105], stage1_41[106], stage1_41[107]},
      {stage1_42[150]},
      {stage1_43[102], stage1_43[103], stage1_43[104], stage1_43[105], stage1_43[106], stage1_43[107]},
      {stage2_45[17],stage2_44[40],stage2_43[40],stage2_42[66],stage2_41[90]}
   );
   gpc615_5 gpc5450 (
      {stage1_41[108], stage1_41[109], stage1_41[110], stage1_41[111], stage1_41[112]},
      {stage1_42[151]},
      {stage1_43[108], stage1_43[109], stage1_43[110], stage1_43[111], stage1_43[112], stage1_43[113]},
      {stage2_45[18],stage2_44[41],stage2_43[41],stage2_42[67],stage2_41[91]}
   );
   gpc615_5 gpc5451 (
      {stage1_41[113], stage1_41[114], stage1_41[115], stage1_41[116], stage1_41[117]},
      {stage1_42[152]},
      {stage1_43[114], stage1_43[115], stage1_43[116], stage1_43[117], stage1_43[118], stage1_43[119]},
      {stage2_45[19],stage2_44[42],stage2_43[42],stage2_42[68],stage2_41[92]}
   );
   gpc615_5 gpc5452 (
      {stage1_41[118], stage1_41[119], stage1_41[120], stage1_41[121], stage1_41[122]},
      {stage1_42[153]},
      {stage1_43[120], stage1_43[121], stage1_43[122], stage1_43[123], stage1_43[124], stage1_43[125]},
      {stage2_45[20],stage2_44[43],stage2_43[43],stage2_42[69],stage2_41[93]}
   );
   gpc615_5 gpc5453 (
      {stage1_41[123], stage1_41[124], stage1_41[125], stage1_41[126], stage1_41[127]},
      {stage1_42[154]},
      {stage1_43[126], stage1_43[127], stage1_43[128], stage1_43[129], stage1_43[130], stage1_43[131]},
      {stage2_45[21],stage2_44[44],stage2_43[44],stage2_42[70],stage2_41[94]}
   );
   gpc615_5 gpc5454 (
      {stage1_41[128], stage1_41[129], stage1_41[130], stage1_41[131], stage1_41[132]},
      {stage1_42[155]},
      {stage1_43[132], stage1_43[133], stage1_43[134], stage1_43[135], stage1_43[136], stage1_43[137]},
      {stage2_45[22],stage2_44[45],stage2_43[45],stage2_42[71],stage2_41[95]}
   );
   gpc615_5 gpc5455 (
      {stage1_41[133], stage1_41[134], stage1_41[135], stage1_41[136], stage1_41[137]},
      {stage1_42[156]},
      {stage1_43[138], stage1_43[139], stage1_43[140], stage1_43[141], stage1_43[142], stage1_43[143]},
      {stage2_45[23],stage2_44[46],stage2_43[46],stage2_42[72],stage2_41[96]}
   );
   gpc615_5 gpc5456 (
      {stage1_41[138], stage1_41[139], stage1_41[140], stage1_41[141], stage1_41[142]},
      {stage1_42[157]},
      {stage1_43[144], stage1_43[145], stage1_43[146], stage1_43[147], stage1_43[148], stage1_43[149]},
      {stage2_45[24],stage2_44[47],stage2_43[47],stage2_42[73],stage2_41[97]}
   );
   gpc615_5 gpc5457 (
      {stage1_41[143], stage1_41[144], stage1_41[145], stage1_41[146], stage1_41[147]},
      {stage1_42[158]},
      {stage1_43[150], stage1_43[151], stage1_43[152], stage1_43[153], stage1_43[154], stage1_43[155]},
      {stage2_45[25],stage2_44[48],stage2_43[48],stage2_42[74],stage2_41[98]}
   );
   gpc615_5 gpc5458 (
      {stage1_41[148], stage1_41[149], stage1_41[150], stage1_41[151], stage1_41[152]},
      {stage1_42[159]},
      {stage1_43[156], stage1_43[157], stage1_43[158], stage1_43[159], stage1_43[160], stage1_43[161]},
      {stage2_45[26],stage2_44[49],stage2_43[49],stage2_42[75],stage2_41[99]}
   );
   gpc615_5 gpc5459 (
      {stage1_41[153], stage1_41[154], stage1_41[155], stage1_41[156], stage1_41[157]},
      {stage1_42[160]},
      {stage1_43[162], stage1_43[163], stage1_43[164], stage1_43[165], stage1_43[166], stage1_43[167]},
      {stage2_45[27],stage2_44[50],stage2_43[50],stage2_42[76],stage2_41[100]}
   );
   gpc615_5 gpc5460 (
      {stage1_41[158], stage1_41[159], stage1_41[160], stage1_41[161], stage1_41[162]},
      {stage1_42[161]},
      {stage1_43[168], stage1_43[169], stage1_43[170], stage1_43[171], stage1_43[172], stage1_43[173]},
      {stage2_45[28],stage2_44[51],stage2_43[51],stage2_42[77],stage2_41[101]}
   );
   gpc615_5 gpc5461 (
      {stage1_41[163], stage1_41[164], stage1_41[165], stage1_41[166], stage1_41[167]},
      {stage1_42[162]},
      {stage1_43[174], stage1_43[175], stage1_43[176], stage1_43[177], stage1_43[178], stage1_43[179]},
      {stage2_45[29],stage2_44[52],stage2_43[52],stage2_42[78],stage2_41[102]}
   );
   gpc615_5 gpc5462 (
      {stage1_42[163], stage1_42[164], stage1_42[165], stage1_42[166], stage1_42[167]},
      {stage1_43[180]},
      {stage1_44[0], stage1_44[1], stage1_44[2], stage1_44[3], stage1_44[4], stage1_44[5]},
      {stage2_46[0],stage2_45[30],stage2_44[53],stage2_43[53],stage2_42[79]}
   );
   gpc615_5 gpc5463 (
      {stage1_43[181], stage1_43[182], stage1_43[183], stage1_43[184], stage1_43[185]},
      {stage1_44[6]},
      {stage1_45[0], stage1_45[1], stage1_45[2], stage1_45[3], stage1_45[4], stage1_45[5]},
      {stage2_47[0],stage2_46[1],stage2_45[31],stage2_44[54],stage2_43[54]}
   );
   gpc615_5 gpc5464 (
      {stage1_43[186], stage1_43[187], stage1_43[188], stage1_43[189], stage1_43[190]},
      {stage1_44[7]},
      {stage1_45[6], stage1_45[7], stage1_45[8], stage1_45[9], stage1_45[10], stage1_45[11]},
      {stage2_47[1],stage2_46[2],stage2_45[32],stage2_44[55],stage2_43[55]}
   );
   gpc615_5 gpc5465 (
      {stage1_43[191], stage1_43[192], stage1_43[193], stage1_43[194], stage1_43[195]},
      {stage1_44[8]},
      {stage1_45[12], stage1_45[13], stage1_45[14], stage1_45[15], stage1_45[16], stage1_45[17]},
      {stage2_47[2],stage2_46[3],stage2_45[33],stage2_44[56],stage2_43[56]}
   );
   gpc615_5 gpc5466 (
      {stage1_43[196], stage1_43[197], stage1_43[198], stage1_43[199], stage1_43[200]},
      {stage1_44[9]},
      {stage1_45[18], stage1_45[19], stage1_45[20], stage1_45[21], stage1_45[22], stage1_45[23]},
      {stage2_47[3],stage2_46[4],stage2_45[34],stage2_44[57],stage2_43[57]}
   );
   gpc615_5 gpc5467 (
      {stage1_43[201], stage1_43[202], stage1_43[203], stage1_43[204], stage1_43[205]},
      {stage1_44[10]},
      {stage1_45[24], stage1_45[25], stage1_45[26], stage1_45[27], stage1_45[28], stage1_45[29]},
      {stage2_47[4],stage2_46[5],stage2_45[35],stage2_44[58],stage2_43[58]}
   );
   gpc615_5 gpc5468 (
      {stage1_43[206], stage1_43[207], stage1_43[208], stage1_43[209], stage1_43[210]},
      {stage1_44[11]},
      {stage1_45[30], stage1_45[31], stage1_45[32], stage1_45[33], stage1_45[34], stage1_45[35]},
      {stage2_47[5],stage2_46[6],stage2_45[36],stage2_44[59],stage2_43[59]}
   );
   gpc615_5 gpc5469 (
      {stage1_43[211], stage1_43[212], stage1_43[213], stage1_43[214], stage1_43[215]},
      {stage1_44[12]},
      {stage1_45[36], stage1_45[37], stage1_45[38], stage1_45[39], stage1_45[40], stage1_45[41]},
      {stage2_47[6],stage2_46[7],stage2_45[37],stage2_44[60],stage2_43[60]}
   );
   gpc615_5 gpc5470 (
      {stage1_43[216], stage1_43[217], stage1_43[218], stage1_43[219], stage1_43[220]},
      {stage1_44[13]},
      {stage1_45[42], stage1_45[43], stage1_45[44], stage1_45[45], stage1_45[46], stage1_45[47]},
      {stage2_47[7],stage2_46[8],stage2_45[38],stage2_44[61],stage2_43[61]}
   );
   gpc615_5 gpc5471 (
      {stage1_43[221], stage1_43[222], stage1_43[223], stage1_43[224], stage1_43[225]},
      {stage1_44[14]},
      {stage1_45[48], stage1_45[49], stage1_45[50], stage1_45[51], stage1_45[52], stage1_45[53]},
      {stage2_47[8],stage2_46[9],stage2_45[39],stage2_44[62],stage2_43[62]}
   );
   gpc615_5 gpc5472 (
      {stage1_43[226], stage1_43[227], stage1_43[228], stage1_43[229], stage1_43[230]},
      {stage1_44[15]},
      {stage1_45[54], stage1_45[55], stage1_45[56], stage1_45[57], stage1_45[58], stage1_45[59]},
      {stage2_47[9],stage2_46[10],stage2_45[40],stage2_44[63],stage2_43[63]}
   );
   gpc615_5 gpc5473 (
      {stage1_43[231], stage1_43[232], stage1_43[233], stage1_43[234], stage1_43[235]},
      {stage1_44[16]},
      {stage1_45[60], stage1_45[61], stage1_45[62], stage1_45[63], stage1_45[64], stage1_45[65]},
      {stage2_47[10],stage2_46[11],stage2_45[41],stage2_44[64],stage2_43[64]}
   );
   gpc615_5 gpc5474 (
      {stage1_43[236], stage1_43[237], stage1_43[238], stage1_43[239], stage1_43[240]},
      {stage1_44[17]},
      {stage1_45[66], stage1_45[67], stage1_45[68], stage1_45[69], stage1_45[70], stage1_45[71]},
      {stage2_47[11],stage2_46[12],stage2_45[42],stage2_44[65],stage2_43[65]}
   );
   gpc606_5 gpc5475 (
      {stage1_44[18], stage1_44[19], stage1_44[20], stage1_44[21], stage1_44[22], stage1_44[23]},
      {stage1_46[0], stage1_46[1], stage1_46[2], stage1_46[3], stage1_46[4], stage1_46[5]},
      {stage2_48[0],stage2_47[12],stage2_46[13],stage2_45[43],stage2_44[66]}
   );
   gpc606_5 gpc5476 (
      {stage1_44[24], stage1_44[25], stage1_44[26], stage1_44[27], stage1_44[28], stage1_44[29]},
      {stage1_46[6], stage1_46[7], stage1_46[8], stage1_46[9], stage1_46[10], stage1_46[11]},
      {stage2_48[1],stage2_47[13],stage2_46[14],stage2_45[44],stage2_44[67]}
   );
   gpc606_5 gpc5477 (
      {stage1_44[30], stage1_44[31], stage1_44[32], stage1_44[33], stage1_44[34], stage1_44[35]},
      {stage1_46[12], stage1_46[13], stage1_46[14], stage1_46[15], stage1_46[16], stage1_46[17]},
      {stage2_48[2],stage2_47[14],stage2_46[15],stage2_45[45],stage2_44[68]}
   );
   gpc606_5 gpc5478 (
      {stage1_44[36], stage1_44[37], stage1_44[38], stage1_44[39], stage1_44[40], stage1_44[41]},
      {stage1_46[18], stage1_46[19], stage1_46[20], stage1_46[21], stage1_46[22], stage1_46[23]},
      {stage2_48[3],stage2_47[15],stage2_46[16],stage2_45[46],stage2_44[69]}
   );
   gpc606_5 gpc5479 (
      {stage1_44[42], stage1_44[43], stage1_44[44], stage1_44[45], stage1_44[46], stage1_44[47]},
      {stage1_46[24], stage1_46[25], stage1_46[26], stage1_46[27], stage1_46[28], stage1_46[29]},
      {stage2_48[4],stage2_47[16],stage2_46[17],stage2_45[47],stage2_44[70]}
   );
   gpc606_5 gpc5480 (
      {stage1_44[48], stage1_44[49], stage1_44[50], stage1_44[51], stage1_44[52], stage1_44[53]},
      {stage1_46[30], stage1_46[31], stage1_46[32], stage1_46[33], stage1_46[34], stage1_46[35]},
      {stage2_48[5],stage2_47[17],stage2_46[18],stage2_45[48],stage2_44[71]}
   );
   gpc606_5 gpc5481 (
      {stage1_44[54], stage1_44[55], stage1_44[56], stage1_44[57], stage1_44[58], stage1_44[59]},
      {stage1_46[36], stage1_46[37], stage1_46[38], stage1_46[39], stage1_46[40], stage1_46[41]},
      {stage2_48[6],stage2_47[18],stage2_46[19],stage2_45[49],stage2_44[72]}
   );
   gpc606_5 gpc5482 (
      {stage1_44[60], stage1_44[61], stage1_44[62], stage1_44[63], stage1_44[64], stage1_44[65]},
      {stage1_46[42], stage1_46[43], stage1_46[44], stage1_46[45], stage1_46[46], stage1_46[47]},
      {stage2_48[7],stage2_47[19],stage2_46[20],stage2_45[50],stage2_44[73]}
   );
   gpc606_5 gpc5483 (
      {stage1_44[66], stage1_44[67], stage1_44[68], stage1_44[69], stage1_44[70], stage1_44[71]},
      {stage1_46[48], stage1_46[49], stage1_46[50], stage1_46[51], stage1_46[52], stage1_46[53]},
      {stage2_48[8],stage2_47[20],stage2_46[21],stage2_45[51],stage2_44[74]}
   );
   gpc606_5 gpc5484 (
      {stage1_44[72], stage1_44[73], stage1_44[74], stage1_44[75], stage1_44[76], stage1_44[77]},
      {stage1_46[54], stage1_46[55], stage1_46[56], stage1_46[57], stage1_46[58], stage1_46[59]},
      {stage2_48[9],stage2_47[21],stage2_46[22],stage2_45[52],stage2_44[75]}
   );
   gpc606_5 gpc5485 (
      {stage1_44[78], stage1_44[79], stage1_44[80], stage1_44[81], stage1_44[82], stage1_44[83]},
      {stage1_46[60], stage1_46[61], stage1_46[62], stage1_46[63], stage1_46[64], stage1_46[65]},
      {stage2_48[10],stage2_47[22],stage2_46[23],stage2_45[53],stage2_44[76]}
   );
   gpc606_5 gpc5486 (
      {stage1_44[84], stage1_44[85], stage1_44[86], stage1_44[87], stage1_44[88], stage1_44[89]},
      {stage1_46[66], stage1_46[67], stage1_46[68], stage1_46[69], stage1_46[70], stage1_46[71]},
      {stage2_48[11],stage2_47[23],stage2_46[24],stage2_45[54],stage2_44[77]}
   );
   gpc606_5 gpc5487 (
      {stage1_44[90], stage1_44[91], stage1_44[92], stage1_44[93], stage1_44[94], stage1_44[95]},
      {stage1_46[72], stage1_46[73], stage1_46[74], stage1_46[75], stage1_46[76], stage1_46[77]},
      {stage2_48[12],stage2_47[24],stage2_46[25],stage2_45[55],stage2_44[78]}
   );
   gpc606_5 gpc5488 (
      {stage1_44[96], stage1_44[97], stage1_44[98], stage1_44[99], stage1_44[100], stage1_44[101]},
      {stage1_46[78], stage1_46[79], stage1_46[80], stage1_46[81], stage1_46[82], stage1_46[83]},
      {stage2_48[13],stage2_47[25],stage2_46[26],stage2_45[56],stage2_44[79]}
   );
   gpc606_5 gpc5489 (
      {stage1_44[102], stage1_44[103], stage1_44[104], stage1_44[105], stage1_44[106], stage1_44[107]},
      {stage1_46[84], stage1_46[85], stage1_46[86], stage1_46[87], stage1_46[88], stage1_46[89]},
      {stage2_48[14],stage2_47[26],stage2_46[27],stage2_45[57],stage2_44[80]}
   );
   gpc606_5 gpc5490 (
      {stage1_44[108], stage1_44[109], stage1_44[110], stage1_44[111], stage1_44[112], stage1_44[113]},
      {stage1_46[90], stage1_46[91], stage1_46[92], stage1_46[93], stage1_46[94], stage1_46[95]},
      {stage2_48[15],stage2_47[27],stage2_46[28],stage2_45[58],stage2_44[81]}
   );
   gpc606_5 gpc5491 (
      {stage1_44[114], stage1_44[115], stage1_44[116], stage1_44[117], stage1_44[118], stage1_44[119]},
      {stage1_46[96], stage1_46[97], stage1_46[98], stage1_46[99], stage1_46[100], stage1_46[101]},
      {stage2_48[16],stage2_47[28],stage2_46[29],stage2_45[59],stage2_44[82]}
   );
   gpc606_5 gpc5492 (
      {stage1_44[120], stage1_44[121], stage1_44[122], stage1_44[123], stage1_44[124], stage1_44[125]},
      {stage1_46[102], stage1_46[103], stage1_46[104], stage1_46[105], stage1_46[106], stage1_46[107]},
      {stage2_48[17],stage2_47[29],stage2_46[30],stage2_45[60],stage2_44[83]}
   );
   gpc606_5 gpc5493 (
      {stage1_44[126], stage1_44[127], stage1_44[128], stage1_44[129], stage1_44[130], stage1_44[131]},
      {stage1_46[108], stage1_46[109], stage1_46[110], stage1_46[111], stage1_46[112], stage1_46[113]},
      {stage2_48[18],stage2_47[30],stage2_46[31],stage2_45[61],stage2_44[84]}
   );
   gpc606_5 gpc5494 (
      {stage1_44[132], stage1_44[133], stage1_44[134], stage1_44[135], stage1_44[136], stage1_44[137]},
      {stage1_46[114], stage1_46[115], stage1_46[116], stage1_46[117], stage1_46[118], stage1_46[119]},
      {stage2_48[19],stage2_47[31],stage2_46[32],stage2_45[62],stage2_44[85]}
   );
   gpc606_5 gpc5495 (
      {stage1_44[138], stage1_44[139], stage1_44[140], stage1_44[141], stage1_44[142], stage1_44[143]},
      {stage1_46[120], stage1_46[121], stage1_46[122], stage1_46[123], stage1_46[124], stage1_46[125]},
      {stage2_48[20],stage2_47[32],stage2_46[33],stage2_45[63],stage2_44[86]}
   );
   gpc606_5 gpc5496 (
      {stage1_44[144], stage1_44[145], stage1_44[146], stage1_44[147], stage1_44[148], stage1_44[149]},
      {stage1_46[126], stage1_46[127], stage1_46[128], stage1_46[129], stage1_46[130], stage1_46[131]},
      {stage2_48[21],stage2_47[33],stage2_46[34],stage2_45[64],stage2_44[87]}
   );
   gpc606_5 gpc5497 (
      {stage1_44[150], stage1_44[151], stage1_44[152], stage1_44[153], stage1_44[154], stage1_44[155]},
      {stage1_46[132], stage1_46[133], stage1_46[134], stage1_46[135], stage1_46[136], stage1_46[137]},
      {stage2_48[22],stage2_47[34],stage2_46[35],stage2_45[65],stage2_44[88]}
   );
   gpc606_5 gpc5498 (
      {stage1_44[156], stage1_44[157], stage1_44[158], stage1_44[159], stage1_44[160], stage1_44[161]},
      {stage1_46[138], stage1_46[139], stage1_46[140], stage1_46[141], stage1_46[142], stage1_46[143]},
      {stage2_48[23],stage2_47[35],stage2_46[36],stage2_45[66],stage2_44[89]}
   );
   gpc606_5 gpc5499 (
      {stage1_44[162], stage1_44[163], stage1_44[164], stage1_44[165], stage1_44[166], stage1_44[167]},
      {stage1_46[144], stage1_46[145], stage1_46[146], stage1_46[147], stage1_46[148], stage1_46[149]},
      {stage2_48[24],stage2_47[36],stage2_46[37],stage2_45[67],stage2_44[90]}
   );
   gpc606_5 gpc5500 (
      {stage1_44[168], stage1_44[169], stage1_44[170], stage1_44[171], stage1_44[172], stage1_44[173]},
      {stage1_46[150], stage1_46[151], stage1_46[152], stage1_46[153], stage1_46[154], stage1_46[155]},
      {stage2_48[25],stage2_47[37],stage2_46[38],stage2_45[68],stage2_44[91]}
   );
   gpc606_5 gpc5501 (
      {stage1_44[174], stage1_44[175], stage1_44[176], stage1_44[177], stage1_44[178], stage1_44[179]},
      {stage1_46[156], stage1_46[157], stage1_46[158], stage1_46[159], stage1_46[160], stage1_46[161]},
      {stage2_48[26],stage2_47[38],stage2_46[39],stage2_45[69],stage2_44[92]}
   );
   gpc606_5 gpc5502 (
      {stage1_44[180], stage1_44[181], stage1_44[182], stage1_44[183], stage1_44[184], stage1_44[185]},
      {stage1_46[162], stage1_46[163], stage1_46[164], stage1_46[165], stage1_46[166], stage1_46[167]},
      {stage2_48[27],stage2_47[39],stage2_46[40],stage2_45[70],stage2_44[93]}
   );
   gpc606_5 gpc5503 (
      {stage1_44[186], stage1_44[187], stage1_44[188], stage1_44[189], stage1_44[190], stage1_44[191]},
      {stage1_46[168], stage1_46[169], stage1_46[170], stage1_46[171], stage1_46[172], stage1_46[173]},
      {stage2_48[28],stage2_47[40],stage2_46[41],stage2_45[71],stage2_44[94]}
   );
   gpc606_5 gpc5504 (
      {stage1_44[192], stage1_44[193], stage1_44[194], stage1_44[195], stage1_44[196], stage1_44[197]},
      {stage1_46[174], stage1_46[175], stage1_46[176], stage1_46[177], stage1_46[178], stage1_46[179]},
      {stage2_48[29],stage2_47[41],stage2_46[42],stage2_45[72],stage2_44[95]}
   );
   gpc606_5 gpc5505 (
      {stage1_44[198], stage1_44[199], stage1_44[200], stage1_44[201], stage1_44[202], stage1_44[203]},
      {stage1_46[180], stage1_46[181], stage1_46[182], stage1_46[183], stage1_46[184], stage1_46[185]},
      {stage2_48[30],stage2_47[42],stage2_46[43],stage2_45[73],stage2_44[96]}
   );
   gpc606_5 gpc5506 (
      {stage1_44[204], stage1_44[205], stage1_44[206], stage1_44[207], stage1_44[208], stage1_44[209]},
      {stage1_46[186], stage1_46[187], stage1_46[188], stage1_46[189], stage1_46[190], stage1_46[191]},
      {stage2_48[31],stage2_47[43],stage2_46[44],stage2_45[74],stage2_44[97]}
   );
   gpc606_5 gpc5507 (
      {stage1_44[210], stage1_44[211], stage1_44[212], stage1_44[213], stage1_44[214], stage1_44[215]},
      {stage1_46[192], stage1_46[193], stage1_46[194], stage1_46[195], stage1_46[196], stage1_46[197]},
      {stage2_48[32],stage2_47[44],stage2_46[45],stage2_45[75],stage2_44[98]}
   );
   gpc606_5 gpc5508 (
      {stage1_44[216], stage1_44[217], stage1_44[218], stage1_44[219], stage1_44[220], stage1_44[221]},
      {stage1_46[198], stage1_46[199], stage1_46[200], stage1_46[201], stage1_46[202], stage1_46[203]},
      {stage2_48[33],stage2_47[45],stage2_46[46],stage2_45[76],stage2_44[99]}
   );
   gpc606_5 gpc5509 (
      {stage1_44[222], stage1_44[223], stage1_44[224], stage1_44[225], stage1_44[226], stage1_44[227]},
      {stage1_46[204], stage1_46[205], stage1_46[206], stage1_46[207], stage1_46[208], stage1_46[209]},
      {stage2_48[34],stage2_47[46],stage2_46[47],stage2_45[77],stage2_44[100]}
   );
   gpc606_5 gpc5510 (
      {stage1_44[228], stage1_44[229], stage1_44[230], stage1_44[231], stage1_44[232], stage1_44[233]},
      {stage1_46[210], stage1_46[211], stage1_46[212], stage1_46[213], stage1_46[214], stage1_46[215]},
      {stage2_48[35],stage2_47[47],stage2_46[48],stage2_45[78],stage2_44[101]}
   );
   gpc606_5 gpc5511 (
      {stage1_44[234], stage1_44[235], stage1_44[236], stage1_44[237], stage1_44[238], stage1_44[239]},
      {stage1_46[216], stage1_46[217], stage1_46[218], stage1_46[219], stage1_46[220], stage1_46[221]},
      {stage2_48[36],stage2_47[48],stage2_46[49],stage2_45[79],stage2_44[102]}
   );
   gpc606_5 gpc5512 (
      {stage1_45[72], stage1_45[73], stage1_45[74], stage1_45[75], stage1_45[76], stage1_45[77]},
      {stage1_47[0], stage1_47[1], stage1_47[2], stage1_47[3], stage1_47[4], stage1_47[5]},
      {stage2_49[0],stage2_48[37],stage2_47[49],stage2_46[50],stage2_45[80]}
   );
   gpc606_5 gpc5513 (
      {stage1_45[78], stage1_45[79], stage1_45[80], stage1_45[81], stage1_45[82], stage1_45[83]},
      {stage1_47[6], stage1_47[7], stage1_47[8], stage1_47[9], stage1_47[10], stage1_47[11]},
      {stage2_49[1],stage2_48[38],stage2_47[50],stage2_46[51],stage2_45[81]}
   );
   gpc615_5 gpc5514 (
      {stage1_45[84], stage1_45[85], stage1_45[86], stage1_45[87], stage1_45[88]},
      {stage1_46[222]},
      {stage1_47[12], stage1_47[13], stage1_47[14], stage1_47[15], stage1_47[16], stage1_47[17]},
      {stage2_49[2],stage2_48[39],stage2_47[51],stage2_46[52],stage2_45[82]}
   );
   gpc615_5 gpc5515 (
      {stage1_45[89], stage1_45[90], stage1_45[91], stage1_45[92], stage1_45[93]},
      {stage1_46[223]},
      {stage1_47[18], stage1_47[19], stage1_47[20], stage1_47[21], stage1_47[22], stage1_47[23]},
      {stage2_49[3],stage2_48[40],stage2_47[52],stage2_46[53],stage2_45[83]}
   );
   gpc615_5 gpc5516 (
      {stage1_45[94], stage1_45[95], stage1_45[96], stage1_45[97], stage1_45[98]},
      {stage1_46[224]},
      {stage1_47[24], stage1_47[25], stage1_47[26], stage1_47[27], stage1_47[28], stage1_47[29]},
      {stage2_49[4],stage2_48[41],stage2_47[53],stage2_46[54],stage2_45[84]}
   );
   gpc615_5 gpc5517 (
      {stage1_45[99], stage1_45[100], stage1_45[101], stage1_45[102], stage1_45[103]},
      {stage1_46[225]},
      {stage1_47[30], stage1_47[31], stage1_47[32], stage1_47[33], stage1_47[34], stage1_47[35]},
      {stage2_49[5],stage2_48[42],stage2_47[54],stage2_46[55],stage2_45[85]}
   );
   gpc615_5 gpc5518 (
      {stage1_45[104], stage1_45[105], stage1_45[106], stage1_45[107], stage1_45[108]},
      {stage1_46[226]},
      {stage1_47[36], stage1_47[37], stage1_47[38], stage1_47[39], stage1_47[40], stage1_47[41]},
      {stage2_49[6],stage2_48[43],stage2_47[55],stage2_46[56],stage2_45[86]}
   );
   gpc615_5 gpc5519 (
      {stage1_45[109], stage1_45[110], stage1_45[111], stage1_45[112], stage1_45[113]},
      {stage1_46[227]},
      {stage1_47[42], stage1_47[43], stage1_47[44], stage1_47[45], stage1_47[46], stage1_47[47]},
      {stage2_49[7],stage2_48[44],stage2_47[56],stage2_46[57],stage2_45[87]}
   );
   gpc615_5 gpc5520 (
      {stage1_45[114], stage1_45[115], stage1_45[116], stage1_45[117], stage1_45[118]},
      {stage1_46[228]},
      {stage1_47[48], stage1_47[49], stage1_47[50], stage1_47[51], stage1_47[52], stage1_47[53]},
      {stage2_49[8],stage2_48[45],stage2_47[57],stage2_46[58],stage2_45[88]}
   );
   gpc615_5 gpc5521 (
      {stage1_45[119], stage1_45[120], stage1_45[121], stage1_45[122], stage1_45[123]},
      {stage1_46[229]},
      {stage1_47[54], stage1_47[55], stage1_47[56], stage1_47[57], stage1_47[58], stage1_47[59]},
      {stage2_49[9],stage2_48[46],stage2_47[58],stage2_46[59],stage2_45[89]}
   );
   gpc615_5 gpc5522 (
      {stage1_45[124], stage1_45[125], stage1_45[126], stage1_45[127], stage1_45[128]},
      {stage1_46[230]},
      {stage1_47[60], stage1_47[61], stage1_47[62], stage1_47[63], stage1_47[64], stage1_47[65]},
      {stage2_49[10],stage2_48[47],stage2_47[59],stage2_46[60],stage2_45[90]}
   );
   gpc615_5 gpc5523 (
      {stage1_45[129], stage1_45[130], stage1_45[131], stage1_45[132], stage1_45[133]},
      {stage1_46[231]},
      {stage1_47[66], stage1_47[67], stage1_47[68], stage1_47[69], stage1_47[70], stage1_47[71]},
      {stage2_49[11],stage2_48[48],stage2_47[60],stage2_46[61],stage2_45[91]}
   );
   gpc615_5 gpc5524 (
      {stage1_45[134], stage1_45[135], stage1_45[136], stage1_45[137], stage1_45[138]},
      {stage1_46[232]},
      {stage1_47[72], stage1_47[73], stage1_47[74], stage1_47[75], stage1_47[76], stage1_47[77]},
      {stage2_49[12],stage2_48[49],stage2_47[61],stage2_46[62],stage2_45[92]}
   );
   gpc615_5 gpc5525 (
      {stage1_45[139], stage1_45[140], stage1_45[141], stage1_45[142], stage1_45[143]},
      {stage1_46[233]},
      {stage1_47[78], stage1_47[79], stage1_47[80], stage1_47[81], stage1_47[82], stage1_47[83]},
      {stage2_49[13],stage2_48[50],stage2_47[62],stage2_46[63],stage2_45[93]}
   );
   gpc615_5 gpc5526 (
      {stage1_45[144], stage1_45[145], stage1_45[146], stage1_45[147], stage1_45[148]},
      {stage1_46[234]},
      {stage1_47[84], stage1_47[85], stage1_47[86], stage1_47[87], stage1_47[88], stage1_47[89]},
      {stage2_49[14],stage2_48[51],stage2_47[63],stage2_46[64],stage2_45[94]}
   );
   gpc615_5 gpc5527 (
      {stage1_45[149], stage1_45[150], stage1_45[151], stage1_45[152], stage1_45[153]},
      {stage1_46[235]},
      {stage1_47[90], stage1_47[91], stage1_47[92], stage1_47[93], stage1_47[94], stage1_47[95]},
      {stage2_49[15],stage2_48[52],stage2_47[64],stage2_46[65],stage2_45[95]}
   );
   gpc615_5 gpc5528 (
      {stage1_45[154], stage1_45[155], stage1_45[156], stage1_45[157], stage1_45[158]},
      {stage1_46[236]},
      {stage1_47[96], stage1_47[97], stage1_47[98], stage1_47[99], stage1_47[100], stage1_47[101]},
      {stage2_49[16],stage2_48[53],stage2_47[65],stage2_46[66],stage2_45[96]}
   );
   gpc615_5 gpc5529 (
      {stage1_45[159], stage1_45[160], stage1_45[161], stage1_45[162], stage1_45[163]},
      {stage1_46[237]},
      {stage1_47[102], stage1_47[103], stage1_47[104], stage1_47[105], stage1_47[106], stage1_47[107]},
      {stage2_49[17],stage2_48[54],stage2_47[66],stage2_46[67],stage2_45[97]}
   );
   gpc615_5 gpc5530 (
      {stage1_45[164], stage1_45[165], stage1_45[166], stage1_45[167], stage1_45[168]},
      {stage1_46[238]},
      {stage1_47[108], stage1_47[109], stage1_47[110], stage1_47[111], stage1_47[112], stage1_47[113]},
      {stage2_49[18],stage2_48[55],stage2_47[67],stage2_46[68],stage2_45[98]}
   );
   gpc615_5 gpc5531 (
      {stage1_45[169], stage1_45[170], stage1_45[171], stage1_45[172], stage1_45[173]},
      {stage1_46[239]},
      {stage1_47[114], stage1_47[115], stage1_47[116], stage1_47[117], stage1_47[118], stage1_47[119]},
      {stage2_49[19],stage2_48[56],stage2_47[68],stage2_46[69],stage2_45[99]}
   );
   gpc615_5 gpc5532 (
      {stage1_45[174], stage1_45[175], stage1_45[176], stage1_45[177], stage1_45[178]},
      {stage1_46[240]},
      {stage1_47[120], stage1_47[121], stage1_47[122], stage1_47[123], stage1_47[124], stage1_47[125]},
      {stage2_49[20],stage2_48[57],stage2_47[69],stage2_46[70],stage2_45[100]}
   );
   gpc615_5 gpc5533 (
      {stage1_45[179], stage1_45[180], stage1_45[181], stage1_45[182], stage1_45[183]},
      {stage1_46[241]},
      {stage1_47[126], stage1_47[127], stage1_47[128], stage1_47[129], stage1_47[130], stage1_47[131]},
      {stage2_49[21],stage2_48[58],stage2_47[70],stage2_46[71],stage2_45[101]}
   );
   gpc615_5 gpc5534 (
      {stage1_45[184], stage1_45[185], stage1_45[186], stage1_45[187], stage1_45[188]},
      {stage1_46[242]},
      {stage1_47[132], stage1_47[133], stage1_47[134], stage1_47[135], stage1_47[136], stage1_47[137]},
      {stage2_49[22],stage2_48[59],stage2_47[71],stage2_46[72],stage2_45[102]}
   );
   gpc615_5 gpc5535 (
      {stage1_45[189], stage1_45[190], stage1_45[191], stage1_45[192], stage1_45[193]},
      {stage1_46[243]},
      {stage1_47[138], stage1_47[139], stage1_47[140], stage1_47[141], stage1_47[142], stage1_47[143]},
      {stage2_49[23],stage2_48[60],stage2_47[72],stage2_46[73],stage2_45[103]}
   );
   gpc615_5 gpc5536 (
      {stage1_45[194], stage1_45[195], stage1_45[196], stage1_45[197], stage1_45[198]},
      {stage1_46[244]},
      {stage1_47[144], stage1_47[145], stage1_47[146], stage1_47[147], stage1_47[148], stage1_47[149]},
      {stage2_49[24],stage2_48[61],stage2_47[73],stage2_46[74],stage2_45[104]}
   );
   gpc615_5 gpc5537 (
      {stage1_46[245], stage1_46[246], stage1_46[247], stage1_46[248], stage1_46[249]},
      {stage1_47[150]},
      {stage1_48[0], stage1_48[1], stage1_48[2], stage1_48[3], stage1_48[4], stage1_48[5]},
      {stage2_50[0],stage2_49[25],stage2_48[62],stage2_47[74],stage2_46[75]}
   );
   gpc615_5 gpc5538 (
      {stage1_46[250], stage1_46[251], stage1_46[252], stage1_46[253], stage1_46[254]},
      {stage1_47[151]},
      {stage1_48[6], stage1_48[7], stage1_48[8], stage1_48[9], stage1_48[10], stage1_48[11]},
      {stage2_50[1],stage2_49[26],stage2_48[63],stage2_47[75],stage2_46[76]}
   );
   gpc615_5 gpc5539 (
      {stage1_46[255], stage1_46[256], stage1_46[257], stage1_46[258], stage1_46[259]},
      {stage1_47[152]},
      {stage1_48[12], stage1_48[13], stage1_48[14], stage1_48[15], stage1_48[16], stage1_48[17]},
      {stage2_50[2],stage2_49[27],stage2_48[64],stage2_47[76],stage2_46[77]}
   );
   gpc615_5 gpc5540 (
      {stage1_46[260], stage1_46[261], stage1_46[262], stage1_46[263], stage1_46[264]},
      {stage1_47[153]},
      {stage1_48[18], stage1_48[19], stage1_48[20], stage1_48[21], stage1_48[22], stage1_48[23]},
      {stage2_50[3],stage2_49[28],stage2_48[65],stage2_47[77],stage2_46[78]}
   );
   gpc615_5 gpc5541 (
      {stage1_46[265], stage1_46[266], stage1_46[267], stage1_46[268], stage1_46[269]},
      {stage1_47[154]},
      {stage1_48[24], stage1_48[25], stage1_48[26], stage1_48[27], stage1_48[28], stage1_48[29]},
      {stage2_50[4],stage2_49[29],stage2_48[66],stage2_47[78],stage2_46[79]}
   );
   gpc615_5 gpc5542 (
      {stage1_46[270], stage1_46[271], stage1_46[272], stage1_46[273], stage1_46[274]},
      {stage1_47[155]},
      {stage1_48[30], stage1_48[31], stage1_48[32], stage1_48[33], stage1_48[34], stage1_48[35]},
      {stage2_50[5],stage2_49[30],stage2_48[67],stage2_47[79],stage2_46[80]}
   );
   gpc615_5 gpc5543 (
      {stage1_46[275], stage1_46[276], stage1_46[277], stage1_46[278], stage1_46[279]},
      {stage1_47[156]},
      {stage1_48[36], stage1_48[37], stage1_48[38], stage1_48[39], stage1_48[40], stage1_48[41]},
      {stage2_50[6],stage2_49[31],stage2_48[68],stage2_47[80],stage2_46[81]}
   );
   gpc615_5 gpc5544 (
      {stage1_46[280], stage1_46[281], stage1_46[282], stage1_46[283], stage1_46[284]},
      {stage1_47[157]},
      {stage1_48[42], stage1_48[43], stage1_48[44], stage1_48[45], stage1_48[46], stage1_48[47]},
      {stage2_50[7],stage2_49[32],stage2_48[69],stage2_47[81],stage2_46[82]}
   );
   gpc615_5 gpc5545 (
      {stage1_46[285], stage1_46[286], stage1_46[287], stage1_46[288], stage1_46[289]},
      {stage1_47[158]},
      {stage1_48[48], stage1_48[49], stage1_48[50], stage1_48[51], stage1_48[52], stage1_48[53]},
      {stage2_50[8],stage2_49[33],stage2_48[70],stage2_47[82],stage2_46[83]}
   );
   gpc615_5 gpc5546 (
      {stage1_46[290], stage1_46[291], stage1_46[292], stage1_46[293], stage1_46[294]},
      {stage1_47[159]},
      {stage1_48[54], stage1_48[55], stage1_48[56], stage1_48[57], stage1_48[58], stage1_48[59]},
      {stage2_50[9],stage2_49[34],stage2_48[71],stage2_47[83],stage2_46[84]}
   );
   gpc615_5 gpc5547 (
      {stage1_47[160], stage1_47[161], stage1_47[162], stage1_47[163], stage1_47[164]},
      {stage1_48[60]},
      {stage1_49[0], stage1_49[1], stage1_49[2], stage1_49[3], stage1_49[4], stage1_49[5]},
      {stage2_51[0],stage2_50[10],stage2_49[35],stage2_48[72],stage2_47[84]}
   );
   gpc615_5 gpc5548 (
      {stage1_47[165], stage1_47[166], stage1_47[167], stage1_47[168], stage1_47[169]},
      {stage1_48[61]},
      {stage1_49[6], stage1_49[7], stage1_49[8], stage1_49[9], stage1_49[10], stage1_49[11]},
      {stage2_51[1],stage2_50[11],stage2_49[36],stage2_48[73],stage2_47[85]}
   );
   gpc615_5 gpc5549 (
      {stage1_47[170], stage1_47[171], stage1_47[172], stage1_47[173], stage1_47[174]},
      {stage1_48[62]},
      {stage1_49[12], stage1_49[13], stage1_49[14], stage1_49[15], stage1_49[16], stage1_49[17]},
      {stage2_51[2],stage2_50[12],stage2_49[37],stage2_48[74],stage2_47[86]}
   );
   gpc615_5 gpc5550 (
      {stage1_47[175], stage1_47[176], stage1_47[177], stage1_47[178], stage1_47[179]},
      {stage1_48[63]},
      {stage1_49[18], stage1_49[19], stage1_49[20], stage1_49[21], stage1_49[22], stage1_49[23]},
      {stage2_51[3],stage2_50[13],stage2_49[38],stage2_48[75],stage2_47[87]}
   );
   gpc615_5 gpc5551 (
      {stage1_47[180], stage1_47[181], stage1_47[182], stage1_47[183], stage1_47[184]},
      {stage1_48[64]},
      {stage1_49[24], stage1_49[25], stage1_49[26], stage1_49[27], stage1_49[28], stage1_49[29]},
      {stage2_51[4],stage2_50[14],stage2_49[39],stage2_48[76],stage2_47[88]}
   );
   gpc615_5 gpc5552 (
      {stage1_47[185], stage1_47[186], stage1_47[187], stage1_47[188], stage1_47[189]},
      {stage1_48[65]},
      {stage1_49[30], stage1_49[31], stage1_49[32], stage1_49[33], stage1_49[34], stage1_49[35]},
      {stage2_51[5],stage2_50[15],stage2_49[40],stage2_48[77],stage2_47[89]}
   );
   gpc615_5 gpc5553 (
      {stage1_47[190], stage1_47[191], stage1_47[192], stage1_47[193], stage1_47[194]},
      {stage1_48[66]},
      {stage1_49[36], stage1_49[37], stage1_49[38], stage1_49[39], stage1_49[40], stage1_49[41]},
      {stage2_51[6],stage2_50[16],stage2_49[41],stage2_48[78],stage2_47[90]}
   );
   gpc615_5 gpc5554 (
      {stage1_47[195], stage1_47[196], stage1_47[197], stage1_47[198], stage1_47[199]},
      {stage1_48[67]},
      {stage1_49[42], stage1_49[43], stage1_49[44], stage1_49[45], stage1_49[46], stage1_49[47]},
      {stage2_51[7],stage2_50[17],stage2_49[42],stage2_48[79],stage2_47[91]}
   );
   gpc615_5 gpc5555 (
      {stage1_47[200], stage1_47[201], stage1_47[202], stage1_47[203], stage1_47[204]},
      {stage1_48[68]},
      {stage1_49[48], stage1_49[49], stage1_49[50], stage1_49[51], stage1_49[52], stage1_49[53]},
      {stage2_51[8],stage2_50[18],stage2_49[43],stage2_48[80],stage2_47[92]}
   );
   gpc615_5 gpc5556 (
      {stage1_47[205], stage1_47[206], stage1_47[207], stage1_47[208], stage1_47[209]},
      {stage1_48[69]},
      {stage1_49[54], stage1_49[55], stage1_49[56], stage1_49[57], stage1_49[58], stage1_49[59]},
      {stage2_51[9],stage2_50[19],stage2_49[44],stage2_48[81],stage2_47[93]}
   );
   gpc615_5 gpc5557 (
      {stage1_47[210], stage1_47[211], stage1_47[212], stage1_47[213], stage1_47[214]},
      {stage1_48[70]},
      {stage1_49[60], stage1_49[61], stage1_49[62], stage1_49[63], stage1_49[64], stage1_49[65]},
      {stage2_51[10],stage2_50[20],stage2_49[45],stage2_48[82],stage2_47[94]}
   );
   gpc615_5 gpc5558 (
      {stage1_47[215], stage1_47[216], stage1_47[217], stage1_47[218], stage1_47[219]},
      {stage1_48[71]},
      {stage1_49[66], stage1_49[67], stage1_49[68], stage1_49[69], stage1_49[70], stage1_49[71]},
      {stage2_51[11],stage2_50[21],stage2_49[46],stage2_48[83],stage2_47[95]}
   );
   gpc615_5 gpc5559 (
      {stage1_47[220], stage1_47[221], stage1_47[222], stage1_47[223], stage1_47[224]},
      {stage1_48[72]},
      {stage1_49[72], stage1_49[73], stage1_49[74], stage1_49[75], stage1_49[76], stage1_49[77]},
      {stage2_51[12],stage2_50[22],stage2_49[47],stage2_48[84],stage2_47[96]}
   );
   gpc615_5 gpc5560 (
      {stage1_47[225], stage1_47[226], stage1_47[227], stage1_47[228], stage1_47[229]},
      {stage1_48[73]},
      {stage1_49[78], stage1_49[79], stage1_49[80], stage1_49[81], stage1_49[82], stage1_49[83]},
      {stage2_51[13],stage2_50[23],stage2_49[48],stage2_48[85],stage2_47[97]}
   );
   gpc606_5 gpc5561 (
      {stage1_48[74], stage1_48[75], stage1_48[76], stage1_48[77], stage1_48[78], stage1_48[79]},
      {stage1_50[0], stage1_50[1], stage1_50[2], stage1_50[3], stage1_50[4], stage1_50[5]},
      {stage2_52[0],stage2_51[14],stage2_50[24],stage2_49[49],stage2_48[86]}
   );
   gpc606_5 gpc5562 (
      {stage1_48[80], stage1_48[81], stage1_48[82], stage1_48[83], stage1_48[84], stage1_48[85]},
      {stage1_50[6], stage1_50[7], stage1_50[8], stage1_50[9], stage1_50[10], stage1_50[11]},
      {stage2_52[1],stage2_51[15],stage2_50[25],stage2_49[50],stage2_48[87]}
   );
   gpc606_5 gpc5563 (
      {stage1_48[86], stage1_48[87], stage1_48[88], stage1_48[89], stage1_48[90], stage1_48[91]},
      {stage1_50[12], stage1_50[13], stage1_50[14], stage1_50[15], stage1_50[16], stage1_50[17]},
      {stage2_52[2],stage2_51[16],stage2_50[26],stage2_49[51],stage2_48[88]}
   );
   gpc606_5 gpc5564 (
      {stage1_48[92], stage1_48[93], stage1_48[94], stage1_48[95], stage1_48[96], stage1_48[97]},
      {stage1_50[18], stage1_50[19], stage1_50[20], stage1_50[21], stage1_50[22], stage1_50[23]},
      {stage2_52[3],stage2_51[17],stage2_50[27],stage2_49[52],stage2_48[89]}
   );
   gpc606_5 gpc5565 (
      {stage1_48[98], stage1_48[99], stage1_48[100], stage1_48[101], stage1_48[102], stage1_48[103]},
      {stage1_50[24], stage1_50[25], stage1_50[26], stage1_50[27], stage1_50[28], stage1_50[29]},
      {stage2_52[4],stage2_51[18],stage2_50[28],stage2_49[53],stage2_48[90]}
   );
   gpc606_5 gpc5566 (
      {stage1_48[104], stage1_48[105], stage1_48[106], stage1_48[107], stage1_48[108], stage1_48[109]},
      {stage1_50[30], stage1_50[31], stage1_50[32], stage1_50[33], stage1_50[34], stage1_50[35]},
      {stage2_52[5],stage2_51[19],stage2_50[29],stage2_49[54],stage2_48[91]}
   );
   gpc606_5 gpc5567 (
      {stage1_48[110], stage1_48[111], stage1_48[112], stage1_48[113], stage1_48[114], stage1_48[115]},
      {stage1_50[36], stage1_50[37], stage1_50[38], stage1_50[39], stage1_50[40], stage1_50[41]},
      {stage2_52[6],stage2_51[20],stage2_50[30],stage2_49[55],stage2_48[92]}
   );
   gpc606_5 gpc5568 (
      {stage1_48[116], stage1_48[117], stage1_48[118], stage1_48[119], stage1_48[120], stage1_48[121]},
      {stage1_50[42], stage1_50[43], stage1_50[44], stage1_50[45], stage1_50[46], stage1_50[47]},
      {stage2_52[7],stage2_51[21],stage2_50[31],stage2_49[56],stage2_48[93]}
   );
   gpc615_5 gpc5569 (
      {stage1_48[122], stage1_48[123], stage1_48[124], stage1_48[125], stage1_48[126]},
      {stage1_49[84]},
      {stage1_50[48], stage1_50[49], stage1_50[50], stage1_50[51], stage1_50[52], stage1_50[53]},
      {stage2_52[8],stage2_51[22],stage2_50[32],stage2_49[57],stage2_48[94]}
   );
   gpc615_5 gpc5570 (
      {stage1_48[127], stage1_48[128], stage1_48[129], stage1_48[130], stage1_48[131]},
      {stage1_49[85]},
      {stage1_50[54], stage1_50[55], stage1_50[56], stage1_50[57], stage1_50[58], stage1_50[59]},
      {stage2_52[9],stage2_51[23],stage2_50[33],stage2_49[58],stage2_48[95]}
   );
   gpc615_5 gpc5571 (
      {stage1_48[132], stage1_48[133], stage1_48[134], stage1_48[135], stage1_48[136]},
      {stage1_49[86]},
      {stage1_50[60], stage1_50[61], stage1_50[62], stage1_50[63], stage1_50[64], stage1_50[65]},
      {stage2_52[10],stage2_51[24],stage2_50[34],stage2_49[59],stage2_48[96]}
   );
   gpc615_5 gpc5572 (
      {stage1_48[137], stage1_48[138], stage1_48[139], stage1_48[140], stage1_48[141]},
      {stage1_49[87]},
      {stage1_50[66], stage1_50[67], stage1_50[68], stage1_50[69], stage1_50[70], stage1_50[71]},
      {stage2_52[11],stage2_51[25],stage2_50[35],stage2_49[60],stage2_48[97]}
   );
   gpc615_5 gpc5573 (
      {stage1_48[142], stage1_48[143], stage1_48[144], stage1_48[145], stage1_48[146]},
      {stage1_49[88]},
      {stage1_50[72], stage1_50[73], stage1_50[74], stage1_50[75], stage1_50[76], stage1_50[77]},
      {stage2_52[12],stage2_51[26],stage2_50[36],stage2_49[61],stage2_48[98]}
   );
   gpc615_5 gpc5574 (
      {stage1_48[147], stage1_48[148], stage1_48[149], stage1_48[150], stage1_48[151]},
      {stage1_49[89]},
      {stage1_50[78], stage1_50[79], stage1_50[80], stage1_50[81], stage1_50[82], stage1_50[83]},
      {stage2_52[13],stage2_51[27],stage2_50[37],stage2_49[62],stage2_48[99]}
   );
   gpc615_5 gpc5575 (
      {stage1_48[152], stage1_48[153], stage1_48[154], stage1_48[155], stage1_48[156]},
      {stage1_49[90]},
      {stage1_50[84], stage1_50[85], stage1_50[86], stage1_50[87], stage1_50[88], stage1_50[89]},
      {stage2_52[14],stage2_51[28],stage2_50[38],stage2_49[63],stage2_48[100]}
   );
   gpc615_5 gpc5576 (
      {stage1_48[157], stage1_48[158], stage1_48[159], stage1_48[160], stage1_48[161]},
      {stage1_49[91]},
      {stage1_50[90], stage1_50[91], stage1_50[92], stage1_50[93], stage1_50[94], stage1_50[95]},
      {stage2_52[15],stage2_51[29],stage2_50[39],stage2_49[64],stage2_48[101]}
   );
   gpc615_5 gpc5577 (
      {stage1_48[162], stage1_48[163], stage1_48[164], stage1_48[165], stage1_48[166]},
      {stage1_49[92]},
      {stage1_50[96], stage1_50[97], stage1_50[98], stage1_50[99], stage1_50[100], stage1_50[101]},
      {stage2_52[16],stage2_51[30],stage2_50[40],stage2_49[65],stage2_48[102]}
   );
   gpc615_5 gpc5578 (
      {stage1_48[167], stage1_48[168], stage1_48[169], stage1_48[170], stage1_48[171]},
      {stage1_49[93]},
      {stage1_50[102], stage1_50[103], stage1_50[104], stage1_50[105], stage1_50[106], stage1_50[107]},
      {stage2_52[17],stage2_51[31],stage2_50[41],stage2_49[66],stage2_48[103]}
   );
   gpc606_5 gpc5579 (
      {stage1_49[94], stage1_49[95], stage1_49[96], stage1_49[97], stage1_49[98], stage1_49[99]},
      {stage1_51[0], stage1_51[1], stage1_51[2], stage1_51[3], stage1_51[4], stage1_51[5]},
      {stage2_53[0],stage2_52[18],stage2_51[32],stage2_50[42],stage2_49[67]}
   );
   gpc606_5 gpc5580 (
      {stage1_49[100], stage1_49[101], stage1_49[102], stage1_49[103], stage1_49[104], stage1_49[105]},
      {stage1_51[6], stage1_51[7], stage1_51[8], stage1_51[9], stage1_51[10], stage1_51[11]},
      {stage2_53[1],stage2_52[19],stage2_51[33],stage2_50[43],stage2_49[68]}
   );
   gpc606_5 gpc5581 (
      {stage1_49[106], stage1_49[107], stage1_49[108], stage1_49[109], stage1_49[110], stage1_49[111]},
      {stage1_51[12], stage1_51[13], stage1_51[14], stage1_51[15], stage1_51[16], stage1_51[17]},
      {stage2_53[2],stage2_52[20],stage2_51[34],stage2_50[44],stage2_49[69]}
   );
   gpc606_5 gpc5582 (
      {stage1_49[112], stage1_49[113], stage1_49[114], stage1_49[115], stage1_49[116], stage1_49[117]},
      {stage1_51[18], stage1_51[19], stage1_51[20], stage1_51[21], stage1_51[22], stage1_51[23]},
      {stage2_53[3],stage2_52[21],stage2_51[35],stage2_50[45],stage2_49[70]}
   );
   gpc606_5 gpc5583 (
      {stage1_49[118], stage1_49[119], stage1_49[120], stage1_49[121], stage1_49[122], stage1_49[123]},
      {stage1_51[24], stage1_51[25], stage1_51[26], stage1_51[27], stage1_51[28], stage1_51[29]},
      {stage2_53[4],stage2_52[22],stage2_51[36],stage2_50[46],stage2_49[71]}
   );
   gpc606_5 gpc5584 (
      {stage1_49[124], stage1_49[125], stage1_49[126], stage1_49[127], stage1_49[128], stage1_49[129]},
      {stage1_51[30], stage1_51[31], stage1_51[32], stage1_51[33], stage1_51[34], stage1_51[35]},
      {stage2_53[5],stage2_52[23],stage2_51[37],stage2_50[47],stage2_49[72]}
   );
   gpc606_5 gpc5585 (
      {stage1_49[130], stage1_49[131], stage1_49[132], stage1_49[133], stage1_49[134], stage1_49[135]},
      {stage1_51[36], stage1_51[37], stage1_51[38], stage1_51[39], stage1_51[40], stage1_51[41]},
      {stage2_53[6],stage2_52[24],stage2_51[38],stage2_50[48],stage2_49[73]}
   );
   gpc606_5 gpc5586 (
      {stage1_49[136], stage1_49[137], stage1_49[138], stage1_49[139], stage1_49[140], stage1_49[141]},
      {stage1_51[42], stage1_51[43], stage1_51[44], stage1_51[45], stage1_51[46], stage1_51[47]},
      {stage2_53[7],stage2_52[25],stage2_51[39],stage2_50[49],stage2_49[74]}
   );
   gpc606_5 gpc5587 (
      {stage1_49[142], stage1_49[143], stage1_49[144], stage1_49[145], stage1_49[146], stage1_49[147]},
      {stage1_51[48], stage1_51[49], stage1_51[50], stage1_51[51], stage1_51[52], stage1_51[53]},
      {stage2_53[8],stage2_52[26],stage2_51[40],stage2_50[50],stage2_49[75]}
   );
   gpc606_5 gpc5588 (
      {stage1_49[148], stage1_49[149], stage1_49[150], stage1_49[151], stage1_49[152], stage1_49[153]},
      {stage1_51[54], stage1_51[55], stage1_51[56], stage1_51[57], stage1_51[58], stage1_51[59]},
      {stage2_53[9],stage2_52[27],stage2_51[41],stage2_50[51],stage2_49[76]}
   );
   gpc2135_5 gpc5589 (
      {stage1_50[108], stage1_50[109], stage1_50[110], stage1_50[111], stage1_50[112]},
      {stage1_51[60], stage1_51[61], stage1_51[62]},
      {stage1_52[0]},
      {stage1_53[0], stage1_53[1]},
      {stage2_54[0],stage2_53[10],stage2_52[28],stage2_51[42],stage2_50[52]}
   );
   gpc1163_5 gpc5590 (
      {stage1_50[113], stage1_50[114], stage1_50[115]},
      {stage1_51[63], stage1_51[64], stage1_51[65], stage1_51[66], stage1_51[67], stage1_51[68]},
      {stage1_52[1]},
      {stage1_53[2]},
      {stage2_54[1],stage2_53[11],stage2_52[29],stage2_51[43],stage2_50[53]}
   );
   gpc1163_5 gpc5591 (
      {stage1_50[116], stage1_50[117], stage1_50[118]},
      {stage1_51[69], stage1_51[70], stage1_51[71], stage1_51[72], stage1_51[73], stage1_51[74]},
      {stage1_52[2]},
      {stage1_53[3]},
      {stage2_54[2],stage2_53[12],stage2_52[30],stage2_51[44],stage2_50[54]}
   );
   gpc1163_5 gpc5592 (
      {stage1_50[119], stage1_50[120], stage1_50[121]},
      {stage1_51[75], stage1_51[76], stage1_51[77], stage1_51[78], stage1_51[79], stage1_51[80]},
      {stage1_52[3]},
      {stage1_53[4]},
      {stage2_54[3],stage2_53[13],stage2_52[31],stage2_51[45],stage2_50[55]}
   );
   gpc1163_5 gpc5593 (
      {stage1_50[122], stage1_50[123], stage1_50[124]},
      {stage1_51[81], stage1_51[82], stage1_51[83], stage1_51[84], stage1_51[85], stage1_51[86]},
      {stage1_52[4]},
      {stage1_53[5]},
      {stage2_54[4],stage2_53[14],stage2_52[32],stage2_51[46],stage2_50[56]}
   );
   gpc1163_5 gpc5594 (
      {stage1_50[125], stage1_50[126], stage1_50[127]},
      {stage1_51[87], stage1_51[88], stage1_51[89], stage1_51[90], stage1_51[91], stage1_51[92]},
      {stage1_52[5]},
      {stage1_53[6]},
      {stage2_54[5],stage2_53[15],stage2_52[33],stage2_51[47],stage2_50[57]}
   );
   gpc1163_5 gpc5595 (
      {stage1_50[128], stage1_50[129], stage1_50[130]},
      {stage1_51[93], stage1_51[94], stage1_51[95], stage1_51[96], stage1_51[97], stage1_51[98]},
      {stage1_52[6]},
      {stage1_53[7]},
      {stage2_54[6],stage2_53[16],stage2_52[34],stage2_51[48],stage2_50[58]}
   );
   gpc1163_5 gpc5596 (
      {stage1_50[131], stage1_50[132], stage1_50[133]},
      {stage1_51[99], stage1_51[100], stage1_51[101], stage1_51[102], stage1_51[103], stage1_51[104]},
      {stage1_52[7]},
      {stage1_53[8]},
      {stage2_54[7],stage2_53[17],stage2_52[35],stage2_51[49],stage2_50[59]}
   );
   gpc1163_5 gpc5597 (
      {stage1_50[134], stage1_50[135], stage1_50[136]},
      {stage1_51[105], stage1_51[106], stage1_51[107], stage1_51[108], stage1_51[109], stage1_51[110]},
      {stage1_52[8]},
      {stage1_53[9]},
      {stage2_54[8],stage2_53[18],stage2_52[36],stage2_51[50],stage2_50[60]}
   );
   gpc1163_5 gpc5598 (
      {stage1_50[137], stage1_50[138], stage1_50[139]},
      {stage1_51[111], stage1_51[112], stage1_51[113], stage1_51[114], stage1_51[115], stage1_51[116]},
      {stage1_52[9]},
      {stage1_53[10]},
      {stage2_54[9],stage2_53[19],stage2_52[37],stage2_51[51],stage2_50[61]}
   );
   gpc1163_5 gpc5599 (
      {stage1_50[140], stage1_50[141], stage1_50[142]},
      {stage1_51[117], stage1_51[118], stage1_51[119], stage1_51[120], stage1_51[121], stage1_51[122]},
      {stage1_52[10]},
      {stage1_53[11]},
      {stage2_54[10],stage2_53[20],stage2_52[38],stage2_51[52],stage2_50[62]}
   );
   gpc1163_5 gpc5600 (
      {stage1_50[143], stage1_50[144], stage1_50[145]},
      {stage1_51[123], stage1_51[124], stage1_51[125], stage1_51[126], stage1_51[127], stage1_51[128]},
      {stage1_52[11]},
      {stage1_53[12]},
      {stage2_54[11],stage2_53[21],stage2_52[39],stage2_51[53],stage2_50[63]}
   );
   gpc1163_5 gpc5601 (
      {stage1_50[146], stage1_50[147], stage1_50[148]},
      {stage1_51[129], stage1_51[130], stage1_51[131], stage1_51[132], stage1_51[133], stage1_51[134]},
      {stage1_52[12]},
      {stage1_53[13]},
      {stage2_54[12],stage2_53[22],stage2_52[40],stage2_51[54],stage2_50[64]}
   );
   gpc1163_5 gpc5602 (
      {stage1_50[149], stage1_50[150], stage1_50[151]},
      {stage1_51[135], stage1_51[136], stage1_51[137], stage1_51[138], stage1_51[139], stage1_51[140]},
      {stage1_52[13]},
      {stage1_53[14]},
      {stage2_54[13],stage2_53[23],stage2_52[41],stage2_51[55],stage2_50[65]}
   );
   gpc1163_5 gpc5603 (
      {stage1_50[152], stage1_50[153], stage1_50[154]},
      {stage1_51[141], stage1_51[142], stage1_51[143], stage1_51[144], stage1_51[145], stage1_51[146]},
      {stage1_52[14]},
      {stage1_53[15]},
      {stage2_54[14],stage2_53[24],stage2_52[42],stage2_51[56],stage2_50[66]}
   );
   gpc1163_5 gpc5604 (
      {stage1_50[155], stage1_50[156], stage1_50[157]},
      {stage1_51[147], stage1_51[148], stage1_51[149], stage1_51[150], stage1_51[151], stage1_51[152]},
      {stage1_52[15]},
      {stage1_53[16]},
      {stage2_54[15],stage2_53[25],stage2_52[43],stage2_51[57],stage2_50[67]}
   );
   gpc1163_5 gpc5605 (
      {stage1_50[158], stage1_50[159], stage1_50[160]},
      {stage1_51[153], stage1_51[154], stage1_51[155], stage1_51[156], stage1_51[157], stage1_51[158]},
      {stage1_52[16]},
      {stage1_53[17]},
      {stage2_54[16],stage2_53[26],stage2_52[44],stage2_51[58],stage2_50[68]}
   );
   gpc1163_5 gpc5606 (
      {stage1_50[161], stage1_50[162], stage1_50[163]},
      {stage1_51[159], stage1_51[160], stage1_51[161], stage1_51[162], stage1_51[163], stage1_51[164]},
      {stage1_52[17]},
      {stage1_53[18]},
      {stage2_54[17],stage2_53[27],stage2_52[45],stage2_51[59],stage2_50[69]}
   );
   gpc1163_5 gpc5607 (
      {stage1_50[164], stage1_50[165], stage1_50[166]},
      {stage1_51[165], stage1_51[166], stage1_51[167], stage1_51[168], stage1_51[169], stage1_51[170]},
      {stage1_52[18]},
      {stage1_53[19]},
      {stage2_54[18],stage2_53[28],stage2_52[46],stage2_51[60],stage2_50[70]}
   );
   gpc1163_5 gpc5608 (
      {stage1_50[167], stage1_50[168], stage1_50[169]},
      {stage1_51[171], stage1_51[172], stage1_51[173], stage1_51[174], stage1_51[175], stage1_51[176]},
      {stage1_52[19]},
      {stage1_53[20]},
      {stage2_54[19],stage2_53[29],stage2_52[47],stage2_51[61],stage2_50[71]}
   );
   gpc1163_5 gpc5609 (
      {stage1_50[170], stage1_50[171], stage1_50[172]},
      {stage1_51[177], stage1_51[178], stage1_51[179], stage1_51[180], stage1_51[181], stage1_51[182]},
      {stage1_52[20]},
      {stage1_53[21]},
      {stage2_54[20],stage2_53[30],stage2_52[48],stage2_51[62],stage2_50[72]}
   );
   gpc1163_5 gpc5610 (
      {stage1_50[173], stage1_50[174], stage1_50[175]},
      {stage1_51[183], stage1_51[184], stage1_51[185], stage1_51[186], stage1_51[187], stage1_51[188]},
      {stage1_52[21]},
      {stage1_53[22]},
      {stage2_54[21],stage2_53[31],stage2_52[49],stage2_51[63],stage2_50[73]}
   );
   gpc1163_5 gpc5611 (
      {stage1_50[176], stage1_50[177], stage1_50[178]},
      {stage1_51[189], stage1_51[190], stage1_51[191], stage1_51[192], stage1_51[193], stage1_51[194]},
      {stage1_52[22]},
      {stage1_53[23]},
      {stage2_54[22],stage2_53[32],stage2_52[50],stage2_51[64],stage2_50[74]}
   );
   gpc606_5 gpc5612 (
      {stage1_51[195], stage1_51[196], stage1_51[197], stage1_51[198], stage1_51[199], stage1_51[200]},
      {stage1_53[24], stage1_53[25], stage1_53[26], stage1_53[27], stage1_53[28], stage1_53[29]},
      {stage2_55[0],stage2_54[23],stage2_53[33],stage2_52[51],stage2_51[65]}
   );
   gpc615_5 gpc5613 (
      {stage1_51[201], stage1_51[202], stage1_51[203], stage1_51[204], stage1_51[205]},
      {stage1_52[23]},
      {stage1_53[30], stage1_53[31], stage1_53[32], stage1_53[33], stage1_53[34], stage1_53[35]},
      {stage2_55[1],stage2_54[24],stage2_53[34],stage2_52[52],stage2_51[66]}
   );
   gpc615_5 gpc5614 (
      {stage1_51[206], stage1_51[207], stage1_51[208], stage1_51[209], stage1_51[210]},
      {stage1_52[24]},
      {stage1_53[36], stage1_53[37], stage1_53[38], stage1_53[39], stage1_53[40], stage1_53[41]},
      {stage2_55[2],stage2_54[25],stage2_53[35],stage2_52[53],stage2_51[67]}
   );
   gpc615_5 gpc5615 (
      {stage1_51[211], stage1_51[212], stage1_51[213], stage1_51[214], stage1_51[215]},
      {stage1_52[25]},
      {stage1_53[42], stage1_53[43], stage1_53[44], stage1_53[45], stage1_53[46], stage1_53[47]},
      {stage2_55[3],stage2_54[26],stage2_53[36],stage2_52[54],stage2_51[68]}
   );
   gpc615_5 gpc5616 (
      {stage1_51[216], stage1_51[217], stage1_51[218], stage1_51[219], stage1_51[220]},
      {stage1_52[26]},
      {stage1_53[48], stage1_53[49], stage1_53[50], stage1_53[51], stage1_53[52], stage1_53[53]},
      {stage2_55[4],stage2_54[27],stage2_53[37],stage2_52[55],stage2_51[69]}
   );
   gpc615_5 gpc5617 (
      {stage1_51[221], stage1_51[222], stage1_51[223], stage1_51[224], stage1_51[225]},
      {stage1_52[27]},
      {stage1_53[54], stage1_53[55], stage1_53[56], stage1_53[57], stage1_53[58], stage1_53[59]},
      {stage2_55[5],stage2_54[28],stage2_53[38],stage2_52[56],stage2_51[70]}
   );
   gpc615_5 gpc5618 (
      {stage1_51[226], stage1_51[227], stage1_51[228], stage1_51[229], stage1_51[230]},
      {stage1_52[28]},
      {stage1_53[60], stage1_53[61], stage1_53[62], stage1_53[63], stage1_53[64], stage1_53[65]},
      {stage2_55[6],stage2_54[29],stage2_53[39],stage2_52[57],stage2_51[71]}
   );
   gpc615_5 gpc5619 (
      {stage1_51[231], stage1_51[232], stage1_51[233], stage1_51[234], stage1_51[235]},
      {stage1_52[29]},
      {stage1_53[66], stage1_53[67], stage1_53[68], stage1_53[69], stage1_53[70], stage1_53[71]},
      {stage2_55[7],stage2_54[30],stage2_53[40],stage2_52[58],stage2_51[72]}
   );
   gpc615_5 gpc5620 (
      {stage1_51[236], stage1_51[237], stage1_51[238], stage1_51[239], stage1_51[240]},
      {stage1_52[30]},
      {stage1_53[72], stage1_53[73], stage1_53[74], stage1_53[75], stage1_53[76], stage1_53[77]},
      {stage2_55[8],stage2_54[31],stage2_53[41],stage2_52[59],stage2_51[73]}
   );
   gpc615_5 gpc5621 (
      {stage1_51[241], stage1_51[242], stage1_51[243], stage1_51[244], stage1_51[245]},
      {stage1_52[31]},
      {stage1_53[78], stage1_53[79], stage1_53[80], stage1_53[81], stage1_53[82], stage1_53[83]},
      {stage2_55[9],stage2_54[32],stage2_53[42],stage2_52[60],stage2_51[74]}
   );
   gpc615_5 gpc5622 (
      {stage1_51[246], stage1_51[247], stage1_51[248], stage1_51[249], stage1_51[250]},
      {stage1_52[32]},
      {stage1_53[84], stage1_53[85], stage1_53[86], stage1_53[87], stage1_53[88], stage1_53[89]},
      {stage2_55[10],stage2_54[33],stage2_53[43],stage2_52[61],stage2_51[75]}
   );
   gpc615_5 gpc5623 (
      {stage1_51[251], stage1_51[252], stage1_51[253], stage1_51[254], stage1_51[255]},
      {stage1_52[33]},
      {stage1_53[90], stage1_53[91], stage1_53[92], stage1_53[93], stage1_53[94], stage1_53[95]},
      {stage2_55[11],stage2_54[34],stage2_53[44],stage2_52[62],stage2_51[76]}
   );
   gpc615_5 gpc5624 (
      {stage1_51[256], stage1_51[257], stage1_51[258], stage1_51[259], stage1_51[260]},
      {stage1_52[34]},
      {stage1_53[96], stage1_53[97], stage1_53[98], stage1_53[99], stage1_53[100], stage1_53[101]},
      {stage2_55[12],stage2_54[35],stage2_53[45],stage2_52[63],stage2_51[77]}
   );
   gpc615_5 gpc5625 (
      {stage1_51[261], stage1_51[262], stage1_51[263], stage1_51[264], stage1_51[265]},
      {stage1_52[35]},
      {stage1_53[102], stage1_53[103], stage1_53[104], stage1_53[105], stage1_53[106], stage1_53[107]},
      {stage2_55[13],stage2_54[36],stage2_53[46],stage2_52[64],stage2_51[78]}
   );
   gpc606_5 gpc5626 (
      {stage1_52[36], stage1_52[37], stage1_52[38], stage1_52[39], stage1_52[40], stage1_52[41]},
      {stage1_54[0], stage1_54[1], stage1_54[2], stage1_54[3], stage1_54[4], stage1_54[5]},
      {stage2_56[0],stage2_55[14],stage2_54[37],stage2_53[47],stage2_52[65]}
   );
   gpc606_5 gpc5627 (
      {stage1_52[42], stage1_52[43], stage1_52[44], stage1_52[45], stage1_52[46], stage1_52[47]},
      {stage1_54[6], stage1_54[7], stage1_54[8], stage1_54[9], stage1_54[10], stage1_54[11]},
      {stage2_56[1],stage2_55[15],stage2_54[38],stage2_53[48],stage2_52[66]}
   );
   gpc606_5 gpc5628 (
      {stage1_52[48], stage1_52[49], stage1_52[50], stage1_52[51], stage1_52[52], stage1_52[53]},
      {stage1_54[12], stage1_54[13], stage1_54[14], stage1_54[15], stage1_54[16], stage1_54[17]},
      {stage2_56[2],stage2_55[16],stage2_54[39],stage2_53[49],stage2_52[67]}
   );
   gpc606_5 gpc5629 (
      {stage1_52[54], stage1_52[55], stage1_52[56], stage1_52[57], stage1_52[58], stage1_52[59]},
      {stage1_54[18], stage1_54[19], stage1_54[20], stage1_54[21], stage1_54[22], stage1_54[23]},
      {stage2_56[3],stage2_55[17],stage2_54[40],stage2_53[50],stage2_52[68]}
   );
   gpc606_5 gpc5630 (
      {stage1_52[60], stage1_52[61], stage1_52[62], stage1_52[63], stage1_52[64], stage1_52[65]},
      {stage1_54[24], stage1_54[25], stage1_54[26], stage1_54[27], stage1_54[28], stage1_54[29]},
      {stage2_56[4],stage2_55[18],stage2_54[41],stage2_53[51],stage2_52[69]}
   );
   gpc606_5 gpc5631 (
      {stage1_52[66], stage1_52[67], stage1_52[68], stage1_52[69], stage1_52[70], stage1_52[71]},
      {stage1_54[30], stage1_54[31], stage1_54[32], stage1_54[33], stage1_54[34], stage1_54[35]},
      {stage2_56[5],stage2_55[19],stage2_54[42],stage2_53[52],stage2_52[70]}
   );
   gpc606_5 gpc5632 (
      {stage1_52[72], stage1_52[73], stage1_52[74], stage1_52[75], stage1_52[76], stage1_52[77]},
      {stage1_54[36], stage1_54[37], stage1_54[38], stage1_54[39], stage1_54[40], stage1_54[41]},
      {stage2_56[6],stage2_55[20],stage2_54[43],stage2_53[53],stage2_52[71]}
   );
   gpc606_5 gpc5633 (
      {stage1_52[78], stage1_52[79], stage1_52[80], stage1_52[81], stage1_52[82], stage1_52[83]},
      {stage1_54[42], stage1_54[43], stage1_54[44], stage1_54[45], stage1_54[46], stage1_54[47]},
      {stage2_56[7],stage2_55[21],stage2_54[44],stage2_53[54],stage2_52[72]}
   );
   gpc606_5 gpc5634 (
      {stage1_52[84], stage1_52[85], stage1_52[86], stage1_52[87], stage1_52[88], stage1_52[89]},
      {stage1_54[48], stage1_54[49], stage1_54[50], stage1_54[51], stage1_54[52], stage1_54[53]},
      {stage2_56[8],stage2_55[22],stage2_54[45],stage2_53[55],stage2_52[73]}
   );
   gpc606_5 gpc5635 (
      {stage1_52[90], stage1_52[91], stage1_52[92], stage1_52[93], stage1_52[94], stage1_52[95]},
      {stage1_54[54], stage1_54[55], stage1_54[56], stage1_54[57], stage1_54[58], stage1_54[59]},
      {stage2_56[9],stage2_55[23],stage2_54[46],stage2_53[56],stage2_52[74]}
   );
   gpc606_5 gpc5636 (
      {stage1_52[96], stage1_52[97], stage1_52[98], stage1_52[99], stage1_52[100], stage1_52[101]},
      {stage1_54[60], stage1_54[61], stage1_54[62], stage1_54[63], stage1_54[64], stage1_54[65]},
      {stage2_56[10],stage2_55[24],stage2_54[47],stage2_53[57],stage2_52[75]}
   );
   gpc615_5 gpc5637 (
      {stage1_52[102], stage1_52[103], stage1_52[104], stage1_52[105], stage1_52[106]},
      {stage1_53[108]},
      {stage1_54[66], stage1_54[67], stage1_54[68], stage1_54[69], stage1_54[70], stage1_54[71]},
      {stage2_56[11],stage2_55[25],stage2_54[48],stage2_53[58],stage2_52[76]}
   );
   gpc615_5 gpc5638 (
      {stage1_52[107], stage1_52[108], stage1_52[109], stage1_52[110], stage1_52[111]},
      {stage1_53[109]},
      {stage1_54[72], stage1_54[73], stage1_54[74], stage1_54[75], stage1_54[76], stage1_54[77]},
      {stage2_56[12],stage2_55[26],stage2_54[49],stage2_53[59],stage2_52[77]}
   );
   gpc615_5 gpc5639 (
      {stage1_52[112], stage1_52[113], stage1_52[114], stage1_52[115], stage1_52[116]},
      {stage1_53[110]},
      {stage1_54[78], stage1_54[79], stage1_54[80], stage1_54[81], stage1_54[82], stage1_54[83]},
      {stage2_56[13],stage2_55[27],stage2_54[50],stage2_53[60],stage2_52[78]}
   );
   gpc615_5 gpc5640 (
      {stage1_52[117], stage1_52[118], stage1_52[119], stage1_52[120], stage1_52[121]},
      {stage1_53[111]},
      {stage1_54[84], stage1_54[85], stage1_54[86], stage1_54[87], stage1_54[88], stage1_54[89]},
      {stage2_56[14],stage2_55[28],stage2_54[51],stage2_53[61],stage2_52[79]}
   );
   gpc615_5 gpc5641 (
      {stage1_52[122], stage1_52[123], stage1_52[124], stage1_52[125], stage1_52[126]},
      {stage1_53[112]},
      {stage1_54[90], stage1_54[91], stage1_54[92], stage1_54[93], stage1_54[94], stage1_54[95]},
      {stage2_56[15],stage2_55[29],stage2_54[52],stage2_53[62],stage2_52[80]}
   );
   gpc615_5 gpc5642 (
      {stage1_52[127], stage1_52[128], stage1_52[129], stage1_52[130], stage1_52[131]},
      {stage1_53[113]},
      {stage1_54[96], stage1_54[97], stage1_54[98], stage1_54[99], stage1_54[100], stage1_54[101]},
      {stage2_56[16],stage2_55[30],stage2_54[53],stage2_53[63],stage2_52[81]}
   );
   gpc615_5 gpc5643 (
      {stage1_52[132], stage1_52[133], stage1_52[134], stage1_52[135], stage1_52[136]},
      {stage1_53[114]},
      {stage1_54[102], stage1_54[103], stage1_54[104], stage1_54[105], stage1_54[106], stage1_54[107]},
      {stage2_56[17],stage2_55[31],stage2_54[54],stage2_53[64],stage2_52[82]}
   );
   gpc615_5 gpc5644 (
      {stage1_52[137], stage1_52[138], stage1_52[139], stage1_52[140], stage1_52[141]},
      {stage1_53[115]},
      {stage1_54[108], stage1_54[109], stage1_54[110], stage1_54[111], stage1_54[112], stage1_54[113]},
      {stage2_56[18],stage2_55[32],stage2_54[55],stage2_53[65],stage2_52[83]}
   );
   gpc615_5 gpc5645 (
      {stage1_52[142], stage1_52[143], stage1_52[144], stage1_52[145], stage1_52[146]},
      {stage1_53[116]},
      {stage1_54[114], stage1_54[115], stage1_54[116], stage1_54[117], stage1_54[118], stage1_54[119]},
      {stage2_56[19],stage2_55[33],stage2_54[56],stage2_53[66],stage2_52[84]}
   );
   gpc615_5 gpc5646 (
      {stage1_52[147], stage1_52[148], stage1_52[149], stage1_52[150], stage1_52[151]},
      {stage1_53[117]},
      {stage1_54[120], stage1_54[121], stage1_54[122], stage1_54[123], stage1_54[124], stage1_54[125]},
      {stage2_56[20],stage2_55[34],stage2_54[57],stage2_53[67],stage2_52[85]}
   );
   gpc615_5 gpc5647 (
      {stage1_52[152], stage1_52[153], stage1_52[154], stage1_52[155], stage1_52[156]},
      {stage1_53[118]},
      {stage1_54[126], stage1_54[127], stage1_54[128], stage1_54[129], stage1_54[130], stage1_54[131]},
      {stage2_56[21],stage2_55[35],stage2_54[58],stage2_53[68],stage2_52[86]}
   );
   gpc615_5 gpc5648 (
      {stage1_52[157], stage1_52[158], stage1_52[159], stage1_52[160], stage1_52[161]},
      {stage1_53[119]},
      {stage1_54[132], stage1_54[133], stage1_54[134], stage1_54[135], stage1_54[136], stage1_54[137]},
      {stage2_56[22],stage2_55[36],stage2_54[59],stage2_53[69],stage2_52[87]}
   );
   gpc615_5 gpc5649 (
      {stage1_52[162], stage1_52[163], stage1_52[164], stage1_52[165], stage1_52[166]},
      {stage1_53[120]},
      {stage1_54[138], stage1_54[139], stage1_54[140], stage1_54[141], stage1_54[142], stage1_54[143]},
      {stage2_56[23],stage2_55[37],stage2_54[60],stage2_53[70],stage2_52[88]}
   );
   gpc615_5 gpc5650 (
      {stage1_52[167], stage1_52[168], stage1_52[169], stage1_52[170], stage1_52[171]},
      {stage1_53[121]},
      {stage1_54[144], stage1_54[145], stage1_54[146], stage1_54[147], stage1_54[148], stage1_54[149]},
      {stage2_56[24],stage2_55[38],stage2_54[61],stage2_53[71],stage2_52[89]}
   );
   gpc615_5 gpc5651 (
      {stage1_52[172], stage1_52[173], stage1_52[174], stage1_52[175], stage1_52[176]},
      {stage1_53[122]},
      {stage1_54[150], stage1_54[151], stage1_54[152], stage1_54[153], stage1_54[154], stage1_54[155]},
      {stage2_56[25],stage2_55[39],stage2_54[62],stage2_53[72],stage2_52[90]}
   );
   gpc615_5 gpc5652 (
      {stage1_52[177], stage1_52[178], stage1_52[179], stage1_52[180], stage1_52[181]},
      {stage1_53[123]},
      {stage1_54[156], stage1_54[157], stage1_54[158], stage1_54[159], stage1_54[160], stage1_54[161]},
      {stage2_56[26],stage2_55[40],stage2_54[63],stage2_53[73],stage2_52[91]}
   );
   gpc615_5 gpc5653 (
      {stage1_52[182], stage1_52[183], stage1_52[184], stage1_52[185], stage1_52[186]},
      {stage1_53[124]},
      {stage1_54[162], stage1_54[163], stage1_54[164], stage1_54[165], stage1_54[166], stage1_54[167]},
      {stage2_56[27],stage2_55[41],stage2_54[64],stage2_53[74],stage2_52[92]}
   );
   gpc615_5 gpc5654 (
      {stage1_53[125], stage1_53[126], stage1_53[127], stage1_53[128], stage1_53[129]},
      {stage1_54[168]},
      {stage1_55[0], stage1_55[1], stage1_55[2], stage1_55[3], stage1_55[4], stage1_55[5]},
      {stage2_57[0],stage2_56[28],stage2_55[42],stage2_54[65],stage2_53[75]}
   );
   gpc606_5 gpc5655 (
      {stage1_54[169], stage1_54[170], stage1_54[171], stage1_54[172], stage1_54[173], stage1_54[174]},
      {stage1_56[0], stage1_56[1], stage1_56[2], stage1_56[3], stage1_56[4], stage1_56[5]},
      {stage2_58[0],stage2_57[1],stage2_56[29],stage2_55[43],stage2_54[66]}
   );
   gpc606_5 gpc5656 (
      {stage1_54[175], stage1_54[176], stage1_54[177], stage1_54[178], stage1_54[179], stage1_54[180]},
      {stage1_56[6], stage1_56[7], stage1_56[8], stage1_56[9], stage1_56[10], stage1_56[11]},
      {stage2_58[1],stage2_57[2],stage2_56[30],stage2_55[44],stage2_54[67]}
   );
   gpc606_5 gpc5657 (
      {stage1_54[181], stage1_54[182], stage1_54[183], stage1_54[184], stage1_54[185], stage1_54[186]},
      {stage1_56[12], stage1_56[13], stage1_56[14], stage1_56[15], stage1_56[16], stage1_56[17]},
      {stage2_58[2],stage2_57[3],stage2_56[31],stage2_55[45],stage2_54[68]}
   );
   gpc606_5 gpc5658 (
      {stage1_54[187], stage1_54[188], stage1_54[189], stage1_54[190], stage1_54[191], stage1_54[192]},
      {stage1_56[18], stage1_56[19], stage1_56[20], stage1_56[21], stage1_56[22], stage1_56[23]},
      {stage2_58[3],stage2_57[4],stage2_56[32],stage2_55[46],stage2_54[69]}
   );
   gpc615_5 gpc5659 (
      {stage1_54[193], stage1_54[194], stage1_54[195], stage1_54[196], stage1_54[197]},
      {stage1_55[6]},
      {stage1_56[24], stage1_56[25], stage1_56[26], stage1_56[27], stage1_56[28], stage1_56[29]},
      {stage2_58[4],stage2_57[5],stage2_56[33],stage2_55[47],stage2_54[70]}
   );
   gpc615_5 gpc5660 (
      {stage1_54[198], stage1_54[199], stage1_54[200], stage1_54[201], stage1_54[202]},
      {stage1_55[7]},
      {stage1_56[30], stage1_56[31], stage1_56[32], stage1_56[33], stage1_56[34], stage1_56[35]},
      {stage2_58[5],stage2_57[6],stage2_56[34],stage2_55[48],stage2_54[71]}
   );
   gpc2135_5 gpc5661 (
      {stage1_55[8], stage1_55[9], stage1_55[10], stage1_55[11], stage1_55[12]},
      {stage1_56[36], stage1_56[37], stage1_56[38]},
      {stage1_57[0]},
      {stage1_58[0], stage1_58[1]},
      {stage2_59[0],stage2_58[6],stage2_57[7],stage2_56[35],stage2_55[49]}
   );
   gpc2135_5 gpc5662 (
      {stage1_55[13], stage1_55[14], stage1_55[15], stage1_55[16], stage1_55[17]},
      {stage1_56[39], stage1_56[40], stage1_56[41]},
      {stage1_57[1]},
      {stage1_58[2], stage1_58[3]},
      {stage2_59[1],stage2_58[7],stage2_57[8],stage2_56[36],stage2_55[50]}
   );
   gpc2135_5 gpc5663 (
      {stage1_55[18], stage1_55[19], stage1_55[20], stage1_55[21], stage1_55[22]},
      {stage1_56[42], stage1_56[43], stage1_56[44]},
      {stage1_57[2]},
      {stage1_58[4], stage1_58[5]},
      {stage2_59[2],stage2_58[8],stage2_57[9],stage2_56[37],stage2_55[51]}
   );
   gpc2135_5 gpc5664 (
      {stage1_55[23], stage1_55[24], stage1_55[25], stage1_55[26], stage1_55[27]},
      {stage1_56[45], stage1_56[46], stage1_56[47]},
      {stage1_57[3]},
      {stage1_58[6], stage1_58[7]},
      {stage2_59[3],stage2_58[9],stage2_57[10],stage2_56[38],stage2_55[52]}
   );
   gpc2135_5 gpc5665 (
      {stage1_55[28], stage1_55[29], stage1_55[30], stage1_55[31], stage1_55[32]},
      {stage1_56[48], stage1_56[49], stage1_56[50]},
      {stage1_57[4]},
      {stage1_58[8], stage1_58[9]},
      {stage2_59[4],stage2_58[10],stage2_57[11],stage2_56[39],stage2_55[53]}
   );
   gpc2135_5 gpc5666 (
      {stage1_55[33], stage1_55[34], stage1_55[35], stage1_55[36], stage1_55[37]},
      {stage1_56[51], stage1_56[52], stage1_56[53]},
      {stage1_57[5]},
      {stage1_58[10], stage1_58[11]},
      {stage2_59[5],stage2_58[11],stage2_57[12],stage2_56[40],stage2_55[54]}
   );
   gpc2135_5 gpc5667 (
      {stage1_55[38], stage1_55[39], stage1_55[40], stage1_55[41], stage1_55[42]},
      {stage1_56[54], stage1_56[55], stage1_56[56]},
      {stage1_57[6]},
      {stage1_58[12], stage1_58[13]},
      {stage2_59[6],stage2_58[12],stage2_57[13],stage2_56[41],stage2_55[55]}
   );
   gpc2135_5 gpc5668 (
      {stage1_55[43], stage1_55[44], stage1_55[45], stage1_55[46], stage1_55[47]},
      {stage1_56[57], stage1_56[58], stage1_56[59]},
      {stage1_57[7]},
      {stage1_58[14], stage1_58[15]},
      {stage2_59[7],stage2_58[13],stage2_57[14],stage2_56[42],stage2_55[56]}
   );
   gpc2135_5 gpc5669 (
      {stage1_55[48], stage1_55[49], stage1_55[50], stage1_55[51], stage1_55[52]},
      {stage1_56[60], stage1_56[61], stage1_56[62]},
      {stage1_57[8]},
      {stage1_58[16], stage1_58[17]},
      {stage2_59[8],stage2_58[14],stage2_57[15],stage2_56[43],stage2_55[57]}
   );
   gpc2135_5 gpc5670 (
      {stage1_55[53], stage1_55[54], stage1_55[55], stage1_55[56], stage1_55[57]},
      {stage1_56[63], stage1_56[64], stage1_56[65]},
      {stage1_57[9]},
      {stage1_58[18], stage1_58[19]},
      {stage2_59[9],stage2_58[15],stage2_57[16],stage2_56[44],stage2_55[58]}
   );
   gpc2135_5 gpc5671 (
      {stage1_55[58], stage1_55[59], stage1_55[60], stage1_55[61], stage1_55[62]},
      {stage1_56[66], stage1_56[67], stage1_56[68]},
      {stage1_57[10]},
      {stage1_58[20], stage1_58[21]},
      {stage2_59[10],stage2_58[16],stage2_57[17],stage2_56[45],stage2_55[59]}
   );
   gpc2135_5 gpc5672 (
      {stage1_55[63], stage1_55[64], stage1_55[65], stage1_55[66], stage1_55[67]},
      {stage1_56[69], stage1_56[70], stage1_56[71]},
      {stage1_57[11]},
      {stage1_58[22], stage1_58[23]},
      {stage2_59[11],stage2_58[17],stage2_57[18],stage2_56[46],stage2_55[60]}
   );
   gpc2135_5 gpc5673 (
      {stage1_55[68], stage1_55[69], stage1_55[70], stage1_55[71], stage1_55[72]},
      {stage1_56[72], stage1_56[73], stage1_56[74]},
      {stage1_57[12]},
      {stage1_58[24], stage1_58[25]},
      {stage2_59[12],stage2_58[18],stage2_57[19],stage2_56[47],stage2_55[61]}
   );
   gpc2135_5 gpc5674 (
      {stage1_55[73], stage1_55[74], stage1_55[75], stage1_55[76], stage1_55[77]},
      {stage1_56[75], stage1_56[76], stage1_56[77]},
      {stage1_57[13]},
      {stage1_58[26], stage1_58[27]},
      {stage2_59[13],stage2_58[19],stage2_57[20],stage2_56[48],stage2_55[62]}
   );
   gpc2135_5 gpc5675 (
      {stage1_55[78], stage1_55[79], stage1_55[80], stage1_55[81], stage1_55[82]},
      {stage1_56[78], stage1_56[79], stage1_56[80]},
      {stage1_57[14]},
      {stage1_58[28], stage1_58[29]},
      {stage2_59[14],stage2_58[20],stage2_57[21],stage2_56[49],stage2_55[63]}
   );
   gpc2135_5 gpc5676 (
      {stage1_55[83], stage1_55[84], stage1_55[85], stage1_55[86], stage1_55[87]},
      {stage1_56[81], stage1_56[82], stage1_56[83]},
      {stage1_57[15]},
      {stage1_58[30], stage1_58[31]},
      {stage2_59[15],stage2_58[21],stage2_57[22],stage2_56[50],stage2_55[64]}
   );
   gpc2135_5 gpc5677 (
      {stage1_55[88], stage1_55[89], stage1_55[90], stage1_55[91], stage1_55[92]},
      {stage1_56[84], stage1_56[85], stage1_56[86]},
      {stage1_57[16]},
      {stage1_58[32], stage1_58[33]},
      {stage2_59[16],stage2_58[22],stage2_57[23],stage2_56[51],stage2_55[65]}
   );
   gpc2135_5 gpc5678 (
      {stage1_55[93], stage1_55[94], stage1_55[95], stage1_55[96], stage1_55[97]},
      {stage1_56[87], stage1_56[88], stage1_56[89]},
      {stage1_57[17]},
      {stage1_58[34], stage1_58[35]},
      {stage2_59[17],stage2_58[23],stage2_57[24],stage2_56[52],stage2_55[66]}
   );
   gpc606_5 gpc5679 (
      {stage1_55[98], stage1_55[99], stage1_55[100], stage1_55[101], stage1_55[102], stage1_55[103]},
      {stage1_57[18], stage1_57[19], stage1_57[20], stage1_57[21], stage1_57[22], stage1_57[23]},
      {stage2_59[18],stage2_58[24],stage2_57[25],stage2_56[53],stage2_55[67]}
   );
   gpc606_5 gpc5680 (
      {stage1_55[104], stage1_55[105], stage1_55[106], stage1_55[107], stage1_55[108], stage1_55[109]},
      {stage1_57[24], stage1_57[25], stage1_57[26], stage1_57[27], stage1_57[28], stage1_57[29]},
      {stage2_59[19],stage2_58[25],stage2_57[26],stage2_56[54],stage2_55[68]}
   );
   gpc606_5 gpc5681 (
      {stage1_55[110], stage1_55[111], stage1_55[112], stage1_55[113], stage1_55[114], stage1_55[115]},
      {stage1_57[30], stage1_57[31], stage1_57[32], stage1_57[33], stage1_57[34], stage1_57[35]},
      {stage2_59[20],stage2_58[26],stage2_57[27],stage2_56[55],stage2_55[69]}
   );
   gpc606_5 gpc5682 (
      {stage1_55[116], stage1_55[117], stage1_55[118], stage1_55[119], stage1_55[120], stage1_55[121]},
      {stage1_57[36], stage1_57[37], stage1_57[38], stage1_57[39], stage1_57[40], stage1_57[41]},
      {stage2_59[21],stage2_58[27],stage2_57[28],stage2_56[56],stage2_55[70]}
   );
   gpc606_5 gpc5683 (
      {stage1_55[122], stage1_55[123], stage1_55[124], stage1_55[125], stage1_55[126], stage1_55[127]},
      {stage1_57[42], stage1_57[43], stage1_57[44], stage1_57[45], stage1_57[46], stage1_57[47]},
      {stage2_59[22],stage2_58[28],stage2_57[29],stage2_56[57],stage2_55[71]}
   );
   gpc606_5 gpc5684 (
      {stage1_55[128], stage1_55[129], stage1_55[130], stage1_55[131], stage1_55[132], stage1_55[133]},
      {stage1_57[48], stage1_57[49], stage1_57[50], stage1_57[51], stage1_57[52], stage1_57[53]},
      {stage2_59[23],stage2_58[29],stage2_57[30],stage2_56[58],stage2_55[72]}
   );
   gpc606_5 gpc5685 (
      {stage1_55[134], stage1_55[135], stage1_55[136], stage1_55[137], stage1_55[138], stage1_55[139]},
      {stage1_57[54], stage1_57[55], stage1_57[56], stage1_57[57], stage1_57[58], stage1_57[59]},
      {stage2_59[24],stage2_58[30],stage2_57[31],stage2_56[59],stage2_55[73]}
   );
   gpc606_5 gpc5686 (
      {stage1_55[140], stage1_55[141], stage1_55[142], stage1_55[143], stage1_55[144], stage1_55[145]},
      {stage1_57[60], stage1_57[61], stage1_57[62], stage1_57[63], stage1_57[64], stage1_57[65]},
      {stage2_59[25],stage2_58[31],stage2_57[32],stage2_56[60],stage2_55[74]}
   );
   gpc606_5 gpc5687 (
      {stage1_55[146], stage1_55[147], stage1_55[148], stage1_55[149], stage1_55[150], stage1_55[151]},
      {stage1_57[66], stage1_57[67], stage1_57[68], stage1_57[69], stage1_57[70], stage1_57[71]},
      {stage2_59[26],stage2_58[32],stage2_57[33],stage2_56[61],stage2_55[75]}
   );
   gpc606_5 gpc5688 (
      {stage1_55[152], stage1_55[153], stage1_55[154], stage1_55[155], stage1_55[156], stage1_55[157]},
      {stage1_57[72], stage1_57[73], stage1_57[74], stage1_57[75], stage1_57[76], stage1_57[77]},
      {stage2_59[27],stage2_58[33],stage2_57[34],stage2_56[62],stage2_55[76]}
   );
   gpc606_5 gpc5689 (
      {stage1_55[158], stage1_55[159], stage1_55[160], stage1_55[161], stage1_55[162], stage1_55[163]},
      {stage1_57[78], stage1_57[79], stage1_57[80], stage1_57[81], stage1_57[82], stage1_57[83]},
      {stage2_59[28],stage2_58[34],stage2_57[35],stage2_56[63],stage2_55[77]}
   );
   gpc606_5 gpc5690 (
      {stage1_55[164], stage1_55[165], stage1_55[166], stage1_55[167], stage1_55[168], stage1_55[169]},
      {stage1_57[84], stage1_57[85], stage1_57[86], stage1_57[87], stage1_57[88], stage1_57[89]},
      {stage2_59[29],stage2_58[35],stage2_57[36],stage2_56[64],stage2_55[78]}
   );
   gpc606_5 gpc5691 (
      {stage1_55[170], stage1_55[171], stage1_55[172], stage1_55[173], stage1_55[174], stage1_55[175]},
      {stage1_57[90], stage1_57[91], stage1_57[92], stage1_57[93], stage1_57[94], stage1_57[95]},
      {stage2_59[30],stage2_58[36],stage2_57[37],stage2_56[65],stage2_55[79]}
   );
   gpc606_5 gpc5692 (
      {stage1_55[176], stage1_55[177], stage1_55[178], stage1_55[179], stage1_55[180], stage1_55[181]},
      {stage1_57[96], stage1_57[97], stage1_57[98], stage1_57[99], stage1_57[100], stage1_57[101]},
      {stage2_59[31],stage2_58[37],stage2_57[38],stage2_56[66],stage2_55[80]}
   );
   gpc606_5 gpc5693 (
      {stage1_55[182], stage1_55[183], stage1_55[184], stage1_55[185], stage1_55[186], stage1_55[187]},
      {stage1_57[102], stage1_57[103], stage1_57[104], stage1_57[105], stage1_57[106], stage1_57[107]},
      {stage2_59[32],stage2_58[38],stage2_57[39],stage2_56[67],stage2_55[81]}
   );
   gpc606_5 gpc5694 (
      {stage1_55[188], stage1_55[189], stage1_55[190], stage1_55[191], stage1_55[192], stage1_55[193]},
      {stage1_57[108], stage1_57[109], stage1_57[110], stage1_57[111], stage1_57[112], stage1_57[113]},
      {stage2_59[33],stage2_58[39],stage2_57[40],stage2_56[68],stage2_55[82]}
   );
   gpc606_5 gpc5695 (
      {stage1_55[194], stage1_55[195], stage1_55[196], stage1_55[197], stage1_55[198], stage1_55[199]},
      {stage1_57[114], stage1_57[115], stage1_57[116], stage1_57[117], stage1_57[118], stage1_57[119]},
      {stage2_59[34],stage2_58[40],stage2_57[41],stage2_56[69],stage2_55[83]}
   );
   gpc606_5 gpc5696 (
      {stage1_55[200], stage1_55[201], stage1_55[202], stage1_55[203], stage1_55[204], stage1_55[205]},
      {stage1_57[120], stage1_57[121], stage1_57[122], stage1_57[123], stage1_57[124], stage1_57[125]},
      {stage2_59[35],stage2_58[41],stage2_57[42],stage2_56[70],stage2_55[84]}
   );
   gpc606_5 gpc5697 (
      {stage1_55[206], stage1_55[207], stage1_55[208], stage1_55[209], stage1_55[210], stage1_55[211]},
      {stage1_57[126], stage1_57[127], stage1_57[128], stage1_57[129], stage1_57[130], stage1_57[131]},
      {stage2_59[36],stage2_58[42],stage2_57[43],stage2_56[71],stage2_55[85]}
   );
   gpc606_5 gpc5698 (
      {stage1_55[212], stage1_55[213], stage1_55[214], stage1_55[215], stage1_55[216], stage1_55[217]},
      {stage1_57[132], stage1_57[133], stage1_57[134], stage1_57[135], stage1_57[136], stage1_57[137]},
      {stage2_59[37],stage2_58[43],stage2_57[44],stage2_56[72],stage2_55[86]}
   );
   gpc606_5 gpc5699 (
      {stage1_55[218], stage1_55[219], stage1_55[220], stage1_55[221], stage1_55[222], stage1_55[223]},
      {stage1_57[138], stage1_57[139], stage1_57[140], stage1_57[141], stage1_57[142], stage1_57[143]},
      {stage2_59[38],stage2_58[44],stage2_57[45],stage2_56[73],stage2_55[87]}
   );
   gpc606_5 gpc5700 (
      {stage1_55[224], stage1_55[225], stage1_55[226], stage1_55[227], stage1_55[228], stage1_55[229]},
      {stage1_57[144], stage1_57[145], stage1_57[146], stage1_57[147], stage1_57[148], stage1_57[149]},
      {stage2_59[39],stage2_58[45],stage2_57[46],stage2_56[74],stage2_55[88]}
   );
   gpc606_5 gpc5701 (
      {stage1_55[230], stage1_55[231], stage1_55[232], stage1_55[233], stage1_55[234], stage1_55[235]},
      {stage1_57[150], stage1_57[151], stage1_57[152], stage1_57[153], stage1_57[154], stage1_57[155]},
      {stage2_59[40],stage2_58[46],stage2_57[47],stage2_56[75],stage2_55[89]}
   );
   gpc606_5 gpc5702 (
      {stage1_55[236], stage1_55[237], stage1_55[238], stage1_55[239], stage1_55[240], stage1_55[241]},
      {stage1_57[156], stage1_57[157], stage1_57[158], stage1_57[159], stage1_57[160], stage1_57[161]},
      {stage2_59[41],stage2_58[47],stage2_57[48],stage2_56[76],stage2_55[90]}
   );
   gpc606_5 gpc5703 (
      {stage1_55[242], stage1_55[243], stage1_55[244], stage1_55[245], stage1_55[246], stage1_55[247]},
      {stage1_57[162], stage1_57[163], stage1_57[164], stage1_57[165], stage1_57[166], stage1_57[167]},
      {stage2_59[42],stage2_58[48],stage2_57[49],stage2_56[77],stage2_55[91]}
   );
   gpc606_5 gpc5704 (
      {stage1_55[248], stage1_55[249], stage1_55[250], stage1_55[251], stage1_55[252], stage1_55[253]},
      {stage1_57[168], stage1_57[169], stage1_57[170], stage1_57[171], stage1_57[172], stage1_57[173]},
      {stage2_59[43],stage2_58[49],stage2_57[50],stage2_56[78],stage2_55[92]}
   );
   gpc606_5 gpc5705 (
      {stage1_56[90], stage1_56[91], stage1_56[92], stage1_56[93], stage1_56[94], stage1_56[95]},
      {stage1_58[36], stage1_58[37], stage1_58[38], stage1_58[39], stage1_58[40], stage1_58[41]},
      {stage2_60[0],stage2_59[44],stage2_58[50],stage2_57[51],stage2_56[79]}
   );
   gpc606_5 gpc5706 (
      {stage1_56[96], stage1_56[97], stage1_56[98], stage1_56[99], stage1_56[100], stage1_56[101]},
      {stage1_58[42], stage1_58[43], stage1_58[44], stage1_58[45], stage1_58[46], stage1_58[47]},
      {stage2_60[1],stage2_59[45],stage2_58[51],stage2_57[52],stage2_56[80]}
   );
   gpc606_5 gpc5707 (
      {stage1_56[102], stage1_56[103], stage1_56[104], stage1_56[105], stage1_56[106], stage1_56[107]},
      {stage1_58[48], stage1_58[49], stage1_58[50], stage1_58[51], stage1_58[52], stage1_58[53]},
      {stage2_60[2],stage2_59[46],stage2_58[52],stage2_57[53],stage2_56[81]}
   );
   gpc606_5 gpc5708 (
      {stage1_56[108], stage1_56[109], stage1_56[110], stage1_56[111], stage1_56[112], stage1_56[113]},
      {stage1_58[54], stage1_58[55], stage1_58[56], stage1_58[57], stage1_58[58], stage1_58[59]},
      {stage2_60[3],stage2_59[47],stage2_58[53],stage2_57[54],stage2_56[82]}
   );
   gpc606_5 gpc5709 (
      {stage1_56[114], stage1_56[115], stage1_56[116], stage1_56[117], stage1_56[118], stage1_56[119]},
      {stage1_58[60], stage1_58[61], stage1_58[62], stage1_58[63], stage1_58[64], stage1_58[65]},
      {stage2_60[4],stage2_59[48],stage2_58[54],stage2_57[55],stage2_56[83]}
   );
   gpc606_5 gpc5710 (
      {stage1_56[120], stage1_56[121], stage1_56[122], stage1_56[123], stage1_56[124], stage1_56[125]},
      {stage1_58[66], stage1_58[67], stage1_58[68], stage1_58[69], stage1_58[70], stage1_58[71]},
      {stage2_60[5],stage2_59[49],stage2_58[55],stage2_57[56],stage2_56[84]}
   );
   gpc606_5 gpc5711 (
      {stage1_56[126], stage1_56[127], stage1_56[128], stage1_56[129], stage1_56[130], stage1_56[131]},
      {stage1_58[72], stage1_58[73], stage1_58[74], stage1_58[75], stage1_58[76], stage1_58[77]},
      {stage2_60[6],stage2_59[50],stage2_58[56],stage2_57[57],stage2_56[85]}
   );
   gpc606_5 gpc5712 (
      {stage1_56[132], stage1_56[133], stage1_56[134], stage1_56[135], stage1_56[136], stage1_56[137]},
      {stage1_58[78], stage1_58[79], stage1_58[80], stage1_58[81], stage1_58[82], stage1_58[83]},
      {stage2_60[7],stage2_59[51],stage2_58[57],stage2_57[58],stage2_56[86]}
   );
   gpc606_5 gpc5713 (
      {stage1_56[138], stage1_56[139], stage1_56[140], stage1_56[141], stage1_56[142], stage1_56[143]},
      {stage1_58[84], stage1_58[85], stage1_58[86], stage1_58[87], stage1_58[88], stage1_58[89]},
      {stage2_60[8],stage2_59[52],stage2_58[58],stage2_57[59],stage2_56[87]}
   );
   gpc615_5 gpc5714 (
      {stage1_56[144], stage1_56[145], stage1_56[146], stage1_56[147], stage1_56[148]},
      {stage1_57[174]},
      {stage1_58[90], stage1_58[91], stage1_58[92], stage1_58[93], stage1_58[94], stage1_58[95]},
      {stage2_60[9],stage2_59[53],stage2_58[59],stage2_57[60],stage2_56[88]}
   );
   gpc615_5 gpc5715 (
      {stage1_56[149], stage1_56[150], stage1_56[151], stage1_56[152], stage1_56[153]},
      {stage1_57[175]},
      {stage1_58[96], stage1_58[97], stage1_58[98], stage1_58[99], stage1_58[100], stage1_58[101]},
      {stage2_60[10],stage2_59[54],stage2_58[60],stage2_57[61],stage2_56[89]}
   );
   gpc615_5 gpc5716 (
      {stage1_56[154], stage1_56[155], stage1_56[156], stage1_56[157], stage1_56[158]},
      {stage1_57[176]},
      {stage1_58[102], stage1_58[103], stage1_58[104], stage1_58[105], stage1_58[106], stage1_58[107]},
      {stage2_60[11],stage2_59[55],stage2_58[61],stage2_57[62],stage2_56[90]}
   );
   gpc615_5 gpc5717 (
      {stage1_56[159], stage1_56[160], stage1_56[161], stage1_56[162], stage1_56[163]},
      {stage1_57[177]},
      {stage1_58[108], stage1_58[109], stage1_58[110], stage1_58[111], stage1_58[112], stage1_58[113]},
      {stage2_60[12],stage2_59[56],stage2_58[62],stage2_57[63],stage2_56[91]}
   );
   gpc606_5 gpc5718 (
      {stage1_57[178], stage1_57[179], stage1_57[180], stage1_57[181], stage1_57[182], stage1_57[183]},
      {stage1_59[0], stage1_59[1], stage1_59[2], stage1_59[3], stage1_59[4], stage1_59[5]},
      {stage2_61[0],stage2_60[13],stage2_59[57],stage2_58[63],stage2_57[64]}
   );
   gpc615_5 gpc5719 (
      {stage1_57[184], stage1_57[185], stage1_57[186], stage1_57[187], stage1_57[188]},
      {stage1_58[114]},
      {stage1_59[6], stage1_59[7], stage1_59[8], stage1_59[9], stage1_59[10], stage1_59[11]},
      {stage2_61[1],stage2_60[14],stage2_59[58],stage2_58[64],stage2_57[65]}
   );
   gpc615_5 gpc5720 (
      {stage1_58[115], stage1_58[116], stage1_58[117], stage1_58[118], stage1_58[119]},
      {stage1_59[12]},
      {stage1_60[0], stage1_60[1], stage1_60[2], stage1_60[3], stage1_60[4], stage1_60[5]},
      {stage2_62[0],stage2_61[2],stage2_60[15],stage2_59[59],stage2_58[65]}
   );
   gpc615_5 gpc5721 (
      {stage1_58[120], stage1_58[121], stage1_58[122], stage1_58[123], stage1_58[124]},
      {stage1_59[13]},
      {stage1_60[6], stage1_60[7], stage1_60[8], stage1_60[9], stage1_60[10], stage1_60[11]},
      {stage2_62[1],stage2_61[3],stage2_60[16],stage2_59[60],stage2_58[66]}
   );
   gpc615_5 gpc5722 (
      {stage1_58[125], stage1_58[126], stage1_58[127], stage1_58[128], stage1_58[129]},
      {stage1_59[14]},
      {stage1_60[12], stage1_60[13], stage1_60[14], stage1_60[15], stage1_60[16], stage1_60[17]},
      {stage2_62[2],stage2_61[4],stage2_60[17],stage2_59[61],stage2_58[67]}
   );
   gpc615_5 gpc5723 (
      {stage1_58[130], stage1_58[131], stage1_58[132], stage1_58[133], stage1_58[134]},
      {stage1_59[15]},
      {stage1_60[18], stage1_60[19], stage1_60[20], stage1_60[21], stage1_60[22], stage1_60[23]},
      {stage2_62[3],stage2_61[5],stage2_60[18],stage2_59[62],stage2_58[68]}
   );
   gpc615_5 gpc5724 (
      {stage1_58[135], stage1_58[136], stage1_58[137], stage1_58[138], stage1_58[139]},
      {stage1_59[16]},
      {stage1_60[24], stage1_60[25], stage1_60[26], stage1_60[27], stage1_60[28], stage1_60[29]},
      {stage2_62[4],stage2_61[6],stage2_60[19],stage2_59[63],stage2_58[69]}
   );
   gpc615_5 gpc5725 (
      {stage1_58[140], stage1_58[141], stage1_58[142], stage1_58[143], stage1_58[144]},
      {stage1_59[17]},
      {stage1_60[30], stage1_60[31], stage1_60[32], stage1_60[33], stage1_60[34], stage1_60[35]},
      {stage2_62[5],stage2_61[7],stage2_60[20],stage2_59[64],stage2_58[70]}
   );
   gpc615_5 gpc5726 (
      {stage1_58[145], stage1_58[146], stage1_58[147], stage1_58[148], stage1_58[149]},
      {stage1_59[18]},
      {stage1_60[36], stage1_60[37], stage1_60[38], stage1_60[39], stage1_60[40], stage1_60[41]},
      {stage2_62[6],stage2_61[8],stage2_60[21],stage2_59[65],stage2_58[71]}
   );
   gpc615_5 gpc5727 (
      {stage1_58[150], stage1_58[151], stage1_58[152], stage1_58[153], stage1_58[154]},
      {stage1_59[19]},
      {stage1_60[42], stage1_60[43], stage1_60[44], stage1_60[45], stage1_60[46], stage1_60[47]},
      {stage2_62[7],stage2_61[9],stage2_60[22],stage2_59[66],stage2_58[72]}
   );
   gpc615_5 gpc5728 (
      {stage1_58[155], stage1_58[156], stage1_58[157], stage1_58[158], stage1_58[159]},
      {stage1_59[20]},
      {stage1_60[48], stage1_60[49], stage1_60[50], stage1_60[51], stage1_60[52], stage1_60[53]},
      {stage2_62[8],stage2_61[10],stage2_60[23],stage2_59[67],stage2_58[73]}
   );
   gpc615_5 gpc5729 (
      {stage1_58[160], stage1_58[161], stage1_58[162], stage1_58[163], stage1_58[164]},
      {stage1_59[21]},
      {stage1_60[54], stage1_60[55], stage1_60[56], stage1_60[57], stage1_60[58], stage1_60[59]},
      {stage2_62[9],stage2_61[11],stage2_60[24],stage2_59[68],stage2_58[74]}
   );
   gpc615_5 gpc5730 (
      {stage1_58[165], stage1_58[166], stage1_58[167], stage1_58[168], stage1_58[169]},
      {stage1_59[22]},
      {stage1_60[60], stage1_60[61], stage1_60[62], stage1_60[63], stage1_60[64], stage1_60[65]},
      {stage2_62[10],stage2_61[12],stage2_60[25],stage2_59[69],stage2_58[75]}
   );
   gpc615_5 gpc5731 (
      {stage1_58[170], stage1_58[171], stage1_58[172], stage1_58[173], stage1_58[174]},
      {stage1_59[23]},
      {stage1_60[66], stage1_60[67], stage1_60[68], stage1_60[69], stage1_60[70], stage1_60[71]},
      {stage2_62[11],stage2_61[13],stage2_60[26],stage2_59[70],stage2_58[76]}
   );
   gpc615_5 gpc5732 (
      {stage1_58[175], stage1_58[176], stage1_58[177], stage1_58[178], stage1_58[179]},
      {stage1_59[24]},
      {stage1_60[72], stage1_60[73], stage1_60[74], stage1_60[75], stage1_60[76], stage1_60[77]},
      {stage2_62[12],stage2_61[14],stage2_60[27],stage2_59[71],stage2_58[77]}
   );
   gpc615_5 gpc5733 (
      {stage1_58[180], stage1_58[181], stage1_58[182], stage1_58[183], stage1_58[184]},
      {stage1_59[25]},
      {stage1_60[78], stage1_60[79], stage1_60[80], stage1_60[81], stage1_60[82], stage1_60[83]},
      {stage2_62[13],stage2_61[15],stage2_60[28],stage2_59[72],stage2_58[78]}
   );
   gpc615_5 gpc5734 (
      {stage1_58[185], stage1_58[186], stage1_58[187], stage1_58[188], stage1_58[189]},
      {stage1_59[26]},
      {stage1_60[84], stage1_60[85], stage1_60[86], stage1_60[87], stage1_60[88], stage1_60[89]},
      {stage2_62[14],stage2_61[16],stage2_60[29],stage2_59[73],stage2_58[79]}
   );
   gpc615_5 gpc5735 (
      {stage1_58[190], stage1_58[191], stage1_58[192], stage1_58[193], stage1_58[194]},
      {stage1_59[27]},
      {stage1_60[90], stage1_60[91], stage1_60[92], stage1_60[93], stage1_60[94], stage1_60[95]},
      {stage2_62[15],stage2_61[17],stage2_60[30],stage2_59[74],stage2_58[80]}
   );
   gpc615_5 gpc5736 (
      {stage1_58[195], stage1_58[196], stage1_58[197], stage1_58[198], stage1_58[199]},
      {stage1_59[28]},
      {stage1_60[96], stage1_60[97], stage1_60[98], stage1_60[99], stage1_60[100], stage1_60[101]},
      {stage2_62[16],stage2_61[18],stage2_60[31],stage2_59[75],stage2_58[81]}
   );
   gpc615_5 gpc5737 (
      {stage1_58[200], stage1_58[201], stage1_58[202], stage1_58[203], stage1_58[204]},
      {stage1_59[29]},
      {stage1_60[102], stage1_60[103], stage1_60[104], stage1_60[105], stage1_60[106], stage1_60[107]},
      {stage2_62[17],stage2_61[19],stage2_60[32],stage2_59[76],stage2_58[82]}
   );
   gpc615_5 gpc5738 (
      {stage1_58[205], stage1_58[206], stage1_58[207], stage1_58[208], stage1_58[209]},
      {stage1_59[30]},
      {stage1_60[108], stage1_60[109], stage1_60[110], stage1_60[111], stage1_60[112], stage1_60[113]},
      {stage2_62[18],stage2_61[20],stage2_60[33],stage2_59[77],stage2_58[83]}
   );
   gpc615_5 gpc5739 (
      {stage1_58[210], stage1_58[211], stage1_58[212], stage1_58[213], stage1_58[214]},
      {stage1_59[31]},
      {stage1_60[114], stage1_60[115], stage1_60[116], stage1_60[117], stage1_60[118], stage1_60[119]},
      {stage2_62[19],stage2_61[21],stage2_60[34],stage2_59[78],stage2_58[84]}
   );
   gpc615_5 gpc5740 (
      {stage1_58[215], stage1_58[216], stage1_58[217], stage1_58[218], stage1_58[219]},
      {stage1_59[32]},
      {stage1_60[120], stage1_60[121], stage1_60[122], stage1_60[123], stage1_60[124], stage1_60[125]},
      {stage2_62[20],stage2_61[22],stage2_60[35],stage2_59[79],stage2_58[85]}
   );
   gpc2135_5 gpc5741 (
      {stage1_59[33], stage1_59[34], stage1_59[35], stage1_59[36], stage1_59[37]},
      {stage1_60[126], stage1_60[127], stage1_60[128]},
      {stage1_61[0]},
      {stage1_62[0], stage1_62[1]},
      {stage2_63[0],stage2_62[21],stage2_61[23],stage2_60[36],stage2_59[80]}
   );
   gpc606_5 gpc5742 (
      {stage1_59[38], stage1_59[39], stage1_59[40], stage1_59[41], stage1_59[42], stage1_59[43]},
      {stage1_61[1], stage1_61[2], stage1_61[3], stage1_61[4], stage1_61[5], stage1_61[6]},
      {stage2_63[1],stage2_62[22],stage2_61[24],stage2_60[37],stage2_59[81]}
   );
   gpc606_5 gpc5743 (
      {stage1_59[44], stage1_59[45], stage1_59[46], stage1_59[47], stage1_59[48], stage1_59[49]},
      {stage1_61[7], stage1_61[8], stage1_61[9], stage1_61[10], stage1_61[11], stage1_61[12]},
      {stage2_63[2],stage2_62[23],stage2_61[25],stage2_60[38],stage2_59[82]}
   );
   gpc606_5 gpc5744 (
      {stage1_59[50], stage1_59[51], stage1_59[52], stage1_59[53], stage1_59[54], stage1_59[55]},
      {stage1_61[13], stage1_61[14], stage1_61[15], stage1_61[16], stage1_61[17], stage1_61[18]},
      {stage2_63[3],stage2_62[24],stage2_61[26],stage2_60[39],stage2_59[83]}
   );
   gpc606_5 gpc5745 (
      {stage1_59[56], stage1_59[57], stage1_59[58], stage1_59[59], stage1_59[60], stage1_59[61]},
      {stage1_61[19], stage1_61[20], stage1_61[21], stage1_61[22], stage1_61[23], stage1_61[24]},
      {stage2_63[4],stage2_62[25],stage2_61[27],stage2_60[40],stage2_59[84]}
   );
   gpc606_5 gpc5746 (
      {stage1_59[62], stage1_59[63], stage1_59[64], stage1_59[65], stage1_59[66], stage1_59[67]},
      {stage1_61[25], stage1_61[26], stage1_61[27], stage1_61[28], stage1_61[29], stage1_61[30]},
      {stage2_63[5],stage2_62[26],stage2_61[28],stage2_60[41],stage2_59[85]}
   );
   gpc606_5 gpc5747 (
      {stage1_59[68], stage1_59[69], stage1_59[70], stage1_59[71], stage1_59[72], stage1_59[73]},
      {stage1_61[31], stage1_61[32], stage1_61[33], stage1_61[34], stage1_61[35], stage1_61[36]},
      {stage2_63[6],stage2_62[27],stage2_61[29],stage2_60[42],stage2_59[86]}
   );
   gpc606_5 gpc5748 (
      {stage1_59[74], stage1_59[75], stage1_59[76], stage1_59[77], stage1_59[78], stage1_59[79]},
      {stage1_61[37], stage1_61[38], stage1_61[39], stage1_61[40], stage1_61[41], stage1_61[42]},
      {stage2_63[7],stage2_62[28],stage2_61[30],stage2_60[43],stage2_59[87]}
   );
   gpc606_5 gpc5749 (
      {stage1_59[80], stage1_59[81], stage1_59[82], stage1_59[83], stage1_59[84], stage1_59[85]},
      {stage1_61[43], stage1_61[44], stage1_61[45], stage1_61[46], stage1_61[47], stage1_61[48]},
      {stage2_63[8],stage2_62[29],stage2_61[31],stage2_60[44],stage2_59[88]}
   );
   gpc606_5 gpc5750 (
      {stage1_59[86], stage1_59[87], stage1_59[88], stage1_59[89], stage1_59[90], stage1_59[91]},
      {stage1_61[49], stage1_61[50], stage1_61[51], stage1_61[52], stage1_61[53], stage1_61[54]},
      {stage2_63[9],stage2_62[30],stage2_61[32],stage2_60[45],stage2_59[89]}
   );
   gpc606_5 gpc5751 (
      {stage1_59[92], stage1_59[93], stage1_59[94], stage1_59[95], stage1_59[96], stage1_59[97]},
      {stage1_61[55], stage1_61[56], stage1_61[57], stage1_61[58], stage1_61[59], stage1_61[60]},
      {stage2_63[10],stage2_62[31],stage2_61[33],stage2_60[46],stage2_59[90]}
   );
   gpc606_5 gpc5752 (
      {stage1_59[98], stage1_59[99], stage1_59[100], stage1_59[101], stage1_59[102], stage1_59[103]},
      {stage1_61[61], stage1_61[62], stage1_61[63], stage1_61[64], stage1_61[65], stage1_61[66]},
      {stage2_63[11],stage2_62[32],stage2_61[34],stage2_60[47],stage2_59[91]}
   );
   gpc606_5 gpc5753 (
      {stage1_59[104], stage1_59[105], stage1_59[106], stage1_59[107], stage1_59[108], stage1_59[109]},
      {stage1_61[67], stage1_61[68], stage1_61[69], stage1_61[70], stage1_61[71], stage1_61[72]},
      {stage2_63[12],stage2_62[33],stage2_61[35],stage2_60[48],stage2_59[92]}
   );
   gpc606_5 gpc5754 (
      {stage1_59[110], stage1_59[111], stage1_59[112], stage1_59[113], stage1_59[114], stage1_59[115]},
      {stage1_61[73], stage1_61[74], stage1_61[75], stage1_61[76], stage1_61[77], stage1_61[78]},
      {stage2_63[13],stage2_62[34],stage2_61[36],stage2_60[49],stage2_59[93]}
   );
   gpc606_5 gpc5755 (
      {stage1_59[116], stage1_59[117], stage1_59[118], stage1_59[119], stage1_59[120], stage1_59[121]},
      {stage1_61[79], stage1_61[80], stage1_61[81], stage1_61[82], stage1_61[83], stage1_61[84]},
      {stage2_63[14],stage2_62[35],stage2_61[37],stage2_60[50],stage2_59[94]}
   );
   gpc606_5 gpc5756 (
      {stage1_59[122], stage1_59[123], stage1_59[124], stage1_59[125], stage1_59[126], stage1_59[127]},
      {stage1_61[85], stage1_61[86], stage1_61[87], stage1_61[88], stage1_61[89], stage1_61[90]},
      {stage2_63[15],stage2_62[36],stage2_61[38],stage2_60[51],stage2_59[95]}
   );
   gpc606_5 gpc5757 (
      {stage1_59[128], stage1_59[129], stage1_59[130], stage1_59[131], stage1_59[132], stage1_59[133]},
      {stage1_61[91], stage1_61[92], stage1_61[93], stage1_61[94], stage1_61[95], stage1_61[96]},
      {stage2_63[16],stage2_62[37],stage2_61[39],stage2_60[52],stage2_59[96]}
   );
   gpc606_5 gpc5758 (
      {stage1_59[134], stage1_59[135], stage1_59[136], stage1_59[137], stage1_59[138], stage1_59[139]},
      {stage1_61[97], stage1_61[98], stage1_61[99], stage1_61[100], stage1_61[101], stage1_61[102]},
      {stage2_63[17],stage2_62[38],stage2_61[40],stage2_60[53],stage2_59[97]}
   );
   gpc606_5 gpc5759 (
      {stage1_59[140], stage1_59[141], stage1_59[142], stage1_59[143], stage1_59[144], stage1_59[145]},
      {stage1_61[103], stage1_61[104], stage1_61[105], stage1_61[106], stage1_61[107], stage1_61[108]},
      {stage2_63[18],stage2_62[39],stage2_61[41],stage2_60[54],stage2_59[98]}
   );
   gpc606_5 gpc5760 (
      {stage1_59[146], stage1_59[147], stage1_59[148], stage1_59[149], stage1_59[150], stage1_59[151]},
      {stage1_61[109], stage1_61[110], stage1_61[111], stage1_61[112], stage1_61[113], stage1_61[114]},
      {stage2_63[19],stage2_62[40],stage2_61[42],stage2_60[55],stage2_59[99]}
   );
   gpc606_5 gpc5761 (
      {stage1_59[152], stage1_59[153], stage1_59[154], stage1_59[155], stage1_59[156], stage1_59[157]},
      {stage1_61[115], stage1_61[116], stage1_61[117], stage1_61[118], stage1_61[119], stage1_61[120]},
      {stage2_63[20],stage2_62[41],stage2_61[43],stage2_60[56],stage2_59[100]}
   );
   gpc606_5 gpc5762 (
      {stage1_59[158], stage1_59[159], stage1_59[160], stage1_59[161], stage1_59[162], stage1_59[163]},
      {stage1_61[121], stage1_61[122], stage1_61[123], stage1_61[124], stage1_61[125], stage1_61[126]},
      {stage2_63[21],stage2_62[42],stage2_61[44],stage2_60[57],stage2_59[101]}
   );
   gpc606_5 gpc5763 (
      {stage1_59[164], stage1_59[165], stage1_59[166], stage1_59[167], stage1_59[168], stage1_59[169]},
      {stage1_61[127], stage1_61[128], stage1_61[129], stage1_61[130], stage1_61[131], stage1_61[132]},
      {stage2_63[22],stage2_62[43],stage2_61[45],stage2_60[58],stage2_59[102]}
   );
   gpc606_5 gpc5764 (
      {stage1_59[170], stage1_59[171], stage1_59[172], stage1_59[173], stage1_59[174], stage1_59[175]},
      {stage1_61[133], stage1_61[134], stage1_61[135], stage1_61[136], stage1_61[137], stage1_61[138]},
      {stage2_63[23],stage2_62[44],stage2_61[46],stage2_60[59],stage2_59[103]}
   );
   gpc606_5 gpc5765 (
      {stage1_59[176], stage1_59[177], stage1_59[178], stage1_59[179], stage1_59[180], stage1_59[181]},
      {stage1_61[139], stage1_61[140], stage1_61[141], stage1_61[142], stage1_61[143], stage1_61[144]},
      {stage2_63[24],stage2_62[45],stage2_61[47],stage2_60[60],stage2_59[104]}
   );
   gpc606_5 gpc5766 (
      {stage1_59[182], stage1_59[183], stage1_59[184], stage1_59[185], stage1_59[186], stage1_59[187]},
      {stage1_61[145], stage1_61[146], stage1_61[147], stage1_61[148], stage1_61[149], stage1_61[150]},
      {stage2_63[25],stage2_62[46],stage2_61[48],stage2_60[61],stage2_59[105]}
   );
   gpc606_5 gpc5767 (
      {stage1_59[188], stage1_59[189], stage1_59[190], stage1_59[191], stage1_59[192], stage1_59[193]},
      {stage1_61[151], stage1_61[152], stage1_61[153], stage1_61[154], stage1_61[155], stage1_61[156]},
      {stage2_63[26],stage2_62[47],stage2_61[49],stage2_60[62],stage2_59[106]}
   );
   gpc606_5 gpc5768 (
      {stage1_59[194], stage1_59[195], stage1_59[196], stage1_59[197], stage1_59[198], stage1_59[199]},
      {stage1_61[157], stage1_61[158], stage1_61[159], stage1_61[160], stage1_61[161], stage1_61[162]},
      {stage2_63[27],stage2_62[48],stage2_61[50],stage2_60[63],stage2_59[107]}
   );
   gpc615_5 gpc5769 (
      {stage1_59[200], stage1_59[201], stage1_59[202], stage1_59[203], stage1_59[204]},
      {stage1_60[129]},
      {stage1_61[163], stage1_61[164], stage1_61[165], stage1_61[166], stage1_61[167], stage1_61[168]},
      {stage2_63[28],stage2_62[49],stage2_61[51],stage2_60[64],stage2_59[108]}
   );
   gpc606_5 gpc5770 (
      {stage1_60[130], stage1_60[131], stage1_60[132], stage1_60[133], stage1_60[134], stage1_60[135]},
      {stage1_62[2], stage1_62[3], stage1_62[4], stage1_62[5], stage1_62[6], stage1_62[7]},
      {stage2_64[0],stage2_63[29],stage2_62[50],stage2_61[52],stage2_60[65]}
   );
   gpc606_5 gpc5771 (
      {stage1_60[136], stage1_60[137], stage1_60[138], stage1_60[139], stage1_60[140], stage1_60[141]},
      {stage1_62[8], stage1_62[9], stage1_62[10], stage1_62[11], stage1_62[12], stage1_62[13]},
      {stage2_64[1],stage2_63[30],stage2_62[51],stage2_61[53],stage2_60[66]}
   );
   gpc606_5 gpc5772 (
      {stage1_60[142], stage1_60[143], stage1_60[144], stage1_60[145], stage1_60[146], stage1_60[147]},
      {stage1_62[14], stage1_62[15], stage1_62[16], stage1_62[17], stage1_62[18], stage1_62[19]},
      {stage2_64[2],stage2_63[31],stage2_62[52],stage2_61[54],stage2_60[67]}
   );
   gpc606_5 gpc5773 (
      {stage1_60[148], stage1_60[149], stage1_60[150], stage1_60[151], stage1_60[152], stage1_60[153]},
      {stage1_62[20], stage1_62[21], stage1_62[22], stage1_62[23], stage1_62[24], stage1_62[25]},
      {stage2_64[3],stage2_63[32],stage2_62[53],stage2_61[55],stage2_60[68]}
   );
   gpc606_5 gpc5774 (
      {stage1_60[154], stage1_60[155], stage1_60[156], stage1_60[157], stage1_60[158], stage1_60[159]},
      {stage1_62[26], stage1_62[27], stage1_62[28], stage1_62[29], stage1_62[30], stage1_62[31]},
      {stage2_64[4],stage2_63[33],stage2_62[54],stage2_61[56],stage2_60[69]}
   );
   gpc606_5 gpc5775 (
      {stage1_60[160], stage1_60[161], stage1_60[162], stage1_60[163], stage1_60[164], stage1_60[165]},
      {stage1_62[32], stage1_62[33], stage1_62[34], stage1_62[35], stage1_62[36], stage1_62[37]},
      {stage2_64[5],stage2_63[34],stage2_62[55],stage2_61[57],stage2_60[70]}
   );
   gpc606_5 gpc5776 (
      {stage1_60[166], stage1_60[167], stage1_60[168], stage1_60[169], stage1_60[170], stage1_60[171]},
      {stage1_62[38], stage1_62[39], stage1_62[40], stage1_62[41], stage1_62[42], stage1_62[43]},
      {stage2_64[6],stage2_63[35],stage2_62[56],stage2_61[58],stage2_60[71]}
   );
   gpc606_5 gpc5777 (
      {stage1_60[172], stage1_60[173], stage1_60[174], stage1_60[175], stage1_60[176], stage1_60[177]},
      {stage1_62[44], stage1_62[45], stage1_62[46], stage1_62[47], stage1_62[48], stage1_62[49]},
      {stage2_64[7],stage2_63[36],stage2_62[57],stage2_61[59],stage2_60[72]}
   );
   gpc606_5 gpc5778 (
      {stage1_60[178], stage1_60[179], stage1_60[180], stage1_60[181], stage1_60[182], stage1_60[183]},
      {stage1_62[50], stage1_62[51], stage1_62[52], stage1_62[53], stage1_62[54], stage1_62[55]},
      {stage2_64[8],stage2_63[37],stage2_62[58],stage2_61[60],stage2_60[73]}
   );
   gpc615_5 gpc5779 (
      {stage1_60[184], stage1_60[185], stage1_60[186], stage1_60[187], stage1_60[188]},
      {stage1_61[169]},
      {stage1_62[56], stage1_62[57], stage1_62[58], stage1_62[59], stage1_62[60], stage1_62[61]},
      {stage2_64[9],stage2_63[38],stage2_62[59],stage2_61[61],stage2_60[74]}
   );
   gpc615_5 gpc5780 (
      {stage1_60[189], stage1_60[190], stage1_60[191], stage1_60[192], stage1_60[193]},
      {stage1_61[170]},
      {stage1_62[62], stage1_62[63], stage1_62[64], stage1_62[65], stage1_62[66], stage1_62[67]},
      {stage2_64[10],stage2_63[39],stage2_62[60],stage2_61[62],stage2_60[75]}
   );
   gpc615_5 gpc5781 (
      {stage1_60[194], stage1_60[195], stage1_60[196], stage1_60[197], stage1_60[198]},
      {stage1_61[171]},
      {stage1_62[68], stage1_62[69], stage1_62[70], stage1_62[71], stage1_62[72], stage1_62[73]},
      {stage2_64[11],stage2_63[40],stage2_62[61],stage2_61[63],stage2_60[76]}
   );
   gpc615_5 gpc5782 (
      {stage1_60[199], stage1_60[200], stage1_60[201], stage1_60[202], stage1_60[203]},
      {stage1_61[172]},
      {stage1_62[74], stage1_62[75], stage1_62[76], stage1_62[77], stage1_62[78], stage1_62[79]},
      {stage2_64[12],stage2_63[41],stage2_62[62],stage2_61[64],stage2_60[77]}
   );
   gpc615_5 gpc5783 (
      {stage1_60[204], stage1_60[205], stage1_60[206], stage1_60[207], stage1_60[208]},
      {stage1_61[173]},
      {stage1_62[80], stage1_62[81], stage1_62[82], stage1_62[83], stage1_62[84], stage1_62[85]},
      {stage2_64[13],stage2_63[42],stage2_62[63],stage2_61[65],stage2_60[78]}
   );
   gpc615_5 gpc5784 (
      {stage1_61[174], stage1_61[175], stage1_61[176], stage1_61[177], stage1_61[178]},
      {stage1_62[86]},
      {stage1_63[0], stage1_63[1], stage1_63[2], stage1_63[3], stage1_63[4], stage1_63[5]},
      {stage2_65[0],stage2_64[14],stage2_63[43],stage2_62[64],stage2_61[66]}
   );
   gpc615_5 gpc5785 (
      {stage1_61[179], stage1_61[180], stage1_61[181], stage1_61[182], stage1_61[183]},
      {stage1_62[87]},
      {stage1_63[6], stage1_63[7], stage1_63[8], stage1_63[9], stage1_63[10], stage1_63[11]},
      {stage2_65[1],stage2_64[15],stage2_63[44],stage2_62[65],stage2_61[67]}
   );
   gpc615_5 gpc5786 (
      {stage1_61[184], stage1_61[185], stage1_61[186], stage1_61[187], stage1_61[188]},
      {stage1_62[88]},
      {stage1_63[12], stage1_63[13], stage1_63[14], stage1_63[15], stage1_63[16], stage1_63[17]},
      {stage2_65[2],stage2_64[16],stage2_63[45],stage2_62[66],stage2_61[68]}
   );
   gpc615_5 gpc5787 (
      {stage1_61[189], stage1_61[190], stage1_61[191], stage1_61[192], stage1_61[193]},
      {stage1_62[89]},
      {stage1_63[18], stage1_63[19], stage1_63[20], stage1_63[21], stage1_63[22], stage1_63[23]},
      {stage2_65[3],stage2_64[17],stage2_63[46],stage2_62[67],stage2_61[69]}
   );
   gpc615_5 gpc5788 (
      {stage1_61[194], stage1_61[195], stage1_61[196], stage1_61[197], stage1_61[198]},
      {stage1_62[90]},
      {stage1_63[24], stage1_63[25], stage1_63[26], stage1_63[27], stage1_63[28], stage1_63[29]},
      {stage2_65[4],stage2_64[18],stage2_63[47],stage2_62[68],stage2_61[70]}
   );
   gpc615_5 gpc5789 (
      {stage1_61[199], stage1_61[200], stage1_61[201], stage1_61[202], stage1_61[203]},
      {stage1_62[91]},
      {stage1_63[30], stage1_63[31], stage1_63[32], stage1_63[33], stage1_63[34], stage1_63[35]},
      {stage2_65[5],stage2_64[19],stage2_63[48],stage2_62[69],stage2_61[71]}
   );
   gpc615_5 gpc5790 (
      {stage1_61[204], stage1_61[205], stage1_61[206], stage1_61[207], stage1_61[208]},
      {stage1_62[92]},
      {stage1_63[36], stage1_63[37], stage1_63[38], stage1_63[39], stage1_63[40], stage1_63[41]},
      {stage2_65[6],stage2_64[20],stage2_63[49],stage2_62[70],stage2_61[72]}
   );
   gpc615_5 gpc5791 (
      {stage1_61[209], stage1_61[210], stage1_61[211], stage1_61[212], stage1_61[213]},
      {stage1_62[93]},
      {stage1_63[42], stage1_63[43], stage1_63[44], stage1_63[45], stage1_63[46], stage1_63[47]},
      {stage2_65[7],stage2_64[21],stage2_63[50],stage2_62[71],stage2_61[73]}
   );
   gpc615_5 gpc5792 (
      {stage1_61[214], stage1_61[215], stage1_61[216], stage1_61[217], stage1_61[218]},
      {stage1_62[94]},
      {stage1_63[48], stage1_63[49], stage1_63[50], stage1_63[51], stage1_63[52], stage1_63[53]},
      {stage2_65[8],stage2_64[22],stage2_63[51],stage2_62[72],stage2_61[74]}
   );
   gpc1163_5 gpc5793 (
      {stage1_62[95], stage1_62[96], stage1_62[97]},
      {stage1_63[54], stage1_63[55], stage1_63[56], stage1_63[57], stage1_63[58], stage1_63[59]},
      {stage1_64[0]},
      {stage1_65[0]},
      {stage2_66[0],stage2_65[9],stage2_64[23],stage2_63[52],stage2_62[73]}
   );
   gpc1163_5 gpc5794 (
      {stage1_62[98], stage1_62[99], stage1_62[100]},
      {stage1_63[60], stage1_63[61], stage1_63[62], stage1_63[63], stage1_63[64], stage1_63[65]},
      {stage1_64[1]},
      {stage1_65[1]},
      {stage2_66[1],stage2_65[10],stage2_64[24],stage2_63[53],stage2_62[74]}
   );
   gpc1163_5 gpc5795 (
      {stage1_62[101], stage1_62[102], stage1_62[103]},
      {stage1_63[66], stage1_63[67], stage1_63[68], stage1_63[69], stage1_63[70], stage1_63[71]},
      {stage1_64[2]},
      {stage1_65[2]},
      {stage2_66[2],stage2_65[11],stage2_64[25],stage2_63[54],stage2_62[75]}
   );
   gpc1163_5 gpc5796 (
      {stage1_62[104], stage1_62[105], stage1_62[106]},
      {stage1_63[72], stage1_63[73], stage1_63[74], stage1_63[75], stage1_63[76], stage1_63[77]},
      {stage1_64[3]},
      {stage1_65[3]},
      {stage2_66[3],stage2_65[12],stage2_64[26],stage2_63[55],stage2_62[76]}
   );
   gpc1163_5 gpc5797 (
      {stage1_62[107], stage1_62[108], stage1_62[109]},
      {stage1_63[78], stage1_63[79], stage1_63[80], stage1_63[81], stage1_63[82], stage1_63[83]},
      {stage1_64[4]},
      {stage1_65[4]},
      {stage2_66[4],stage2_65[13],stage2_64[27],stage2_63[56],stage2_62[77]}
   );
   gpc1163_5 gpc5798 (
      {stage1_62[110], stage1_62[111], stage1_62[112]},
      {stage1_63[84], stage1_63[85], stage1_63[86], stage1_63[87], stage1_63[88], stage1_63[89]},
      {stage1_64[5]},
      {stage1_65[5]},
      {stage2_66[5],stage2_65[14],stage2_64[28],stage2_63[57],stage2_62[78]}
   );
   gpc1163_5 gpc5799 (
      {stage1_62[113], stage1_62[114], stage1_62[115]},
      {stage1_63[90], stage1_63[91], stage1_63[92], stage1_63[93], stage1_63[94], stage1_63[95]},
      {stage1_64[6]},
      {stage1_65[6]},
      {stage2_66[6],stage2_65[15],stage2_64[29],stage2_63[58],stage2_62[79]}
   );
   gpc1163_5 gpc5800 (
      {stage1_62[116], stage1_62[117], stage1_62[118]},
      {stage1_63[96], stage1_63[97], stage1_63[98], stage1_63[99], stage1_63[100], stage1_63[101]},
      {stage1_64[7]},
      {stage1_65[7]},
      {stage2_66[7],stage2_65[16],stage2_64[30],stage2_63[59],stage2_62[80]}
   );
   gpc1163_5 gpc5801 (
      {stage1_62[119], stage1_62[120], stage1_62[121]},
      {stage1_63[102], stage1_63[103], stage1_63[104], stage1_63[105], stage1_63[106], stage1_63[107]},
      {stage1_64[8]},
      {stage1_65[8]},
      {stage2_66[8],stage2_65[17],stage2_64[31],stage2_63[60],stage2_62[81]}
   );
   gpc1163_5 gpc5802 (
      {stage1_62[122], stage1_62[123], stage1_62[124]},
      {stage1_63[108], stage1_63[109], stage1_63[110], stage1_63[111], stage1_63[112], stage1_63[113]},
      {stage1_64[9]},
      {stage1_65[9]},
      {stage2_66[9],stage2_65[18],stage2_64[32],stage2_63[61],stage2_62[82]}
   );
   gpc1163_5 gpc5803 (
      {stage1_62[125], stage1_62[126], stage1_62[127]},
      {stage1_63[114], stage1_63[115], stage1_63[116], stage1_63[117], stage1_63[118], stage1_63[119]},
      {stage1_64[10]},
      {stage1_65[10]},
      {stage2_66[10],stage2_65[19],stage2_64[33],stage2_63[62],stage2_62[83]}
   );
   gpc1163_5 gpc5804 (
      {stage1_62[128], stage1_62[129], stage1_62[130]},
      {stage1_63[120], stage1_63[121], stage1_63[122], stage1_63[123], stage1_63[124], stage1_63[125]},
      {stage1_64[11]},
      {stage1_65[11]},
      {stage2_66[11],stage2_65[20],stage2_64[34],stage2_63[63],stage2_62[84]}
   );
   gpc1163_5 gpc5805 (
      {stage1_62[131], stage1_62[132], stage1_62[133]},
      {stage1_63[126], stage1_63[127], stage1_63[128], stage1_63[129], stage1_63[130], stage1_63[131]},
      {stage1_64[12]},
      {stage1_65[12]},
      {stage2_66[12],stage2_65[21],stage2_64[35],stage2_63[64],stage2_62[85]}
   );
   gpc1163_5 gpc5806 (
      {stage1_62[134], stage1_62[135], stage1_62[136]},
      {stage1_63[132], stage1_63[133], stage1_63[134], stage1_63[135], stage1_63[136], stage1_63[137]},
      {stage1_64[13]},
      {stage1_65[13]},
      {stage2_66[13],stage2_65[22],stage2_64[36],stage2_63[65],stage2_62[86]}
   );
   gpc1163_5 gpc5807 (
      {stage1_62[137], stage1_62[138], stage1_62[139]},
      {stage1_63[138], stage1_63[139], stage1_63[140], stage1_63[141], stage1_63[142], stage1_63[143]},
      {stage1_64[14]},
      {stage1_65[14]},
      {stage2_66[14],stage2_65[23],stage2_64[37],stage2_63[66],stage2_62[87]}
   );
   gpc1163_5 gpc5808 (
      {stage1_62[140], stage1_62[141], stage1_62[142]},
      {stage1_63[144], stage1_63[145], stage1_63[146], stage1_63[147], stage1_63[148], stage1_63[149]},
      {stage1_64[15]},
      {stage1_65[15]},
      {stage2_66[15],stage2_65[24],stage2_64[38],stage2_63[67],stage2_62[88]}
   );
   gpc1163_5 gpc5809 (
      {stage1_62[143], stage1_62[144], stage1_62[145]},
      {stage1_63[150], stage1_63[151], stage1_63[152], stage1_63[153], stage1_63[154], stage1_63[155]},
      {stage1_64[16]},
      {stage1_65[16]},
      {stage2_66[16],stage2_65[25],stage2_64[39],stage2_63[68],stage2_62[89]}
   );
   gpc1163_5 gpc5810 (
      {stage1_62[146], stage1_62[147], stage1_62[148]},
      {stage1_63[156], stage1_63[157], stage1_63[158], stage1_63[159], stage1_63[160], stage1_63[161]},
      {stage1_64[17]},
      {stage1_65[17]},
      {stage2_66[17],stage2_65[26],stage2_64[40],stage2_63[69],stage2_62[90]}
   );
   gpc1163_5 gpc5811 (
      {stage1_62[149], stage1_62[150], stage1_62[151]},
      {stage1_63[162], stage1_63[163], stage1_63[164], stage1_63[165], stage1_63[166], stage1_63[167]},
      {stage1_64[18]},
      {stage1_65[18]},
      {stage2_66[18],stage2_65[27],stage2_64[41],stage2_63[70],stage2_62[91]}
   );
   gpc1163_5 gpc5812 (
      {stage1_62[152], stage1_62[153], stage1_62[154]},
      {stage1_63[168], stage1_63[169], stage1_63[170], stage1_63[171], stage1_63[172], stage1_63[173]},
      {stage1_64[19]},
      {stage1_65[19]},
      {stage2_66[19],stage2_65[28],stage2_64[42],stage2_63[71],stage2_62[92]}
   );
   gpc1163_5 gpc5813 (
      {stage1_62[155], stage1_62[156], stage1_62[157]},
      {stage1_63[174], stage1_63[175], stage1_63[176], stage1_63[177], stage1_63[178], stage1_63[179]},
      {stage1_64[20]},
      {stage1_65[20]},
      {stage2_66[20],stage2_65[29],stage2_64[43],stage2_63[72],stage2_62[93]}
   );
   gpc1163_5 gpc5814 (
      {stage1_62[158], stage1_62[159], stage1_62[160]},
      {stage1_63[180], stage1_63[181], stage1_63[182], stage1_63[183], stage1_63[184], stage1_63[185]},
      {stage1_64[21]},
      {stage1_65[21]},
      {stage2_66[21],stage2_65[30],stage2_64[44],stage2_63[73],stage2_62[94]}
   );
   gpc1163_5 gpc5815 (
      {stage1_62[161], stage1_62[162], stage1_62[163]},
      {stage1_63[186], stage1_63[187], stage1_63[188], stage1_63[189], stage1_63[190], stage1_63[191]},
      {stage1_64[22]},
      {stage1_65[22]},
      {stage2_66[22],stage2_65[31],stage2_64[45],stage2_63[74],stage2_62[95]}
   );
   gpc1163_5 gpc5816 (
      {stage1_62[164], stage1_62[165], stage1_62[166]},
      {stage1_63[192], stage1_63[193], stage1_63[194], stage1_63[195], stage1_63[196], stage1_63[197]},
      {stage1_64[23]},
      {stage1_65[23]},
      {stage2_66[23],stage2_65[32],stage2_64[46],stage2_63[75],stage2_62[96]}
   );
   gpc1163_5 gpc5817 (
      {stage1_62[167], stage1_62[168], stage1_62[169]},
      {stage1_63[198], stage1_63[199], stage1_63[200], stage1_63[201], stage1_63[202], stage1_63[203]},
      {stage1_64[24]},
      {stage1_65[24]},
      {stage2_66[24],stage2_65[33],stage2_64[47],stage2_63[76],stage2_62[97]}
   );
   gpc1163_5 gpc5818 (
      {stage1_62[170], stage1_62[171], stage1_62[172]},
      {stage1_63[204], stage1_63[205], stage1_63[206], stage1_63[207], stage1_63[208], stage1_63[209]},
      {stage1_64[25]},
      {stage1_65[25]},
      {stage2_66[25],stage2_65[34],stage2_64[48],stage2_63[77],stage2_62[98]}
   );
   gpc1163_5 gpc5819 (
      {stage1_62[173], stage1_62[174], stage1_62[175]},
      {stage1_63[210], stage1_63[211], stage1_63[212], stage1_63[213], stage1_63[214], stage1_63[215]},
      {stage1_64[26]},
      {stage1_65[26]},
      {stage2_66[26],stage2_65[35],stage2_64[49],stage2_63[78],stage2_62[99]}
   );
   gpc1163_5 gpc5820 (
      {stage1_62[176], stage1_62[177], stage1_62[178]},
      {stage1_63[216], stage1_63[217], stage1_63[218], stage1_63[219], stage1_63[220], stage1_63[221]},
      {stage1_64[27]},
      {stage1_65[27]},
      {stage2_66[27],stage2_65[36],stage2_64[50],stage2_63[79],stage2_62[100]}
   );
   gpc1163_5 gpc5821 (
      {stage1_62[179], stage1_62[180], stage1_62[181]},
      {stage1_63[222], stage1_63[223], stage1_63[224], stage1_63[225], stage1_63[226], stage1_63[227]},
      {stage1_64[28]},
      {stage1_65[28]},
      {stage2_66[28],stage2_65[37],stage2_64[51],stage2_63[80],stage2_62[101]}
   );
   gpc615_5 gpc5822 (
      {stage1_62[182], stage1_62[183], stage1_62[184], stage1_62[185], stage1_62[186]},
      {stage1_63[228]},
      {stage1_64[29], stage1_64[30], stage1_64[31], stage1_64[32], stage1_64[33], stage1_64[34]},
      {stage2_66[29],stage2_65[38],stage2_64[52],stage2_63[81],stage2_62[102]}
   );
   gpc615_5 gpc5823 (
      {stage1_62[187], stage1_62[188], stage1_62[189], stage1_62[190], stage1_62[191]},
      {stage1_63[229]},
      {stage1_64[35], stage1_64[36], stage1_64[37], stage1_64[38], stage1_64[39], stage1_64[40]},
      {stage2_66[30],stage2_65[39],stage2_64[53],stage2_63[82],stage2_62[103]}
   );
   gpc135_4 gpc5824 (
      {stage1_63[230], stage1_63[231], stage1_63[232], stage1_63[233], stage1_63[234]},
      {stage1_64[41], stage1_64[42], stage1_64[43]},
      {stage1_65[29]},
      {stage2_66[31],stage2_65[40],stage2_64[54],stage2_63[83]}
   );
   gpc135_4 gpc5825 (
      {stage1_63[235], stage1_63[236], stage1_63[237], stage1_63[238], stage1_63[239]},
      {stage1_64[44], stage1_64[45], stage1_64[46]},
      {stage1_65[30]},
      {stage2_66[32],stage2_65[41],stage2_64[55],stage2_63[84]}
   );
   gpc207_4 gpc5826 (
      {stage1_63[240], stage1_63[241], stage1_63[242], stage1_63[243], stage1_63[244], stage1_63[245], stage1_63[246]},
      {stage1_65[31], stage1_65[32]},
      {stage2_66[33],stage2_65[42],stage2_64[56],stage2_63[85]}
   );
   gpc207_4 gpc5827 (
      {stage1_63[247], stage1_63[248], stage1_63[249], stage1_63[250], stage1_63[251], stage1_63[252], stage1_63[253]},
      {stage1_65[33], stage1_65[34]},
      {stage2_66[34],stage2_65[43],stage2_64[57],stage2_63[86]}
   );
   gpc207_4 gpc5828 (
      {stage1_63[254], stage1_63[255], stage1_63[256], stage1_63[257], stage1_63[258], stage1_63[259], stage1_63[260]},
      {stage1_65[35], stage1_65[36]},
      {stage2_66[35],stage2_65[44],stage2_64[58],stage2_63[87]}
   );
   gpc207_4 gpc5829 (
      {stage1_63[261], stage1_63[262], stage1_63[263], stage1_63[264], stage1_63[265], stage1_63[266], stage1_63[267]},
      {stage1_65[37], stage1_65[38]},
      {stage2_66[36],stage2_65[45],stage2_64[59],stage2_63[88]}
   );
   gpc207_4 gpc5830 (
      {stage1_63[268], stage1_63[269], stage1_63[270], stage1_63[271], stage1_63[272], stage1_63[273], stage1_63[274]},
      {stage1_65[39], stage1_65[40]},
      {stage2_66[37],stage2_65[46],stage2_64[60],stage2_63[89]}
   );
   gpc207_4 gpc5831 (
      {stage1_63[275], stage1_63[276], stage1_63[277], stage1_63[278], stage1_63[279], stage1_63[280], stage1_63[281]},
      {stage1_65[41], stage1_65[42]},
      {stage2_66[38],stage2_65[47],stage2_64[61],stage2_63[90]}
   );
   gpc207_4 gpc5832 (
      {stage1_63[282], stage1_63[283], stage1_63[284], stage1_63[285], stage1_63[286], stage1_63[287], stage1_63[288]},
      {stage1_65[43], stage1_65[44]},
      {stage2_66[39],stage2_65[48],stage2_64[62],stage2_63[91]}
   );
   gpc207_4 gpc5833 (
      {stage1_63[289], stage1_63[290], stage1_63[291], stage1_63[292], stage1_63[293], stage1_63[294], stage1_63[295]},
      {stage1_65[45], stage1_65[46]},
      {stage2_66[40],stage2_65[49],stage2_64[63],stage2_63[92]}
   );
   gpc207_4 gpc5834 (
      {stage1_63[296], stage1_63[297], stage1_63[298], stage1_63[299], stage1_63[300], stage1_63[301], stage1_63[302]},
      {stage1_65[47], stage1_65[48]},
      {stage2_66[41],stage2_65[50],stage2_64[64],stage2_63[93]}
   );
   gpc1_1 gpc5835 (
      {stage1_0[108]},
      {stage2_0[21]}
   );
   gpc1_1 gpc5836 (
      {stage1_0[109]},
      {stage2_0[22]}
   );
   gpc1_1 gpc5837 (
      {stage1_0[110]},
      {stage2_0[23]}
   );
   gpc1_1 gpc5838 (
      {stage1_0[111]},
      {stage2_0[24]}
   );
   gpc1_1 gpc5839 (
      {stage1_0[112]},
      {stage2_0[25]}
   );
   gpc1_1 gpc5840 (
      {stage1_0[113]},
      {stage2_0[26]}
   );
   gpc1_1 gpc5841 (
      {stage1_0[114]},
      {stage2_0[27]}
   );
   gpc1_1 gpc5842 (
      {stage1_0[115]},
      {stage2_0[28]}
   );
   gpc1_1 gpc5843 (
      {stage1_0[116]},
      {stage2_0[29]}
   );
   gpc1_1 gpc5844 (
      {stage1_0[117]},
      {stage2_0[30]}
   );
   gpc1_1 gpc5845 (
      {stage1_0[118]},
      {stage2_0[31]}
   );
   gpc1_1 gpc5846 (
      {stage1_0[119]},
      {stage2_0[32]}
   );
   gpc1_1 gpc5847 (
      {stage1_0[120]},
      {stage2_0[33]}
   );
   gpc1_1 gpc5848 (
      {stage1_0[121]},
      {stage2_0[34]}
   );
   gpc1_1 gpc5849 (
      {stage1_0[122]},
      {stage2_0[35]}
   );
   gpc1_1 gpc5850 (
      {stage1_0[123]},
      {stage2_0[36]}
   );
   gpc1_1 gpc5851 (
      {stage1_0[124]},
      {stage2_0[37]}
   );
   gpc1_1 gpc5852 (
      {stage1_1[168]},
      {stage2_1[46]}
   );
   gpc1_1 gpc5853 (
      {stage1_1[169]},
      {stage2_1[47]}
   );
   gpc1_1 gpc5854 (
      {stage1_1[170]},
      {stage2_1[48]}
   );
   gpc1_1 gpc5855 (
      {stage1_1[171]},
      {stage2_1[49]}
   );
   gpc1_1 gpc5856 (
      {stage1_1[172]},
      {stage2_1[50]}
   );
   gpc1_1 gpc5857 (
      {stage1_1[173]},
      {stage2_1[51]}
   );
   gpc1_1 gpc5858 (
      {stage1_1[174]},
      {stage2_1[52]}
   );
   gpc1_1 gpc5859 (
      {stage1_1[175]},
      {stage2_1[53]}
   );
   gpc1_1 gpc5860 (
      {stage1_2[144]},
      {stage2_2[49]}
   );
   gpc1_1 gpc5861 (
      {stage1_2[145]},
      {stage2_2[50]}
   );
   gpc1_1 gpc5862 (
      {stage1_2[146]},
      {stage2_2[51]}
   );
   gpc1_1 gpc5863 (
      {stage1_2[147]},
      {stage2_2[52]}
   );
   gpc1_1 gpc5864 (
      {stage1_2[148]},
      {stage2_2[53]}
   );
   gpc1_1 gpc5865 (
      {stage1_2[149]},
      {stage2_2[54]}
   );
   gpc1_1 gpc5866 (
      {stage1_2[150]},
      {stage2_2[55]}
   );
   gpc1_1 gpc5867 (
      {stage1_2[151]},
      {stage2_2[56]}
   );
   gpc1_1 gpc5868 (
      {stage1_2[152]},
      {stage2_2[57]}
   );
   gpc1_1 gpc5869 (
      {stage1_2[153]},
      {stage2_2[58]}
   );
   gpc1_1 gpc5870 (
      {stage1_2[154]},
      {stage2_2[59]}
   );
   gpc1_1 gpc5871 (
      {stage1_2[155]},
      {stage2_2[60]}
   );
   gpc1_1 gpc5872 (
      {stage1_2[156]},
      {stage2_2[61]}
   );
   gpc1_1 gpc5873 (
      {stage1_2[157]},
      {stage2_2[62]}
   );
   gpc1_1 gpc5874 (
      {stage1_3[150]},
      {stage2_3[49]}
   );
   gpc1_1 gpc5875 (
      {stage1_3[151]},
      {stage2_3[50]}
   );
   gpc1_1 gpc5876 (
      {stage1_3[152]},
      {stage2_3[51]}
   );
   gpc1_1 gpc5877 (
      {stage1_3[153]},
      {stage2_3[52]}
   );
   gpc1_1 gpc5878 (
      {stage1_3[154]},
      {stage2_3[53]}
   );
   gpc1_1 gpc5879 (
      {stage1_3[155]},
      {stage2_3[54]}
   );
   gpc1_1 gpc5880 (
      {stage1_3[156]},
      {stage2_3[55]}
   );
   gpc1_1 gpc5881 (
      {stage1_3[157]},
      {stage2_3[56]}
   );
   gpc1_1 gpc5882 (
      {stage1_3[158]},
      {stage2_3[57]}
   );
   gpc1_1 gpc5883 (
      {stage1_3[159]},
      {stage2_3[58]}
   );
   gpc1_1 gpc5884 (
      {stage1_3[160]},
      {stage2_3[59]}
   );
   gpc1_1 gpc5885 (
      {stage1_3[161]},
      {stage2_3[60]}
   );
   gpc1_1 gpc5886 (
      {stage1_3[162]},
      {stage2_3[61]}
   );
   gpc1_1 gpc5887 (
      {stage1_3[163]},
      {stage2_3[62]}
   );
   gpc1_1 gpc5888 (
      {stage1_3[164]},
      {stage2_3[63]}
   );
   gpc1_1 gpc5889 (
      {stage1_3[165]},
      {stage2_3[64]}
   );
   gpc1_1 gpc5890 (
      {stage1_3[166]},
      {stage2_3[65]}
   );
   gpc1_1 gpc5891 (
      {stage1_3[167]},
      {stage2_3[66]}
   );
   gpc1_1 gpc5892 (
      {stage1_3[168]},
      {stage2_3[67]}
   );
   gpc1_1 gpc5893 (
      {stage1_3[169]},
      {stage2_3[68]}
   );
   gpc1_1 gpc5894 (
      {stage1_3[170]},
      {stage2_3[69]}
   );
   gpc1_1 gpc5895 (
      {stage1_3[171]},
      {stage2_3[70]}
   );
   gpc1_1 gpc5896 (
      {stage1_3[172]},
      {stage2_3[71]}
   );
   gpc1_1 gpc5897 (
      {stage1_3[173]},
      {stage2_3[72]}
   );
   gpc1_1 gpc5898 (
      {stage1_3[174]},
      {stage2_3[73]}
   );
   gpc1_1 gpc5899 (
      {stage1_3[175]},
      {stage2_3[74]}
   );
   gpc1_1 gpc5900 (
      {stage1_3[176]},
      {stage2_3[75]}
   );
   gpc1_1 gpc5901 (
      {stage1_3[177]},
      {stage2_3[76]}
   );
   gpc1_1 gpc5902 (
      {stage1_3[178]},
      {stage2_3[77]}
   );
   gpc1_1 gpc5903 (
      {stage1_3[179]},
      {stage2_3[78]}
   );
   gpc1_1 gpc5904 (
      {stage1_3[180]},
      {stage2_3[79]}
   );
   gpc1_1 gpc5905 (
      {stage1_3[181]},
      {stage2_3[80]}
   );
   gpc1_1 gpc5906 (
      {stage1_3[182]},
      {stage2_3[81]}
   );
   gpc1_1 gpc5907 (
      {stage1_3[183]},
      {stage2_3[82]}
   );
   gpc1_1 gpc5908 (
      {stage1_3[184]},
      {stage2_3[83]}
   );
   gpc1_1 gpc5909 (
      {stage1_3[185]},
      {stage2_3[84]}
   );
   gpc1_1 gpc5910 (
      {stage1_3[186]},
      {stage2_3[85]}
   );
   gpc1_1 gpc5911 (
      {stage1_3[187]},
      {stage2_3[86]}
   );
   gpc1_1 gpc5912 (
      {stage1_3[188]},
      {stage2_3[87]}
   );
   gpc1_1 gpc5913 (
      {stage1_3[189]},
      {stage2_3[88]}
   );
   gpc1_1 gpc5914 (
      {stage1_3[190]},
      {stage2_3[89]}
   );
   gpc1_1 gpc5915 (
      {stage1_3[191]},
      {stage2_3[90]}
   );
   gpc1_1 gpc5916 (
      {stage1_3[192]},
      {stage2_3[91]}
   );
   gpc1_1 gpc5917 (
      {stage1_3[193]},
      {stage2_3[92]}
   );
   gpc1_1 gpc5918 (
      {stage1_3[194]},
      {stage2_3[93]}
   );
   gpc1_1 gpc5919 (
      {stage1_3[195]},
      {stage2_3[94]}
   );
   gpc1_1 gpc5920 (
      {stage1_3[196]},
      {stage2_3[95]}
   );
   gpc1_1 gpc5921 (
      {stage1_3[197]},
      {stage2_3[96]}
   );
   gpc1_1 gpc5922 (
      {stage1_3[198]},
      {stage2_3[97]}
   );
   gpc1_1 gpc5923 (
      {stage1_3[199]},
      {stage2_3[98]}
   );
   gpc1_1 gpc5924 (
      {stage1_3[200]},
      {stage2_3[99]}
   );
   gpc1_1 gpc5925 (
      {stage1_3[201]},
      {stage2_3[100]}
   );
   gpc1_1 gpc5926 (
      {stage1_3[202]},
      {stage2_3[101]}
   );
   gpc1_1 gpc5927 (
      {stage1_3[203]},
      {stage2_3[102]}
   );
   gpc1_1 gpc5928 (
      {stage1_3[204]},
      {stage2_3[103]}
   );
   gpc1_1 gpc5929 (
      {stage1_3[205]},
      {stage2_3[104]}
   );
   gpc1_1 gpc5930 (
      {stage1_3[206]},
      {stage2_3[105]}
   );
   gpc1_1 gpc5931 (
      {stage1_3[207]},
      {stage2_3[106]}
   );
   gpc1_1 gpc5932 (
      {stage1_3[208]},
      {stage2_3[107]}
   );
   gpc1_1 gpc5933 (
      {stage1_3[209]},
      {stage2_3[108]}
   );
   gpc1_1 gpc5934 (
      {stage1_3[210]},
      {stage2_3[109]}
   );
   gpc1_1 gpc5935 (
      {stage1_3[211]},
      {stage2_3[110]}
   );
   gpc1_1 gpc5936 (
      {stage1_3[212]},
      {stage2_3[111]}
   );
   gpc1_1 gpc5937 (
      {stage1_3[213]},
      {stage2_3[112]}
   );
   gpc1_1 gpc5938 (
      {stage1_3[214]},
      {stage2_3[113]}
   );
   gpc1_1 gpc5939 (
      {stage1_4[195]},
      {stage2_4[79]}
   );
   gpc1_1 gpc5940 (
      {stage1_4[196]},
      {stage2_4[80]}
   );
   gpc1_1 gpc5941 (
      {stage1_4[197]},
      {stage2_4[81]}
   );
   gpc1_1 gpc5942 (
      {stage1_4[198]},
      {stage2_4[82]}
   );
   gpc1_1 gpc5943 (
      {stage1_4[199]},
      {stage2_4[83]}
   );
   gpc1_1 gpc5944 (
      {stage1_4[200]},
      {stage2_4[84]}
   );
   gpc1_1 gpc5945 (
      {stage1_4[201]},
      {stage2_4[85]}
   );
   gpc1_1 gpc5946 (
      {stage1_4[202]},
      {stage2_4[86]}
   );
   gpc1_1 gpc5947 (
      {stage1_4[203]},
      {stage2_4[87]}
   );
   gpc1_1 gpc5948 (
      {stage1_4[204]},
      {stage2_4[88]}
   );
   gpc1_1 gpc5949 (
      {stage1_4[205]},
      {stage2_4[89]}
   );
   gpc1_1 gpc5950 (
      {stage1_4[206]},
      {stage2_4[90]}
   );
   gpc1_1 gpc5951 (
      {stage1_4[207]},
      {stage2_4[91]}
   );
   gpc1_1 gpc5952 (
      {stage1_4[208]},
      {stage2_4[92]}
   );
   gpc1_1 gpc5953 (
      {stage1_4[209]},
      {stage2_4[93]}
   );
   gpc1_1 gpc5954 (
      {stage1_4[210]},
      {stage2_4[94]}
   );
   gpc1_1 gpc5955 (
      {stage1_4[211]},
      {stage2_4[95]}
   );
   gpc1_1 gpc5956 (
      {stage1_4[212]},
      {stage2_4[96]}
   );
   gpc1_1 gpc5957 (
      {stage1_4[213]},
      {stage2_4[97]}
   );
   gpc1_1 gpc5958 (
      {stage1_4[214]},
      {stage2_4[98]}
   );
   gpc1_1 gpc5959 (
      {stage1_4[215]},
      {stage2_4[99]}
   );
   gpc1_1 gpc5960 (
      {stage1_4[216]},
      {stage2_4[100]}
   );
   gpc1_1 gpc5961 (
      {stage1_4[217]},
      {stage2_4[101]}
   );
   gpc1_1 gpc5962 (
      {stage1_4[218]},
      {stage2_4[102]}
   );
   gpc1_1 gpc5963 (
      {stage1_4[219]},
      {stage2_4[103]}
   );
   gpc1_1 gpc5964 (
      {stage1_4[220]},
      {stage2_4[104]}
   );
   gpc1_1 gpc5965 (
      {stage1_4[221]},
      {stage2_4[105]}
   );
   gpc1_1 gpc5966 (
      {stage1_4[222]},
      {stage2_4[106]}
   );
   gpc1_1 gpc5967 (
      {stage1_4[223]},
      {stage2_4[107]}
   );
   gpc1_1 gpc5968 (
      {stage1_4[224]},
      {stage2_4[108]}
   );
   gpc1_1 gpc5969 (
      {stage1_4[225]},
      {stage2_4[109]}
   );
   gpc1_1 gpc5970 (
      {stage1_4[226]},
      {stage2_4[110]}
   );
   gpc1_1 gpc5971 (
      {stage1_4[227]},
      {stage2_4[111]}
   );
   gpc1_1 gpc5972 (
      {stage1_5[124]},
      {stage2_5[78]}
   );
   gpc1_1 gpc5973 (
      {stage1_5[125]},
      {stage2_5[79]}
   );
   gpc1_1 gpc5974 (
      {stage1_5[126]},
      {stage2_5[80]}
   );
   gpc1_1 gpc5975 (
      {stage1_5[127]},
      {stage2_5[81]}
   );
   gpc1_1 gpc5976 (
      {stage1_5[128]},
      {stage2_5[82]}
   );
   gpc1_1 gpc5977 (
      {stage1_5[129]},
      {stage2_5[83]}
   );
   gpc1_1 gpc5978 (
      {stage1_5[130]},
      {stage2_5[84]}
   );
   gpc1_1 gpc5979 (
      {stage1_5[131]},
      {stage2_5[85]}
   );
   gpc1_1 gpc5980 (
      {stage1_5[132]},
      {stage2_5[86]}
   );
   gpc1_1 gpc5981 (
      {stage1_5[133]},
      {stage2_5[87]}
   );
   gpc1_1 gpc5982 (
      {stage1_5[134]},
      {stage2_5[88]}
   );
   gpc1_1 gpc5983 (
      {stage1_5[135]},
      {stage2_5[89]}
   );
   gpc1_1 gpc5984 (
      {stage1_5[136]},
      {stage2_5[90]}
   );
   gpc1_1 gpc5985 (
      {stage1_5[137]},
      {stage2_5[91]}
   );
   gpc1_1 gpc5986 (
      {stage1_5[138]},
      {stage2_5[92]}
   );
   gpc1_1 gpc5987 (
      {stage1_5[139]},
      {stage2_5[93]}
   );
   gpc1_1 gpc5988 (
      {stage1_5[140]},
      {stage2_5[94]}
   );
   gpc1_1 gpc5989 (
      {stage1_5[141]},
      {stage2_5[95]}
   );
   gpc1_1 gpc5990 (
      {stage1_5[142]},
      {stage2_5[96]}
   );
   gpc1_1 gpc5991 (
      {stage1_5[143]},
      {stage2_5[97]}
   );
   gpc1_1 gpc5992 (
      {stage1_5[144]},
      {stage2_5[98]}
   );
   gpc1_1 gpc5993 (
      {stage1_5[145]},
      {stage2_5[99]}
   );
   gpc1_1 gpc5994 (
      {stage1_5[146]},
      {stage2_5[100]}
   );
   gpc1_1 gpc5995 (
      {stage1_5[147]},
      {stage2_5[101]}
   );
   gpc1_1 gpc5996 (
      {stage1_5[148]},
      {stage2_5[102]}
   );
   gpc1_1 gpc5997 (
      {stage1_5[149]},
      {stage2_5[103]}
   );
   gpc1_1 gpc5998 (
      {stage1_5[150]},
      {stage2_5[104]}
   );
   gpc1_1 gpc5999 (
      {stage1_5[151]},
      {stage2_5[105]}
   );
   gpc1_1 gpc6000 (
      {stage1_5[152]},
      {stage2_5[106]}
   );
   gpc1_1 gpc6001 (
      {stage1_5[153]},
      {stage2_5[107]}
   );
   gpc1_1 gpc6002 (
      {stage1_5[154]},
      {stage2_5[108]}
   );
   gpc1_1 gpc6003 (
      {stage1_5[155]},
      {stage2_5[109]}
   );
   gpc1_1 gpc6004 (
      {stage1_5[156]},
      {stage2_5[110]}
   );
   gpc1_1 gpc6005 (
      {stage1_5[157]},
      {stage2_5[111]}
   );
   gpc1_1 gpc6006 (
      {stage1_5[158]},
      {stage2_5[112]}
   );
   gpc1_1 gpc6007 (
      {stage1_5[159]},
      {stage2_5[113]}
   );
   gpc1_1 gpc6008 (
      {stage1_5[160]},
      {stage2_5[114]}
   );
   gpc1_1 gpc6009 (
      {stage1_5[161]},
      {stage2_5[115]}
   );
   gpc1_1 gpc6010 (
      {stage1_5[162]},
      {stage2_5[116]}
   );
   gpc1_1 gpc6011 (
      {stage1_5[163]},
      {stage2_5[117]}
   );
   gpc1_1 gpc6012 (
      {stage1_5[164]},
      {stage2_5[118]}
   );
   gpc1_1 gpc6013 (
      {stage1_5[165]},
      {stage2_5[119]}
   );
   gpc1_1 gpc6014 (
      {stage1_5[166]},
      {stage2_5[120]}
   );
   gpc1_1 gpc6015 (
      {stage1_5[167]},
      {stage2_5[121]}
   );
   gpc1_1 gpc6016 (
      {stage1_5[168]},
      {stage2_5[122]}
   );
   gpc1_1 gpc6017 (
      {stage1_5[169]},
      {stage2_5[123]}
   );
   gpc1_1 gpc6018 (
      {stage1_5[170]},
      {stage2_5[124]}
   );
   gpc1_1 gpc6019 (
      {stage1_5[171]},
      {stage2_5[125]}
   );
   gpc1_1 gpc6020 (
      {stage1_5[172]},
      {stage2_5[126]}
   );
   gpc1_1 gpc6021 (
      {stage1_5[173]},
      {stage2_5[127]}
   );
   gpc1_1 gpc6022 (
      {stage1_5[174]},
      {stage2_5[128]}
   );
   gpc1_1 gpc6023 (
      {stage1_5[175]},
      {stage2_5[129]}
   );
   gpc1_1 gpc6024 (
      {stage1_5[176]},
      {stage2_5[130]}
   );
   gpc1_1 gpc6025 (
      {stage1_5[177]},
      {stage2_5[131]}
   );
   gpc1_1 gpc6026 (
      {stage1_5[178]},
      {stage2_5[132]}
   );
   gpc1_1 gpc6027 (
      {stage1_5[179]},
      {stage2_5[133]}
   );
   gpc1_1 gpc6028 (
      {stage1_5[180]},
      {stage2_5[134]}
   );
   gpc1_1 gpc6029 (
      {stage1_5[181]},
      {stage2_5[135]}
   );
   gpc1_1 gpc6030 (
      {stage1_5[182]},
      {stage2_5[136]}
   );
   gpc1_1 gpc6031 (
      {stage1_5[183]},
      {stage2_5[137]}
   );
   gpc1_1 gpc6032 (
      {stage1_5[184]},
      {stage2_5[138]}
   );
   gpc1_1 gpc6033 (
      {stage1_5[185]},
      {stage2_5[139]}
   );
   gpc1_1 gpc6034 (
      {stage1_5[186]},
      {stage2_5[140]}
   );
   gpc1_1 gpc6035 (
      {stage1_5[187]},
      {stage2_5[141]}
   );
   gpc1_1 gpc6036 (
      {stage1_5[188]},
      {stage2_5[142]}
   );
   gpc1_1 gpc6037 (
      {stage1_5[189]},
      {stage2_5[143]}
   );
   gpc1_1 gpc6038 (
      {stage1_5[190]},
      {stage2_5[144]}
   );
   gpc1_1 gpc6039 (
      {stage1_5[191]},
      {stage2_5[145]}
   );
   gpc1_1 gpc6040 (
      {stage1_5[192]},
      {stage2_5[146]}
   );
   gpc1_1 gpc6041 (
      {stage1_5[193]},
      {stage2_5[147]}
   );
   gpc1_1 gpc6042 (
      {stage1_5[194]},
      {stage2_5[148]}
   );
   gpc1_1 gpc6043 (
      {stage1_5[195]},
      {stage2_5[149]}
   );
   gpc1_1 gpc6044 (
      {stage1_5[196]},
      {stage2_5[150]}
   );
   gpc1_1 gpc6045 (
      {stage1_5[197]},
      {stage2_5[151]}
   );
   gpc1_1 gpc6046 (
      {stage1_6[175]},
      {stage2_6[53]}
   );
   gpc1_1 gpc6047 (
      {stage1_6[176]},
      {stage2_6[54]}
   );
   gpc1_1 gpc6048 (
      {stage1_6[177]},
      {stage2_6[55]}
   );
   gpc1_1 gpc6049 (
      {stage1_6[178]},
      {stage2_6[56]}
   );
   gpc1_1 gpc6050 (
      {stage1_6[179]},
      {stage2_6[57]}
   );
   gpc1_1 gpc6051 (
      {stage1_6[180]},
      {stage2_6[58]}
   );
   gpc1_1 gpc6052 (
      {stage1_6[181]},
      {stage2_6[59]}
   );
   gpc1_1 gpc6053 (
      {stage1_6[182]},
      {stage2_6[60]}
   );
   gpc1_1 gpc6054 (
      {stage1_6[183]},
      {stage2_6[61]}
   );
   gpc1_1 gpc6055 (
      {stage1_6[184]},
      {stage2_6[62]}
   );
   gpc1_1 gpc6056 (
      {stage1_6[185]},
      {stage2_6[63]}
   );
   gpc1_1 gpc6057 (
      {stage1_6[186]},
      {stage2_6[64]}
   );
   gpc1_1 gpc6058 (
      {stage1_6[187]},
      {stage2_6[65]}
   );
   gpc1_1 gpc6059 (
      {stage1_6[188]},
      {stage2_6[66]}
   );
   gpc1_1 gpc6060 (
      {stage1_6[189]},
      {stage2_6[67]}
   );
   gpc1_1 gpc6061 (
      {stage1_6[190]},
      {stage2_6[68]}
   );
   gpc1_1 gpc6062 (
      {stage1_6[191]},
      {stage2_6[69]}
   );
   gpc1_1 gpc6063 (
      {stage1_6[192]},
      {stage2_6[70]}
   );
   gpc1_1 gpc6064 (
      {stage1_6[193]},
      {stage2_6[71]}
   );
   gpc1_1 gpc6065 (
      {stage1_6[194]},
      {stage2_6[72]}
   );
   gpc1_1 gpc6066 (
      {stage1_6[195]},
      {stage2_6[73]}
   );
   gpc1_1 gpc6067 (
      {stage1_6[196]},
      {stage2_6[74]}
   );
   gpc1_1 gpc6068 (
      {stage1_6[197]},
      {stage2_6[75]}
   );
   gpc1_1 gpc6069 (
      {stage1_6[198]},
      {stage2_6[76]}
   );
   gpc1_1 gpc6070 (
      {stage1_6[199]},
      {stage2_6[77]}
   );
   gpc1_1 gpc6071 (
      {stage1_6[200]},
      {stage2_6[78]}
   );
   gpc1_1 gpc6072 (
      {stage1_6[201]},
      {stage2_6[79]}
   );
   gpc1_1 gpc6073 (
      {stage1_6[202]},
      {stage2_6[80]}
   );
   gpc1_1 gpc6074 (
      {stage1_6[203]},
      {stage2_6[81]}
   );
   gpc1_1 gpc6075 (
      {stage1_6[204]},
      {stage2_6[82]}
   );
   gpc1_1 gpc6076 (
      {stage1_6[205]},
      {stage2_6[83]}
   );
   gpc1_1 gpc6077 (
      {stage1_6[206]},
      {stage2_6[84]}
   );
   gpc1_1 gpc6078 (
      {stage1_6[207]},
      {stage2_6[85]}
   );
   gpc1_1 gpc6079 (
      {stage1_6[208]},
      {stage2_6[86]}
   );
   gpc1_1 gpc6080 (
      {stage1_6[209]},
      {stage2_6[87]}
   );
   gpc1_1 gpc6081 (
      {stage1_6[210]},
      {stage2_6[88]}
   );
   gpc1_1 gpc6082 (
      {stage1_6[211]},
      {stage2_6[89]}
   );
   gpc1_1 gpc6083 (
      {stage1_6[212]},
      {stage2_6[90]}
   );
   gpc1_1 gpc6084 (
      {stage1_6[213]},
      {stage2_6[91]}
   );
   gpc1_1 gpc6085 (
      {stage1_7[217]},
      {stage2_7[69]}
   );
   gpc1_1 gpc6086 (
      {stage1_7[218]},
      {stage2_7[70]}
   );
   gpc1_1 gpc6087 (
      {stage1_7[219]},
      {stage2_7[71]}
   );
   gpc1_1 gpc6088 (
      {stage1_7[220]},
      {stage2_7[72]}
   );
   gpc1_1 gpc6089 (
      {stage1_8[134]},
      {stage2_8[88]}
   );
   gpc1_1 gpc6090 (
      {stage1_8[135]},
      {stage2_8[89]}
   );
   gpc1_1 gpc6091 (
      {stage1_8[136]},
      {stage2_8[90]}
   );
   gpc1_1 gpc6092 (
      {stage1_8[137]},
      {stage2_8[91]}
   );
   gpc1_1 gpc6093 (
      {stage1_8[138]},
      {stage2_8[92]}
   );
   gpc1_1 gpc6094 (
      {stage1_8[139]},
      {stage2_8[93]}
   );
   gpc1_1 gpc6095 (
      {stage1_8[140]},
      {stage2_8[94]}
   );
   gpc1_1 gpc6096 (
      {stage1_8[141]},
      {stage2_8[95]}
   );
   gpc1_1 gpc6097 (
      {stage1_8[142]},
      {stage2_8[96]}
   );
   gpc1_1 gpc6098 (
      {stage1_8[143]},
      {stage2_8[97]}
   );
   gpc1_1 gpc6099 (
      {stage1_8[144]},
      {stage2_8[98]}
   );
   gpc1_1 gpc6100 (
      {stage1_8[145]},
      {stage2_8[99]}
   );
   gpc1_1 gpc6101 (
      {stage1_8[146]},
      {stage2_8[100]}
   );
   gpc1_1 gpc6102 (
      {stage1_8[147]},
      {stage2_8[101]}
   );
   gpc1_1 gpc6103 (
      {stage1_8[148]},
      {stage2_8[102]}
   );
   gpc1_1 gpc6104 (
      {stage1_8[149]},
      {stage2_8[103]}
   );
   gpc1_1 gpc6105 (
      {stage1_8[150]},
      {stage2_8[104]}
   );
   gpc1_1 gpc6106 (
      {stage1_8[151]},
      {stage2_8[105]}
   );
   gpc1_1 gpc6107 (
      {stage1_8[152]},
      {stage2_8[106]}
   );
   gpc1_1 gpc6108 (
      {stage1_8[153]},
      {stage2_8[107]}
   );
   gpc1_1 gpc6109 (
      {stage1_8[154]},
      {stage2_8[108]}
   );
   gpc1_1 gpc6110 (
      {stage1_8[155]},
      {stage2_8[109]}
   );
   gpc1_1 gpc6111 (
      {stage1_8[156]},
      {stage2_8[110]}
   );
   gpc1_1 gpc6112 (
      {stage1_8[157]},
      {stage2_8[111]}
   );
   gpc1_1 gpc6113 (
      {stage1_8[158]},
      {stage2_8[112]}
   );
   gpc1_1 gpc6114 (
      {stage1_8[159]},
      {stage2_8[113]}
   );
   gpc1_1 gpc6115 (
      {stage1_8[160]},
      {stage2_8[114]}
   );
   gpc1_1 gpc6116 (
      {stage1_8[161]},
      {stage2_8[115]}
   );
   gpc1_1 gpc6117 (
      {stage1_8[162]},
      {stage2_8[116]}
   );
   gpc1_1 gpc6118 (
      {stage1_8[163]},
      {stage2_8[117]}
   );
   gpc1_1 gpc6119 (
      {stage1_8[164]},
      {stage2_8[118]}
   );
   gpc1_1 gpc6120 (
      {stage1_8[165]},
      {stage2_8[119]}
   );
   gpc1_1 gpc6121 (
      {stage1_8[166]},
      {stage2_8[120]}
   );
   gpc1_1 gpc6122 (
      {stage1_8[167]},
      {stage2_8[121]}
   );
   gpc1_1 gpc6123 (
      {stage1_8[168]},
      {stage2_8[122]}
   );
   gpc1_1 gpc6124 (
      {stage1_8[169]},
      {stage2_8[123]}
   );
   gpc1_1 gpc6125 (
      {stage1_8[170]},
      {stage2_8[124]}
   );
   gpc1_1 gpc6126 (
      {stage1_8[171]},
      {stage2_8[125]}
   );
   gpc1_1 gpc6127 (
      {stage1_8[172]},
      {stage2_8[126]}
   );
   gpc1_1 gpc6128 (
      {stage1_8[173]},
      {stage2_8[127]}
   );
   gpc1_1 gpc6129 (
      {stage1_8[174]},
      {stage2_8[128]}
   );
   gpc1_1 gpc6130 (
      {stage1_8[175]},
      {stage2_8[129]}
   );
   gpc1_1 gpc6131 (
      {stage1_8[176]},
      {stage2_8[130]}
   );
   gpc1_1 gpc6132 (
      {stage1_8[177]},
      {stage2_8[131]}
   );
   gpc1_1 gpc6133 (
      {stage1_8[178]},
      {stage2_8[132]}
   );
   gpc1_1 gpc6134 (
      {stage1_8[179]},
      {stage2_8[133]}
   );
   gpc1_1 gpc6135 (
      {stage1_8[180]},
      {stage2_8[134]}
   );
   gpc1_1 gpc6136 (
      {stage1_8[181]},
      {stage2_8[135]}
   );
   gpc1_1 gpc6137 (
      {stage1_8[182]},
      {stage2_8[136]}
   );
   gpc1_1 gpc6138 (
      {stage1_8[183]},
      {stage2_8[137]}
   );
   gpc1_1 gpc6139 (
      {stage1_8[184]},
      {stage2_8[138]}
   );
   gpc1_1 gpc6140 (
      {stage1_8[185]},
      {stage2_8[139]}
   );
   gpc1_1 gpc6141 (
      {stage1_8[186]},
      {stage2_8[140]}
   );
   gpc1_1 gpc6142 (
      {stage1_8[187]},
      {stage2_8[141]}
   );
   gpc1_1 gpc6143 (
      {stage1_8[188]},
      {stage2_8[142]}
   );
   gpc1_1 gpc6144 (
      {stage1_8[189]},
      {stage2_8[143]}
   );
   gpc1_1 gpc6145 (
      {stage1_8[190]},
      {stage2_8[144]}
   );
   gpc1_1 gpc6146 (
      {stage1_8[191]},
      {stage2_8[145]}
   );
   gpc1_1 gpc6147 (
      {stage1_8[192]},
      {stage2_8[146]}
   );
   gpc1_1 gpc6148 (
      {stage1_8[193]},
      {stage2_8[147]}
   );
   gpc1_1 gpc6149 (
      {stage1_8[194]},
      {stage2_8[148]}
   );
   gpc1_1 gpc6150 (
      {stage1_8[195]},
      {stage2_8[149]}
   );
   gpc1_1 gpc6151 (
      {stage1_8[196]},
      {stage2_8[150]}
   );
   gpc1_1 gpc6152 (
      {stage1_8[197]},
      {stage2_8[151]}
   );
   gpc1_1 gpc6153 (
      {stage1_8[198]},
      {stage2_8[152]}
   );
   gpc1_1 gpc6154 (
      {stage1_8[199]},
      {stage2_8[153]}
   );
   gpc1_1 gpc6155 (
      {stage1_8[200]},
      {stage2_8[154]}
   );
   gpc1_1 gpc6156 (
      {stage1_8[201]},
      {stage2_8[155]}
   );
   gpc1_1 gpc6157 (
      {stage1_8[202]},
      {stage2_8[156]}
   );
   gpc1_1 gpc6158 (
      {stage1_8[203]},
      {stage2_8[157]}
   );
   gpc1_1 gpc6159 (
      {stage1_8[204]},
      {stage2_8[158]}
   );
   gpc1_1 gpc6160 (
      {stage1_8[205]},
      {stage2_8[159]}
   );
   gpc1_1 gpc6161 (
      {stage1_9[132]},
      {stage2_9[61]}
   );
   gpc1_1 gpc6162 (
      {stage1_9[133]},
      {stage2_9[62]}
   );
   gpc1_1 gpc6163 (
      {stage1_9[134]},
      {stage2_9[63]}
   );
   gpc1_1 gpc6164 (
      {stage1_9[135]},
      {stage2_9[64]}
   );
   gpc1_1 gpc6165 (
      {stage1_9[136]},
      {stage2_9[65]}
   );
   gpc1_1 gpc6166 (
      {stage1_9[137]},
      {stage2_9[66]}
   );
   gpc1_1 gpc6167 (
      {stage1_9[138]},
      {stage2_9[67]}
   );
   gpc1_1 gpc6168 (
      {stage1_9[139]},
      {stage2_9[68]}
   );
   gpc1_1 gpc6169 (
      {stage1_9[140]},
      {stage2_9[69]}
   );
   gpc1_1 gpc6170 (
      {stage1_9[141]},
      {stage2_9[70]}
   );
   gpc1_1 gpc6171 (
      {stage1_9[142]},
      {stage2_9[71]}
   );
   gpc1_1 gpc6172 (
      {stage1_9[143]},
      {stage2_9[72]}
   );
   gpc1_1 gpc6173 (
      {stage1_9[144]},
      {stage2_9[73]}
   );
   gpc1_1 gpc6174 (
      {stage1_9[145]},
      {stage2_9[74]}
   );
   gpc1_1 gpc6175 (
      {stage1_9[146]},
      {stage2_9[75]}
   );
   gpc1_1 gpc6176 (
      {stage1_9[147]},
      {stage2_9[76]}
   );
   gpc1_1 gpc6177 (
      {stage1_9[148]},
      {stage2_9[77]}
   );
   gpc1_1 gpc6178 (
      {stage1_9[149]},
      {stage2_9[78]}
   );
   gpc1_1 gpc6179 (
      {stage1_9[150]},
      {stage2_9[79]}
   );
   gpc1_1 gpc6180 (
      {stage1_9[151]},
      {stage2_9[80]}
   );
   gpc1_1 gpc6181 (
      {stage1_9[152]},
      {stage2_9[81]}
   );
   gpc1_1 gpc6182 (
      {stage1_9[153]},
      {stage2_9[82]}
   );
   gpc1_1 gpc6183 (
      {stage1_9[154]},
      {stage2_9[83]}
   );
   gpc1_1 gpc6184 (
      {stage1_9[155]},
      {stage2_9[84]}
   );
   gpc1_1 gpc6185 (
      {stage1_9[156]},
      {stage2_9[85]}
   );
   gpc1_1 gpc6186 (
      {stage1_9[157]},
      {stage2_9[86]}
   );
   gpc1_1 gpc6187 (
      {stage1_9[158]},
      {stage2_9[87]}
   );
   gpc1_1 gpc6188 (
      {stage1_9[159]},
      {stage2_9[88]}
   );
   gpc1_1 gpc6189 (
      {stage1_9[160]},
      {stage2_9[89]}
   );
   gpc1_1 gpc6190 (
      {stage1_9[161]},
      {stage2_9[90]}
   );
   gpc1_1 gpc6191 (
      {stage1_9[162]},
      {stage2_9[91]}
   );
   gpc1_1 gpc6192 (
      {stage1_9[163]},
      {stage2_9[92]}
   );
   gpc1_1 gpc6193 (
      {stage1_9[164]},
      {stage2_9[93]}
   );
   gpc1_1 gpc6194 (
      {stage1_9[165]},
      {stage2_9[94]}
   );
   gpc1_1 gpc6195 (
      {stage1_9[166]},
      {stage2_9[95]}
   );
   gpc1_1 gpc6196 (
      {stage1_9[167]},
      {stage2_9[96]}
   );
   gpc1_1 gpc6197 (
      {stage1_9[168]},
      {stage2_9[97]}
   );
   gpc1_1 gpc6198 (
      {stage1_9[169]},
      {stage2_9[98]}
   );
   gpc1_1 gpc6199 (
      {stage1_9[170]},
      {stage2_9[99]}
   );
   gpc1_1 gpc6200 (
      {stage1_9[171]},
      {stage2_9[100]}
   );
   gpc1_1 gpc6201 (
      {stage1_9[172]},
      {stage2_9[101]}
   );
   gpc1_1 gpc6202 (
      {stage1_9[173]},
      {stage2_9[102]}
   );
   gpc1_1 gpc6203 (
      {stage1_9[174]},
      {stage2_9[103]}
   );
   gpc1_1 gpc6204 (
      {stage1_9[175]},
      {stage2_9[104]}
   );
   gpc1_1 gpc6205 (
      {stage1_9[176]},
      {stage2_9[105]}
   );
   gpc1_1 gpc6206 (
      {stage1_9[177]},
      {stage2_9[106]}
   );
   gpc1_1 gpc6207 (
      {stage1_9[178]},
      {stage2_9[107]}
   );
   gpc1_1 gpc6208 (
      {stage1_9[179]},
      {stage2_9[108]}
   );
   gpc1_1 gpc6209 (
      {stage1_9[180]},
      {stage2_9[109]}
   );
   gpc1_1 gpc6210 (
      {stage1_9[181]},
      {stage2_9[110]}
   );
   gpc1_1 gpc6211 (
      {stage1_9[182]},
      {stage2_9[111]}
   );
   gpc1_1 gpc6212 (
      {stage1_9[183]},
      {stage2_9[112]}
   );
   gpc1_1 gpc6213 (
      {stage1_9[184]},
      {stage2_9[113]}
   );
   gpc1_1 gpc6214 (
      {stage1_9[185]},
      {stage2_9[114]}
   );
   gpc1_1 gpc6215 (
      {stage1_9[186]},
      {stage2_9[115]}
   );
   gpc1_1 gpc6216 (
      {stage1_9[187]},
      {stage2_9[116]}
   );
   gpc1_1 gpc6217 (
      {stage1_9[188]},
      {stage2_9[117]}
   );
   gpc1_1 gpc6218 (
      {stage1_9[189]},
      {stage2_9[118]}
   );
   gpc1_1 gpc6219 (
      {stage1_9[190]},
      {stage2_9[119]}
   );
   gpc1_1 gpc6220 (
      {stage1_9[191]},
      {stage2_9[120]}
   );
   gpc1_1 gpc6221 (
      {stage1_9[192]},
      {stage2_9[121]}
   );
   gpc1_1 gpc6222 (
      {stage1_9[193]},
      {stage2_9[122]}
   );
   gpc1_1 gpc6223 (
      {stage1_9[194]},
      {stage2_9[123]}
   );
   gpc1_1 gpc6224 (
      {stage1_9[195]},
      {stage2_9[124]}
   );
   gpc1_1 gpc6225 (
      {stage1_9[196]},
      {stage2_9[125]}
   );
   gpc1_1 gpc6226 (
      {stage1_9[197]},
      {stage2_9[126]}
   );
   gpc1_1 gpc6227 (
      {stage1_9[198]},
      {stage2_9[127]}
   );
   gpc1_1 gpc6228 (
      {stage1_9[199]},
      {stage2_9[128]}
   );
   gpc1_1 gpc6229 (
      {stage1_9[200]},
      {stage2_9[129]}
   );
   gpc1_1 gpc6230 (
      {stage1_9[201]},
      {stage2_9[130]}
   );
   gpc1_1 gpc6231 (
      {stage1_9[202]},
      {stage2_9[131]}
   );
   gpc1_1 gpc6232 (
      {stage1_9[203]},
      {stage2_9[132]}
   );
   gpc1_1 gpc6233 (
      {stage1_9[204]},
      {stage2_9[133]}
   );
   gpc1_1 gpc6234 (
      {stage1_9[205]},
      {stage2_9[134]}
   );
   gpc1_1 gpc6235 (
      {stage1_9[206]},
      {stage2_9[135]}
   );
   gpc1_1 gpc6236 (
      {stage1_9[207]},
      {stage2_9[136]}
   );
   gpc1_1 gpc6237 (
      {stage1_9[208]},
      {stage2_9[137]}
   );
   gpc1_1 gpc6238 (
      {stage1_9[209]},
      {stage2_9[138]}
   );
   gpc1_1 gpc6239 (
      {stage1_9[210]},
      {stage2_9[139]}
   );
   gpc1_1 gpc6240 (
      {stage1_9[211]},
      {stage2_9[140]}
   );
   gpc1_1 gpc6241 (
      {stage1_9[212]},
      {stage2_9[141]}
   );
   gpc1_1 gpc6242 (
      {stage1_9[213]},
      {stage2_9[142]}
   );
   gpc1_1 gpc6243 (
      {stage1_10[175]},
      {stage2_10[54]}
   );
   gpc1_1 gpc6244 (
      {stage1_10[176]},
      {stage2_10[55]}
   );
   gpc1_1 gpc6245 (
      {stage1_10[177]},
      {stage2_10[56]}
   );
   gpc1_1 gpc6246 (
      {stage1_10[178]},
      {stage2_10[57]}
   );
   gpc1_1 gpc6247 (
      {stage1_10[179]},
      {stage2_10[58]}
   );
   gpc1_1 gpc6248 (
      {stage1_10[180]},
      {stage2_10[59]}
   );
   gpc1_1 gpc6249 (
      {stage1_10[181]},
      {stage2_10[60]}
   );
   gpc1_1 gpc6250 (
      {stage1_10[182]},
      {stage2_10[61]}
   );
   gpc1_1 gpc6251 (
      {stage1_10[183]},
      {stage2_10[62]}
   );
   gpc1_1 gpc6252 (
      {stage1_10[184]},
      {stage2_10[63]}
   );
   gpc1_1 gpc6253 (
      {stage1_10[185]},
      {stage2_10[64]}
   );
   gpc1_1 gpc6254 (
      {stage1_10[186]},
      {stage2_10[65]}
   );
   gpc1_1 gpc6255 (
      {stage1_10[187]},
      {stage2_10[66]}
   );
   gpc1_1 gpc6256 (
      {stage1_10[188]},
      {stage2_10[67]}
   );
   gpc1_1 gpc6257 (
      {stage1_10[189]},
      {stage2_10[68]}
   );
   gpc1_1 gpc6258 (
      {stage1_10[190]},
      {stage2_10[69]}
   );
   gpc1_1 gpc6259 (
      {stage1_10[191]},
      {stage2_10[70]}
   );
   gpc1_1 gpc6260 (
      {stage1_10[192]},
      {stage2_10[71]}
   );
   gpc1_1 gpc6261 (
      {stage1_10[193]},
      {stage2_10[72]}
   );
   gpc1_1 gpc6262 (
      {stage1_10[194]},
      {stage2_10[73]}
   );
   gpc1_1 gpc6263 (
      {stage1_10[195]},
      {stage2_10[74]}
   );
   gpc1_1 gpc6264 (
      {stage1_10[196]},
      {stage2_10[75]}
   );
   gpc1_1 gpc6265 (
      {stage1_10[197]},
      {stage2_10[76]}
   );
   gpc1_1 gpc6266 (
      {stage1_10[198]},
      {stage2_10[77]}
   );
   gpc1_1 gpc6267 (
      {stage1_10[199]},
      {stage2_10[78]}
   );
   gpc1_1 gpc6268 (
      {stage1_10[200]},
      {stage2_10[79]}
   );
   gpc1_1 gpc6269 (
      {stage1_10[201]},
      {stage2_10[80]}
   );
   gpc1_1 gpc6270 (
      {stage1_10[202]},
      {stage2_10[81]}
   );
   gpc1_1 gpc6271 (
      {stage1_10[203]},
      {stage2_10[82]}
   );
   gpc1_1 gpc6272 (
      {stage1_10[204]},
      {stage2_10[83]}
   );
   gpc1_1 gpc6273 (
      {stage1_10[205]},
      {stage2_10[84]}
   );
   gpc1_1 gpc6274 (
      {stage1_10[206]},
      {stage2_10[85]}
   );
   gpc1_1 gpc6275 (
      {stage1_10[207]},
      {stage2_10[86]}
   );
   gpc1_1 gpc6276 (
      {stage1_10[208]},
      {stage2_10[87]}
   );
   gpc1_1 gpc6277 (
      {stage1_10[209]},
      {stage2_10[88]}
   );
   gpc1_1 gpc6278 (
      {stage1_10[210]},
      {stage2_10[89]}
   );
   gpc1_1 gpc6279 (
      {stage1_10[211]},
      {stage2_10[90]}
   );
   gpc1_1 gpc6280 (
      {stage1_10[212]},
      {stage2_10[91]}
   );
   gpc1_1 gpc6281 (
      {stage1_10[213]},
      {stage2_10[92]}
   );
   gpc1_1 gpc6282 (
      {stage1_10[214]},
      {stage2_10[93]}
   );
   gpc1_1 gpc6283 (
      {stage1_10[215]},
      {stage2_10[94]}
   );
   gpc1_1 gpc6284 (
      {stage1_10[216]},
      {stage2_10[95]}
   );
   gpc1_1 gpc6285 (
      {stage1_10[217]},
      {stage2_10[96]}
   );
   gpc1_1 gpc6286 (
      {stage1_10[218]},
      {stage2_10[97]}
   );
   gpc1_1 gpc6287 (
      {stage1_10[219]},
      {stage2_10[98]}
   );
   gpc1_1 gpc6288 (
      {stage1_10[220]},
      {stage2_10[99]}
   );
   gpc1_1 gpc6289 (
      {stage1_10[221]},
      {stage2_10[100]}
   );
   gpc1_1 gpc6290 (
      {stage1_10[222]},
      {stage2_10[101]}
   );
   gpc1_1 gpc6291 (
      {stage1_10[223]},
      {stage2_10[102]}
   );
   gpc1_1 gpc6292 (
      {stage1_10[224]},
      {stage2_10[103]}
   );
   gpc1_1 gpc6293 (
      {stage1_10[225]},
      {stage2_10[104]}
   );
   gpc1_1 gpc6294 (
      {stage1_10[226]},
      {stage2_10[105]}
   );
   gpc1_1 gpc6295 (
      {stage1_10[227]},
      {stage2_10[106]}
   );
   gpc1_1 gpc6296 (
      {stage1_10[228]},
      {stage2_10[107]}
   );
   gpc1_1 gpc6297 (
      {stage1_10[229]},
      {stage2_10[108]}
   );
   gpc1_1 gpc6298 (
      {stage1_10[230]},
      {stage2_10[109]}
   );
   gpc1_1 gpc6299 (
      {stage1_10[231]},
      {stage2_10[110]}
   );
   gpc1_1 gpc6300 (
      {stage1_10[232]},
      {stage2_10[111]}
   );
   gpc1_1 gpc6301 (
      {stage1_10[233]},
      {stage2_10[112]}
   );
   gpc1_1 gpc6302 (
      {stage1_10[234]},
      {stage2_10[113]}
   );
   gpc1_1 gpc6303 (
      {stage1_10[235]},
      {stage2_10[114]}
   );
   gpc1_1 gpc6304 (
      {stage1_10[236]},
      {stage2_10[115]}
   );
   gpc1_1 gpc6305 (
      {stage1_10[237]},
      {stage2_10[116]}
   );
   gpc1_1 gpc6306 (
      {stage1_10[238]},
      {stage2_10[117]}
   );
   gpc1_1 gpc6307 (
      {stage1_10[239]},
      {stage2_10[118]}
   );
   gpc1_1 gpc6308 (
      {stage1_10[240]},
      {stage2_10[119]}
   );
   gpc1_1 gpc6309 (
      {stage1_10[241]},
      {stage2_10[120]}
   );
   gpc1_1 gpc6310 (
      {stage1_10[242]},
      {stage2_10[121]}
   );
   gpc1_1 gpc6311 (
      {stage1_10[243]},
      {stage2_10[122]}
   );
   gpc1_1 gpc6312 (
      {stage1_10[244]},
      {stage2_10[123]}
   );
   gpc1_1 gpc6313 (
      {stage1_10[245]},
      {stage2_10[124]}
   );
   gpc1_1 gpc6314 (
      {stage1_10[246]},
      {stage2_10[125]}
   );
   gpc1_1 gpc6315 (
      {stage1_10[247]},
      {stage2_10[126]}
   );
   gpc1_1 gpc6316 (
      {stage1_10[248]},
      {stage2_10[127]}
   );
   gpc1_1 gpc6317 (
      {stage1_10[249]},
      {stage2_10[128]}
   );
   gpc1_1 gpc6318 (
      {stage1_10[250]},
      {stage2_10[129]}
   );
   gpc1_1 gpc6319 (
      {stage1_10[251]},
      {stage2_10[130]}
   );
   gpc1_1 gpc6320 (
      {stage1_10[252]},
      {stage2_10[131]}
   );
   gpc1_1 gpc6321 (
      {stage1_10[253]},
      {stage2_10[132]}
   );
   gpc1_1 gpc6322 (
      {stage1_10[254]},
      {stage2_10[133]}
   );
   gpc1_1 gpc6323 (
      {stage1_10[255]},
      {stage2_10[134]}
   );
   gpc1_1 gpc6324 (
      {stage1_10[256]},
      {stage2_10[135]}
   );
   gpc1_1 gpc6325 (
      {stage1_10[257]},
      {stage2_10[136]}
   );
   gpc1_1 gpc6326 (
      {stage1_10[258]},
      {stage2_10[137]}
   );
   gpc1_1 gpc6327 (
      {stage1_10[259]},
      {stage2_10[138]}
   );
   gpc1_1 gpc6328 (
      {stage1_10[260]},
      {stage2_10[139]}
   );
   gpc1_1 gpc6329 (
      {stage1_10[261]},
      {stage2_10[140]}
   );
   gpc1_1 gpc6330 (
      {stage1_10[262]},
      {stage2_10[141]}
   );
   gpc1_1 gpc6331 (
      {stage1_10[263]},
      {stage2_10[142]}
   );
   gpc1_1 gpc6332 (
      {stage1_10[264]},
      {stage2_10[143]}
   );
   gpc1_1 gpc6333 (
      {stage1_10[265]},
      {stage2_10[144]}
   );
   gpc1_1 gpc6334 (
      {stage1_10[266]},
      {stage2_10[145]}
   );
   gpc1_1 gpc6335 (
      {stage1_10[267]},
      {stage2_10[146]}
   );
   gpc1_1 gpc6336 (
      {stage1_10[268]},
      {stage2_10[147]}
   );
   gpc1_1 gpc6337 (
      {stage1_10[269]},
      {stage2_10[148]}
   );
   gpc1_1 gpc6338 (
      {stage1_10[270]},
      {stage2_10[149]}
   );
   gpc1_1 gpc6339 (
      {stage1_10[271]},
      {stage2_10[150]}
   );
   gpc1_1 gpc6340 (
      {stage1_10[272]},
      {stage2_10[151]}
   );
   gpc1_1 gpc6341 (
      {stage1_10[273]},
      {stage2_10[152]}
   );
   gpc1_1 gpc6342 (
      {stage1_10[274]},
      {stage2_10[153]}
   );
   gpc1_1 gpc6343 (
      {stage1_10[275]},
      {stage2_10[154]}
   );
   gpc1_1 gpc6344 (
      {stage1_10[276]},
      {stage2_10[155]}
   );
   gpc1_1 gpc6345 (
      {stage1_10[277]},
      {stage2_10[156]}
   );
   gpc1_1 gpc6346 (
      {stage1_10[278]},
      {stage2_10[157]}
   );
   gpc1_1 gpc6347 (
      {stage1_10[279]},
      {stage2_10[158]}
   );
   gpc1_1 gpc6348 (
      {stage1_10[280]},
      {stage2_10[159]}
   );
   gpc1_1 gpc6349 (
      {stage1_10[281]},
      {stage2_10[160]}
   );
   gpc1_1 gpc6350 (
      {stage1_10[282]},
      {stage2_10[161]}
   );
   gpc1_1 gpc6351 (
      {stage1_10[283]},
      {stage2_10[162]}
   );
   gpc1_1 gpc6352 (
      {stage1_10[284]},
      {stage2_10[163]}
   );
   gpc1_1 gpc6353 (
      {stage1_11[228]},
      {stage2_11[90]}
   );
   gpc1_1 gpc6354 (
      {stage1_11[229]},
      {stage2_11[91]}
   );
   gpc1_1 gpc6355 (
      {stage1_11[230]},
      {stage2_11[92]}
   );
   gpc1_1 gpc6356 (
      {stage1_11[231]},
      {stage2_11[93]}
   );
   gpc1_1 gpc6357 (
      {stage1_11[232]},
      {stage2_11[94]}
   );
   gpc1_1 gpc6358 (
      {stage1_11[233]},
      {stage2_11[95]}
   );
   gpc1_1 gpc6359 (
      {stage1_11[234]},
      {stage2_11[96]}
   );
   gpc1_1 gpc6360 (
      {stage1_11[235]},
      {stage2_11[97]}
   );
   gpc1_1 gpc6361 (
      {stage1_11[236]},
      {stage2_11[98]}
   );
   gpc1_1 gpc6362 (
      {stage1_11[237]},
      {stage2_11[99]}
   );
   gpc1_1 gpc6363 (
      {stage1_11[238]},
      {stage2_11[100]}
   );
   gpc1_1 gpc6364 (
      {stage1_11[239]},
      {stage2_11[101]}
   );
   gpc1_1 gpc6365 (
      {stage1_11[240]},
      {stage2_11[102]}
   );
   gpc1_1 gpc6366 (
      {stage1_11[241]},
      {stage2_11[103]}
   );
   gpc1_1 gpc6367 (
      {stage1_11[242]},
      {stage2_11[104]}
   );
   gpc1_1 gpc6368 (
      {stage1_11[243]},
      {stage2_11[105]}
   );
   gpc1_1 gpc6369 (
      {stage1_11[244]},
      {stage2_11[106]}
   );
   gpc1_1 gpc6370 (
      {stage1_11[245]},
      {stage2_11[107]}
   );
   gpc1_1 gpc6371 (
      {stage1_11[246]},
      {stage2_11[108]}
   );
   gpc1_1 gpc6372 (
      {stage1_11[247]},
      {stage2_11[109]}
   );
   gpc1_1 gpc6373 (
      {stage1_11[248]},
      {stage2_11[110]}
   );
   gpc1_1 gpc6374 (
      {stage1_11[249]},
      {stage2_11[111]}
   );
   gpc1_1 gpc6375 (
      {stage1_11[250]},
      {stage2_11[112]}
   );
   gpc1_1 gpc6376 (
      {stage1_11[251]},
      {stage2_11[113]}
   );
   gpc1_1 gpc6377 (
      {stage1_11[252]},
      {stage2_11[114]}
   );
   gpc1_1 gpc6378 (
      {stage1_11[253]},
      {stage2_11[115]}
   );
   gpc1_1 gpc6379 (
      {stage1_11[254]},
      {stage2_11[116]}
   );
   gpc1_1 gpc6380 (
      {stage1_11[255]},
      {stage2_11[117]}
   );
   gpc1_1 gpc6381 (
      {stage1_11[256]},
      {stage2_11[118]}
   );
   gpc1_1 gpc6382 (
      {stage1_11[257]},
      {stage2_11[119]}
   );
   gpc1_1 gpc6383 (
      {stage1_11[258]},
      {stage2_11[120]}
   );
   gpc1_1 gpc6384 (
      {stage1_11[259]},
      {stage2_11[121]}
   );
   gpc1_1 gpc6385 (
      {stage1_11[260]},
      {stage2_11[122]}
   );
   gpc1_1 gpc6386 (
      {stage1_11[261]},
      {stage2_11[123]}
   );
   gpc1_1 gpc6387 (
      {stage1_11[262]},
      {stage2_11[124]}
   );
   gpc1_1 gpc6388 (
      {stage1_11[263]},
      {stage2_11[125]}
   );
   gpc1_1 gpc6389 (
      {stage1_11[264]},
      {stage2_11[126]}
   );
   gpc1_1 gpc6390 (
      {stage1_11[265]},
      {stage2_11[127]}
   );
   gpc1_1 gpc6391 (
      {stage1_11[266]},
      {stage2_11[128]}
   );
   gpc1_1 gpc6392 (
      {stage1_11[267]},
      {stage2_11[129]}
   );
   gpc1_1 gpc6393 (
      {stage1_11[268]},
      {stage2_11[130]}
   );
   gpc1_1 gpc6394 (
      {stage1_11[269]},
      {stage2_11[131]}
   );
   gpc1_1 gpc6395 (
      {stage1_11[270]},
      {stage2_11[132]}
   );
   gpc1_1 gpc6396 (
      {stage1_11[271]},
      {stage2_11[133]}
   );
   gpc1_1 gpc6397 (
      {stage1_11[272]},
      {stage2_11[134]}
   );
   gpc1_1 gpc6398 (
      {stage1_11[273]},
      {stage2_11[135]}
   );
   gpc1_1 gpc6399 (
      {stage1_11[274]},
      {stage2_11[136]}
   );
   gpc1_1 gpc6400 (
      {stage1_11[275]},
      {stage2_11[137]}
   );
   gpc1_1 gpc6401 (
      {stage1_11[276]},
      {stage2_11[138]}
   );
   gpc1_1 gpc6402 (
      {stage1_12[163]},
      {stage2_12[81]}
   );
   gpc1_1 gpc6403 (
      {stage1_12[164]},
      {stage2_12[82]}
   );
   gpc1_1 gpc6404 (
      {stage1_12[165]},
      {stage2_12[83]}
   );
   gpc1_1 gpc6405 (
      {stage1_12[166]},
      {stage2_12[84]}
   );
   gpc1_1 gpc6406 (
      {stage1_12[167]},
      {stage2_12[85]}
   );
   gpc1_1 gpc6407 (
      {stage1_12[168]},
      {stage2_12[86]}
   );
   gpc1_1 gpc6408 (
      {stage1_12[169]},
      {stage2_12[87]}
   );
   gpc1_1 gpc6409 (
      {stage1_12[170]},
      {stage2_12[88]}
   );
   gpc1_1 gpc6410 (
      {stage1_12[171]},
      {stage2_12[89]}
   );
   gpc1_1 gpc6411 (
      {stage1_12[172]},
      {stage2_12[90]}
   );
   gpc1_1 gpc6412 (
      {stage1_12[173]},
      {stage2_12[91]}
   );
   gpc1_1 gpc6413 (
      {stage1_12[174]},
      {stage2_12[92]}
   );
   gpc1_1 gpc6414 (
      {stage1_12[175]},
      {stage2_12[93]}
   );
   gpc1_1 gpc6415 (
      {stage1_12[176]},
      {stage2_12[94]}
   );
   gpc1_1 gpc6416 (
      {stage1_12[177]},
      {stage2_12[95]}
   );
   gpc1_1 gpc6417 (
      {stage1_12[178]},
      {stage2_12[96]}
   );
   gpc1_1 gpc6418 (
      {stage1_12[179]},
      {stage2_12[97]}
   );
   gpc1_1 gpc6419 (
      {stage1_12[180]},
      {stage2_12[98]}
   );
   gpc1_1 gpc6420 (
      {stage1_12[181]},
      {stage2_12[99]}
   );
   gpc1_1 gpc6421 (
      {stage1_12[182]},
      {stage2_12[100]}
   );
   gpc1_1 gpc6422 (
      {stage1_12[183]},
      {stage2_12[101]}
   );
   gpc1_1 gpc6423 (
      {stage1_12[184]},
      {stage2_12[102]}
   );
   gpc1_1 gpc6424 (
      {stage1_12[185]},
      {stage2_12[103]}
   );
   gpc1_1 gpc6425 (
      {stage1_12[186]},
      {stage2_12[104]}
   );
   gpc1_1 gpc6426 (
      {stage1_12[187]},
      {stage2_12[105]}
   );
   gpc1_1 gpc6427 (
      {stage1_12[188]},
      {stage2_12[106]}
   );
   gpc1_1 gpc6428 (
      {stage1_14[217]},
      {stage2_14[106]}
   );
   gpc1_1 gpc6429 (
      {stage1_14[218]},
      {stage2_14[107]}
   );
   gpc1_1 gpc6430 (
      {stage1_15[123]},
      {stage2_15[93]}
   );
   gpc1_1 gpc6431 (
      {stage1_15[124]},
      {stage2_15[94]}
   );
   gpc1_1 gpc6432 (
      {stage1_15[125]},
      {stage2_15[95]}
   );
   gpc1_1 gpc6433 (
      {stage1_15[126]},
      {stage2_15[96]}
   );
   gpc1_1 gpc6434 (
      {stage1_15[127]},
      {stage2_15[97]}
   );
   gpc1_1 gpc6435 (
      {stage1_15[128]},
      {stage2_15[98]}
   );
   gpc1_1 gpc6436 (
      {stage1_15[129]},
      {stage2_15[99]}
   );
   gpc1_1 gpc6437 (
      {stage1_15[130]},
      {stage2_15[100]}
   );
   gpc1_1 gpc6438 (
      {stage1_15[131]},
      {stage2_15[101]}
   );
   gpc1_1 gpc6439 (
      {stage1_15[132]},
      {stage2_15[102]}
   );
   gpc1_1 gpc6440 (
      {stage1_15[133]},
      {stage2_15[103]}
   );
   gpc1_1 gpc6441 (
      {stage1_15[134]},
      {stage2_15[104]}
   );
   gpc1_1 gpc6442 (
      {stage1_15[135]},
      {stage2_15[105]}
   );
   gpc1_1 gpc6443 (
      {stage1_15[136]},
      {stage2_15[106]}
   );
   gpc1_1 gpc6444 (
      {stage1_15[137]},
      {stage2_15[107]}
   );
   gpc1_1 gpc6445 (
      {stage1_15[138]},
      {stage2_15[108]}
   );
   gpc1_1 gpc6446 (
      {stage1_15[139]},
      {stage2_15[109]}
   );
   gpc1_1 gpc6447 (
      {stage1_15[140]},
      {stage2_15[110]}
   );
   gpc1_1 gpc6448 (
      {stage1_15[141]},
      {stage2_15[111]}
   );
   gpc1_1 gpc6449 (
      {stage1_15[142]},
      {stage2_15[112]}
   );
   gpc1_1 gpc6450 (
      {stage1_15[143]},
      {stage2_15[113]}
   );
   gpc1_1 gpc6451 (
      {stage1_15[144]},
      {stage2_15[114]}
   );
   gpc1_1 gpc6452 (
      {stage1_15[145]},
      {stage2_15[115]}
   );
   gpc1_1 gpc6453 (
      {stage1_15[146]},
      {stage2_15[116]}
   );
   gpc1_1 gpc6454 (
      {stage1_15[147]},
      {stage2_15[117]}
   );
   gpc1_1 gpc6455 (
      {stage1_15[148]},
      {stage2_15[118]}
   );
   gpc1_1 gpc6456 (
      {stage1_15[149]},
      {stage2_15[119]}
   );
   gpc1_1 gpc6457 (
      {stage1_15[150]},
      {stage2_15[120]}
   );
   gpc1_1 gpc6458 (
      {stage1_15[151]},
      {stage2_15[121]}
   );
   gpc1_1 gpc6459 (
      {stage1_15[152]},
      {stage2_15[122]}
   );
   gpc1_1 gpc6460 (
      {stage1_15[153]},
      {stage2_15[123]}
   );
   gpc1_1 gpc6461 (
      {stage1_15[154]},
      {stage2_15[124]}
   );
   gpc1_1 gpc6462 (
      {stage1_15[155]},
      {stage2_15[125]}
   );
   gpc1_1 gpc6463 (
      {stage1_15[156]},
      {stage2_15[126]}
   );
   gpc1_1 gpc6464 (
      {stage1_15[157]},
      {stage2_15[127]}
   );
   gpc1_1 gpc6465 (
      {stage1_15[158]},
      {stage2_15[128]}
   );
   gpc1_1 gpc6466 (
      {stage1_15[159]},
      {stage2_15[129]}
   );
   gpc1_1 gpc6467 (
      {stage1_15[160]},
      {stage2_15[130]}
   );
   gpc1_1 gpc6468 (
      {stage1_15[161]},
      {stage2_15[131]}
   );
   gpc1_1 gpc6469 (
      {stage1_15[162]},
      {stage2_15[132]}
   );
   gpc1_1 gpc6470 (
      {stage1_15[163]},
      {stage2_15[133]}
   );
   gpc1_1 gpc6471 (
      {stage1_15[164]},
      {stage2_15[134]}
   );
   gpc1_1 gpc6472 (
      {stage1_15[165]},
      {stage2_15[135]}
   );
   gpc1_1 gpc6473 (
      {stage1_15[166]},
      {stage2_15[136]}
   );
   gpc1_1 gpc6474 (
      {stage1_15[167]},
      {stage2_15[137]}
   );
   gpc1_1 gpc6475 (
      {stage1_15[168]},
      {stage2_15[138]}
   );
   gpc1_1 gpc6476 (
      {stage1_15[169]},
      {stage2_15[139]}
   );
   gpc1_1 gpc6477 (
      {stage1_15[170]},
      {stage2_15[140]}
   );
   gpc1_1 gpc6478 (
      {stage1_16[198]},
      {stage2_16[59]}
   );
   gpc1_1 gpc6479 (
      {stage1_16[199]},
      {stage2_16[60]}
   );
   gpc1_1 gpc6480 (
      {stage1_16[200]},
      {stage2_16[61]}
   );
   gpc1_1 gpc6481 (
      {stage1_16[201]},
      {stage2_16[62]}
   );
   gpc1_1 gpc6482 (
      {stage1_16[202]},
      {stage2_16[63]}
   );
   gpc1_1 gpc6483 (
      {stage1_16[203]},
      {stage2_16[64]}
   );
   gpc1_1 gpc6484 (
      {stage1_16[204]},
      {stage2_16[65]}
   );
   gpc1_1 gpc6485 (
      {stage1_16[205]},
      {stage2_16[66]}
   );
   gpc1_1 gpc6486 (
      {stage1_16[206]},
      {stage2_16[67]}
   );
   gpc1_1 gpc6487 (
      {stage1_16[207]},
      {stage2_16[68]}
   );
   gpc1_1 gpc6488 (
      {stage1_16[208]},
      {stage2_16[69]}
   );
   gpc1_1 gpc6489 (
      {stage1_16[209]},
      {stage2_16[70]}
   );
   gpc1_1 gpc6490 (
      {stage1_16[210]},
      {stage2_16[71]}
   );
   gpc1_1 gpc6491 (
      {stage1_16[211]},
      {stage2_16[72]}
   );
   gpc1_1 gpc6492 (
      {stage1_16[212]},
      {stage2_16[73]}
   );
   gpc1_1 gpc6493 (
      {stage1_16[213]},
      {stage2_16[74]}
   );
   gpc1_1 gpc6494 (
      {stage1_16[214]},
      {stage2_16[75]}
   );
   gpc1_1 gpc6495 (
      {stage1_16[215]},
      {stage2_16[76]}
   );
   gpc1_1 gpc6496 (
      {stage1_16[216]},
      {stage2_16[77]}
   );
   gpc1_1 gpc6497 (
      {stage1_16[217]},
      {stage2_16[78]}
   );
   gpc1_1 gpc6498 (
      {stage1_16[218]},
      {stage2_16[79]}
   );
   gpc1_1 gpc6499 (
      {stage1_16[219]},
      {stage2_16[80]}
   );
   gpc1_1 gpc6500 (
      {stage1_16[220]},
      {stage2_16[81]}
   );
   gpc1_1 gpc6501 (
      {stage1_16[221]},
      {stage2_16[82]}
   );
   gpc1_1 gpc6502 (
      {stage1_17[228]},
      {stage2_17[86]}
   );
   gpc1_1 gpc6503 (
      {stage1_18[191]},
      {stage2_18[101]}
   );
   gpc1_1 gpc6504 (
      {stage1_18[192]},
      {stage2_18[102]}
   );
   gpc1_1 gpc6505 (
      {stage1_18[193]},
      {stage2_18[103]}
   );
   gpc1_1 gpc6506 (
      {stage1_18[194]},
      {stage2_18[104]}
   );
   gpc1_1 gpc6507 (
      {stage1_18[195]},
      {stage2_18[105]}
   );
   gpc1_1 gpc6508 (
      {stage1_18[196]},
      {stage2_18[106]}
   );
   gpc1_1 gpc6509 (
      {stage1_18[197]},
      {stage2_18[107]}
   );
   gpc1_1 gpc6510 (
      {stage1_18[198]},
      {stage2_18[108]}
   );
   gpc1_1 gpc6511 (
      {stage1_18[199]},
      {stage2_18[109]}
   );
   gpc1_1 gpc6512 (
      {stage1_18[200]},
      {stage2_18[110]}
   );
   gpc1_1 gpc6513 (
      {stage1_18[201]},
      {stage2_18[111]}
   );
   gpc1_1 gpc6514 (
      {stage1_18[202]},
      {stage2_18[112]}
   );
   gpc1_1 gpc6515 (
      {stage1_18[203]},
      {stage2_18[113]}
   );
   gpc1_1 gpc6516 (
      {stage1_18[204]},
      {stage2_18[114]}
   );
   gpc1_1 gpc6517 (
      {stage1_18[205]},
      {stage2_18[115]}
   );
   gpc1_1 gpc6518 (
      {stage1_18[206]},
      {stage2_18[116]}
   );
   gpc1_1 gpc6519 (
      {stage1_18[207]},
      {stage2_18[117]}
   );
   gpc1_1 gpc6520 (
      {stage1_18[208]},
      {stage2_18[118]}
   );
   gpc1_1 gpc6521 (
      {stage1_19[234]},
      {stage2_19[71]}
   );
   gpc1_1 gpc6522 (
      {stage1_19[235]},
      {stage2_19[72]}
   );
   gpc1_1 gpc6523 (
      {stage1_19[236]},
      {stage2_19[73]}
   );
   gpc1_1 gpc6524 (
      {stage1_19[237]},
      {stage2_19[74]}
   );
   gpc1_1 gpc6525 (
      {stage1_19[238]},
      {stage2_19[75]}
   );
   gpc1_1 gpc6526 (
      {stage1_19[239]},
      {stage2_19[76]}
   );
   gpc1_1 gpc6527 (
      {stage1_19[240]},
      {stage2_19[77]}
   );
   gpc1_1 gpc6528 (
      {stage1_19[241]},
      {stage2_19[78]}
   );
   gpc1_1 gpc6529 (
      {stage1_19[242]},
      {stage2_19[79]}
   );
   gpc1_1 gpc6530 (
      {stage1_19[243]},
      {stage2_19[80]}
   );
   gpc1_1 gpc6531 (
      {stage1_19[244]},
      {stage2_19[81]}
   );
   gpc1_1 gpc6532 (
      {stage1_19[245]},
      {stage2_19[82]}
   );
   gpc1_1 gpc6533 (
      {stage1_19[246]},
      {stage2_19[83]}
   );
   gpc1_1 gpc6534 (
      {stage1_19[247]},
      {stage2_19[84]}
   );
   gpc1_1 gpc6535 (
      {stage1_19[248]},
      {stage2_19[85]}
   );
   gpc1_1 gpc6536 (
      {stage1_19[249]},
      {stage2_19[86]}
   );
   gpc1_1 gpc6537 (
      {stage1_19[250]},
      {stage2_19[87]}
   );
   gpc1_1 gpc6538 (
      {stage1_19[251]},
      {stage2_19[88]}
   );
   gpc1_1 gpc6539 (
      {stage1_19[252]},
      {stage2_19[89]}
   );
   gpc1_1 gpc6540 (
      {stage1_19[253]},
      {stage2_19[90]}
   );
   gpc1_1 gpc6541 (
      {stage1_19[254]},
      {stage2_19[91]}
   );
   gpc1_1 gpc6542 (
      {stage1_19[255]},
      {stage2_19[92]}
   );
   gpc1_1 gpc6543 (
      {stage1_19[256]},
      {stage2_19[93]}
   );
   gpc1_1 gpc6544 (
      {stage1_19[257]},
      {stage2_19[94]}
   );
   gpc1_1 gpc6545 (
      {stage1_19[258]},
      {stage2_19[95]}
   );
   gpc1_1 gpc6546 (
      {stage1_19[259]},
      {stage2_19[96]}
   );
   gpc1_1 gpc6547 (
      {stage1_19[260]},
      {stage2_19[97]}
   );
   gpc1_1 gpc6548 (
      {stage1_19[261]},
      {stage2_19[98]}
   );
   gpc1_1 gpc6549 (
      {stage1_19[262]},
      {stage2_19[99]}
   );
   gpc1_1 gpc6550 (
      {stage1_19[263]},
      {stage2_19[100]}
   );
   gpc1_1 gpc6551 (
      {stage1_19[264]},
      {stage2_19[101]}
   );
   gpc1_1 gpc6552 (
      {stage1_19[265]},
      {stage2_19[102]}
   );
   gpc1_1 gpc6553 (
      {stage1_19[266]},
      {stage2_19[103]}
   );
   gpc1_1 gpc6554 (
      {stage1_19[267]},
      {stage2_19[104]}
   );
   gpc1_1 gpc6555 (
      {stage1_19[268]},
      {stage2_19[105]}
   );
   gpc1_1 gpc6556 (
      {stage1_19[269]},
      {stage2_19[106]}
   );
   gpc1_1 gpc6557 (
      {stage1_19[270]},
      {stage2_19[107]}
   );
   gpc1_1 gpc6558 (
      {stage1_19[271]},
      {stage2_19[108]}
   );
   gpc1_1 gpc6559 (
      {stage1_19[272]},
      {stage2_19[109]}
   );
   gpc1_1 gpc6560 (
      {stage1_19[273]},
      {stage2_19[110]}
   );
   gpc1_1 gpc6561 (
      {stage1_19[274]},
      {stage2_19[111]}
   );
   gpc1_1 gpc6562 (
      {stage1_19[275]},
      {stage2_19[112]}
   );
   gpc1_1 gpc6563 (
      {stage1_20[262]},
      {stage2_20[87]}
   );
   gpc1_1 gpc6564 (
      {stage1_20[263]},
      {stage2_20[88]}
   );
   gpc1_1 gpc6565 (
      {stage1_20[264]},
      {stage2_20[89]}
   );
   gpc1_1 gpc6566 (
      {stage1_20[265]},
      {stage2_20[90]}
   );
   gpc1_1 gpc6567 (
      {stage1_20[266]},
      {stage2_20[91]}
   );
   gpc1_1 gpc6568 (
      {stage1_20[267]},
      {stage2_20[92]}
   );
   gpc1_1 gpc6569 (
      {stage1_21[174]},
      {stage2_21[112]}
   );
   gpc1_1 gpc6570 (
      {stage1_21[175]},
      {stage2_21[113]}
   );
   gpc1_1 gpc6571 (
      {stage1_21[176]},
      {stage2_21[114]}
   );
   gpc1_1 gpc6572 (
      {stage1_21[177]},
      {stage2_21[115]}
   );
   gpc1_1 gpc6573 (
      {stage1_21[178]},
      {stage2_21[116]}
   );
   gpc1_1 gpc6574 (
      {stage1_21[179]},
      {stage2_21[117]}
   );
   gpc1_1 gpc6575 (
      {stage1_21[180]},
      {stage2_21[118]}
   );
   gpc1_1 gpc6576 (
      {stage1_21[181]},
      {stage2_21[119]}
   );
   gpc1_1 gpc6577 (
      {stage1_21[182]},
      {stage2_21[120]}
   );
   gpc1_1 gpc6578 (
      {stage1_21[183]},
      {stage2_21[121]}
   );
   gpc1_1 gpc6579 (
      {stage1_21[184]},
      {stage2_21[122]}
   );
   gpc1_1 gpc6580 (
      {stage1_21[185]},
      {stage2_21[123]}
   );
   gpc1_1 gpc6581 (
      {stage1_21[186]},
      {stage2_21[124]}
   );
   gpc1_1 gpc6582 (
      {stage1_21[187]},
      {stage2_21[125]}
   );
   gpc1_1 gpc6583 (
      {stage1_21[188]},
      {stage2_21[126]}
   );
   gpc1_1 gpc6584 (
      {stage1_21[189]},
      {stage2_21[127]}
   );
   gpc1_1 gpc6585 (
      {stage1_22[145]},
      {stage2_22[82]}
   );
   gpc1_1 gpc6586 (
      {stage1_22[146]},
      {stage2_22[83]}
   );
   gpc1_1 gpc6587 (
      {stage1_22[147]},
      {stage2_22[84]}
   );
   gpc1_1 gpc6588 (
      {stage1_22[148]},
      {stage2_22[85]}
   );
   gpc1_1 gpc6589 (
      {stage1_22[149]},
      {stage2_22[86]}
   );
   gpc1_1 gpc6590 (
      {stage1_22[150]},
      {stage2_22[87]}
   );
   gpc1_1 gpc6591 (
      {stage1_22[151]},
      {stage2_22[88]}
   );
   gpc1_1 gpc6592 (
      {stage1_22[152]},
      {stage2_22[89]}
   );
   gpc1_1 gpc6593 (
      {stage1_22[153]},
      {stage2_22[90]}
   );
   gpc1_1 gpc6594 (
      {stage1_22[154]},
      {stage2_22[91]}
   );
   gpc1_1 gpc6595 (
      {stage1_22[155]},
      {stage2_22[92]}
   );
   gpc1_1 gpc6596 (
      {stage1_22[156]},
      {stage2_22[93]}
   );
   gpc1_1 gpc6597 (
      {stage1_22[157]},
      {stage2_22[94]}
   );
   gpc1_1 gpc6598 (
      {stage1_22[158]},
      {stage2_22[95]}
   );
   gpc1_1 gpc6599 (
      {stage1_22[159]},
      {stage2_22[96]}
   );
   gpc1_1 gpc6600 (
      {stage1_22[160]},
      {stage2_22[97]}
   );
   gpc1_1 gpc6601 (
      {stage1_22[161]},
      {stage2_22[98]}
   );
   gpc1_1 gpc6602 (
      {stage1_22[162]},
      {stage2_22[99]}
   );
   gpc1_1 gpc6603 (
      {stage1_22[163]},
      {stage2_22[100]}
   );
   gpc1_1 gpc6604 (
      {stage1_22[164]},
      {stage2_22[101]}
   );
   gpc1_1 gpc6605 (
      {stage1_22[165]},
      {stage2_22[102]}
   );
   gpc1_1 gpc6606 (
      {stage1_22[166]},
      {stage2_22[103]}
   );
   gpc1_1 gpc6607 (
      {stage1_22[167]},
      {stage2_22[104]}
   );
   gpc1_1 gpc6608 (
      {stage1_22[168]},
      {stage2_22[105]}
   );
   gpc1_1 gpc6609 (
      {stage1_22[169]},
      {stage2_22[106]}
   );
   gpc1_1 gpc6610 (
      {stage1_22[170]},
      {stage2_22[107]}
   );
   gpc1_1 gpc6611 (
      {stage1_24[210]},
      {stage2_24[98]}
   );
   gpc1_1 gpc6612 (
      {stage1_24[211]},
      {stage2_24[99]}
   );
   gpc1_1 gpc6613 (
      {stage1_24[212]},
      {stage2_24[100]}
   );
   gpc1_1 gpc6614 (
      {stage1_24[213]},
      {stage2_24[101]}
   );
   gpc1_1 gpc6615 (
      {stage1_25[175]},
      {stage2_25[87]}
   );
   gpc1_1 gpc6616 (
      {stage1_25[176]},
      {stage2_25[88]}
   );
   gpc1_1 gpc6617 (
      {stage1_25[177]},
      {stage2_25[89]}
   );
   gpc1_1 gpc6618 (
      {stage1_25[178]},
      {stage2_25[90]}
   );
   gpc1_1 gpc6619 (
      {stage1_25[179]},
      {stage2_25[91]}
   );
   gpc1_1 gpc6620 (
      {stage1_25[180]},
      {stage2_25[92]}
   );
   gpc1_1 gpc6621 (
      {stage1_25[181]},
      {stage2_25[93]}
   );
   gpc1_1 gpc6622 (
      {stage1_25[182]},
      {stage2_25[94]}
   );
   gpc1_1 gpc6623 (
      {stage1_25[183]},
      {stage2_25[95]}
   );
   gpc1_1 gpc6624 (
      {stage1_26[248]},
      {stage2_26[82]}
   );
   gpc1_1 gpc6625 (
      {stage1_26[249]},
      {stage2_26[83]}
   );
   gpc1_1 gpc6626 (
      {stage1_26[250]},
      {stage2_26[84]}
   );
   gpc1_1 gpc6627 (
      {stage1_29[216]},
      {stage2_29[74]}
   );
   gpc1_1 gpc6628 (
      {stage1_29[217]},
      {stage2_29[75]}
   );
   gpc1_1 gpc6629 (
      {stage1_29[218]},
      {stage2_29[76]}
   );
   gpc1_1 gpc6630 (
      {stage1_29[219]},
      {stage2_29[77]}
   );
   gpc1_1 gpc6631 (
      {stage1_29[220]},
      {stage2_29[78]}
   );
   gpc1_1 gpc6632 (
      {stage1_29[221]},
      {stage2_29[79]}
   );
   gpc1_1 gpc6633 (
      {stage1_29[222]},
      {stage2_29[80]}
   );
   gpc1_1 gpc6634 (
      {stage1_29[223]},
      {stage2_29[81]}
   );
   gpc1_1 gpc6635 (
      {stage1_29[224]},
      {stage2_29[82]}
   );
   gpc1_1 gpc6636 (
      {stage1_29[225]},
      {stage2_29[83]}
   );
   gpc1_1 gpc6637 (
      {stage1_29[226]},
      {stage2_29[84]}
   );
   gpc1_1 gpc6638 (
      {stage1_29[227]},
      {stage2_29[85]}
   );
   gpc1_1 gpc6639 (
      {stage1_29[228]},
      {stage2_29[86]}
   );
   gpc1_1 gpc6640 (
      {stage1_30[160]},
      {stage2_30[85]}
   );
   gpc1_1 gpc6641 (
      {stage1_30[161]},
      {stage2_30[86]}
   );
   gpc1_1 gpc6642 (
      {stage1_30[162]},
      {stage2_30[87]}
   );
   gpc1_1 gpc6643 (
      {stage1_30[163]},
      {stage2_30[88]}
   );
   gpc1_1 gpc6644 (
      {stage1_30[164]},
      {stage2_30[89]}
   );
   gpc1_1 gpc6645 (
      {stage1_30[165]},
      {stage2_30[90]}
   );
   gpc1_1 gpc6646 (
      {stage1_30[166]},
      {stage2_30[91]}
   );
   gpc1_1 gpc6647 (
      {stage1_30[167]},
      {stage2_30[92]}
   );
   gpc1_1 gpc6648 (
      {stage1_30[168]},
      {stage2_30[93]}
   );
   gpc1_1 gpc6649 (
      {stage1_30[169]},
      {stage2_30[94]}
   );
   gpc1_1 gpc6650 (
      {stage1_30[170]},
      {stage2_30[95]}
   );
   gpc1_1 gpc6651 (
      {stage1_30[171]},
      {stage2_30[96]}
   );
   gpc1_1 gpc6652 (
      {stage1_30[172]},
      {stage2_30[97]}
   );
   gpc1_1 gpc6653 (
      {stage1_30[173]},
      {stage2_30[98]}
   );
   gpc1_1 gpc6654 (
      {stage1_30[174]},
      {stage2_30[99]}
   );
   gpc1_1 gpc6655 (
      {stage1_30[175]},
      {stage2_30[100]}
   );
   gpc1_1 gpc6656 (
      {stage1_30[176]},
      {stage2_30[101]}
   );
   gpc1_1 gpc6657 (
      {stage1_30[177]},
      {stage2_30[102]}
   );
   gpc1_1 gpc6658 (
      {stage1_30[178]},
      {stage2_30[103]}
   );
   gpc1_1 gpc6659 (
      {stage1_30[179]},
      {stage2_30[104]}
   );
   gpc1_1 gpc6660 (
      {stage1_30[180]},
      {stage2_30[105]}
   );
   gpc1_1 gpc6661 (
      {stage1_30[181]},
      {stage2_30[106]}
   );
   gpc1_1 gpc6662 (
      {stage1_30[182]},
      {stage2_30[107]}
   );
   gpc1_1 gpc6663 (
      {stage1_30[183]},
      {stage2_30[108]}
   );
   gpc1_1 gpc6664 (
      {stage1_30[184]},
      {stage2_30[109]}
   );
   gpc1_1 gpc6665 (
      {stage1_30[185]},
      {stage2_30[110]}
   );
   gpc1_1 gpc6666 (
      {stage1_30[186]},
      {stage2_30[111]}
   );
   gpc1_1 gpc6667 (
      {stage1_30[187]},
      {stage2_30[112]}
   );
   gpc1_1 gpc6668 (
      {stage1_30[188]},
      {stage2_30[113]}
   );
   gpc1_1 gpc6669 (
      {stage1_30[189]},
      {stage2_30[114]}
   );
   gpc1_1 gpc6670 (
      {stage1_30[190]},
      {stage2_30[115]}
   );
   gpc1_1 gpc6671 (
      {stage1_30[191]},
      {stage2_30[116]}
   );
   gpc1_1 gpc6672 (
      {stage1_32[189]},
      {stage2_32[78]}
   );
   gpc1_1 gpc6673 (
      {stage1_32[190]},
      {stage2_32[79]}
   );
   gpc1_1 gpc6674 (
      {stage1_32[191]},
      {stage2_32[80]}
   );
   gpc1_1 gpc6675 (
      {stage1_32[192]},
      {stage2_32[81]}
   );
   gpc1_1 gpc6676 (
      {stage1_32[193]},
      {stage2_32[82]}
   );
   gpc1_1 gpc6677 (
      {stage1_32[194]},
      {stage2_32[83]}
   );
   gpc1_1 gpc6678 (
      {stage1_32[195]},
      {stage2_32[84]}
   );
   gpc1_1 gpc6679 (
      {stage1_32[196]},
      {stage2_32[85]}
   );
   gpc1_1 gpc6680 (
      {stage1_32[197]},
      {stage2_32[86]}
   );
   gpc1_1 gpc6681 (
      {stage1_32[198]},
      {stage2_32[87]}
   );
   gpc1_1 gpc6682 (
      {stage1_32[199]},
      {stage2_32[88]}
   );
   gpc1_1 gpc6683 (
      {stage1_32[200]},
      {stage2_32[89]}
   );
   gpc1_1 gpc6684 (
      {stage1_32[201]},
      {stage2_32[90]}
   );
   gpc1_1 gpc6685 (
      {stage1_32[202]},
      {stage2_32[91]}
   );
   gpc1_1 gpc6686 (
      {stage1_32[203]},
      {stage2_32[92]}
   );
   gpc1_1 gpc6687 (
      {stage1_32[204]},
      {stage2_32[93]}
   );
   gpc1_1 gpc6688 (
      {stage1_32[205]},
      {stage2_32[94]}
   );
   gpc1_1 gpc6689 (
      {stage1_32[206]},
      {stage2_32[95]}
   );
   gpc1_1 gpc6690 (
      {stage1_32[207]},
      {stage2_32[96]}
   );
   gpc1_1 gpc6691 (
      {stage1_32[208]},
      {stage2_32[97]}
   );
   gpc1_1 gpc6692 (
      {stage1_32[209]},
      {stage2_32[98]}
   );
   gpc1_1 gpc6693 (
      {stage1_32[210]},
      {stage2_32[99]}
   );
   gpc1_1 gpc6694 (
      {stage1_32[211]},
      {stage2_32[100]}
   );
   gpc1_1 gpc6695 (
      {stage1_32[212]},
      {stage2_32[101]}
   );
   gpc1_1 gpc6696 (
      {stage1_32[213]},
      {stage2_32[102]}
   );
   gpc1_1 gpc6697 (
      {stage1_32[214]},
      {stage2_32[103]}
   );
   gpc1_1 gpc6698 (
      {stage1_32[215]},
      {stage2_32[104]}
   );
   gpc1_1 gpc6699 (
      {stage1_32[216]},
      {stage2_32[105]}
   );
   gpc1_1 gpc6700 (
      {stage1_34[140]},
      {stage2_34[82]}
   );
   gpc1_1 gpc6701 (
      {stage1_34[141]},
      {stage2_34[83]}
   );
   gpc1_1 gpc6702 (
      {stage1_34[142]},
      {stage2_34[84]}
   );
   gpc1_1 gpc6703 (
      {stage1_34[143]},
      {stage2_34[85]}
   );
   gpc1_1 gpc6704 (
      {stage1_34[144]},
      {stage2_34[86]}
   );
   gpc1_1 gpc6705 (
      {stage1_34[145]},
      {stage2_34[87]}
   );
   gpc1_1 gpc6706 (
      {stage1_34[146]},
      {stage2_34[88]}
   );
   gpc1_1 gpc6707 (
      {stage1_34[147]},
      {stage2_34[89]}
   );
   gpc1_1 gpc6708 (
      {stage1_34[148]},
      {stage2_34[90]}
   );
   gpc1_1 gpc6709 (
      {stage1_34[149]},
      {stage2_34[91]}
   );
   gpc1_1 gpc6710 (
      {stage1_34[150]},
      {stage2_34[92]}
   );
   gpc1_1 gpc6711 (
      {stage1_34[151]},
      {stage2_34[93]}
   );
   gpc1_1 gpc6712 (
      {stage1_34[152]},
      {stage2_34[94]}
   );
   gpc1_1 gpc6713 (
      {stage1_34[153]},
      {stage2_34[95]}
   );
   gpc1_1 gpc6714 (
      {stage1_34[154]},
      {stage2_34[96]}
   );
   gpc1_1 gpc6715 (
      {stage1_34[155]},
      {stage2_34[97]}
   );
   gpc1_1 gpc6716 (
      {stage1_34[156]},
      {stage2_34[98]}
   );
   gpc1_1 gpc6717 (
      {stage1_34[157]},
      {stage2_34[99]}
   );
   gpc1_1 gpc6718 (
      {stage1_34[158]},
      {stage2_34[100]}
   );
   gpc1_1 gpc6719 (
      {stage1_34[159]},
      {stage2_34[101]}
   );
   gpc1_1 gpc6720 (
      {stage1_34[160]},
      {stage2_34[102]}
   );
   gpc1_1 gpc6721 (
      {stage1_34[161]},
      {stage2_34[103]}
   );
   gpc1_1 gpc6722 (
      {stage1_34[162]},
      {stage2_34[104]}
   );
   gpc1_1 gpc6723 (
      {stage1_34[163]},
      {stage2_34[105]}
   );
   gpc1_1 gpc6724 (
      {stage1_34[164]},
      {stage2_34[106]}
   );
   gpc1_1 gpc6725 (
      {stage1_34[165]},
      {stage2_34[107]}
   );
   gpc1_1 gpc6726 (
      {stage1_34[166]},
      {stage2_34[108]}
   );
   gpc1_1 gpc6727 (
      {stage1_34[167]},
      {stage2_34[109]}
   );
   gpc1_1 gpc6728 (
      {stage1_34[168]},
      {stage2_34[110]}
   );
   gpc1_1 gpc6729 (
      {stage1_34[169]},
      {stage2_34[111]}
   );
   gpc1_1 gpc6730 (
      {stage1_34[170]},
      {stage2_34[112]}
   );
   gpc1_1 gpc6731 (
      {stage1_34[171]},
      {stage2_34[113]}
   );
   gpc1_1 gpc6732 (
      {stage1_34[172]},
      {stage2_34[114]}
   );
   gpc1_1 gpc6733 (
      {stage1_34[173]},
      {stage2_34[115]}
   );
   gpc1_1 gpc6734 (
      {stage1_34[174]},
      {stage2_34[116]}
   );
   gpc1_1 gpc6735 (
      {stage1_34[175]},
      {stage2_34[117]}
   );
   gpc1_1 gpc6736 (
      {stage1_34[176]},
      {stage2_34[118]}
   );
   gpc1_1 gpc6737 (
      {stage1_34[177]},
      {stage2_34[119]}
   );
   gpc1_1 gpc6738 (
      {stage1_34[178]},
      {stage2_34[120]}
   );
   gpc1_1 gpc6739 (
      {stage1_34[179]},
      {stage2_34[121]}
   );
   gpc1_1 gpc6740 (
      {stage1_34[180]},
      {stage2_34[122]}
   );
   gpc1_1 gpc6741 (
      {stage1_34[181]},
      {stage2_34[123]}
   );
   gpc1_1 gpc6742 (
      {stage1_34[182]},
      {stage2_34[124]}
   );
   gpc1_1 gpc6743 (
      {stage1_34[183]},
      {stage2_34[125]}
   );
   gpc1_1 gpc6744 (
      {stage1_34[184]},
      {stage2_34[126]}
   );
   gpc1_1 gpc6745 (
      {stage1_34[185]},
      {stage2_34[127]}
   );
   gpc1_1 gpc6746 (
      {stage1_34[186]},
      {stage2_34[128]}
   );
   gpc1_1 gpc6747 (
      {stage1_34[187]},
      {stage2_34[129]}
   );
   gpc1_1 gpc6748 (
      {stage1_34[188]},
      {stage2_34[130]}
   );
   gpc1_1 gpc6749 (
      {stage1_34[189]},
      {stage2_34[131]}
   );
   gpc1_1 gpc6750 (
      {stage1_35[178]},
      {stage2_35[94]}
   );
   gpc1_1 gpc6751 (
      {stage1_35[179]},
      {stage2_35[95]}
   );
   gpc1_1 gpc6752 (
      {stage1_35[180]},
      {stage2_35[96]}
   );
   gpc1_1 gpc6753 (
      {stage1_35[181]},
      {stage2_35[97]}
   );
   gpc1_1 gpc6754 (
      {stage1_35[182]},
      {stage2_35[98]}
   );
   gpc1_1 gpc6755 (
      {stage1_35[183]},
      {stage2_35[99]}
   );
   gpc1_1 gpc6756 (
      {stage1_35[184]},
      {stage2_35[100]}
   );
   gpc1_1 gpc6757 (
      {stage1_35[185]},
      {stage2_35[101]}
   );
   gpc1_1 gpc6758 (
      {stage1_35[186]},
      {stage2_35[102]}
   );
   gpc1_1 gpc6759 (
      {stage1_35[187]},
      {stage2_35[103]}
   );
   gpc1_1 gpc6760 (
      {stage1_35[188]},
      {stage2_35[104]}
   );
   gpc1_1 gpc6761 (
      {stage1_35[189]},
      {stage2_35[105]}
   );
   gpc1_1 gpc6762 (
      {stage1_35[190]},
      {stage2_35[106]}
   );
   gpc1_1 gpc6763 (
      {stage1_35[191]},
      {stage2_35[107]}
   );
   gpc1_1 gpc6764 (
      {stage1_35[192]},
      {stage2_35[108]}
   );
   gpc1_1 gpc6765 (
      {stage1_35[193]},
      {stage2_35[109]}
   );
   gpc1_1 gpc6766 (
      {stage1_35[194]},
      {stage2_35[110]}
   );
   gpc1_1 gpc6767 (
      {stage1_35[195]},
      {stage2_35[111]}
   );
   gpc1_1 gpc6768 (
      {stage1_35[196]},
      {stage2_35[112]}
   );
   gpc1_1 gpc6769 (
      {stage1_35[197]},
      {stage2_35[113]}
   );
   gpc1_1 gpc6770 (
      {stage1_35[198]},
      {stage2_35[114]}
   );
   gpc1_1 gpc6771 (
      {stage1_35[199]},
      {stage2_35[115]}
   );
   gpc1_1 gpc6772 (
      {stage1_35[200]},
      {stage2_35[116]}
   );
   gpc1_1 gpc6773 (
      {stage1_35[201]},
      {stage2_35[117]}
   );
   gpc1_1 gpc6774 (
      {stage1_35[202]},
      {stage2_35[118]}
   );
   gpc1_1 gpc6775 (
      {stage1_35[203]},
      {stage2_35[119]}
   );
   gpc1_1 gpc6776 (
      {stage1_35[204]},
      {stage2_35[120]}
   );
   gpc1_1 gpc6777 (
      {stage1_35[205]},
      {stage2_35[121]}
   );
   gpc1_1 gpc6778 (
      {stage1_35[206]},
      {stage2_35[122]}
   );
   gpc1_1 gpc6779 (
      {stage1_35[207]},
      {stage2_35[123]}
   );
   gpc1_1 gpc6780 (
      {stage1_35[208]},
      {stage2_35[124]}
   );
   gpc1_1 gpc6781 (
      {stage1_35[209]},
      {stage2_35[125]}
   );
   gpc1_1 gpc6782 (
      {stage1_35[210]},
      {stage2_35[126]}
   );
   gpc1_1 gpc6783 (
      {stage1_35[211]},
      {stage2_35[127]}
   );
   gpc1_1 gpc6784 (
      {stage1_35[212]},
      {stage2_35[128]}
   );
   gpc1_1 gpc6785 (
      {stage1_35[213]},
      {stage2_35[129]}
   );
   gpc1_1 gpc6786 (
      {stage1_35[214]},
      {stage2_35[130]}
   );
   gpc1_1 gpc6787 (
      {stage1_35[215]},
      {stage2_35[131]}
   );
   gpc1_1 gpc6788 (
      {stage1_35[216]},
      {stage2_35[132]}
   );
   gpc1_1 gpc6789 (
      {stage1_37[306]},
      {stage2_37[88]}
   );
   gpc1_1 gpc6790 (
      {stage1_37[307]},
      {stage2_37[89]}
   );
   gpc1_1 gpc6791 (
      {stage1_38[231]},
      {stage2_38[106]}
   );
   gpc1_1 gpc6792 (
      {stage1_38[232]},
      {stage2_38[107]}
   );
   gpc1_1 gpc6793 (
      {stage1_38[233]},
      {stage2_38[108]}
   );
   gpc1_1 gpc6794 (
      {stage1_38[234]},
      {stage2_38[109]}
   );
   gpc1_1 gpc6795 (
      {stage1_38[235]},
      {stage2_38[110]}
   );
   gpc1_1 gpc6796 (
      {stage1_38[236]},
      {stage2_38[111]}
   );
   gpc1_1 gpc6797 (
      {stage1_38[237]},
      {stage2_38[112]}
   );
   gpc1_1 gpc6798 (
      {stage1_38[238]},
      {stage2_38[113]}
   );
   gpc1_1 gpc6799 (
      {stage1_38[239]},
      {stage2_38[114]}
   );
   gpc1_1 gpc6800 (
      {stage1_38[240]},
      {stage2_38[115]}
   );
   gpc1_1 gpc6801 (
      {stage1_38[241]},
      {stage2_38[116]}
   );
   gpc1_1 gpc6802 (
      {stage1_38[242]},
      {stage2_38[117]}
   );
   gpc1_1 gpc6803 (
      {stage1_38[243]},
      {stage2_38[118]}
   );
   gpc1_1 gpc6804 (
      {stage1_38[244]},
      {stage2_38[119]}
   );
   gpc1_1 gpc6805 (
      {stage1_38[245]},
      {stage2_38[120]}
   );
   gpc1_1 gpc6806 (
      {stage1_38[246]},
      {stage2_38[121]}
   );
   gpc1_1 gpc6807 (
      {stage1_38[247]},
      {stage2_38[122]}
   );
   gpc1_1 gpc6808 (
      {stage1_38[248]},
      {stage2_38[123]}
   );
   gpc1_1 gpc6809 (
      {stage1_38[249]},
      {stage2_38[124]}
   );
   gpc1_1 gpc6810 (
      {stage1_38[250]},
      {stage2_38[125]}
   );
   gpc1_1 gpc6811 (
      {stage1_38[251]},
      {stage2_38[126]}
   );
   gpc1_1 gpc6812 (
      {stage1_38[252]},
      {stage2_38[127]}
   );
   gpc1_1 gpc6813 (
      {stage1_38[253]},
      {stage2_38[128]}
   );
   gpc1_1 gpc6814 (
      {stage1_38[254]},
      {stage2_38[129]}
   );
   gpc1_1 gpc6815 (
      {stage1_38[255]},
      {stage2_38[130]}
   );
   gpc1_1 gpc6816 (
      {stage1_38[256]},
      {stage2_38[131]}
   );
   gpc1_1 gpc6817 (
      {stage1_38[257]},
      {stage2_38[132]}
   );
   gpc1_1 gpc6818 (
      {stage1_38[258]},
      {stage2_38[133]}
   );
   gpc1_1 gpc6819 (
      {stage1_38[259]},
      {stage2_38[134]}
   );
   gpc1_1 gpc6820 (
      {stage1_38[260]},
      {stage2_38[135]}
   );
   gpc1_1 gpc6821 (
      {stage1_38[261]},
      {stage2_38[136]}
   );
   gpc1_1 gpc6822 (
      {stage1_38[262]},
      {stage2_38[137]}
   );
   gpc1_1 gpc6823 (
      {stage1_38[263]},
      {stage2_38[138]}
   );
   gpc1_1 gpc6824 (
      {stage1_38[264]},
      {stage2_38[139]}
   );
   gpc1_1 gpc6825 (
      {stage1_39[170]},
      {stage2_39[94]}
   );
   gpc1_1 gpc6826 (
      {stage1_39[171]},
      {stage2_39[95]}
   );
   gpc1_1 gpc6827 (
      {stage1_39[172]},
      {stage2_39[96]}
   );
   gpc1_1 gpc6828 (
      {stage1_39[173]},
      {stage2_39[97]}
   );
   gpc1_1 gpc6829 (
      {stage1_39[174]},
      {stage2_39[98]}
   );
   gpc1_1 gpc6830 (
      {stage1_39[175]},
      {stage2_39[99]}
   );
   gpc1_1 gpc6831 (
      {stage1_39[176]},
      {stage2_39[100]}
   );
   gpc1_1 gpc6832 (
      {stage1_39[177]},
      {stage2_39[101]}
   );
   gpc1_1 gpc6833 (
      {stage1_39[178]},
      {stage2_39[102]}
   );
   gpc1_1 gpc6834 (
      {stage1_39[179]},
      {stage2_39[103]}
   );
   gpc1_1 gpc6835 (
      {stage1_39[180]},
      {stage2_39[104]}
   );
   gpc1_1 gpc6836 (
      {stage1_39[181]},
      {stage2_39[105]}
   );
   gpc1_1 gpc6837 (
      {stage1_39[182]},
      {stage2_39[106]}
   );
   gpc1_1 gpc6838 (
      {stage1_39[183]},
      {stage2_39[107]}
   );
   gpc1_1 gpc6839 (
      {stage1_39[184]},
      {stage2_39[108]}
   );
   gpc1_1 gpc6840 (
      {stage1_39[185]},
      {stage2_39[109]}
   );
   gpc1_1 gpc6841 (
      {stage1_39[186]},
      {stage2_39[110]}
   );
   gpc1_1 gpc6842 (
      {stage1_39[187]},
      {stage2_39[111]}
   );
   gpc1_1 gpc6843 (
      {stage1_39[188]},
      {stage2_39[112]}
   );
   gpc1_1 gpc6844 (
      {stage1_39[189]},
      {stage2_39[113]}
   );
   gpc1_1 gpc6845 (
      {stage1_39[190]},
      {stage2_39[114]}
   );
   gpc1_1 gpc6846 (
      {stage1_39[191]},
      {stage2_39[115]}
   );
   gpc1_1 gpc6847 (
      {stage1_39[192]},
      {stage2_39[116]}
   );
   gpc1_1 gpc6848 (
      {stage1_39[193]},
      {stage2_39[117]}
   );
   gpc1_1 gpc6849 (
      {stage1_39[194]},
      {stage2_39[118]}
   );
   gpc1_1 gpc6850 (
      {stage1_39[195]},
      {stage2_39[119]}
   );
   gpc1_1 gpc6851 (
      {stage1_39[196]},
      {stage2_39[120]}
   );
   gpc1_1 gpc6852 (
      {stage1_39[197]},
      {stage2_39[121]}
   );
   gpc1_1 gpc6853 (
      {stage1_39[198]},
      {stage2_39[122]}
   );
   gpc1_1 gpc6854 (
      {stage1_39[199]},
      {stage2_39[123]}
   );
   gpc1_1 gpc6855 (
      {stage1_39[200]},
      {stage2_39[124]}
   );
   gpc1_1 gpc6856 (
      {stage1_39[201]},
      {stage2_39[125]}
   );
   gpc1_1 gpc6857 (
      {stage1_39[202]},
      {stage2_39[126]}
   );
   gpc1_1 gpc6858 (
      {stage1_39[203]},
      {stage2_39[127]}
   );
   gpc1_1 gpc6859 (
      {stage1_39[204]},
      {stage2_39[128]}
   );
   gpc1_1 gpc6860 (
      {stage1_39[205]},
      {stage2_39[129]}
   );
   gpc1_1 gpc6861 (
      {stage1_39[206]},
      {stage2_39[130]}
   );
   gpc1_1 gpc6862 (
      {stage1_39[207]},
      {stage2_39[131]}
   );
   gpc1_1 gpc6863 (
      {stage1_39[208]},
      {stage2_39[132]}
   );
   gpc1_1 gpc6864 (
      {stage1_39[209]},
      {stage2_39[133]}
   );
   gpc1_1 gpc6865 (
      {stage1_39[210]},
      {stage2_39[134]}
   );
   gpc1_1 gpc6866 (
      {stage1_39[211]},
      {stage2_39[135]}
   );
   gpc1_1 gpc6867 (
      {stage1_39[212]},
      {stage2_39[136]}
   );
   gpc1_1 gpc6868 (
      {stage1_40[281]},
      {stage2_40[90]}
   );
   gpc1_1 gpc6869 (
      {stage1_40[282]},
      {stage2_40[91]}
   );
   gpc1_1 gpc6870 (
      {stage1_40[283]},
      {stage2_40[92]}
   );
   gpc1_1 gpc6871 (
      {stage1_40[284]},
      {stage2_40[93]}
   );
   gpc1_1 gpc6872 (
      {stage1_40[285]},
      {stage2_40[94]}
   );
   gpc1_1 gpc6873 (
      {stage1_40[286]},
      {stage2_40[95]}
   );
   gpc1_1 gpc6874 (
      {stage1_40[287]},
      {stage2_40[96]}
   );
   gpc1_1 gpc6875 (
      {stage1_40[288]},
      {stage2_40[97]}
   );
   gpc1_1 gpc6876 (
      {stage1_40[289]},
      {stage2_40[98]}
   );
   gpc1_1 gpc6877 (
      {stage1_40[290]},
      {stage2_40[99]}
   );
   gpc1_1 gpc6878 (
      {stage1_40[291]},
      {stage2_40[100]}
   );
   gpc1_1 gpc6879 (
      {stage1_40[292]},
      {stage2_40[101]}
   );
   gpc1_1 gpc6880 (
      {stage1_40[293]},
      {stage2_40[102]}
   );
   gpc1_1 gpc6881 (
      {stage1_40[294]},
      {stage2_40[103]}
   );
   gpc1_1 gpc6882 (
      {stage1_40[295]},
      {stage2_40[104]}
   );
   gpc1_1 gpc6883 (
      {stage1_40[296]},
      {stage2_40[105]}
   );
   gpc1_1 gpc6884 (
      {stage1_40[297]},
      {stage2_40[106]}
   );
   gpc1_1 gpc6885 (
      {stage1_40[298]},
      {stage2_40[107]}
   );
   gpc1_1 gpc6886 (
      {stage1_40[299]},
      {stage2_40[108]}
   );
   gpc1_1 gpc6887 (
      {stage1_40[300]},
      {stage2_40[109]}
   );
   gpc1_1 gpc6888 (
      {stage1_40[301]},
      {stage2_40[110]}
   );
   gpc1_1 gpc6889 (
      {stage1_40[302]},
      {stage2_40[111]}
   );
   gpc1_1 gpc6890 (
      {stage1_40[303]},
      {stage2_40[112]}
   );
   gpc1_1 gpc6891 (
      {stage1_41[168]},
      {stage2_41[103]}
   );
   gpc1_1 gpc6892 (
      {stage1_41[169]},
      {stage2_41[104]}
   );
   gpc1_1 gpc6893 (
      {stage1_41[170]},
      {stage2_41[105]}
   );
   gpc1_1 gpc6894 (
      {stage1_42[168]},
      {stage2_42[80]}
   );
   gpc1_1 gpc6895 (
      {stage1_42[169]},
      {stage2_42[81]}
   );
   gpc1_1 gpc6896 (
      {stage1_42[170]},
      {stage2_42[82]}
   );
   gpc1_1 gpc6897 (
      {stage1_42[171]},
      {stage2_42[83]}
   );
   gpc1_1 gpc6898 (
      {stage1_42[172]},
      {stage2_42[84]}
   );
   gpc1_1 gpc6899 (
      {stage1_42[173]},
      {stage2_42[85]}
   );
   gpc1_1 gpc6900 (
      {stage1_43[241]},
      {stage2_43[66]}
   );
   gpc1_1 gpc6901 (
      {stage1_43[242]},
      {stage2_43[67]}
   );
   gpc1_1 gpc6902 (
      {stage1_43[243]},
      {stage2_43[68]}
   );
   gpc1_1 gpc6903 (
      {stage1_43[244]},
      {stage2_43[69]}
   );
   gpc1_1 gpc6904 (
      {stage1_43[245]},
      {stage2_43[70]}
   );
   gpc1_1 gpc6905 (
      {stage1_43[246]},
      {stage2_43[71]}
   );
   gpc1_1 gpc6906 (
      {stage1_43[247]},
      {stage2_43[72]}
   );
   gpc1_1 gpc6907 (
      {stage1_43[248]},
      {stage2_43[73]}
   );
   gpc1_1 gpc6908 (
      {stage1_43[249]},
      {stage2_43[74]}
   );
   gpc1_1 gpc6909 (
      {stage1_43[250]},
      {stage2_43[75]}
   );
   gpc1_1 gpc6910 (
      {stage1_43[251]},
      {stage2_43[76]}
   );
   gpc1_1 gpc6911 (
      {stage1_43[252]},
      {stage2_43[77]}
   );
   gpc1_1 gpc6912 (
      {stage1_43[253]},
      {stage2_43[78]}
   );
   gpc1_1 gpc6913 (
      {stage1_44[240]},
      {stage2_44[103]}
   );
   gpc1_1 gpc6914 (
      {stage1_44[241]},
      {stage2_44[104]}
   );
   gpc1_1 gpc6915 (
      {stage1_44[242]},
      {stage2_44[105]}
   );
   gpc1_1 gpc6916 (
      {stage1_44[243]},
      {stage2_44[106]}
   );
   gpc1_1 gpc6917 (
      {stage1_44[244]},
      {stage2_44[107]}
   );
   gpc1_1 gpc6918 (
      {stage1_44[245]},
      {stage2_44[108]}
   );
   gpc1_1 gpc6919 (
      {stage1_44[246]},
      {stage2_44[109]}
   );
   gpc1_1 gpc6920 (
      {stage1_44[247]},
      {stage2_44[110]}
   );
   gpc1_1 gpc6921 (
      {stage1_44[248]},
      {stage2_44[111]}
   );
   gpc1_1 gpc6922 (
      {stage1_44[249]},
      {stage2_44[112]}
   );
   gpc1_1 gpc6923 (
      {stage1_44[250]},
      {stage2_44[113]}
   );
   gpc1_1 gpc6924 (
      {stage1_44[251]},
      {stage2_44[114]}
   );
   gpc1_1 gpc6925 (
      {stage1_44[252]},
      {stage2_44[115]}
   );
   gpc1_1 gpc6926 (
      {stage1_44[253]},
      {stage2_44[116]}
   );
   gpc1_1 gpc6927 (
      {stage1_44[254]},
      {stage2_44[117]}
   );
   gpc1_1 gpc6928 (
      {stage1_44[255]},
      {stage2_44[118]}
   );
   gpc1_1 gpc6929 (
      {stage1_45[199]},
      {stage2_45[105]}
   );
   gpc1_1 gpc6930 (
      {stage1_45[200]},
      {stage2_45[106]}
   );
   gpc1_1 gpc6931 (
      {stage1_45[201]},
      {stage2_45[107]}
   );
   gpc1_1 gpc6932 (
      {stage1_45[202]},
      {stage2_45[108]}
   );
   gpc1_1 gpc6933 (
      {stage1_45[203]},
      {stage2_45[109]}
   );
   gpc1_1 gpc6934 (
      {stage1_45[204]},
      {stage2_45[110]}
   );
   gpc1_1 gpc6935 (
      {stage1_45[205]},
      {stage2_45[111]}
   );
   gpc1_1 gpc6936 (
      {stage1_45[206]},
      {stage2_45[112]}
   );
   gpc1_1 gpc6937 (
      {stage1_45[207]},
      {stage2_45[113]}
   );
   gpc1_1 gpc6938 (
      {stage1_45[208]},
      {stage2_45[114]}
   );
   gpc1_1 gpc6939 (
      {stage1_45[209]},
      {stage2_45[115]}
   );
   gpc1_1 gpc6940 (
      {stage1_45[210]},
      {stage2_45[116]}
   );
   gpc1_1 gpc6941 (
      {stage1_45[211]},
      {stage2_45[117]}
   );
   gpc1_1 gpc6942 (
      {stage1_46[295]},
      {stage2_46[85]}
   );
   gpc1_1 gpc6943 (
      {stage1_46[296]},
      {stage2_46[86]}
   );
   gpc1_1 gpc6944 (
      {stage1_46[297]},
      {stage2_46[87]}
   );
   gpc1_1 gpc6945 (
      {stage1_47[230]},
      {stage2_47[98]}
   );
   gpc1_1 gpc6946 (
      {stage1_47[231]},
      {stage2_47[99]}
   );
   gpc1_1 gpc6947 (
      {stage1_47[232]},
      {stage2_47[100]}
   );
   gpc1_1 gpc6948 (
      {stage1_47[233]},
      {stage2_47[101]}
   );
   gpc1_1 gpc6949 (
      {stage1_47[234]},
      {stage2_47[102]}
   );
   gpc1_1 gpc6950 (
      {stage1_47[235]},
      {stage2_47[103]}
   );
   gpc1_1 gpc6951 (
      {stage1_48[172]},
      {stage2_48[104]}
   );
   gpc1_1 gpc6952 (
      {stage1_48[173]},
      {stage2_48[105]}
   );
   gpc1_1 gpc6953 (
      {stage1_48[174]},
      {stage2_48[106]}
   );
   gpc1_1 gpc6954 (
      {stage1_48[175]},
      {stage2_48[107]}
   );
   gpc1_1 gpc6955 (
      {stage1_48[176]},
      {stage2_48[108]}
   );
   gpc1_1 gpc6956 (
      {stage1_48[177]},
      {stage2_48[109]}
   );
   gpc1_1 gpc6957 (
      {stage1_48[178]},
      {stage2_48[110]}
   );
   gpc1_1 gpc6958 (
      {stage1_48[179]},
      {stage2_48[111]}
   );
   gpc1_1 gpc6959 (
      {stage1_48[180]},
      {stage2_48[112]}
   );
   gpc1_1 gpc6960 (
      {stage1_48[181]},
      {stage2_48[113]}
   );
   gpc1_1 gpc6961 (
      {stage1_48[182]},
      {stage2_48[114]}
   );
   gpc1_1 gpc6962 (
      {stage1_48[183]},
      {stage2_48[115]}
   );
   gpc1_1 gpc6963 (
      {stage1_48[184]},
      {stage2_48[116]}
   );
   gpc1_1 gpc6964 (
      {stage1_48[185]},
      {stage2_48[117]}
   );
   gpc1_1 gpc6965 (
      {stage1_48[186]},
      {stage2_48[118]}
   );
   gpc1_1 gpc6966 (
      {stage1_48[187]},
      {stage2_48[119]}
   );
   gpc1_1 gpc6967 (
      {stage1_48[188]},
      {stage2_48[120]}
   );
   gpc1_1 gpc6968 (
      {stage1_48[189]},
      {stage2_48[121]}
   );
   gpc1_1 gpc6969 (
      {stage1_48[190]},
      {stage2_48[122]}
   );
   gpc1_1 gpc6970 (
      {stage1_48[191]},
      {stage2_48[123]}
   );
   gpc1_1 gpc6971 (
      {stage1_48[192]},
      {stage2_48[124]}
   );
   gpc1_1 gpc6972 (
      {stage1_48[193]},
      {stage2_48[125]}
   );
   gpc1_1 gpc6973 (
      {stage1_48[194]},
      {stage2_48[126]}
   );
   gpc1_1 gpc6974 (
      {stage1_48[195]},
      {stage2_48[127]}
   );
   gpc1_1 gpc6975 (
      {stage1_48[196]},
      {stage2_48[128]}
   );
   gpc1_1 gpc6976 (
      {stage1_48[197]},
      {stage2_48[129]}
   );
   gpc1_1 gpc6977 (
      {stage1_49[154]},
      {stage2_49[77]}
   );
   gpc1_1 gpc6978 (
      {stage1_49[155]},
      {stage2_49[78]}
   );
   gpc1_1 gpc6979 (
      {stage1_49[156]},
      {stage2_49[79]}
   );
   gpc1_1 gpc6980 (
      {stage1_49[157]},
      {stage2_49[80]}
   );
   gpc1_1 gpc6981 (
      {stage1_49[158]},
      {stage2_49[81]}
   );
   gpc1_1 gpc6982 (
      {stage1_49[159]},
      {stage2_49[82]}
   );
   gpc1_1 gpc6983 (
      {stage1_49[160]},
      {stage2_49[83]}
   );
   gpc1_1 gpc6984 (
      {stage1_49[161]},
      {stage2_49[84]}
   );
   gpc1_1 gpc6985 (
      {stage1_49[162]},
      {stage2_49[85]}
   );
   gpc1_1 gpc6986 (
      {stage1_49[163]},
      {stage2_49[86]}
   );
   gpc1_1 gpc6987 (
      {stage1_49[164]},
      {stage2_49[87]}
   );
   gpc1_1 gpc6988 (
      {stage1_49[165]},
      {stage2_49[88]}
   );
   gpc1_1 gpc6989 (
      {stage1_49[166]},
      {stage2_49[89]}
   );
   gpc1_1 gpc6990 (
      {stage1_49[167]},
      {stage2_49[90]}
   );
   gpc1_1 gpc6991 (
      {stage1_49[168]},
      {stage2_49[91]}
   );
   gpc1_1 gpc6992 (
      {stage1_49[169]},
      {stage2_49[92]}
   );
   gpc1_1 gpc6993 (
      {stage1_49[170]},
      {stage2_49[93]}
   );
   gpc1_1 gpc6994 (
      {stage1_49[171]},
      {stage2_49[94]}
   );
   gpc1_1 gpc6995 (
      {stage1_49[172]},
      {stage2_49[95]}
   );
   gpc1_1 gpc6996 (
      {stage1_50[179]},
      {stage2_50[75]}
   );
   gpc1_1 gpc6997 (
      {stage1_50[180]},
      {stage2_50[76]}
   );
   gpc1_1 gpc6998 (
      {stage1_50[181]},
      {stage2_50[77]}
   );
   gpc1_1 gpc6999 (
      {stage1_50[182]},
      {stage2_50[78]}
   );
   gpc1_1 gpc7000 (
      {stage1_50[183]},
      {stage2_50[79]}
   );
   gpc1_1 gpc7001 (
      {stage1_50[184]},
      {stage2_50[80]}
   );
   gpc1_1 gpc7002 (
      {stage1_50[185]},
      {stage2_50[81]}
   );
   gpc1_1 gpc7003 (
      {stage1_50[186]},
      {stage2_50[82]}
   );
   gpc1_1 gpc7004 (
      {stage1_50[187]},
      {stage2_50[83]}
   );
   gpc1_1 gpc7005 (
      {stage1_50[188]},
      {stage2_50[84]}
   );
   gpc1_1 gpc7006 (
      {stage1_50[189]},
      {stage2_50[85]}
   );
   gpc1_1 gpc7007 (
      {stage1_51[266]},
      {stage2_51[79]}
   );
   gpc1_1 gpc7008 (
      {stage1_51[267]},
      {stage2_51[80]}
   );
   gpc1_1 gpc7009 (
      {stage1_51[268]},
      {stage2_51[81]}
   );
   gpc1_1 gpc7010 (
      {stage1_51[269]},
      {stage2_51[82]}
   );
   gpc1_1 gpc7011 (
      {stage1_51[270]},
      {stage2_51[83]}
   );
   gpc1_1 gpc7012 (
      {stage1_51[271]},
      {stage2_51[84]}
   );
   gpc1_1 gpc7013 (
      {stage1_51[272]},
      {stage2_51[85]}
   );
   gpc1_1 gpc7014 (
      {stage1_51[273]},
      {stage2_51[86]}
   );
   gpc1_1 gpc7015 (
      {stage1_51[274]},
      {stage2_51[87]}
   );
   gpc1_1 gpc7016 (
      {stage1_52[187]},
      {stage2_52[93]}
   );
   gpc1_1 gpc7017 (
      {stage1_52[188]},
      {stage2_52[94]}
   );
   gpc1_1 gpc7018 (
      {stage1_52[189]},
      {stage2_52[95]}
   );
   gpc1_1 gpc7019 (
      {stage1_52[190]},
      {stage2_52[96]}
   );
   gpc1_1 gpc7020 (
      {stage1_52[191]},
      {stage2_52[97]}
   );
   gpc1_1 gpc7021 (
      {stage1_52[192]},
      {stage2_52[98]}
   );
   gpc1_1 gpc7022 (
      {stage1_52[193]},
      {stage2_52[99]}
   );
   gpc1_1 gpc7023 (
      {stage1_52[194]},
      {stage2_52[100]}
   );
   gpc1_1 gpc7024 (
      {stage1_52[195]},
      {stage2_52[101]}
   );
   gpc1_1 gpc7025 (
      {stage1_52[196]},
      {stage2_52[102]}
   );
   gpc1_1 gpc7026 (
      {stage1_52[197]},
      {stage2_52[103]}
   );
   gpc1_1 gpc7027 (
      {stage1_52[198]},
      {stage2_52[104]}
   );
   gpc1_1 gpc7028 (
      {stage1_53[130]},
      {stage2_53[76]}
   );
   gpc1_1 gpc7029 (
      {stage1_53[131]},
      {stage2_53[77]}
   );
   gpc1_1 gpc7030 (
      {stage1_53[132]},
      {stage2_53[78]}
   );
   gpc1_1 gpc7031 (
      {stage1_53[133]},
      {stage2_53[79]}
   );
   gpc1_1 gpc7032 (
      {stage1_53[134]},
      {stage2_53[80]}
   );
   gpc1_1 gpc7033 (
      {stage1_53[135]},
      {stage2_53[81]}
   );
   gpc1_1 gpc7034 (
      {stage1_53[136]},
      {stage2_53[82]}
   );
   gpc1_1 gpc7035 (
      {stage1_53[137]},
      {stage2_53[83]}
   );
   gpc1_1 gpc7036 (
      {stage1_53[138]},
      {stage2_53[84]}
   );
   gpc1_1 gpc7037 (
      {stage1_53[139]},
      {stage2_53[85]}
   );
   gpc1_1 gpc7038 (
      {stage1_53[140]},
      {stage2_53[86]}
   );
   gpc1_1 gpc7039 (
      {stage1_53[141]},
      {stage2_53[87]}
   );
   gpc1_1 gpc7040 (
      {stage1_53[142]},
      {stage2_53[88]}
   );
   gpc1_1 gpc7041 (
      {stage1_53[143]},
      {stage2_53[89]}
   );
   gpc1_1 gpc7042 (
      {stage1_53[144]},
      {stage2_53[90]}
   );
   gpc1_1 gpc7043 (
      {stage1_53[145]},
      {stage2_53[91]}
   );
   gpc1_1 gpc7044 (
      {stage1_53[146]},
      {stage2_53[92]}
   );
   gpc1_1 gpc7045 (
      {stage1_53[147]},
      {stage2_53[93]}
   );
   gpc1_1 gpc7046 (
      {stage1_53[148]},
      {stage2_53[94]}
   );
   gpc1_1 gpc7047 (
      {stage1_53[149]},
      {stage2_53[95]}
   );
   gpc1_1 gpc7048 (
      {stage1_53[150]},
      {stage2_53[96]}
   );
   gpc1_1 gpc7049 (
      {stage1_53[151]},
      {stage2_53[97]}
   );
   gpc1_1 gpc7050 (
      {stage1_53[152]},
      {stage2_53[98]}
   );
   gpc1_1 gpc7051 (
      {stage1_53[153]},
      {stage2_53[99]}
   );
   gpc1_1 gpc7052 (
      {stage1_53[154]},
      {stage2_53[100]}
   );
   gpc1_1 gpc7053 (
      {stage1_53[155]},
      {stage2_53[101]}
   );
   gpc1_1 gpc7054 (
      {stage1_53[156]},
      {stage2_53[102]}
   );
   gpc1_1 gpc7055 (
      {stage1_53[157]},
      {stage2_53[103]}
   );
   gpc1_1 gpc7056 (
      {stage1_53[158]},
      {stage2_53[104]}
   );
   gpc1_1 gpc7057 (
      {stage1_53[159]},
      {stage2_53[105]}
   );
   gpc1_1 gpc7058 (
      {stage1_53[160]},
      {stage2_53[106]}
   );
   gpc1_1 gpc7059 (
      {stage1_53[161]},
      {stage2_53[107]}
   );
   gpc1_1 gpc7060 (
      {stage1_53[162]},
      {stage2_53[108]}
   );
   gpc1_1 gpc7061 (
      {stage1_53[163]},
      {stage2_53[109]}
   );
   gpc1_1 gpc7062 (
      {stage1_53[164]},
      {stage2_53[110]}
   );
   gpc1_1 gpc7063 (
      {stage1_53[165]},
      {stage2_53[111]}
   );
   gpc1_1 gpc7064 (
      {stage1_53[166]},
      {stage2_53[112]}
   );
   gpc1_1 gpc7065 (
      {stage1_53[167]},
      {stage2_53[113]}
   );
   gpc1_1 gpc7066 (
      {stage1_53[168]},
      {stage2_53[114]}
   );
   gpc1_1 gpc7067 (
      {stage1_54[203]},
      {stage2_54[72]}
   );
   gpc1_1 gpc7068 (
      {stage1_54[204]},
      {stage2_54[73]}
   );
   gpc1_1 gpc7069 (
      {stage1_54[205]},
      {stage2_54[74]}
   );
   gpc1_1 gpc7070 (
      {stage1_54[206]},
      {stage2_54[75]}
   );
   gpc1_1 gpc7071 (
      {stage1_54[207]},
      {stage2_54[76]}
   );
   gpc1_1 gpc7072 (
      {stage1_54[208]},
      {stage2_54[77]}
   );
   gpc1_1 gpc7073 (
      {stage1_54[209]},
      {stage2_54[78]}
   );
   gpc1_1 gpc7074 (
      {stage1_54[210]},
      {stage2_54[79]}
   );
   gpc1_1 gpc7075 (
      {stage1_54[211]},
      {stage2_54[80]}
   );
   gpc1_1 gpc7076 (
      {stage1_54[212]},
      {stage2_54[81]}
   );
   gpc1_1 gpc7077 (
      {stage1_54[213]},
      {stage2_54[82]}
   );
   gpc1_1 gpc7078 (
      {stage1_54[214]},
      {stage2_54[83]}
   );
   gpc1_1 gpc7079 (
      {stage1_54[215]},
      {stage2_54[84]}
   );
   gpc1_1 gpc7080 (
      {stage1_54[216]},
      {stage2_54[85]}
   );
   gpc1_1 gpc7081 (
      {stage1_54[217]},
      {stage2_54[86]}
   );
   gpc1_1 gpc7082 (
      {stage1_54[218]},
      {stage2_54[87]}
   );
   gpc1_1 gpc7083 (
      {stage1_54[219]},
      {stage2_54[88]}
   );
   gpc1_1 gpc7084 (
      {stage1_54[220]},
      {stage2_54[89]}
   );
   gpc1_1 gpc7085 (
      {stage1_54[221]},
      {stage2_54[90]}
   );
   gpc1_1 gpc7086 (
      {stage1_54[222]},
      {stage2_54[91]}
   );
   gpc1_1 gpc7087 (
      {stage1_54[223]},
      {stage2_54[92]}
   );
   gpc1_1 gpc7088 (
      {stage1_54[224]},
      {stage2_54[93]}
   );
   gpc1_1 gpc7089 (
      {stage1_54[225]},
      {stage2_54[94]}
   );
   gpc1_1 gpc7090 (
      {stage1_54[226]},
      {stage2_54[95]}
   );
   gpc1_1 gpc7091 (
      {stage1_54[227]},
      {stage2_54[96]}
   );
   gpc1_1 gpc7092 (
      {stage1_54[228]},
      {stage2_54[97]}
   );
   gpc1_1 gpc7093 (
      {stage1_54[229]},
      {stage2_54[98]}
   );
   gpc1_1 gpc7094 (
      {stage1_54[230]},
      {stage2_54[99]}
   );
   gpc1_1 gpc7095 (
      {stage1_55[254]},
      {stage2_55[93]}
   );
   gpc1_1 gpc7096 (
      {stage1_55[255]},
      {stage2_55[94]}
   );
   gpc1_1 gpc7097 (
      {stage1_55[256]},
      {stage2_55[95]}
   );
   gpc1_1 gpc7098 (
      {stage1_55[257]},
      {stage2_55[96]}
   );
   gpc1_1 gpc7099 (
      {stage1_55[258]},
      {stage2_55[97]}
   );
   gpc1_1 gpc7100 (
      {stage1_55[259]},
      {stage2_55[98]}
   );
   gpc1_1 gpc7101 (
      {stage1_55[260]},
      {stage2_55[99]}
   );
   gpc1_1 gpc7102 (
      {stage1_55[261]},
      {stage2_55[100]}
   );
   gpc1_1 gpc7103 (
      {stage1_55[262]},
      {stage2_55[101]}
   );
   gpc1_1 gpc7104 (
      {stage1_55[263]},
      {stage2_55[102]}
   );
   gpc1_1 gpc7105 (
      {stage1_55[264]},
      {stage2_55[103]}
   );
   gpc1_1 gpc7106 (
      {stage1_55[265]},
      {stage2_55[104]}
   );
   gpc1_1 gpc7107 (
      {stage1_55[266]},
      {stage2_55[105]}
   );
   gpc1_1 gpc7108 (
      {stage1_56[164]},
      {stage2_56[92]}
   );
   gpc1_1 gpc7109 (
      {stage1_56[165]},
      {stage2_56[93]}
   );
   gpc1_1 gpc7110 (
      {stage1_56[166]},
      {stage2_56[94]}
   );
   gpc1_1 gpc7111 (
      {stage1_56[167]},
      {stage2_56[95]}
   );
   gpc1_1 gpc7112 (
      {stage1_56[168]},
      {stage2_56[96]}
   );
   gpc1_1 gpc7113 (
      {stage1_56[169]},
      {stage2_56[97]}
   );
   gpc1_1 gpc7114 (
      {stage1_56[170]},
      {stage2_56[98]}
   );
   gpc1_1 gpc7115 (
      {stage1_56[171]},
      {stage2_56[99]}
   );
   gpc1_1 gpc7116 (
      {stage1_56[172]},
      {stage2_56[100]}
   );
   gpc1_1 gpc7117 (
      {stage1_56[173]},
      {stage2_56[101]}
   );
   gpc1_1 gpc7118 (
      {stage1_56[174]},
      {stage2_56[102]}
   );
   gpc1_1 gpc7119 (
      {stage1_56[175]},
      {stage2_56[103]}
   );
   gpc1_1 gpc7120 (
      {stage1_56[176]},
      {stage2_56[104]}
   );
   gpc1_1 gpc7121 (
      {stage1_56[177]},
      {stage2_56[105]}
   );
   gpc1_1 gpc7122 (
      {stage1_56[178]},
      {stage2_56[106]}
   );
   gpc1_1 gpc7123 (
      {stage1_56[179]},
      {stage2_56[107]}
   );
   gpc1_1 gpc7124 (
      {stage1_56[180]},
      {stage2_56[108]}
   );
   gpc1_1 gpc7125 (
      {stage1_56[181]},
      {stage2_56[109]}
   );
   gpc1_1 gpc7126 (
      {stage1_56[182]},
      {stage2_56[110]}
   );
   gpc1_1 gpc7127 (
      {stage1_56[183]},
      {stage2_56[111]}
   );
   gpc1_1 gpc7128 (
      {stage1_56[184]},
      {stage2_56[112]}
   );
   gpc1_1 gpc7129 (
      {stage1_56[185]},
      {stage2_56[113]}
   );
   gpc1_1 gpc7130 (
      {stage1_56[186]},
      {stage2_56[114]}
   );
   gpc1_1 gpc7131 (
      {stage1_59[205]},
      {stage2_59[109]}
   );
   gpc1_1 gpc7132 (
      {stage1_60[209]},
      {stage2_60[79]}
   );
   gpc1_1 gpc7133 (
      {stage1_60[210]},
      {stage2_60[80]}
   );
   gpc1_1 gpc7134 (
      {stage1_60[211]},
      {stage2_60[81]}
   );
   gpc1_1 gpc7135 (
      {stage1_60[212]},
      {stage2_60[82]}
   );
   gpc1_1 gpc7136 (
      {stage1_60[213]},
      {stage2_60[83]}
   );
   gpc1_1 gpc7137 (
      {stage1_60[214]},
      {stage2_60[84]}
   );
   gpc1_1 gpc7138 (
      {stage1_62[192]},
      {stage2_62[104]}
   );
   gpc1_1 gpc7139 (
      {stage1_63[303]},
      {stage2_63[94]}
   );
   gpc1_1 gpc7140 (
      {stage1_63[304]},
      {stage2_63[95]}
   );
   gpc1_1 gpc7141 (
      {stage1_63[305]},
      {stage2_63[96]}
   );
   gpc1_1 gpc7142 (
      {stage1_63[306]},
      {stage2_63[97]}
   );
   gpc1_1 gpc7143 (
      {stage1_63[307]},
      {stage2_63[98]}
   );
   gpc1_1 gpc7144 (
      {stage1_64[47]},
      {stage2_64[65]}
   );
   gpc1_1 gpc7145 (
      {stage1_64[48]},
      {stage2_64[66]}
   );
   gpc1_1 gpc7146 (
      {stage1_64[49]},
      {stage2_64[67]}
   );
   gpc1_1 gpc7147 (
      {stage1_64[50]},
      {stage2_64[68]}
   );
   gpc1_1 gpc7148 (
      {stage1_64[51]},
      {stage2_64[69]}
   );
   gpc1_1 gpc7149 (
      {stage1_64[52]},
      {stage2_64[70]}
   );
   gpc1_1 gpc7150 (
      {stage1_64[53]},
      {stage2_64[71]}
   );
   gpc1_1 gpc7151 (
      {stage1_64[54]},
      {stage2_64[72]}
   );
   gpc1_1 gpc7152 (
      {stage1_64[55]},
      {stage2_64[73]}
   );
   gpc1_1 gpc7153 (
      {stage1_64[56]},
      {stage2_64[74]}
   );
   gpc1_1 gpc7154 (
      {stage1_64[57]},
      {stage2_64[75]}
   );
   gpc1_1 gpc7155 (
      {stage1_64[58]},
      {stage2_64[76]}
   );
   gpc1_1 gpc7156 (
      {stage1_64[59]},
      {stage2_64[77]}
   );
   gpc1_1 gpc7157 (
      {stage1_64[60]},
      {stage2_64[78]}
   );
   gpc1_1 gpc7158 (
      {stage1_64[61]},
      {stage2_64[79]}
   );
   gpc1_1 gpc7159 (
      {stage1_64[62]},
      {stage2_64[80]}
   );
   gpc1_1 gpc7160 (
      {stage1_64[63]},
      {stage2_64[81]}
   );
   gpc1_1 gpc7161 (
      {stage1_64[64]},
      {stage2_64[82]}
   );
   gpc1_1 gpc7162 (
      {stage1_64[65]},
      {stage2_64[83]}
   );
   gpc1_1 gpc7163 (
      {stage1_64[66]},
      {stage2_64[84]}
   );
   gpc1_1 gpc7164 (
      {stage1_64[67]},
      {stage2_64[85]}
   );
   gpc1_1 gpc7165 (
      {stage1_64[68]},
      {stage2_64[86]}
   );
   gpc1_1 gpc7166 (
      {stage1_64[69]},
      {stage2_64[87]}
   );
   gpc1_1 gpc7167 (
      {stage1_64[70]},
      {stage2_64[88]}
   );
   gpc1_1 gpc7168 (
      {stage1_64[71]},
      {stage2_64[89]}
   );
   gpc1_1 gpc7169 (
      {stage1_64[72]},
      {stage2_64[90]}
   );
   gpc1_1 gpc7170 (
      {stage1_64[73]},
      {stage2_64[91]}
   );
   gpc1_1 gpc7171 (
      {stage1_64[74]},
      {stage2_64[92]}
   );
   gpc1_1 gpc7172 (
      {stage1_64[75]},
      {stage2_64[93]}
   );
   gpc1_1 gpc7173 (
      {stage1_64[76]},
      {stage2_64[94]}
   );
   gpc1_1 gpc7174 (
      {stage1_64[77]},
      {stage2_64[95]}
   );
   gpc1_1 gpc7175 (
      {stage1_64[78]},
      {stage2_64[96]}
   );
   gpc1_1 gpc7176 (
      {stage1_64[79]},
      {stage2_64[97]}
   );
   gpc1_1 gpc7177 (
      {stage1_64[80]},
      {stage2_64[98]}
   );
   gpc1_1 gpc7178 (
      {stage1_64[81]},
      {stage2_64[99]}
   );
   gpc1_1 gpc7179 (
      {stage1_64[82]},
      {stage2_64[100]}
   );
   gpc1_1 gpc7180 (
      {stage1_64[83]},
      {stage2_64[101]}
   );
   gpc1_1 gpc7181 (
      {stage1_64[84]},
      {stage2_64[102]}
   );
   gpc1_1 gpc7182 (
      {stage1_64[85]},
      {stage2_64[103]}
   );
   gpc1_1 gpc7183 (
      {stage1_64[86]},
      {stage2_64[104]}
   );
   gpc1_1 gpc7184 (
      {stage1_64[87]},
      {stage2_64[105]}
   );
   gpc1_1 gpc7185 (
      {stage1_64[88]},
      {stage2_64[106]}
   );
   gpc1_1 gpc7186 (
      {stage1_64[89]},
      {stage2_64[107]}
   );
   gpc1_1 gpc7187 (
      {stage1_64[90]},
      {stage2_64[108]}
   );
   gpc1_1 gpc7188 (
      {stage1_64[91]},
      {stage2_64[109]}
   );
   gpc1_1 gpc7189 (
      {stage1_64[92]},
      {stage2_64[110]}
   );
   gpc1_1 gpc7190 (
      {stage1_64[93]},
      {stage2_64[111]}
   );
   gpc1_1 gpc7191 (
      {stage1_64[94]},
      {stage2_64[112]}
   );
   gpc1_1 gpc7192 (
      {stage1_64[95]},
      {stage2_64[113]}
   );
   gpc1_1 gpc7193 (
      {stage1_64[96]},
      {stage2_64[114]}
   );
   gpc1_1 gpc7194 (
      {stage1_64[97]},
      {stage2_64[115]}
   );
   gpc1_1 gpc7195 (
      {stage1_64[98]},
      {stage2_64[116]}
   );
   gpc1_1 gpc7196 (
      {stage1_64[99]},
      {stage2_64[117]}
   );
   gpc1_1 gpc7197 (
      {stage1_64[100]},
      {stage2_64[118]}
   );
   gpc1_1 gpc7198 (
      {stage1_64[101]},
      {stage2_64[119]}
   );
   gpc1_1 gpc7199 (
      {stage1_64[102]},
      {stage2_64[120]}
   );
   gpc1_1 gpc7200 (
      {stage1_64[103]},
      {stage2_64[121]}
   );
   gpc1_1 gpc7201 (
      {stage1_64[104]},
      {stage2_64[122]}
   );
   gpc1_1 gpc7202 (
      {stage1_64[105]},
      {stage2_64[123]}
   );
   gpc1_1 gpc7203 (
      {stage1_64[106]},
      {stage2_64[124]}
   );
   gpc1_1 gpc7204 (
      {stage1_64[107]},
      {stage2_64[125]}
   );
   gpc1_1 gpc7205 (
      {stage1_64[108]},
      {stage2_64[126]}
   );
   gpc1_1 gpc7206 (
      {stage1_64[109]},
      {stage2_64[127]}
   );
   gpc1_1 gpc7207 (
      {stage1_64[110]},
      {stage2_64[128]}
   );
   gpc1_1 gpc7208 (
      {stage1_64[111]},
      {stage2_64[129]}
   );
   gpc1_1 gpc7209 (
      {stage1_64[112]},
      {stage2_64[130]}
   );
   gpc1_1 gpc7210 (
      {stage1_64[113]},
      {stage2_64[131]}
   );
   gpc1_1 gpc7211 (
      {stage1_64[114]},
      {stage2_64[132]}
   );
   gpc1_1 gpc7212 (
      {stage1_64[115]},
      {stage2_64[133]}
   );
   gpc1_1 gpc7213 (
      {stage1_64[116]},
      {stage2_64[134]}
   );
   gpc1_1 gpc7214 (
      {stage1_64[117]},
      {stage2_64[135]}
   );
   gpc1_1 gpc7215 (
      {stage1_64[118]},
      {stage2_64[136]}
   );
   gpc1_1 gpc7216 (
      {stage1_64[119]},
      {stage2_64[137]}
   );
   gpc1_1 gpc7217 (
      {stage1_64[120]},
      {stage2_64[138]}
   );
   gpc1_1 gpc7218 (
      {stage1_64[121]},
      {stage2_64[139]}
   );
   gpc1_1 gpc7219 (
      {stage1_64[122]},
      {stage2_64[140]}
   );
   gpc1_1 gpc7220 (
      {stage1_64[123]},
      {stage2_64[141]}
   );
   gpc1_1 gpc7221 (
      {stage1_65[49]},
      {stage2_65[51]}
   );
   gpc1_1 gpc7222 (
      {stage1_65[50]},
      {stage2_65[52]}
   );
   gpc1_1 gpc7223 (
      {stage1_65[51]},
      {stage2_65[53]}
   );
   gpc1_1 gpc7224 (
      {stage1_65[52]},
      {stage2_65[54]}
   );
   gpc1_1 gpc7225 (
      {stage1_65[53]},
      {stage2_65[55]}
   );
   gpc1343_5 gpc7226 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3]},
      {stage2_2[0], stage2_2[1], stage2_2[2]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc1343_5 gpc7227 (
      {stage2_0[3], stage2_0[4], stage2_0[5]},
      {stage2_1[4], stage2_1[5], stage2_1[6], stage2_1[7]},
      {stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage2_3[1]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc1343_5 gpc7228 (
      {stage2_0[6], stage2_0[7], stage2_0[8]},
      {stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_2[6], stage2_2[7], stage2_2[8]},
      {stage2_3[2]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc1343_5 gpc7229 (
      {stage2_0[9], stage2_0[10], stage2_0[11]},
      {stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15]},
      {stage2_2[9], stage2_2[10], stage2_2[11]},
      {stage2_3[3]},
      {stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3],stage3_0[3]}
   );
   gpc2135_5 gpc7230 (
      {stage2_0[12], stage2_0[13], stage2_0[14], stage2_0[15], stage2_0[16]},
      {stage2_1[16], stage2_1[17], stage2_1[18]},
      {stage2_2[12]},
      {stage2_3[4], stage2_3[5]},
      {stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4],stage3_0[4]}
   );
   gpc606_5 gpc7231 (
      {stage2_0[17], stage2_0[18], stage2_0[19], stage2_0[20], stage2_0[21], stage2_0[22]},
      {stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17], stage2_2[18]},
      {stage3_4[5],stage3_3[5],stage3_2[5],stage3_1[5],stage3_0[5]}
   );
   gpc606_5 gpc7232 (
      {stage2_1[19], stage2_1[20], stage2_1[21], stage2_1[22], stage2_1[23], stage2_1[24]},
      {stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11]},
      {stage3_5[0],stage3_4[6],stage3_3[6],stage3_2[6],stage3_1[6]}
   );
   gpc606_5 gpc7233 (
      {stage2_1[25], stage2_1[26], stage2_1[27], stage2_1[28], stage2_1[29], stage2_1[30]},
      {stage2_3[12], stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17]},
      {stage3_5[1],stage3_4[7],stage3_3[7],stage3_2[7],stage3_1[7]}
   );
   gpc606_5 gpc7234 (
      {stage2_1[31], stage2_1[32], stage2_1[33], stage2_1[34], stage2_1[35], stage2_1[36]},
      {stage2_3[18], stage2_3[19], stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23]},
      {stage3_5[2],stage3_4[8],stage3_3[8],stage3_2[8],stage3_1[8]}
   );
   gpc615_5 gpc7235 (
      {stage2_1[37], stage2_1[38], stage2_1[39], stage2_1[40], stage2_1[41]},
      {stage2_2[19]},
      {stage2_3[24], stage2_3[25], stage2_3[26], stage2_3[27], stage2_3[28], stage2_3[29]},
      {stage3_5[3],stage3_4[9],stage3_3[9],stage3_2[9],stage3_1[9]}
   );
   gpc606_5 gpc7236 (
      {stage2_2[20], stage2_2[21], stage2_2[22], stage2_2[23], stage2_2[24], stage2_2[25]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[4],stage3_4[10],stage3_3[10],stage3_2[10]}
   );
   gpc606_5 gpc7237 (
      {stage2_2[26], stage2_2[27], stage2_2[28], stage2_2[29], stage2_2[30], stage2_2[31]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[5],stage3_4[11],stage3_3[11],stage3_2[11]}
   );
   gpc615_5 gpc7238 (
      {stage2_3[30], stage2_3[31], stage2_3[32], stage2_3[33], stage2_3[34]},
      {stage2_4[12]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[2],stage3_5[6],stage3_4[12],stage3_3[12]}
   );
   gpc615_5 gpc7239 (
      {stage2_3[35], stage2_3[36], stage2_3[37], stage2_3[38], stage2_3[39]},
      {stage2_4[13]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[3],stage3_5[7],stage3_4[13],stage3_3[13]}
   );
   gpc615_5 gpc7240 (
      {stage2_3[40], stage2_3[41], stage2_3[42], stage2_3[43], stage2_3[44]},
      {stage2_4[14]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[4],stage3_5[8],stage3_4[14],stage3_3[14]}
   );
   gpc615_5 gpc7241 (
      {stage2_3[45], stage2_3[46], stage2_3[47], stage2_3[48], stage2_3[49]},
      {stage2_4[15]},
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage3_7[3],stage3_6[5],stage3_5[9],stage3_4[15],stage3_3[15]}
   );
   gpc615_5 gpc7242 (
      {stage2_3[50], stage2_3[51], stage2_3[52], stage2_3[53], stage2_3[54]},
      {stage2_4[16]},
      {stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29]},
      {stage3_7[4],stage3_6[6],stage3_5[10],stage3_4[16],stage3_3[16]}
   );
   gpc615_5 gpc7243 (
      {stage2_3[55], stage2_3[56], stage2_3[57], stage2_3[58], stage2_3[59]},
      {stage2_4[17]},
      {stage2_5[30], stage2_5[31], stage2_5[32], stage2_5[33], stage2_5[34], stage2_5[35]},
      {stage3_7[5],stage3_6[7],stage3_5[11],stage3_4[17],stage3_3[17]}
   );
   gpc615_5 gpc7244 (
      {stage2_3[60], stage2_3[61], stage2_3[62], stage2_3[63], stage2_3[64]},
      {stage2_4[18]},
      {stage2_5[36], stage2_5[37], stage2_5[38], stage2_5[39], stage2_5[40], stage2_5[41]},
      {stage3_7[6],stage3_6[8],stage3_5[12],stage3_4[18],stage3_3[18]}
   );
   gpc615_5 gpc7245 (
      {stage2_3[65], stage2_3[66], stage2_3[67], stage2_3[68], stage2_3[69]},
      {stage2_4[19]},
      {stage2_5[42], stage2_5[43], stage2_5[44], stage2_5[45], stage2_5[46], stage2_5[47]},
      {stage3_7[7],stage3_6[9],stage3_5[13],stage3_4[19],stage3_3[19]}
   );
   gpc615_5 gpc7246 (
      {stage2_3[70], stage2_3[71], stage2_3[72], stage2_3[73], stage2_3[74]},
      {stage2_4[20]},
      {stage2_5[48], stage2_5[49], stage2_5[50], stage2_5[51], stage2_5[52], stage2_5[53]},
      {stage3_7[8],stage3_6[10],stage3_5[14],stage3_4[20],stage3_3[20]}
   );
   gpc615_5 gpc7247 (
      {stage2_3[75], stage2_3[76], stage2_3[77], stage2_3[78], stage2_3[79]},
      {stage2_4[21]},
      {stage2_5[54], stage2_5[55], stage2_5[56], stage2_5[57], stage2_5[58], stage2_5[59]},
      {stage3_7[9],stage3_6[11],stage3_5[15],stage3_4[21],stage3_3[21]}
   );
   gpc615_5 gpc7248 (
      {stage2_3[80], stage2_3[81], stage2_3[82], stage2_3[83], stage2_3[84]},
      {stage2_4[22]},
      {stage2_5[60], stage2_5[61], stage2_5[62], stage2_5[63], stage2_5[64], stage2_5[65]},
      {stage3_7[10],stage3_6[12],stage3_5[16],stage3_4[22],stage3_3[22]}
   );
   gpc615_5 gpc7249 (
      {stage2_3[85], stage2_3[86], stage2_3[87], stage2_3[88], stage2_3[89]},
      {stage2_4[23]},
      {stage2_5[66], stage2_5[67], stage2_5[68], stage2_5[69], stage2_5[70], stage2_5[71]},
      {stage3_7[11],stage3_6[13],stage3_5[17],stage3_4[23],stage3_3[23]}
   );
   gpc615_5 gpc7250 (
      {stage2_3[90], stage2_3[91], stage2_3[92], stage2_3[93], stage2_3[94]},
      {stage2_4[24]},
      {stage2_5[72], stage2_5[73], stage2_5[74], stage2_5[75], stage2_5[76], stage2_5[77]},
      {stage3_7[12],stage3_6[14],stage3_5[18],stage3_4[24],stage3_3[24]}
   );
   gpc615_5 gpc7251 (
      {stage2_3[95], stage2_3[96], stage2_3[97], stage2_3[98], stage2_3[99]},
      {stage2_4[25]},
      {stage2_5[78], stage2_5[79], stage2_5[80], stage2_5[81], stage2_5[82], stage2_5[83]},
      {stage3_7[13],stage3_6[15],stage3_5[19],stage3_4[25],stage3_3[25]}
   );
   gpc615_5 gpc7252 (
      {stage2_3[100], stage2_3[101], stage2_3[102], stage2_3[103], stage2_3[104]},
      {stage2_4[26]},
      {stage2_5[84], stage2_5[85], stage2_5[86], stage2_5[87], stage2_5[88], stage2_5[89]},
      {stage3_7[14],stage3_6[16],stage3_5[20],stage3_4[26],stage3_3[26]}
   );
   gpc615_5 gpc7253 (
      {stage2_3[105], stage2_3[106], stage2_3[107], stage2_3[108], stage2_3[109]},
      {stage2_4[27]},
      {stage2_5[90], stage2_5[91], stage2_5[92], stage2_5[93], stage2_5[94], stage2_5[95]},
      {stage3_7[15],stage3_6[17],stage3_5[21],stage3_4[27],stage3_3[27]}
   );
   gpc615_5 gpc7254 (
      {stage2_3[110], stage2_3[111], stage2_3[112], stage2_3[113], 1'b0},
      {stage2_4[28]},
      {stage2_5[96], stage2_5[97], stage2_5[98], stage2_5[99], stage2_5[100], stage2_5[101]},
      {stage3_7[16],stage3_6[18],stage3_5[22],stage3_4[28],stage3_3[28]}
   );
   gpc606_5 gpc7255 (
      {stage2_5[102], stage2_5[103], stage2_5[104], stage2_5[105], stage2_5[106], stage2_5[107]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[0],stage3_7[17],stage3_6[19],stage3_5[23]}
   );
   gpc606_5 gpc7256 (
      {stage2_5[108], stage2_5[109], stage2_5[110], stage2_5[111], stage2_5[112], stage2_5[113]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[1],stage3_7[18],stage3_6[20],stage3_5[24]}
   );
   gpc606_5 gpc7257 (
      {stage2_5[114], stage2_5[115], stage2_5[116], stage2_5[117], stage2_5[118], stage2_5[119]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[2],stage3_7[19],stage3_6[21],stage3_5[25]}
   );
   gpc606_5 gpc7258 (
      {stage2_5[120], stage2_5[121], stage2_5[122], stage2_5[123], stage2_5[124], stage2_5[125]},
      {stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage3_9[3],stage3_8[3],stage3_7[20],stage3_6[22],stage3_5[26]}
   );
   gpc606_5 gpc7259 (
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[4],stage3_8[4],stage3_7[21],stage3_6[23]}
   );
   gpc615_5 gpc7260 (
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10]},
      {stage2_7[24]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[5],stage3_8[5],stage3_7[22],stage3_6[24]}
   );
   gpc615_5 gpc7261 (
      {stage2_6[11], stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15]},
      {stage2_7[25]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[6],stage3_8[6],stage3_7[23],stage3_6[25]}
   );
   gpc615_5 gpc7262 (
      {stage2_6[16], stage2_6[17], stage2_6[18], stage2_6[19], stage2_6[20]},
      {stage2_7[26]},
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23]},
      {stage3_10[3],stage3_9[7],stage3_8[7],stage3_7[24],stage3_6[26]}
   );
   gpc615_5 gpc7263 (
      {stage2_6[21], stage2_6[22], stage2_6[23], stage2_6[24], stage2_6[25]},
      {stage2_7[27]},
      {stage2_8[24], stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29]},
      {stage3_10[4],stage3_9[8],stage3_8[8],stage3_7[25],stage3_6[27]}
   );
   gpc615_5 gpc7264 (
      {stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29], stage2_6[30]},
      {stage2_7[28]},
      {stage2_8[30], stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35]},
      {stage3_10[5],stage3_9[9],stage3_8[9],stage3_7[26],stage3_6[28]}
   );
   gpc615_5 gpc7265 (
      {stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage2_7[29]},
      {stage2_8[36], stage2_8[37], stage2_8[38], stage2_8[39], stage2_8[40], stage2_8[41]},
      {stage3_10[6],stage3_9[10],stage3_8[10],stage3_7[27],stage3_6[29]}
   );
   gpc615_5 gpc7266 (
      {stage2_6[36], stage2_6[37], stage2_6[38], stage2_6[39], stage2_6[40]},
      {stage2_7[30]},
      {stage2_8[42], stage2_8[43], stage2_8[44], stage2_8[45], stage2_8[46], stage2_8[47]},
      {stage3_10[7],stage3_9[11],stage3_8[11],stage3_7[28],stage3_6[30]}
   );
   gpc615_5 gpc7267 (
      {stage2_6[41], stage2_6[42], stage2_6[43], stage2_6[44], stage2_6[45]},
      {stage2_7[31]},
      {stage2_8[48], stage2_8[49], stage2_8[50], stage2_8[51], stage2_8[52], stage2_8[53]},
      {stage3_10[8],stage3_9[12],stage3_8[12],stage3_7[29],stage3_6[31]}
   );
   gpc615_5 gpc7268 (
      {stage2_7[32], stage2_7[33], stage2_7[34], stage2_7[35], stage2_7[36]},
      {stage2_8[54]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[9],stage3_9[13],stage3_8[13],stage3_7[30]}
   );
   gpc615_5 gpc7269 (
      {stage2_7[37], stage2_7[38], stage2_7[39], stage2_7[40], stage2_7[41]},
      {stage2_8[55]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[10],stage3_9[14],stage3_8[14],stage3_7[31]}
   );
   gpc615_5 gpc7270 (
      {stage2_7[42], stage2_7[43], stage2_7[44], stage2_7[45], stage2_7[46]},
      {stage2_8[56]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[11],stage3_9[15],stage3_8[15],stage3_7[32]}
   );
   gpc615_5 gpc7271 (
      {stage2_7[47], stage2_7[48], stage2_7[49], stage2_7[50], stage2_7[51]},
      {stage2_8[57]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[12],stage3_9[16],stage3_8[16],stage3_7[33]}
   );
   gpc615_5 gpc7272 (
      {stage2_7[52], stage2_7[53], stage2_7[54], stage2_7[55], stage2_7[56]},
      {stage2_8[58]},
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage3_11[4],stage3_10[13],stage3_9[17],stage3_8[17],stage3_7[34]}
   );
   gpc606_5 gpc7273 (
      {stage2_8[59], stage2_8[60], stage2_8[61], stage2_8[62], stage2_8[63], stage2_8[64]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[5],stage3_10[14],stage3_9[18],stage3_8[18]}
   );
   gpc606_5 gpc7274 (
      {stage2_8[65], stage2_8[66], stage2_8[67], stage2_8[68], stage2_8[69], stage2_8[70]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[6],stage3_10[15],stage3_9[19],stage3_8[19]}
   );
   gpc606_5 gpc7275 (
      {stage2_8[71], stage2_8[72], stage2_8[73], stage2_8[74], stage2_8[75], stage2_8[76]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[7],stage3_10[16],stage3_9[20],stage3_8[20]}
   );
   gpc606_5 gpc7276 (
      {stage2_8[77], stage2_8[78], stage2_8[79], stage2_8[80], stage2_8[81], stage2_8[82]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage3_12[3],stage3_11[8],stage3_10[17],stage3_9[21],stage3_8[21]}
   );
   gpc606_5 gpc7277 (
      {stage2_8[83], stage2_8[84], stage2_8[85], stage2_8[86], stage2_8[87], stage2_8[88]},
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage3_12[4],stage3_11[9],stage3_10[18],stage3_9[22],stage3_8[22]}
   );
   gpc606_5 gpc7278 (
      {stage2_8[89], stage2_8[90], stage2_8[91], stage2_8[92], stage2_8[93], stage2_8[94]},
      {stage2_10[30], stage2_10[31], stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35]},
      {stage3_12[5],stage3_11[10],stage3_10[19],stage3_9[23],stage3_8[23]}
   );
   gpc606_5 gpc7279 (
      {stage2_8[95], stage2_8[96], stage2_8[97], stage2_8[98], stage2_8[99], stage2_8[100]},
      {stage2_10[36], stage2_10[37], stage2_10[38], stage2_10[39], stage2_10[40], stage2_10[41]},
      {stage3_12[6],stage3_11[11],stage3_10[20],stage3_9[24],stage3_8[24]}
   );
   gpc606_5 gpc7280 (
      {stage2_8[101], stage2_8[102], stage2_8[103], stage2_8[104], stage2_8[105], stage2_8[106]},
      {stage2_10[42], stage2_10[43], stage2_10[44], stage2_10[45], stage2_10[46], stage2_10[47]},
      {stage3_12[7],stage3_11[12],stage3_10[21],stage3_9[25],stage3_8[25]}
   );
   gpc606_5 gpc7281 (
      {stage2_8[107], stage2_8[108], stage2_8[109], stage2_8[110], stage2_8[111], stage2_8[112]},
      {stage2_10[48], stage2_10[49], stage2_10[50], stage2_10[51], stage2_10[52], stage2_10[53]},
      {stage3_12[8],stage3_11[13],stage3_10[22],stage3_9[26],stage3_8[26]}
   );
   gpc606_5 gpc7282 (
      {stage2_8[113], stage2_8[114], stage2_8[115], stage2_8[116], stage2_8[117], stage2_8[118]},
      {stage2_10[54], stage2_10[55], stage2_10[56], stage2_10[57], stage2_10[58], stage2_10[59]},
      {stage3_12[9],stage3_11[14],stage3_10[23],stage3_9[27],stage3_8[27]}
   );
   gpc606_5 gpc7283 (
      {stage2_8[119], stage2_8[120], stage2_8[121], stage2_8[122], stage2_8[123], stage2_8[124]},
      {stage2_10[60], stage2_10[61], stage2_10[62], stage2_10[63], stage2_10[64], stage2_10[65]},
      {stage3_12[10],stage3_11[15],stage3_10[24],stage3_9[28],stage3_8[28]}
   );
   gpc606_5 gpc7284 (
      {stage2_8[125], stage2_8[126], stage2_8[127], stage2_8[128], stage2_8[129], stage2_8[130]},
      {stage2_10[66], stage2_10[67], stage2_10[68], stage2_10[69], stage2_10[70], stage2_10[71]},
      {stage3_12[11],stage3_11[16],stage3_10[25],stage3_9[29],stage3_8[29]}
   );
   gpc606_5 gpc7285 (
      {stage2_8[131], stage2_8[132], stage2_8[133], stage2_8[134], stage2_8[135], stage2_8[136]},
      {stage2_10[72], stage2_10[73], stage2_10[74], stage2_10[75], stage2_10[76], stage2_10[77]},
      {stage3_12[12],stage3_11[17],stage3_10[26],stage3_9[30],stage3_8[30]}
   );
   gpc606_5 gpc7286 (
      {stage2_8[137], stage2_8[138], stage2_8[139], stage2_8[140], stage2_8[141], stage2_8[142]},
      {stage2_10[78], stage2_10[79], stage2_10[80], stage2_10[81], stage2_10[82], stage2_10[83]},
      {stage3_12[13],stage3_11[18],stage3_10[27],stage3_9[31],stage3_8[31]}
   );
   gpc606_5 gpc7287 (
      {stage2_8[143], stage2_8[144], stage2_8[145], stage2_8[146], stage2_8[147], stage2_8[148]},
      {stage2_10[84], stage2_10[85], stage2_10[86], stage2_10[87], stage2_10[88], stage2_10[89]},
      {stage3_12[14],stage3_11[19],stage3_10[28],stage3_9[32],stage3_8[32]}
   );
   gpc606_5 gpc7288 (
      {stage2_8[149], stage2_8[150], stage2_8[151], stage2_8[152], stage2_8[153], stage2_8[154]},
      {stage2_10[90], stage2_10[91], stage2_10[92], stage2_10[93], stage2_10[94], stage2_10[95]},
      {stage3_12[15],stage3_11[20],stage3_10[29],stage3_9[33],stage3_8[33]}
   );
   gpc606_5 gpc7289 (
      {stage2_8[155], stage2_8[156], stage2_8[157], stage2_8[158], stage2_8[159], 1'b0},
      {stage2_10[96], stage2_10[97], stage2_10[98], stage2_10[99], stage2_10[100], stage2_10[101]},
      {stage3_12[16],stage3_11[21],stage3_10[30],stage3_9[34],stage3_8[34]}
   );
   gpc606_5 gpc7290 (
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[17],stage3_11[22],stage3_10[31],stage3_9[35]}
   );
   gpc606_5 gpc7291 (
      {stage2_9[36], stage2_9[37], stage2_9[38], stage2_9[39], stage2_9[40], stage2_9[41]},
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage3_13[1],stage3_12[18],stage3_11[23],stage3_10[32],stage3_9[36]}
   );
   gpc606_5 gpc7292 (
      {stage2_9[42], stage2_9[43], stage2_9[44], stage2_9[45], stage2_9[46], stage2_9[47]},
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17]},
      {stage3_13[2],stage3_12[19],stage3_11[24],stage3_10[33],stage3_9[37]}
   );
   gpc606_5 gpc7293 (
      {stage2_9[48], stage2_9[49], stage2_9[50], stage2_9[51], stage2_9[52], stage2_9[53]},
      {stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23]},
      {stage3_13[3],stage3_12[20],stage3_11[25],stage3_10[34],stage3_9[38]}
   );
   gpc606_5 gpc7294 (
      {stage2_9[54], stage2_9[55], stage2_9[56], stage2_9[57], stage2_9[58], stage2_9[59]},
      {stage2_11[24], stage2_11[25], stage2_11[26], stage2_11[27], stage2_11[28], stage2_11[29]},
      {stage3_13[4],stage3_12[21],stage3_11[26],stage3_10[35],stage3_9[39]}
   );
   gpc606_5 gpc7295 (
      {stage2_9[60], stage2_9[61], stage2_9[62], stage2_9[63], stage2_9[64], stage2_9[65]},
      {stage2_11[30], stage2_11[31], stage2_11[32], stage2_11[33], stage2_11[34], stage2_11[35]},
      {stage3_13[5],stage3_12[22],stage3_11[27],stage3_10[36],stage3_9[40]}
   );
   gpc606_5 gpc7296 (
      {stage2_9[66], stage2_9[67], stage2_9[68], stage2_9[69], stage2_9[70], stage2_9[71]},
      {stage2_11[36], stage2_11[37], stage2_11[38], stage2_11[39], stage2_11[40], stage2_11[41]},
      {stage3_13[6],stage3_12[23],stage3_11[28],stage3_10[37],stage3_9[41]}
   );
   gpc606_5 gpc7297 (
      {stage2_9[72], stage2_9[73], stage2_9[74], stage2_9[75], stage2_9[76], stage2_9[77]},
      {stage2_11[42], stage2_11[43], stage2_11[44], stage2_11[45], stage2_11[46], stage2_11[47]},
      {stage3_13[7],stage3_12[24],stage3_11[29],stage3_10[38],stage3_9[42]}
   );
   gpc606_5 gpc7298 (
      {stage2_9[78], stage2_9[79], stage2_9[80], stage2_9[81], stage2_9[82], stage2_9[83]},
      {stage2_11[48], stage2_11[49], stage2_11[50], stage2_11[51], stage2_11[52], stage2_11[53]},
      {stage3_13[8],stage3_12[25],stage3_11[30],stage3_10[39],stage3_9[43]}
   );
   gpc606_5 gpc7299 (
      {stage2_9[84], stage2_9[85], stage2_9[86], stage2_9[87], stage2_9[88], stage2_9[89]},
      {stage2_11[54], stage2_11[55], stage2_11[56], stage2_11[57], stage2_11[58], stage2_11[59]},
      {stage3_13[9],stage3_12[26],stage3_11[31],stage3_10[40],stage3_9[44]}
   );
   gpc606_5 gpc7300 (
      {stage2_9[90], stage2_9[91], stage2_9[92], stage2_9[93], stage2_9[94], stage2_9[95]},
      {stage2_11[60], stage2_11[61], stage2_11[62], stage2_11[63], stage2_11[64], stage2_11[65]},
      {stage3_13[10],stage3_12[27],stage3_11[32],stage3_10[41],stage3_9[45]}
   );
   gpc606_5 gpc7301 (
      {stage2_9[96], stage2_9[97], stage2_9[98], stage2_9[99], stage2_9[100], stage2_9[101]},
      {stage2_11[66], stage2_11[67], stage2_11[68], stage2_11[69], stage2_11[70], stage2_11[71]},
      {stage3_13[11],stage3_12[28],stage3_11[33],stage3_10[42],stage3_9[46]}
   );
   gpc606_5 gpc7302 (
      {stage2_9[102], stage2_9[103], stage2_9[104], stage2_9[105], stage2_9[106], stage2_9[107]},
      {stage2_11[72], stage2_11[73], stage2_11[74], stage2_11[75], stage2_11[76], stage2_11[77]},
      {stage3_13[12],stage3_12[29],stage3_11[34],stage3_10[43],stage3_9[47]}
   );
   gpc606_5 gpc7303 (
      {stage2_9[108], stage2_9[109], stage2_9[110], stage2_9[111], stage2_9[112], stage2_9[113]},
      {stage2_11[78], stage2_11[79], stage2_11[80], stage2_11[81], stage2_11[82], stage2_11[83]},
      {stage3_13[13],stage3_12[30],stage3_11[35],stage3_10[44],stage3_9[48]}
   );
   gpc606_5 gpc7304 (
      {stage2_9[114], stage2_9[115], stage2_9[116], stage2_9[117], stage2_9[118], stage2_9[119]},
      {stage2_11[84], stage2_11[85], stage2_11[86], stage2_11[87], stage2_11[88], stage2_11[89]},
      {stage3_13[14],stage3_12[31],stage3_11[36],stage3_10[45],stage3_9[49]}
   );
   gpc606_5 gpc7305 (
      {stage2_9[120], stage2_9[121], stage2_9[122], stage2_9[123], stage2_9[124], stage2_9[125]},
      {stage2_11[90], stage2_11[91], stage2_11[92], stage2_11[93], stage2_11[94], stage2_11[95]},
      {stage3_13[15],stage3_12[32],stage3_11[37],stage3_10[46],stage3_9[50]}
   );
   gpc606_5 gpc7306 (
      {stage2_9[126], stage2_9[127], stage2_9[128], stage2_9[129], stage2_9[130], stage2_9[131]},
      {stage2_11[96], stage2_11[97], stage2_11[98], stage2_11[99], stage2_11[100], stage2_11[101]},
      {stage3_13[16],stage3_12[33],stage3_11[38],stage3_10[47],stage3_9[51]}
   );
   gpc606_5 gpc7307 (
      {stage2_9[132], stage2_9[133], stage2_9[134], stage2_9[135], stage2_9[136], stage2_9[137]},
      {stage2_11[102], stage2_11[103], stage2_11[104], stage2_11[105], stage2_11[106], stage2_11[107]},
      {stage3_13[17],stage3_12[34],stage3_11[39],stage3_10[48],stage3_9[52]}
   );
   gpc606_5 gpc7308 (
      {stage2_9[138], stage2_9[139], stage2_9[140], stage2_9[141], stage2_9[142], 1'b0},
      {stage2_11[108], stage2_11[109], stage2_11[110], stage2_11[111], stage2_11[112], stage2_11[113]},
      {stage3_13[18],stage3_12[35],stage3_11[40],stage3_10[49],stage3_9[53]}
   );
   gpc615_5 gpc7309 (
      {stage2_10[102], stage2_10[103], stage2_10[104], stage2_10[105], stage2_10[106]},
      {stage2_11[114]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[19],stage3_12[36],stage3_11[41],stage3_10[50]}
   );
   gpc615_5 gpc7310 (
      {stage2_10[107], stage2_10[108], stage2_10[109], stage2_10[110], stage2_10[111]},
      {stage2_11[115]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[20],stage3_12[37],stage3_11[42],stage3_10[51]}
   );
   gpc615_5 gpc7311 (
      {stage2_10[112], stage2_10[113], stage2_10[114], stage2_10[115], stage2_10[116]},
      {stage2_11[116]},
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage3_14[2],stage3_13[21],stage3_12[38],stage3_11[43],stage3_10[52]}
   );
   gpc615_5 gpc7312 (
      {stage2_11[117], stage2_11[118], stage2_11[119], stage2_11[120], stage2_11[121]},
      {stage2_12[18]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[3],stage3_13[22],stage3_12[39],stage3_11[44]}
   );
   gpc615_5 gpc7313 (
      {stage2_11[122], stage2_11[123], stage2_11[124], stage2_11[125], stage2_11[126]},
      {stage2_12[19]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[4],stage3_13[23],stage3_12[40],stage3_11[45]}
   );
   gpc606_5 gpc7314 (
      {stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23], stage2_12[24], stage2_12[25]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[2],stage3_14[5],stage3_13[24],stage3_12[41]}
   );
   gpc606_5 gpc7315 (
      {stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29], stage2_12[30], stage2_12[31]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[3],stage3_14[6],stage3_13[25],stage3_12[42]}
   );
   gpc606_5 gpc7316 (
      {stage2_12[32], stage2_12[33], stage2_12[34], stage2_12[35], stage2_12[36], stage2_12[37]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[4],stage3_14[7],stage3_13[26],stage3_12[43]}
   );
   gpc606_5 gpc7317 (
      {stage2_12[38], stage2_12[39], stage2_12[40], stage2_12[41], stage2_12[42], stage2_12[43]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[5],stage3_14[8],stage3_13[27],stage3_12[44]}
   );
   gpc606_5 gpc7318 (
      {stage2_12[44], stage2_12[45], stage2_12[46], stage2_12[47], stage2_12[48], stage2_12[49]},
      {stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29]},
      {stage3_16[4],stage3_15[6],stage3_14[9],stage3_13[28],stage3_12[45]}
   );
   gpc606_5 gpc7319 (
      {stage2_12[50], stage2_12[51], stage2_12[52], stage2_12[53], stage2_12[54], stage2_12[55]},
      {stage2_14[30], stage2_14[31], stage2_14[32], stage2_14[33], stage2_14[34], stage2_14[35]},
      {stage3_16[5],stage3_15[7],stage3_14[10],stage3_13[29],stage3_12[46]}
   );
   gpc606_5 gpc7320 (
      {stage2_12[56], stage2_12[57], stage2_12[58], stage2_12[59], stage2_12[60], stage2_12[61]},
      {stage2_14[36], stage2_14[37], stage2_14[38], stage2_14[39], stage2_14[40], stage2_14[41]},
      {stage3_16[6],stage3_15[8],stage3_14[11],stage3_13[30],stage3_12[47]}
   );
   gpc606_5 gpc7321 (
      {stage2_12[62], stage2_12[63], stage2_12[64], stage2_12[65], stage2_12[66], stage2_12[67]},
      {stage2_14[42], stage2_14[43], stage2_14[44], stage2_14[45], stage2_14[46], stage2_14[47]},
      {stage3_16[7],stage3_15[9],stage3_14[12],stage3_13[31],stage3_12[48]}
   );
   gpc606_5 gpc7322 (
      {stage2_12[68], stage2_12[69], stage2_12[70], stage2_12[71], stage2_12[72], stage2_12[73]},
      {stage2_14[48], stage2_14[49], stage2_14[50], stage2_14[51], stage2_14[52], stage2_14[53]},
      {stage3_16[8],stage3_15[10],stage3_14[13],stage3_13[32],stage3_12[49]}
   );
   gpc606_5 gpc7323 (
      {stage2_12[74], stage2_12[75], stage2_12[76], stage2_12[77], stage2_12[78], stage2_12[79]},
      {stage2_14[54], stage2_14[55], stage2_14[56], stage2_14[57], stage2_14[58], stage2_14[59]},
      {stage3_16[9],stage3_15[11],stage3_14[14],stage3_13[33],stage3_12[50]}
   );
   gpc606_5 gpc7324 (
      {stage2_12[80], stage2_12[81], stage2_12[82], stage2_12[83], stage2_12[84], stage2_12[85]},
      {stage2_14[60], stage2_14[61], stage2_14[62], stage2_14[63], stage2_14[64], stage2_14[65]},
      {stage3_16[10],stage3_15[12],stage3_14[15],stage3_13[34],stage3_12[51]}
   );
   gpc606_5 gpc7325 (
      {stage2_12[86], stage2_12[87], stage2_12[88], stage2_12[89], stage2_12[90], stage2_12[91]},
      {stage2_14[66], stage2_14[67], stage2_14[68], stage2_14[69], stage2_14[70], stage2_14[71]},
      {stage3_16[11],stage3_15[13],stage3_14[16],stage3_13[35],stage3_12[52]}
   );
   gpc606_5 gpc7326 (
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[12],stage3_15[14],stage3_14[17],stage3_13[36]}
   );
   gpc606_5 gpc7327 (
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage3_17[1],stage3_16[13],stage3_15[15],stage3_14[18],stage3_13[37]}
   );
   gpc606_5 gpc7328 (
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17]},
      {stage3_17[2],stage3_16[14],stage3_15[16],stage3_14[19],stage3_13[38]}
   );
   gpc606_5 gpc7329 (
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage2_15[18], stage2_15[19], stage2_15[20], stage2_15[21], stage2_15[22], stage2_15[23]},
      {stage3_17[3],stage3_16[15],stage3_15[17],stage3_14[20],stage3_13[39]}
   );
   gpc606_5 gpc7330 (
      {stage2_13[36], stage2_13[37], stage2_13[38], stage2_13[39], stage2_13[40], stage2_13[41]},
      {stage2_15[24], stage2_15[25], stage2_15[26], stage2_15[27], stage2_15[28], stage2_15[29]},
      {stage3_17[4],stage3_16[16],stage3_15[18],stage3_14[21],stage3_13[40]}
   );
   gpc606_5 gpc7331 (
      {stage2_13[42], stage2_13[43], stage2_13[44], stage2_13[45], stage2_13[46], stage2_13[47]},
      {stage2_15[30], stage2_15[31], stage2_15[32], stage2_15[33], stage2_15[34], stage2_15[35]},
      {stage3_17[5],stage3_16[17],stage3_15[19],stage3_14[22],stage3_13[41]}
   );
   gpc606_5 gpc7332 (
      {stage2_13[48], stage2_13[49], stage2_13[50], stage2_13[51], stage2_13[52], stage2_13[53]},
      {stage2_15[36], stage2_15[37], stage2_15[38], stage2_15[39], stage2_15[40], stage2_15[41]},
      {stage3_17[6],stage3_16[18],stage3_15[20],stage3_14[23],stage3_13[42]}
   );
   gpc606_5 gpc7333 (
      {stage2_13[54], stage2_13[55], stage2_13[56], stage2_13[57], stage2_13[58], stage2_13[59]},
      {stage2_15[42], stage2_15[43], stage2_15[44], stage2_15[45], stage2_15[46], stage2_15[47]},
      {stage3_17[7],stage3_16[19],stage3_15[21],stage3_14[24],stage3_13[43]}
   );
   gpc606_5 gpc7334 (
      {stage2_13[60], stage2_13[61], stage2_13[62], stage2_13[63], stage2_13[64], stage2_13[65]},
      {stage2_15[48], stage2_15[49], stage2_15[50], stage2_15[51], stage2_15[52], stage2_15[53]},
      {stage3_17[8],stage3_16[20],stage3_15[22],stage3_14[25],stage3_13[44]}
   );
   gpc606_5 gpc7335 (
      {stage2_14[72], stage2_14[73], stage2_14[74], stage2_14[75], stage2_14[76], stage2_14[77]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[9],stage3_16[21],stage3_15[23],stage3_14[26]}
   );
   gpc606_5 gpc7336 (
      {stage2_14[78], stage2_14[79], stage2_14[80], stage2_14[81], stage2_14[82], stage2_14[83]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[10],stage3_16[22],stage3_15[24],stage3_14[27]}
   );
   gpc606_5 gpc7337 (
      {stage2_14[84], stage2_14[85], stage2_14[86], stage2_14[87], stage2_14[88], stage2_14[89]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[11],stage3_16[23],stage3_15[25],stage3_14[28]}
   );
   gpc606_5 gpc7338 (
      {stage2_14[90], stage2_14[91], stage2_14[92], stage2_14[93], stage2_14[94], stage2_14[95]},
      {stage2_16[18], stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23]},
      {stage3_18[3],stage3_17[12],stage3_16[24],stage3_15[26],stage3_14[29]}
   );
   gpc606_5 gpc7339 (
      {stage2_14[96], stage2_14[97], stage2_14[98], stage2_14[99], stage2_14[100], stage2_14[101]},
      {stage2_16[24], stage2_16[25], stage2_16[26], stage2_16[27], stage2_16[28], stage2_16[29]},
      {stage3_18[4],stage3_17[13],stage3_16[25],stage3_15[27],stage3_14[30]}
   );
   gpc606_5 gpc7340 (
      {stage2_14[102], stage2_14[103], stage2_14[104], stage2_14[105], stage2_14[106], stage2_14[107]},
      {stage2_16[30], stage2_16[31], stage2_16[32], stage2_16[33], stage2_16[34], stage2_16[35]},
      {stage3_18[5],stage3_17[14],stage3_16[26],stage3_15[28],stage3_14[31]}
   );
   gpc207_4 gpc7341 (
      {stage2_15[54], stage2_15[55], stage2_15[56], stage2_15[57], stage2_15[58], stage2_15[59], stage2_15[60]},
      {stage2_17[0], stage2_17[1]},
      {stage3_18[6],stage3_17[15],stage3_16[27],stage3_15[29]}
   );
   gpc207_4 gpc7342 (
      {stage2_15[61], stage2_15[62], stage2_15[63], stage2_15[64], stage2_15[65], stage2_15[66], stage2_15[67]},
      {stage2_17[2], stage2_17[3]},
      {stage3_18[7],stage3_17[16],stage3_16[28],stage3_15[30]}
   );
   gpc615_5 gpc7343 (
      {stage2_15[68], stage2_15[69], stage2_15[70], stage2_15[71], stage2_15[72]},
      {stage2_16[36]},
      {stage2_17[4], stage2_17[5], stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9]},
      {stage3_19[0],stage3_18[8],stage3_17[17],stage3_16[29],stage3_15[31]}
   );
   gpc615_5 gpc7344 (
      {stage2_15[73], stage2_15[74], stage2_15[75], stage2_15[76], stage2_15[77]},
      {stage2_16[37]},
      {stage2_17[10], stage2_17[11], stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15]},
      {stage3_19[1],stage3_18[9],stage3_17[18],stage3_16[30],stage3_15[32]}
   );
   gpc615_5 gpc7345 (
      {stage2_15[78], stage2_15[79], stage2_15[80], stage2_15[81], stage2_15[82]},
      {stage2_16[38]},
      {stage2_17[16], stage2_17[17], stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21]},
      {stage3_19[2],stage3_18[10],stage3_17[19],stage3_16[31],stage3_15[33]}
   );
   gpc615_5 gpc7346 (
      {stage2_15[83], stage2_15[84], stage2_15[85], stage2_15[86], stage2_15[87]},
      {stage2_16[39]},
      {stage2_17[22], stage2_17[23], stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27]},
      {stage3_19[3],stage3_18[11],stage3_17[20],stage3_16[32],stage3_15[34]}
   );
   gpc615_5 gpc7347 (
      {stage2_15[88], stage2_15[89], stage2_15[90], stage2_15[91], stage2_15[92]},
      {stage2_16[40]},
      {stage2_17[28], stage2_17[29], stage2_17[30], stage2_17[31], stage2_17[32], stage2_17[33]},
      {stage3_19[4],stage3_18[12],stage3_17[21],stage3_16[33],stage3_15[35]}
   );
   gpc615_5 gpc7348 (
      {stage2_15[93], stage2_15[94], stage2_15[95], stage2_15[96], stage2_15[97]},
      {stage2_16[41]},
      {stage2_17[34], stage2_17[35], stage2_17[36], stage2_17[37], stage2_17[38], stage2_17[39]},
      {stage3_19[5],stage3_18[13],stage3_17[22],stage3_16[34],stage3_15[36]}
   );
   gpc615_5 gpc7349 (
      {stage2_15[98], stage2_15[99], stage2_15[100], stage2_15[101], stage2_15[102]},
      {stage2_16[42]},
      {stage2_17[40], stage2_17[41], stage2_17[42], stage2_17[43], stage2_17[44], stage2_17[45]},
      {stage3_19[6],stage3_18[14],stage3_17[23],stage3_16[35],stage3_15[37]}
   );
   gpc615_5 gpc7350 (
      {stage2_15[103], stage2_15[104], stage2_15[105], stage2_15[106], stage2_15[107]},
      {stage2_16[43]},
      {stage2_17[46], stage2_17[47], stage2_17[48], stage2_17[49], stage2_17[50], stage2_17[51]},
      {stage3_19[7],stage3_18[15],stage3_17[24],stage3_16[36],stage3_15[38]}
   );
   gpc615_5 gpc7351 (
      {stage2_15[108], stage2_15[109], stage2_15[110], stage2_15[111], stage2_15[112]},
      {stage2_16[44]},
      {stage2_17[52], stage2_17[53], stage2_17[54], stage2_17[55], stage2_17[56], stage2_17[57]},
      {stage3_19[8],stage3_18[16],stage3_17[25],stage3_16[37],stage3_15[39]}
   );
   gpc615_5 gpc7352 (
      {stage2_15[113], stage2_15[114], stage2_15[115], stage2_15[116], stage2_15[117]},
      {stage2_16[45]},
      {stage2_17[58], stage2_17[59], stage2_17[60], stage2_17[61], stage2_17[62], stage2_17[63]},
      {stage3_19[9],stage3_18[17],stage3_17[26],stage3_16[38],stage3_15[40]}
   );
   gpc615_5 gpc7353 (
      {stage2_15[118], stage2_15[119], stage2_15[120], stage2_15[121], stage2_15[122]},
      {stage2_16[46]},
      {stage2_17[64], stage2_17[65], stage2_17[66], stage2_17[67], stage2_17[68], stage2_17[69]},
      {stage3_19[10],stage3_18[18],stage3_17[27],stage3_16[39],stage3_15[41]}
   );
   gpc615_5 gpc7354 (
      {stage2_15[123], stage2_15[124], stage2_15[125], stage2_15[126], stage2_15[127]},
      {stage2_16[47]},
      {stage2_17[70], stage2_17[71], stage2_17[72], stage2_17[73], stage2_17[74], stage2_17[75]},
      {stage3_19[11],stage3_18[19],stage3_17[28],stage3_16[40],stage3_15[42]}
   );
   gpc615_5 gpc7355 (
      {stage2_15[128], stage2_15[129], stage2_15[130], stage2_15[131], stage2_15[132]},
      {stage2_16[48]},
      {stage2_17[76], stage2_17[77], stage2_17[78], stage2_17[79], stage2_17[80], stage2_17[81]},
      {stage3_19[12],stage3_18[20],stage3_17[29],stage3_16[41],stage3_15[43]}
   );
   gpc615_5 gpc7356 (
      {stage2_15[133], stage2_15[134], stage2_15[135], stage2_15[136], stage2_15[137]},
      {stage2_16[49]},
      {stage2_17[82], stage2_17[83], stage2_17[84], stage2_17[85], stage2_17[86], 1'b0},
      {stage3_19[13],stage3_18[21],stage3_17[30],stage3_16[42],stage3_15[44]}
   );
   gpc606_5 gpc7357 (
      {stage2_16[50], stage2_16[51], stage2_16[52], stage2_16[53], stage2_16[54], stage2_16[55]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[14],stage3_18[22],stage3_17[31],stage3_16[43]}
   );
   gpc606_5 gpc7358 (
      {stage2_16[56], stage2_16[57], stage2_16[58], stage2_16[59], stage2_16[60], stage2_16[61]},
      {stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10], stage2_18[11]},
      {stage3_20[1],stage3_19[15],stage3_18[23],stage3_17[32],stage3_16[44]}
   );
   gpc606_5 gpc7359 (
      {stage2_16[62], stage2_16[63], stage2_16[64], stage2_16[65], stage2_16[66], stage2_16[67]},
      {stage2_18[12], stage2_18[13], stage2_18[14], stage2_18[15], stage2_18[16], stage2_18[17]},
      {stage3_20[2],stage3_19[16],stage3_18[24],stage3_17[33],stage3_16[45]}
   );
   gpc606_5 gpc7360 (
      {stage2_16[68], stage2_16[69], stage2_16[70], stage2_16[71], stage2_16[72], stage2_16[73]},
      {stage2_18[18], stage2_18[19], stage2_18[20], stage2_18[21], stage2_18[22], stage2_18[23]},
      {stage3_20[3],stage3_19[17],stage3_18[25],stage3_17[34],stage3_16[46]}
   );
   gpc606_5 gpc7361 (
      {stage2_16[74], stage2_16[75], stage2_16[76], stage2_16[77], stage2_16[78], stage2_16[79]},
      {stage2_18[24], stage2_18[25], stage2_18[26], stage2_18[27], stage2_18[28], stage2_18[29]},
      {stage3_20[4],stage3_19[18],stage3_18[26],stage3_17[35],stage3_16[47]}
   );
   gpc2135_5 gpc7362 (
      {stage2_18[30], stage2_18[31], stage2_18[32], stage2_18[33], stage2_18[34]},
      {stage2_19[0], stage2_19[1], stage2_19[2]},
      {stage2_20[0]},
      {stage2_21[0], stage2_21[1]},
      {stage3_22[0],stage3_21[0],stage3_20[5],stage3_19[19],stage3_18[27]}
   );
   gpc2135_5 gpc7363 (
      {stage2_18[35], stage2_18[36], stage2_18[37], stage2_18[38], stage2_18[39]},
      {stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage2_20[1]},
      {stage2_21[2], stage2_21[3]},
      {stage3_22[1],stage3_21[1],stage3_20[6],stage3_19[20],stage3_18[28]}
   );
   gpc2135_5 gpc7364 (
      {stage2_18[40], stage2_18[41], stage2_18[42], stage2_18[43], stage2_18[44]},
      {stage2_19[6], stage2_19[7], stage2_19[8]},
      {stage2_20[2]},
      {stage2_21[4], stage2_21[5]},
      {stage3_22[2],stage3_21[2],stage3_20[7],stage3_19[21],stage3_18[29]}
   );
   gpc2135_5 gpc7365 (
      {stage2_18[45], stage2_18[46], stage2_18[47], stage2_18[48], stage2_18[49]},
      {stage2_19[9], stage2_19[10], stage2_19[11]},
      {stage2_20[3]},
      {stage2_21[6], stage2_21[7]},
      {stage3_22[3],stage3_21[3],stage3_20[8],stage3_19[22],stage3_18[30]}
   );
   gpc2135_5 gpc7366 (
      {stage2_18[50], stage2_18[51], stage2_18[52], stage2_18[53], stage2_18[54]},
      {stage2_19[12], stage2_19[13], stage2_19[14]},
      {stage2_20[4]},
      {stage2_21[8], stage2_21[9]},
      {stage3_22[4],stage3_21[4],stage3_20[9],stage3_19[23],stage3_18[31]}
   );
   gpc2135_5 gpc7367 (
      {stage2_18[55], stage2_18[56], stage2_18[57], stage2_18[58], stage2_18[59]},
      {stage2_19[15], stage2_19[16], stage2_19[17]},
      {stage2_20[5]},
      {stage2_21[10], stage2_21[11]},
      {stage3_22[5],stage3_21[5],stage3_20[10],stage3_19[24],stage3_18[32]}
   );
   gpc2135_5 gpc7368 (
      {stage2_18[60], stage2_18[61], stage2_18[62], stage2_18[63], stage2_18[64]},
      {stage2_19[18], stage2_19[19], stage2_19[20]},
      {stage2_20[6]},
      {stage2_21[12], stage2_21[13]},
      {stage3_22[6],stage3_21[6],stage3_20[11],stage3_19[25],stage3_18[33]}
   );
   gpc2135_5 gpc7369 (
      {stage2_18[65], stage2_18[66], stage2_18[67], stage2_18[68], stage2_18[69]},
      {stage2_19[21], stage2_19[22], stage2_19[23]},
      {stage2_20[7]},
      {stage2_21[14], stage2_21[15]},
      {stage3_22[7],stage3_21[7],stage3_20[12],stage3_19[26],stage3_18[34]}
   );
   gpc2135_5 gpc7370 (
      {stage2_18[70], stage2_18[71], stage2_18[72], stage2_18[73], stage2_18[74]},
      {stage2_19[24], stage2_19[25], stage2_19[26]},
      {stage2_20[8]},
      {stage2_21[16], stage2_21[17]},
      {stage3_22[8],stage3_21[8],stage3_20[13],stage3_19[27],stage3_18[35]}
   );
   gpc2135_5 gpc7371 (
      {stage2_18[75], stage2_18[76], stage2_18[77], stage2_18[78], stage2_18[79]},
      {stage2_19[27], stage2_19[28], stage2_19[29]},
      {stage2_20[9]},
      {stage2_21[18], stage2_21[19]},
      {stage3_22[9],stage3_21[9],stage3_20[14],stage3_19[28],stage3_18[36]}
   );
   gpc2135_5 gpc7372 (
      {stage2_18[80], stage2_18[81], stage2_18[82], stage2_18[83], stage2_18[84]},
      {stage2_19[30], stage2_19[31], stage2_19[32]},
      {stage2_20[10]},
      {stage2_21[20], stage2_21[21]},
      {stage3_22[10],stage3_21[10],stage3_20[15],stage3_19[29],stage3_18[37]}
   );
   gpc2135_5 gpc7373 (
      {stage2_18[85], stage2_18[86], stage2_18[87], stage2_18[88], stage2_18[89]},
      {stage2_19[33], stage2_19[34], stage2_19[35]},
      {stage2_20[11]},
      {stage2_21[22], stage2_21[23]},
      {stage3_22[11],stage3_21[11],stage3_20[16],stage3_19[30],stage3_18[38]}
   );
   gpc615_5 gpc7374 (
      {stage2_18[90], stage2_18[91], stage2_18[92], stage2_18[93], stage2_18[94]},
      {stage2_19[36]},
      {stage2_20[12], stage2_20[13], stage2_20[14], stage2_20[15], stage2_20[16], stage2_20[17]},
      {stage3_22[12],stage3_21[12],stage3_20[17],stage3_19[31],stage3_18[39]}
   );
   gpc615_5 gpc7375 (
      {stage2_18[95], stage2_18[96], stage2_18[97], stage2_18[98], stage2_18[99]},
      {stage2_19[37]},
      {stage2_20[18], stage2_20[19], stage2_20[20], stage2_20[21], stage2_20[22], stage2_20[23]},
      {stage3_22[13],stage3_21[13],stage3_20[18],stage3_19[32],stage3_18[40]}
   );
   gpc615_5 gpc7376 (
      {stage2_19[38], stage2_19[39], stage2_19[40], stage2_19[41], stage2_19[42]},
      {stage2_20[24]},
      {stage2_21[24], stage2_21[25], stage2_21[26], stage2_21[27], stage2_21[28], stage2_21[29]},
      {stage3_23[0],stage3_22[14],stage3_21[14],stage3_20[19],stage3_19[33]}
   );
   gpc615_5 gpc7377 (
      {stage2_19[43], stage2_19[44], stage2_19[45], stage2_19[46], stage2_19[47]},
      {stage2_20[25]},
      {stage2_21[30], stage2_21[31], stage2_21[32], stage2_21[33], stage2_21[34], stage2_21[35]},
      {stage3_23[1],stage3_22[15],stage3_21[15],stage3_20[20],stage3_19[34]}
   );
   gpc615_5 gpc7378 (
      {stage2_19[48], stage2_19[49], stage2_19[50], stage2_19[51], stage2_19[52]},
      {stage2_20[26]},
      {stage2_21[36], stage2_21[37], stage2_21[38], stage2_21[39], stage2_21[40], stage2_21[41]},
      {stage3_23[2],stage3_22[16],stage3_21[16],stage3_20[21],stage3_19[35]}
   );
   gpc615_5 gpc7379 (
      {stage2_19[53], stage2_19[54], stage2_19[55], stage2_19[56], stage2_19[57]},
      {stage2_20[27]},
      {stage2_21[42], stage2_21[43], stage2_21[44], stage2_21[45], stage2_21[46], stage2_21[47]},
      {stage3_23[3],stage3_22[17],stage3_21[17],stage3_20[22],stage3_19[36]}
   );
   gpc615_5 gpc7380 (
      {stage2_19[58], stage2_19[59], stage2_19[60], stage2_19[61], stage2_19[62]},
      {stage2_20[28]},
      {stage2_21[48], stage2_21[49], stage2_21[50], stage2_21[51], stage2_21[52], stage2_21[53]},
      {stage3_23[4],stage3_22[18],stage3_21[18],stage3_20[23],stage3_19[37]}
   );
   gpc615_5 gpc7381 (
      {stage2_19[63], stage2_19[64], stage2_19[65], stage2_19[66], stage2_19[67]},
      {stage2_20[29]},
      {stage2_21[54], stage2_21[55], stage2_21[56], stage2_21[57], stage2_21[58], stage2_21[59]},
      {stage3_23[5],stage3_22[19],stage3_21[19],stage3_20[24],stage3_19[38]}
   );
   gpc615_5 gpc7382 (
      {stage2_19[68], stage2_19[69], stage2_19[70], stage2_19[71], stage2_19[72]},
      {stage2_20[30]},
      {stage2_21[60], stage2_21[61], stage2_21[62], stage2_21[63], stage2_21[64], stage2_21[65]},
      {stage3_23[6],stage3_22[20],stage3_21[20],stage3_20[25],stage3_19[39]}
   );
   gpc615_5 gpc7383 (
      {stage2_19[73], stage2_19[74], stage2_19[75], stage2_19[76], stage2_19[77]},
      {stage2_20[31]},
      {stage2_21[66], stage2_21[67], stage2_21[68], stage2_21[69], stage2_21[70], stage2_21[71]},
      {stage3_23[7],stage3_22[21],stage3_21[21],stage3_20[26],stage3_19[40]}
   );
   gpc615_5 gpc7384 (
      {stage2_19[78], stage2_19[79], stage2_19[80], stage2_19[81], stage2_19[82]},
      {stage2_20[32]},
      {stage2_21[72], stage2_21[73], stage2_21[74], stage2_21[75], stage2_21[76], stage2_21[77]},
      {stage3_23[8],stage3_22[22],stage3_21[22],stage3_20[27],stage3_19[41]}
   );
   gpc615_5 gpc7385 (
      {stage2_19[83], stage2_19[84], stage2_19[85], stage2_19[86], stage2_19[87]},
      {stage2_20[33]},
      {stage2_21[78], stage2_21[79], stage2_21[80], stage2_21[81], stage2_21[82], stage2_21[83]},
      {stage3_23[9],stage3_22[23],stage3_21[23],stage3_20[28],stage3_19[42]}
   );
   gpc615_5 gpc7386 (
      {stage2_19[88], stage2_19[89], stage2_19[90], stage2_19[91], stage2_19[92]},
      {stage2_20[34]},
      {stage2_21[84], stage2_21[85], stage2_21[86], stage2_21[87], stage2_21[88], stage2_21[89]},
      {stage3_23[10],stage3_22[24],stage3_21[24],stage3_20[29],stage3_19[43]}
   );
   gpc615_5 gpc7387 (
      {stage2_19[93], stage2_19[94], stage2_19[95], stage2_19[96], stage2_19[97]},
      {stage2_20[35]},
      {stage2_21[90], stage2_21[91], stage2_21[92], stage2_21[93], stage2_21[94], stage2_21[95]},
      {stage3_23[11],stage3_22[25],stage3_21[25],stage3_20[30],stage3_19[44]}
   );
   gpc615_5 gpc7388 (
      {stage2_19[98], stage2_19[99], stage2_19[100], stage2_19[101], stage2_19[102]},
      {stage2_20[36]},
      {stage2_21[96], stage2_21[97], stage2_21[98], stage2_21[99], stage2_21[100], stage2_21[101]},
      {stage3_23[12],stage3_22[26],stage3_21[26],stage3_20[31],stage3_19[45]}
   );
   gpc615_5 gpc7389 (
      {stage2_19[103], stage2_19[104], stage2_19[105], stage2_19[106], stage2_19[107]},
      {stage2_20[37]},
      {stage2_21[102], stage2_21[103], stage2_21[104], stage2_21[105], stage2_21[106], stage2_21[107]},
      {stage3_23[13],stage3_22[27],stage3_21[27],stage3_20[32],stage3_19[46]}
   );
   gpc615_5 gpc7390 (
      {stage2_19[108], stage2_19[109], stage2_19[110], stage2_19[111], stage2_19[112]},
      {stage2_20[38]},
      {stage2_21[108], stage2_21[109], stage2_21[110], stage2_21[111], stage2_21[112], stage2_21[113]},
      {stage3_23[14],stage3_22[28],stage3_21[28],stage3_20[33],stage3_19[47]}
   );
   gpc606_5 gpc7391 (
      {stage2_20[39], stage2_20[40], stage2_20[41], stage2_20[42], stage2_20[43], stage2_20[44]},
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage3_24[0],stage3_23[15],stage3_22[29],stage3_21[29],stage3_20[34]}
   );
   gpc606_5 gpc7392 (
      {stage2_21[114], stage2_21[115], stage2_21[116], stage2_21[117], stage2_21[118], stage2_21[119]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[1],stage3_23[16],stage3_22[30],stage3_21[30]}
   );
   gpc606_5 gpc7393 (
      {stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10], stage2_22[11]},
      {stage2_24[0], stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5]},
      {stage3_26[0],stage3_25[1],stage3_24[2],stage3_23[17],stage3_22[31]}
   );
   gpc606_5 gpc7394 (
      {stage2_22[12], stage2_22[13], stage2_22[14], stage2_22[15], stage2_22[16], stage2_22[17]},
      {stage2_24[6], stage2_24[7], stage2_24[8], stage2_24[9], stage2_24[10], stage2_24[11]},
      {stage3_26[1],stage3_25[2],stage3_24[3],stage3_23[18],stage3_22[32]}
   );
   gpc606_5 gpc7395 (
      {stage2_22[18], stage2_22[19], stage2_22[20], stage2_22[21], stage2_22[22], stage2_22[23]},
      {stage2_24[12], stage2_24[13], stage2_24[14], stage2_24[15], stage2_24[16], stage2_24[17]},
      {stage3_26[2],stage3_25[3],stage3_24[4],stage3_23[19],stage3_22[33]}
   );
   gpc606_5 gpc7396 (
      {stage2_22[24], stage2_22[25], stage2_22[26], stage2_22[27], stage2_22[28], stage2_22[29]},
      {stage2_24[18], stage2_24[19], stage2_24[20], stage2_24[21], stage2_24[22], stage2_24[23]},
      {stage3_26[3],stage3_25[4],stage3_24[5],stage3_23[20],stage3_22[34]}
   );
   gpc615_5 gpc7397 (
      {stage2_22[30], stage2_22[31], stage2_22[32], stage2_22[33], stage2_22[34]},
      {stage2_23[6]},
      {stage2_24[24], stage2_24[25], stage2_24[26], stage2_24[27], stage2_24[28], stage2_24[29]},
      {stage3_26[4],stage3_25[5],stage3_24[6],stage3_23[21],stage3_22[35]}
   );
   gpc615_5 gpc7398 (
      {stage2_22[35], stage2_22[36], stage2_22[37], stage2_22[38], stage2_22[39]},
      {stage2_23[7]},
      {stage2_24[30], stage2_24[31], stage2_24[32], stage2_24[33], stage2_24[34], stage2_24[35]},
      {stage3_26[5],stage3_25[6],stage3_24[7],stage3_23[22],stage3_22[36]}
   );
   gpc615_5 gpc7399 (
      {stage2_22[40], stage2_22[41], stage2_22[42], stage2_22[43], stage2_22[44]},
      {stage2_23[8]},
      {stage2_24[36], stage2_24[37], stage2_24[38], stage2_24[39], stage2_24[40], stage2_24[41]},
      {stage3_26[6],stage3_25[7],stage3_24[8],stage3_23[23],stage3_22[37]}
   );
   gpc615_5 gpc7400 (
      {stage2_22[45], stage2_22[46], stage2_22[47], stage2_22[48], stage2_22[49]},
      {stage2_23[9]},
      {stage2_24[42], stage2_24[43], stage2_24[44], stage2_24[45], stage2_24[46], stage2_24[47]},
      {stage3_26[7],stage3_25[8],stage3_24[9],stage3_23[24],stage3_22[38]}
   );
   gpc615_5 gpc7401 (
      {stage2_22[50], stage2_22[51], stage2_22[52], stage2_22[53], stage2_22[54]},
      {stage2_23[10]},
      {stage2_24[48], stage2_24[49], stage2_24[50], stage2_24[51], stage2_24[52], stage2_24[53]},
      {stage3_26[8],stage3_25[9],stage3_24[10],stage3_23[25],stage3_22[39]}
   );
   gpc615_5 gpc7402 (
      {stage2_22[55], stage2_22[56], stage2_22[57], stage2_22[58], stage2_22[59]},
      {stage2_23[11]},
      {stage2_24[54], stage2_24[55], stage2_24[56], stage2_24[57], stage2_24[58], stage2_24[59]},
      {stage3_26[9],stage3_25[10],stage3_24[11],stage3_23[26],stage3_22[40]}
   );
   gpc615_5 gpc7403 (
      {stage2_22[60], stage2_22[61], stage2_22[62], stage2_22[63], stage2_22[64]},
      {stage2_23[12]},
      {stage2_24[60], stage2_24[61], stage2_24[62], stage2_24[63], stage2_24[64], stage2_24[65]},
      {stage3_26[10],stage3_25[11],stage3_24[12],stage3_23[27],stage3_22[41]}
   );
   gpc615_5 gpc7404 (
      {stage2_22[65], stage2_22[66], stage2_22[67], stage2_22[68], stage2_22[69]},
      {stage2_23[13]},
      {stage2_24[66], stage2_24[67], stage2_24[68], stage2_24[69], stage2_24[70], stage2_24[71]},
      {stage3_26[11],stage3_25[12],stage3_24[13],stage3_23[28],stage3_22[42]}
   );
   gpc615_5 gpc7405 (
      {stage2_22[70], stage2_22[71], stage2_22[72], stage2_22[73], stage2_22[74]},
      {stage2_23[14]},
      {stage2_24[72], stage2_24[73], stage2_24[74], stage2_24[75], stage2_24[76], stage2_24[77]},
      {stage3_26[12],stage3_25[13],stage3_24[14],stage3_23[29],stage3_22[43]}
   );
   gpc615_5 gpc7406 (
      {stage2_22[75], stage2_22[76], stage2_22[77], stage2_22[78], stage2_22[79]},
      {stage2_23[15]},
      {stage2_24[78], stage2_24[79], stage2_24[80], stage2_24[81], stage2_24[82], stage2_24[83]},
      {stage3_26[13],stage3_25[14],stage3_24[15],stage3_23[30],stage3_22[44]}
   );
   gpc2116_5 gpc7407 (
      {stage2_23[16], stage2_23[17], stage2_23[18], stage2_23[19], stage2_23[20], stage2_23[21]},
      {stage2_24[84]},
      {stage2_25[0]},
      {stage2_26[0], stage2_26[1]},
      {stage3_27[0],stage3_26[14],stage3_25[15],stage3_24[16],stage3_23[31]}
   );
   gpc615_5 gpc7408 (
      {stage2_23[22], stage2_23[23], stage2_23[24], stage2_23[25], stage2_23[26]},
      {stage2_24[85]},
      {stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5], stage2_25[6]},
      {stage3_27[1],stage3_26[15],stage3_25[16],stage3_24[17],stage3_23[32]}
   );
   gpc615_5 gpc7409 (
      {stage2_23[27], stage2_23[28], stage2_23[29], stage2_23[30], stage2_23[31]},
      {stage2_24[86]},
      {stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11], stage2_25[12]},
      {stage3_27[2],stage3_26[16],stage3_25[17],stage3_24[18],stage3_23[33]}
   );
   gpc615_5 gpc7410 (
      {stage2_23[32], stage2_23[33], stage2_23[34], stage2_23[35], stage2_23[36]},
      {stage2_24[87]},
      {stage2_25[13], stage2_25[14], stage2_25[15], stage2_25[16], stage2_25[17], stage2_25[18]},
      {stage3_27[3],stage3_26[17],stage3_25[18],stage3_24[19],stage3_23[34]}
   );
   gpc615_5 gpc7411 (
      {stage2_23[37], stage2_23[38], stage2_23[39], stage2_23[40], stage2_23[41]},
      {stage2_24[88]},
      {stage2_25[19], stage2_25[20], stage2_25[21], stage2_25[22], stage2_25[23], stage2_25[24]},
      {stage3_27[4],stage3_26[18],stage3_25[19],stage3_24[20],stage3_23[35]}
   );
   gpc615_5 gpc7412 (
      {stage2_23[42], stage2_23[43], stage2_23[44], stage2_23[45], stage2_23[46]},
      {stage2_24[89]},
      {stage2_25[25], stage2_25[26], stage2_25[27], stage2_25[28], stage2_25[29], stage2_25[30]},
      {stage3_27[5],stage3_26[19],stage3_25[20],stage3_24[21],stage3_23[36]}
   );
   gpc615_5 gpc7413 (
      {stage2_23[47], stage2_23[48], stage2_23[49], stage2_23[50], stage2_23[51]},
      {stage2_24[90]},
      {stage2_25[31], stage2_25[32], stage2_25[33], stage2_25[34], stage2_25[35], stage2_25[36]},
      {stage3_27[6],stage3_26[20],stage3_25[21],stage3_24[22],stage3_23[37]}
   );
   gpc615_5 gpc7414 (
      {stage2_23[52], stage2_23[53], stage2_23[54], stage2_23[55], stage2_23[56]},
      {stage2_24[91]},
      {stage2_25[37], stage2_25[38], stage2_25[39], stage2_25[40], stage2_25[41], stage2_25[42]},
      {stage3_27[7],stage3_26[21],stage3_25[22],stage3_24[23],stage3_23[38]}
   );
   gpc615_5 gpc7415 (
      {stage2_23[57], stage2_23[58], stage2_23[59], stage2_23[60], stage2_23[61]},
      {stage2_24[92]},
      {stage2_25[43], stage2_25[44], stage2_25[45], stage2_25[46], stage2_25[47], stage2_25[48]},
      {stage3_27[8],stage3_26[22],stage3_25[23],stage3_24[24],stage3_23[39]}
   );
   gpc615_5 gpc7416 (
      {stage2_23[62], stage2_23[63], stage2_23[64], stage2_23[65], stage2_23[66]},
      {stage2_24[93]},
      {stage2_25[49], stage2_25[50], stage2_25[51], stage2_25[52], stage2_25[53], stage2_25[54]},
      {stage3_27[9],stage3_26[23],stage3_25[24],stage3_24[25],stage3_23[40]}
   );
   gpc615_5 gpc7417 (
      {stage2_23[67], stage2_23[68], stage2_23[69], stage2_23[70], stage2_23[71]},
      {stage2_24[94]},
      {stage2_25[55], stage2_25[56], stage2_25[57], stage2_25[58], stage2_25[59], stage2_25[60]},
      {stage3_27[10],stage3_26[24],stage3_25[25],stage3_24[26],stage3_23[41]}
   );
   gpc615_5 gpc7418 (
      {stage2_23[72], stage2_23[73], stage2_23[74], stage2_23[75], 1'b0},
      {stage2_24[95]},
      {stage2_25[61], stage2_25[62], stage2_25[63], stage2_25[64], stage2_25[65], stage2_25[66]},
      {stage3_27[11],stage3_26[25],stage3_25[26],stage3_24[27],stage3_23[42]}
   );
   gpc606_5 gpc7419 (
      {stage2_24[96], stage2_24[97], stage2_24[98], stage2_24[99], stage2_24[100], stage2_24[101]},
      {stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5], stage2_26[6], stage2_26[7]},
      {stage3_28[0],stage3_27[12],stage3_26[26],stage3_25[27],stage3_24[28]}
   );
   gpc606_5 gpc7420 (
      {stage2_25[67], stage2_25[68], stage2_25[69], stage2_25[70], stage2_25[71], stage2_25[72]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage3_29[0],stage3_28[1],stage3_27[13],stage3_26[27],stage3_25[28]}
   );
   gpc606_5 gpc7421 (
      {stage2_25[73], stage2_25[74], stage2_25[75], stage2_25[76], stage2_25[77], stage2_25[78]},
      {stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11]},
      {stage3_29[1],stage3_28[2],stage3_27[14],stage3_26[28],stage3_25[29]}
   );
   gpc606_5 gpc7422 (
      {stage2_25[79], stage2_25[80], stage2_25[81], stage2_25[82], stage2_25[83], stage2_25[84]},
      {stage2_27[12], stage2_27[13], stage2_27[14], stage2_27[15], stage2_27[16], stage2_27[17]},
      {stage3_29[2],stage3_28[3],stage3_27[15],stage3_26[29],stage3_25[30]}
   );
   gpc606_5 gpc7423 (
      {stage2_25[85], stage2_25[86], stage2_25[87], stage2_25[88], stage2_25[89], stage2_25[90]},
      {stage2_27[18], stage2_27[19], stage2_27[20], stage2_27[21], stage2_27[22], stage2_27[23]},
      {stage3_29[3],stage3_28[4],stage3_27[16],stage3_26[30],stage3_25[31]}
   );
   gpc606_5 gpc7424 (
      {stage2_25[91], stage2_25[92], stage2_25[93], stage2_25[94], stage2_25[95], 1'b0},
      {stage2_27[24], stage2_27[25], stage2_27[26], stage2_27[27], stage2_27[28], stage2_27[29]},
      {stage3_29[4],stage3_28[5],stage3_27[17],stage3_26[31],stage3_25[32]}
   );
   gpc135_4 gpc7425 (
      {stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11], stage2_26[12]},
      {stage2_27[30], stage2_27[31], stage2_27[32]},
      {stage2_28[0]},
      {stage3_29[5],stage3_28[6],stage3_27[18],stage3_26[32]}
   );
   gpc135_4 gpc7426 (
      {stage2_26[13], stage2_26[14], stage2_26[15], stage2_26[16], stage2_26[17]},
      {stage2_27[33], stage2_27[34], stage2_27[35]},
      {stage2_28[1]},
      {stage3_29[6],stage3_28[7],stage3_27[19],stage3_26[33]}
   );
   gpc135_4 gpc7427 (
      {stage2_26[18], stage2_26[19], stage2_26[20], stage2_26[21], stage2_26[22]},
      {stage2_27[36], stage2_27[37], stage2_27[38]},
      {stage2_28[2]},
      {stage3_29[7],stage3_28[8],stage3_27[20],stage3_26[34]}
   );
   gpc135_4 gpc7428 (
      {stage2_26[23], stage2_26[24], stage2_26[25], stage2_26[26], stage2_26[27]},
      {stage2_27[39], stage2_27[40], stage2_27[41]},
      {stage2_28[3]},
      {stage3_29[8],stage3_28[9],stage3_27[21],stage3_26[35]}
   );
   gpc135_4 gpc7429 (
      {stage2_26[28], stage2_26[29], stage2_26[30], stage2_26[31], stage2_26[32]},
      {stage2_27[42], stage2_27[43], stage2_27[44]},
      {stage2_28[4]},
      {stage3_29[9],stage3_28[10],stage3_27[22],stage3_26[36]}
   );
   gpc135_4 gpc7430 (
      {stage2_26[33], stage2_26[34], stage2_26[35], stage2_26[36], stage2_26[37]},
      {stage2_27[45], stage2_27[46], stage2_27[47]},
      {stage2_28[5]},
      {stage3_29[10],stage3_28[11],stage3_27[23],stage3_26[37]}
   );
   gpc135_4 gpc7431 (
      {stage2_26[38], stage2_26[39], stage2_26[40], stage2_26[41], stage2_26[42]},
      {stage2_27[48], stage2_27[49], stage2_27[50]},
      {stage2_28[6]},
      {stage3_29[11],stage3_28[12],stage3_27[24],stage3_26[38]}
   );
   gpc135_4 gpc7432 (
      {stage2_26[43], stage2_26[44], stage2_26[45], stage2_26[46], stage2_26[47]},
      {stage2_27[51], stage2_27[52], stage2_27[53]},
      {stage2_28[7]},
      {stage3_29[12],stage3_28[13],stage3_27[25],stage3_26[39]}
   );
   gpc135_4 gpc7433 (
      {stage2_26[48], stage2_26[49], stage2_26[50], stage2_26[51], stage2_26[52]},
      {stage2_27[54], stage2_27[55], stage2_27[56]},
      {stage2_28[8]},
      {stage3_29[13],stage3_28[14],stage3_27[26],stage3_26[40]}
   );
   gpc135_4 gpc7434 (
      {stage2_26[53], stage2_26[54], stage2_26[55], stage2_26[56], stage2_26[57]},
      {stage2_27[57], stage2_27[58], stage2_27[59]},
      {stage2_28[9]},
      {stage3_29[14],stage3_28[15],stage3_27[27],stage3_26[41]}
   );
   gpc135_4 gpc7435 (
      {stage2_26[58], stage2_26[59], stage2_26[60], stage2_26[61], stage2_26[62]},
      {stage2_27[60], stage2_27[61], stage2_27[62]},
      {stage2_28[10]},
      {stage3_29[15],stage3_28[16],stage3_27[28],stage3_26[42]}
   );
   gpc135_4 gpc7436 (
      {stage2_26[63], stage2_26[64], stage2_26[65], stage2_26[66], stage2_26[67]},
      {stage2_27[63], stage2_27[64], stage2_27[65]},
      {stage2_28[11]},
      {stage3_29[16],stage3_28[17],stage3_27[29],stage3_26[43]}
   );
   gpc135_4 gpc7437 (
      {stage2_26[68], stage2_26[69], stage2_26[70], stage2_26[71], stage2_26[72]},
      {stage2_27[66], stage2_27[67], stage2_27[68]},
      {stage2_28[12]},
      {stage3_29[17],stage3_28[18],stage3_27[30],stage3_26[44]}
   );
   gpc1343_5 gpc7438 (
      {stage2_26[73], stage2_26[74], stage2_26[75]},
      {stage2_27[69], stage2_27[70], stage2_27[71], stage2_27[72]},
      {stage2_28[13], stage2_28[14], stage2_28[15]},
      {stage2_29[0]},
      {stage3_30[0],stage3_29[18],stage3_28[19],stage3_27[31],stage3_26[45]}
   );
   gpc117_4 gpc7439 (
      {stage2_26[76], stage2_26[77], stage2_26[78], stage2_26[79], stage2_26[80], stage2_26[81], stage2_26[82]},
      {stage2_27[73]},
      {stage2_28[16]},
      {stage3_29[19],stage3_28[20],stage3_27[32],stage3_26[46]}
   );
   gpc7_3 gpc7440 (
      {stage2_27[74], stage2_27[75], stage2_27[76], stage2_27[77], stage2_27[78], stage2_27[79], stage2_27[80]},
      {stage3_29[20],stage3_28[21],stage3_27[33]}
   );
   gpc7_3 gpc7441 (
      {stage2_27[81], stage2_27[82], stage2_27[83], stage2_27[84], stage2_27[85], stage2_27[86], stage2_27[87]},
      {stage3_29[21],stage3_28[22],stage3_27[34]}
   );
   gpc615_5 gpc7442 (
      {stage2_27[88], stage2_27[89], stage2_27[90], stage2_27[91], stage2_27[92]},
      {stage2_28[17]},
      {stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5], stage2_29[6]},
      {stage3_31[0],stage3_30[1],stage3_29[22],stage3_28[23],stage3_27[35]}
   );
   gpc606_5 gpc7443 (
      {stage2_28[18], stage2_28[19], stage2_28[20], stage2_28[21], stage2_28[22], stage2_28[23]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[1],stage3_30[2],stage3_29[23],stage3_28[24]}
   );
   gpc615_5 gpc7444 (
      {stage2_28[24], stage2_28[25], stage2_28[26], stage2_28[27], stage2_28[28]},
      {stage2_29[7]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage3_32[1],stage3_31[2],stage3_30[3],stage3_29[24],stage3_28[25]}
   );
   gpc615_5 gpc7445 (
      {stage2_28[29], stage2_28[30], stage2_28[31], stage2_28[32], stage2_28[33]},
      {stage2_29[8]},
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16], stage2_30[17]},
      {stage3_32[2],stage3_31[3],stage3_30[4],stage3_29[25],stage3_28[26]}
   );
   gpc615_5 gpc7446 (
      {stage2_28[34], stage2_28[35], stage2_28[36], stage2_28[37], stage2_28[38]},
      {stage2_29[9]},
      {stage2_30[18], stage2_30[19], stage2_30[20], stage2_30[21], stage2_30[22], stage2_30[23]},
      {stage3_32[3],stage3_31[4],stage3_30[5],stage3_29[26],stage3_28[27]}
   );
   gpc615_5 gpc7447 (
      {stage2_28[39], stage2_28[40], stage2_28[41], stage2_28[42], stage2_28[43]},
      {stage2_29[10]},
      {stage2_30[24], stage2_30[25], stage2_30[26], stage2_30[27], stage2_30[28], stage2_30[29]},
      {stage3_32[4],stage3_31[5],stage3_30[6],stage3_29[27],stage3_28[28]}
   );
   gpc615_5 gpc7448 (
      {stage2_28[44], stage2_28[45], stage2_28[46], stage2_28[47], stage2_28[48]},
      {stage2_29[11]},
      {stage2_30[30], stage2_30[31], stage2_30[32], stage2_30[33], stage2_30[34], stage2_30[35]},
      {stage3_32[5],stage3_31[6],stage3_30[7],stage3_29[28],stage3_28[29]}
   );
   gpc615_5 gpc7449 (
      {stage2_28[49], stage2_28[50], stage2_28[51], stage2_28[52], stage2_28[53]},
      {stage2_29[12]},
      {stage2_30[36], stage2_30[37], stage2_30[38], stage2_30[39], stage2_30[40], stage2_30[41]},
      {stage3_32[6],stage3_31[7],stage3_30[8],stage3_29[29],stage3_28[30]}
   );
   gpc615_5 gpc7450 (
      {stage2_28[54], stage2_28[55], stage2_28[56], stage2_28[57], stage2_28[58]},
      {stage2_29[13]},
      {stage2_30[42], stage2_30[43], stage2_30[44], stage2_30[45], stage2_30[46], stage2_30[47]},
      {stage3_32[7],stage3_31[8],stage3_30[9],stage3_29[30],stage3_28[31]}
   );
   gpc615_5 gpc7451 (
      {stage2_28[59], stage2_28[60], stage2_28[61], stage2_28[62], stage2_28[63]},
      {stage2_29[14]},
      {stage2_30[48], stage2_30[49], stage2_30[50], stage2_30[51], stage2_30[52], stage2_30[53]},
      {stage3_32[8],stage3_31[9],stage3_30[10],stage3_29[31],stage3_28[32]}
   );
   gpc615_5 gpc7452 (
      {stage2_28[64], stage2_28[65], stage2_28[66], stage2_28[67], stage2_28[68]},
      {stage2_29[15]},
      {stage2_30[54], stage2_30[55], stage2_30[56], stage2_30[57], stage2_30[58], stage2_30[59]},
      {stage3_32[9],stage3_31[10],stage3_30[11],stage3_29[32],stage3_28[33]}
   );
   gpc1163_5 gpc7453 (
      {stage2_29[16], stage2_29[17], stage2_29[18]},
      {stage2_30[60], stage2_30[61], stage2_30[62], stage2_30[63], stage2_30[64], stage2_30[65]},
      {stage2_31[0]},
      {stage2_32[0]},
      {stage3_33[0],stage3_32[10],stage3_31[11],stage3_30[12],stage3_29[33]}
   );
   gpc1163_5 gpc7454 (
      {stage2_29[19], stage2_29[20], stage2_29[21]},
      {stage2_30[66], stage2_30[67], stage2_30[68], stage2_30[69], stage2_30[70], stage2_30[71]},
      {stage2_31[1]},
      {stage2_32[1]},
      {stage3_33[1],stage3_32[11],stage3_31[12],stage3_30[13],stage3_29[34]}
   );
   gpc1163_5 gpc7455 (
      {stage2_29[22], stage2_29[23], stage2_29[24]},
      {stage2_30[72], stage2_30[73], stage2_30[74], stage2_30[75], stage2_30[76], stage2_30[77]},
      {stage2_31[2]},
      {stage2_32[2]},
      {stage3_33[2],stage3_32[12],stage3_31[13],stage3_30[14],stage3_29[35]}
   );
   gpc1163_5 gpc7456 (
      {stage2_29[25], stage2_29[26], stage2_29[27]},
      {stage2_30[78], stage2_30[79], stage2_30[80], stage2_30[81], stage2_30[82], stage2_30[83]},
      {stage2_31[3]},
      {stage2_32[3]},
      {stage3_33[3],stage3_32[13],stage3_31[14],stage3_30[15],stage3_29[36]}
   );
   gpc1163_5 gpc7457 (
      {stage2_29[28], stage2_29[29], stage2_29[30]},
      {stage2_30[84], stage2_30[85], stage2_30[86], stage2_30[87], stage2_30[88], stage2_30[89]},
      {stage2_31[4]},
      {stage2_32[4]},
      {stage3_33[4],stage3_32[14],stage3_31[15],stage3_30[16],stage3_29[37]}
   );
   gpc1163_5 gpc7458 (
      {stage2_29[31], stage2_29[32], stage2_29[33]},
      {stage2_30[90], stage2_30[91], stage2_30[92], stage2_30[93], stage2_30[94], stage2_30[95]},
      {stage2_31[5]},
      {stage2_32[5]},
      {stage3_33[5],stage3_32[15],stage3_31[16],stage3_30[17],stage3_29[38]}
   );
   gpc606_5 gpc7459 (
      {stage2_29[34], stage2_29[35], stage2_29[36], stage2_29[37], stage2_29[38], stage2_29[39]},
      {stage2_31[6], stage2_31[7], stage2_31[8], stage2_31[9], stage2_31[10], stage2_31[11]},
      {stage3_33[6],stage3_32[16],stage3_31[17],stage3_30[18],stage3_29[39]}
   );
   gpc606_5 gpc7460 (
      {stage2_29[40], stage2_29[41], stage2_29[42], stage2_29[43], stage2_29[44], stage2_29[45]},
      {stage2_31[12], stage2_31[13], stage2_31[14], stage2_31[15], stage2_31[16], stage2_31[17]},
      {stage3_33[7],stage3_32[17],stage3_31[18],stage3_30[19],stage3_29[40]}
   );
   gpc606_5 gpc7461 (
      {stage2_29[46], stage2_29[47], stage2_29[48], stage2_29[49], stage2_29[50], stage2_29[51]},
      {stage2_31[18], stage2_31[19], stage2_31[20], stage2_31[21], stage2_31[22], stage2_31[23]},
      {stage3_33[8],stage3_32[18],stage3_31[19],stage3_30[20],stage3_29[41]}
   );
   gpc606_5 gpc7462 (
      {stage2_29[52], stage2_29[53], stage2_29[54], stage2_29[55], stage2_29[56], stage2_29[57]},
      {stage2_31[24], stage2_31[25], stage2_31[26], stage2_31[27], stage2_31[28], stage2_31[29]},
      {stage3_33[9],stage3_32[19],stage3_31[20],stage3_30[21],stage3_29[42]}
   );
   gpc606_5 gpc7463 (
      {stage2_29[58], stage2_29[59], stage2_29[60], stage2_29[61], stage2_29[62], stage2_29[63]},
      {stage2_31[30], stage2_31[31], stage2_31[32], stage2_31[33], stage2_31[34], stage2_31[35]},
      {stage3_33[10],stage3_32[20],stage3_31[21],stage3_30[22],stage3_29[43]}
   );
   gpc606_5 gpc7464 (
      {stage2_29[64], stage2_29[65], stage2_29[66], stage2_29[67], stage2_29[68], stage2_29[69]},
      {stage2_31[36], stage2_31[37], stage2_31[38], stage2_31[39], stage2_31[40], stage2_31[41]},
      {stage3_33[11],stage3_32[21],stage3_31[22],stage3_30[23],stage3_29[44]}
   );
   gpc606_5 gpc7465 (
      {stage2_29[70], stage2_29[71], stage2_29[72], stage2_29[73], stage2_29[74], stage2_29[75]},
      {stage2_31[42], stage2_31[43], stage2_31[44], stage2_31[45], stage2_31[46], stage2_31[47]},
      {stage3_33[12],stage3_32[22],stage3_31[23],stage3_30[24],stage3_29[45]}
   );
   gpc606_5 gpc7466 (
      {stage2_29[76], stage2_29[77], stage2_29[78], stage2_29[79], stage2_29[80], stage2_29[81]},
      {stage2_31[48], stage2_31[49], stage2_31[50], stage2_31[51], stage2_31[52], stage2_31[53]},
      {stage3_33[13],stage3_32[23],stage3_31[24],stage3_30[25],stage3_29[46]}
   );
   gpc606_5 gpc7467 (
      {stage2_29[82], stage2_29[83], stage2_29[84], stage2_29[85], stage2_29[86], 1'b0},
      {stage2_31[54], stage2_31[55], stage2_31[56], stage2_31[57], stage2_31[58], stage2_31[59]},
      {stage3_33[14],stage3_32[24],stage3_31[25],stage3_30[26],stage3_29[47]}
   );
   gpc207_4 gpc7468 (
      {stage2_30[96], stage2_30[97], stage2_30[98], stage2_30[99], stage2_30[100], stage2_30[101], stage2_30[102]},
      {stage2_32[6], stage2_32[7]},
      {stage3_33[15],stage3_32[25],stage3_31[26],stage3_30[27]}
   );
   gpc615_5 gpc7469 (
      {stage2_31[60], stage2_31[61], stage2_31[62], stage2_31[63], stage2_31[64]},
      {stage2_32[8]},
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5]},
      {stage3_35[0],stage3_34[0],stage3_33[16],stage3_32[26],stage3_31[27]}
   );
   gpc615_5 gpc7470 (
      {stage2_31[65], stage2_31[66], stage2_31[67], stage2_31[68], stage2_31[69]},
      {stage2_32[9]},
      {stage2_33[6], stage2_33[7], stage2_33[8], stage2_33[9], stage2_33[10], stage2_33[11]},
      {stage3_35[1],stage3_34[1],stage3_33[17],stage3_32[27],stage3_31[28]}
   );
   gpc615_5 gpc7471 (
      {stage2_31[70], stage2_31[71], stage2_31[72], stage2_31[73], stage2_31[74]},
      {stage2_32[10]},
      {stage2_33[12], stage2_33[13], stage2_33[14], stage2_33[15], stage2_33[16], stage2_33[17]},
      {stage3_35[2],stage3_34[2],stage3_33[18],stage3_32[28],stage3_31[29]}
   );
   gpc615_5 gpc7472 (
      {stage2_31[75], stage2_31[76], stage2_31[77], stage2_31[78], stage2_31[79]},
      {stage2_32[11]},
      {stage2_33[18], stage2_33[19], stage2_33[20], stage2_33[21], stage2_33[22], stage2_33[23]},
      {stage3_35[3],stage3_34[3],stage3_33[19],stage3_32[29],stage3_31[30]}
   );
   gpc615_5 gpc7473 (
      {stage2_31[80], stage2_31[81], stage2_31[82], stage2_31[83], stage2_31[84]},
      {stage2_32[12]},
      {stage2_33[24], stage2_33[25], stage2_33[26], stage2_33[27], stage2_33[28], stage2_33[29]},
      {stage3_35[4],stage3_34[4],stage3_33[20],stage3_32[30],stage3_31[31]}
   );
   gpc615_5 gpc7474 (
      {stage2_31[85], stage2_31[86], stage2_31[87], stage2_31[88], stage2_31[89]},
      {stage2_32[13]},
      {stage2_33[30], stage2_33[31], stage2_33[32], stage2_33[33], stage2_33[34], stage2_33[35]},
      {stage3_35[5],stage3_34[5],stage3_33[21],stage3_32[31],stage3_31[32]}
   );
   gpc615_5 gpc7475 (
      {stage2_31[90], stage2_31[91], stage2_31[92], stage2_31[93], stage2_31[94]},
      {stage2_32[14]},
      {stage2_33[36], stage2_33[37], stage2_33[38], stage2_33[39], stage2_33[40], stage2_33[41]},
      {stage3_35[6],stage3_34[6],stage3_33[22],stage3_32[32],stage3_31[33]}
   );
   gpc606_5 gpc7476 (
      {stage2_32[15], stage2_32[16], stage2_32[17], stage2_32[18], stage2_32[19], stage2_32[20]},
      {stage2_34[0], stage2_34[1], stage2_34[2], stage2_34[3], stage2_34[4], stage2_34[5]},
      {stage3_36[0],stage3_35[7],stage3_34[7],stage3_33[23],stage3_32[33]}
   );
   gpc606_5 gpc7477 (
      {stage2_32[21], stage2_32[22], stage2_32[23], stage2_32[24], stage2_32[25], stage2_32[26]},
      {stage2_34[6], stage2_34[7], stage2_34[8], stage2_34[9], stage2_34[10], stage2_34[11]},
      {stage3_36[1],stage3_35[8],stage3_34[8],stage3_33[24],stage3_32[34]}
   );
   gpc606_5 gpc7478 (
      {stage2_32[27], stage2_32[28], stage2_32[29], stage2_32[30], stage2_32[31], stage2_32[32]},
      {stage2_34[12], stage2_34[13], stage2_34[14], stage2_34[15], stage2_34[16], stage2_34[17]},
      {stage3_36[2],stage3_35[9],stage3_34[9],stage3_33[25],stage3_32[35]}
   );
   gpc606_5 gpc7479 (
      {stage2_32[33], stage2_32[34], stage2_32[35], stage2_32[36], stage2_32[37], stage2_32[38]},
      {stage2_34[18], stage2_34[19], stage2_34[20], stage2_34[21], stage2_34[22], stage2_34[23]},
      {stage3_36[3],stage3_35[10],stage3_34[10],stage3_33[26],stage3_32[36]}
   );
   gpc606_5 gpc7480 (
      {stage2_32[39], stage2_32[40], stage2_32[41], stage2_32[42], stage2_32[43], stage2_32[44]},
      {stage2_34[24], stage2_34[25], stage2_34[26], stage2_34[27], stage2_34[28], stage2_34[29]},
      {stage3_36[4],stage3_35[11],stage3_34[11],stage3_33[27],stage3_32[37]}
   );
   gpc606_5 gpc7481 (
      {stage2_32[45], stage2_32[46], stage2_32[47], stage2_32[48], stage2_32[49], stage2_32[50]},
      {stage2_34[30], stage2_34[31], stage2_34[32], stage2_34[33], stage2_34[34], stage2_34[35]},
      {stage3_36[5],stage3_35[12],stage3_34[12],stage3_33[28],stage3_32[38]}
   );
   gpc606_5 gpc7482 (
      {stage2_32[51], stage2_32[52], stage2_32[53], stage2_32[54], stage2_32[55], stage2_32[56]},
      {stage2_34[36], stage2_34[37], stage2_34[38], stage2_34[39], stage2_34[40], stage2_34[41]},
      {stage3_36[6],stage3_35[13],stage3_34[13],stage3_33[29],stage3_32[39]}
   );
   gpc606_5 gpc7483 (
      {stage2_32[57], stage2_32[58], stage2_32[59], stage2_32[60], stage2_32[61], stage2_32[62]},
      {stage2_34[42], stage2_34[43], stage2_34[44], stage2_34[45], stage2_34[46], stage2_34[47]},
      {stage3_36[7],stage3_35[14],stage3_34[14],stage3_33[30],stage3_32[40]}
   );
   gpc606_5 gpc7484 (
      {stage2_32[63], stage2_32[64], stage2_32[65], stage2_32[66], stage2_32[67], stage2_32[68]},
      {stage2_34[48], stage2_34[49], stage2_34[50], stage2_34[51], stage2_34[52], stage2_34[53]},
      {stage3_36[8],stage3_35[15],stage3_34[15],stage3_33[31],stage3_32[41]}
   );
   gpc606_5 gpc7485 (
      {stage2_32[69], stage2_32[70], stage2_32[71], stage2_32[72], stage2_32[73], stage2_32[74]},
      {stage2_34[54], stage2_34[55], stage2_34[56], stage2_34[57], stage2_34[58], stage2_34[59]},
      {stage3_36[9],stage3_35[16],stage3_34[16],stage3_33[32],stage3_32[42]}
   );
   gpc606_5 gpc7486 (
      {stage2_32[75], stage2_32[76], stage2_32[77], stage2_32[78], stage2_32[79], stage2_32[80]},
      {stage2_34[60], stage2_34[61], stage2_34[62], stage2_34[63], stage2_34[64], stage2_34[65]},
      {stage3_36[10],stage3_35[17],stage3_34[17],stage3_33[33],stage3_32[43]}
   );
   gpc606_5 gpc7487 (
      {stage2_32[81], stage2_32[82], stage2_32[83], stage2_32[84], stage2_32[85], stage2_32[86]},
      {stage2_34[66], stage2_34[67], stage2_34[68], stage2_34[69], stage2_34[70], stage2_34[71]},
      {stage3_36[11],stage3_35[18],stage3_34[18],stage3_33[34],stage3_32[44]}
   );
   gpc606_5 gpc7488 (
      {stage2_32[87], stage2_32[88], stage2_32[89], stage2_32[90], stage2_32[91], stage2_32[92]},
      {stage2_34[72], stage2_34[73], stage2_34[74], stage2_34[75], stage2_34[76], stage2_34[77]},
      {stage3_36[12],stage3_35[19],stage3_34[19],stage3_33[35],stage3_32[45]}
   );
   gpc606_5 gpc7489 (
      {stage2_32[93], stage2_32[94], stage2_32[95], stage2_32[96], stage2_32[97], stage2_32[98]},
      {stage2_34[78], stage2_34[79], stage2_34[80], stage2_34[81], stage2_34[82], stage2_34[83]},
      {stage3_36[13],stage3_35[20],stage3_34[20],stage3_33[36],stage3_32[46]}
   );
   gpc606_5 gpc7490 (
      {stage2_33[42], stage2_33[43], stage2_33[44], stage2_33[45], stage2_33[46], stage2_33[47]},
      {stage2_35[0], stage2_35[1], stage2_35[2], stage2_35[3], stage2_35[4], stage2_35[5]},
      {stage3_37[0],stage3_36[14],stage3_35[21],stage3_34[21],stage3_33[37]}
   );
   gpc606_5 gpc7491 (
      {stage2_33[48], stage2_33[49], stage2_33[50], stage2_33[51], stage2_33[52], stage2_33[53]},
      {stage2_35[6], stage2_35[7], stage2_35[8], stage2_35[9], stage2_35[10], stage2_35[11]},
      {stage3_37[1],stage3_36[15],stage3_35[22],stage3_34[22],stage3_33[38]}
   );
   gpc606_5 gpc7492 (
      {stage2_33[54], stage2_33[55], stage2_33[56], stage2_33[57], stage2_33[58], stage2_33[59]},
      {stage2_35[12], stage2_35[13], stage2_35[14], stage2_35[15], stage2_35[16], stage2_35[17]},
      {stage3_37[2],stage3_36[16],stage3_35[23],stage3_34[23],stage3_33[39]}
   );
   gpc606_5 gpc7493 (
      {stage2_33[60], stage2_33[61], stage2_33[62], stage2_33[63], stage2_33[64], stage2_33[65]},
      {stage2_35[18], stage2_35[19], stage2_35[20], stage2_35[21], stage2_35[22], stage2_35[23]},
      {stage3_37[3],stage3_36[17],stage3_35[24],stage3_34[24],stage3_33[40]}
   );
   gpc606_5 gpc7494 (
      {stage2_33[66], stage2_33[67], stage2_33[68], stage2_33[69], stage2_33[70], stage2_33[71]},
      {stage2_35[24], stage2_35[25], stage2_35[26], stage2_35[27], stage2_35[28], stage2_35[29]},
      {stage3_37[4],stage3_36[18],stage3_35[25],stage3_34[25],stage3_33[41]}
   );
   gpc1163_5 gpc7495 (
      {stage2_34[84], stage2_34[85], stage2_34[86]},
      {stage2_35[30], stage2_35[31], stage2_35[32], stage2_35[33], stage2_35[34], stage2_35[35]},
      {stage2_36[0]},
      {stage2_37[0]},
      {stage3_38[0],stage3_37[5],stage3_36[19],stage3_35[26],stage3_34[26]}
   );
   gpc1163_5 gpc7496 (
      {stage2_34[87], stage2_34[88], stage2_34[89]},
      {stage2_35[36], stage2_35[37], stage2_35[38], stage2_35[39], stage2_35[40], stage2_35[41]},
      {stage2_36[1]},
      {stage2_37[1]},
      {stage3_38[1],stage3_37[6],stage3_36[20],stage3_35[27],stage3_34[27]}
   );
   gpc1163_5 gpc7497 (
      {stage2_34[90], stage2_34[91], stage2_34[92]},
      {stage2_35[42], stage2_35[43], stage2_35[44], stage2_35[45], stage2_35[46], stage2_35[47]},
      {stage2_36[2]},
      {stage2_37[2]},
      {stage3_38[2],stage3_37[7],stage3_36[21],stage3_35[28],stage3_34[28]}
   );
   gpc1163_5 gpc7498 (
      {stage2_34[93], stage2_34[94], stage2_34[95]},
      {stage2_35[48], stage2_35[49], stage2_35[50], stage2_35[51], stage2_35[52], stage2_35[53]},
      {stage2_36[3]},
      {stage2_37[3]},
      {stage3_38[3],stage3_37[8],stage3_36[22],stage3_35[29],stage3_34[29]}
   );
   gpc1163_5 gpc7499 (
      {stage2_34[96], stage2_34[97], stage2_34[98]},
      {stage2_35[54], stage2_35[55], stage2_35[56], stage2_35[57], stage2_35[58], stage2_35[59]},
      {stage2_36[4]},
      {stage2_37[4]},
      {stage3_38[4],stage3_37[9],stage3_36[23],stage3_35[30],stage3_34[30]}
   );
   gpc1163_5 gpc7500 (
      {stage2_34[99], stage2_34[100], stage2_34[101]},
      {stage2_35[60], stage2_35[61], stage2_35[62], stage2_35[63], stage2_35[64], stage2_35[65]},
      {stage2_36[5]},
      {stage2_37[5]},
      {stage3_38[5],stage3_37[10],stage3_36[24],stage3_35[31],stage3_34[31]}
   );
   gpc1163_5 gpc7501 (
      {stage2_34[102], stage2_34[103], stage2_34[104]},
      {stage2_35[66], stage2_35[67], stage2_35[68], stage2_35[69], stage2_35[70], stage2_35[71]},
      {stage2_36[6]},
      {stage2_37[6]},
      {stage3_38[6],stage3_37[11],stage3_36[25],stage3_35[32],stage3_34[32]}
   );
   gpc1163_5 gpc7502 (
      {stage2_34[105], stage2_34[106], stage2_34[107]},
      {stage2_35[72], stage2_35[73], stage2_35[74], stage2_35[75], stage2_35[76], stage2_35[77]},
      {stage2_36[7]},
      {stage2_37[7]},
      {stage3_38[7],stage3_37[12],stage3_36[26],stage3_35[33],stage3_34[33]}
   );
   gpc1163_5 gpc7503 (
      {stage2_34[108], stage2_34[109], stage2_34[110]},
      {stage2_35[78], stage2_35[79], stage2_35[80], stage2_35[81], stage2_35[82], stage2_35[83]},
      {stage2_36[8]},
      {stage2_37[8]},
      {stage3_38[8],stage3_37[13],stage3_36[27],stage3_35[34],stage3_34[34]}
   );
   gpc1163_5 gpc7504 (
      {stage2_34[111], stage2_34[112], stage2_34[113]},
      {stage2_35[84], stage2_35[85], stage2_35[86], stage2_35[87], stage2_35[88], stage2_35[89]},
      {stage2_36[9]},
      {stage2_37[9]},
      {stage3_38[9],stage3_37[14],stage3_36[28],stage3_35[35],stage3_34[35]}
   );
   gpc615_5 gpc7505 (
      {stage2_34[114], stage2_34[115], stage2_34[116], stage2_34[117], stage2_34[118]},
      {stage2_35[90]},
      {stage2_36[10], stage2_36[11], stage2_36[12], stage2_36[13], stage2_36[14], stage2_36[15]},
      {stage3_38[10],stage3_37[15],stage3_36[29],stage3_35[36],stage3_34[36]}
   );
   gpc615_5 gpc7506 (
      {stage2_34[119], stage2_34[120], stage2_34[121], stage2_34[122], stage2_34[123]},
      {stage2_35[91]},
      {stage2_36[16], stage2_36[17], stage2_36[18], stage2_36[19], stage2_36[20], stage2_36[21]},
      {stage3_38[11],stage3_37[16],stage3_36[30],stage3_35[37],stage3_34[37]}
   );
   gpc615_5 gpc7507 (
      {stage2_34[124], stage2_34[125], stage2_34[126], stage2_34[127], stage2_34[128]},
      {stage2_35[92]},
      {stage2_36[22], stage2_36[23], stage2_36[24], stage2_36[25], stage2_36[26], stage2_36[27]},
      {stage3_38[12],stage3_37[17],stage3_36[31],stage3_35[38],stage3_34[38]}
   );
   gpc1406_5 gpc7508 (
      {stage2_35[93], stage2_35[94], stage2_35[95], stage2_35[96], stage2_35[97], stage2_35[98]},
      {stage2_37[10], stage2_37[11], stage2_37[12], stage2_37[13]},
      {stage2_38[0]},
      {stage3_39[0],stage3_38[13],stage3_37[18],stage3_36[32],stage3_35[39]}
   );
   gpc1406_5 gpc7509 (
      {stage2_35[99], stage2_35[100], stage2_35[101], stage2_35[102], stage2_35[103], stage2_35[104]},
      {stage2_37[14], stage2_37[15], stage2_37[16], stage2_37[17]},
      {stage2_38[1]},
      {stage3_39[1],stage3_38[14],stage3_37[19],stage3_36[33],stage3_35[40]}
   );
   gpc615_5 gpc7510 (
      {stage2_35[105], stage2_35[106], stage2_35[107], stage2_35[108], stage2_35[109]},
      {stage2_36[28]},
      {stage2_37[18], stage2_37[19], stage2_37[20], stage2_37[21], stage2_37[22], stage2_37[23]},
      {stage3_39[2],stage3_38[15],stage3_37[20],stage3_36[34],stage3_35[41]}
   );
   gpc615_5 gpc7511 (
      {stage2_35[110], stage2_35[111], stage2_35[112], stage2_35[113], stage2_35[114]},
      {stage2_36[29]},
      {stage2_37[24], stage2_37[25], stage2_37[26], stage2_37[27], stage2_37[28], stage2_37[29]},
      {stage3_39[3],stage3_38[16],stage3_37[21],stage3_36[35],stage3_35[42]}
   );
   gpc615_5 gpc7512 (
      {stage2_35[115], stage2_35[116], stage2_35[117], stage2_35[118], stage2_35[119]},
      {stage2_36[30]},
      {stage2_37[30], stage2_37[31], stage2_37[32], stage2_37[33], stage2_37[34], stage2_37[35]},
      {stage3_39[4],stage3_38[17],stage3_37[22],stage3_36[36],stage3_35[43]}
   );
   gpc606_5 gpc7513 (
      {stage2_36[31], stage2_36[32], stage2_36[33], stage2_36[34], stage2_36[35], stage2_36[36]},
      {stage2_38[2], stage2_38[3], stage2_38[4], stage2_38[5], stage2_38[6], stage2_38[7]},
      {stage3_40[0],stage3_39[5],stage3_38[18],stage3_37[23],stage3_36[37]}
   );
   gpc606_5 gpc7514 (
      {stage2_36[37], stage2_36[38], stage2_36[39], stage2_36[40], stage2_36[41], stage2_36[42]},
      {stage2_38[8], stage2_38[9], stage2_38[10], stage2_38[11], stage2_38[12], stage2_38[13]},
      {stage3_40[1],stage3_39[6],stage3_38[19],stage3_37[24],stage3_36[38]}
   );
   gpc606_5 gpc7515 (
      {stage2_36[43], stage2_36[44], stage2_36[45], stage2_36[46], stage2_36[47], stage2_36[48]},
      {stage2_38[14], stage2_38[15], stage2_38[16], stage2_38[17], stage2_38[18], stage2_38[19]},
      {stage3_40[2],stage3_39[7],stage3_38[20],stage3_37[25],stage3_36[39]}
   );
   gpc606_5 gpc7516 (
      {stage2_36[49], stage2_36[50], stage2_36[51], stage2_36[52], stage2_36[53], stage2_36[54]},
      {stage2_38[20], stage2_38[21], stage2_38[22], stage2_38[23], stage2_38[24], stage2_38[25]},
      {stage3_40[3],stage3_39[8],stage3_38[21],stage3_37[26],stage3_36[40]}
   );
   gpc606_5 gpc7517 (
      {stage2_36[55], stage2_36[56], stage2_36[57], stage2_36[58], stage2_36[59], stage2_36[60]},
      {stage2_38[26], stage2_38[27], stage2_38[28], stage2_38[29], stage2_38[30], stage2_38[31]},
      {stage3_40[4],stage3_39[9],stage3_38[22],stage3_37[27],stage3_36[41]}
   );
   gpc606_5 gpc7518 (
      {stage2_36[61], stage2_36[62], stage2_36[63], stage2_36[64], stage2_36[65], stage2_36[66]},
      {stage2_38[32], stage2_38[33], stage2_38[34], stage2_38[35], stage2_38[36], stage2_38[37]},
      {stage3_40[5],stage3_39[10],stage3_38[23],stage3_37[28],stage3_36[42]}
   );
   gpc606_5 gpc7519 (
      {stage2_36[67], stage2_36[68], stage2_36[69], stage2_36[70], stage2_36[71], stage2_36[72]},
      {stage2_38[38], stage2_38[39], stage2_38[40], stage2_38[41], stage2_38[42], stage2_38[43]},
      {stage3_40[6],stage3_39[11],stage3_38[24],stage3_37[29],stage3_36[43]}
   );
   gpc606_5 gpc7520 (
      {stage2_37[36], stage2_37[37], stage2_37[38], stage2_37[39], stage2_37[40], stage2_37[41]},
      {stage2_39[0], stage2_39[1], stage2_39[2], stage2_39[3], stage2_39[4], stage2_39[5]},
      {stage3_41[0],stage3_40[7],stage3_39[12],stage3_38[25],stage3_37[30]}
   );
   gpc606_5 gpc7521 (
      {stage2_37[42], stage2_37[43], stage2_37[44], stage2_37[45], stage2_37[46], stage2_37[47]},
      {stage2_39[6], stage2_39[7], stage2_39[8], stage2_39[9], stage2_39[10], stage2_39[11]},
      {stage3_41[1],stage3_40[8],stage3_39[13],stage3_38[26],stage3_37[31]}
   );
   gpc606_5 gpc7522 (
      {stage2_37[48], stage2_37[49], stage2_37[50], stage2_37[51], stage2_37[52], stage2_37[53]},
      {stage2_39[12], stage2_39[13], stage2_39[14], stage2_39[15], stage2_39[16], stage2_39[17]},
      {stage3_41[2],stage3_40[9],stage3_39[14],stage3_38[27],stage3_37[32]}
   );
   gpc615_5 gpc7523 (
      {stage2_37[54], stage2_37[55], stage2_37[56], stage2_37[57], stage2_37[58]},
      {stage2_38[44]},
      {stage2_39[18], stage2_39[19], stage2_39[20], stage2_39[21], stage2_39[22], stage2_39[23]},
      {stage3_41[3],stage3_40[10],stage3_39[15],stage3_38[28],stage3_37[33]}
   );
   gpc615_5 gpc7524 (
      {stage2_37[59], stage2_37[60], stage2_37[61], stage2_37[62], stage2_37[63]},
      {stage2_38[45]},
      {stage2_39[24], stage2_39[25], stage2_39[26], stage2_39[27], stage2_39[28], stage2_39[29]},
      {stage3_41[4],stage3_40[11],stage3_39[16],stage3_38[29],stage3_37[34]}
   );
   gpc615_5 gpc7525 (
      {stage2_37[64], stage2_37[65], stage2_37[66], stage2_37[67], stage2_37[68]},
      {stage2_38[46]},
      {stage2_39[30], stage2_39[31], stage2_39[32], stage2_39[33], stage2_39[34], stage2_39[35]},
      {stage3_41[5],stage3_40[12],stage3_39[17],stage3_38[30],stage3_37[35]}
   );
   gpc615_5 gpc7526 (
      {stage2_37[69], stage2_37[70], stage2_37[71], stage2_37[72], stage2_37[73]},
      {stage2_38[47]},
      {stage2_39[36], stage2_39[37], stage2_39[38], stage2_39[39], stage2_39[40], stage2_39[41]},
      {stage3_41[6],stage3_40[13],stage3_39[18],stage3_38[31],stage3_37[36]}
   );
   gpc606_5 gpc7527 (
      {stage2_38[48], stage2_38[49], stage2_38[50], stage2_38[51], stage2_38[52], stage2_38[53]},
      {stage2_40[0], stage2_40[1], stage2_40[2], stage2_40[3], stage2_40[4], stage2_40[5]},
      {stage3_42[0],stage3_41[7],stage3_40[14],stage3_39[19],stage3_38[32]}
   );
   gpc606_5 gpc7528 (
      {stage2_38[54], stage2_38[55], stage2_38[56], stage2_38[57], stage2_38[58], stage2_38[59]},
      {stage2_40[6], stage2_40[7], stage2_40[8], stage2_40[9], stage2_40[10], stage2_40[11]},
      {stage3_42[1],stage3_41[8],stage3_40[15],stage3_39[20],stage3_38[33]}
   );
   gpc606_5 gpc7529 (
      {stage2_38[60], stage2_38[61], stage2_38[62], stage2_38[63], stage2_38[64], stage2_38[65]},
      {stage2_40[12], stage2_40[13], stage2_40[14], stage2_40[15], stage2_40[16], stage2_40[17]},
      {stage3_42[2],stage3_41[9],stage3_40[16],stage3_39[21],stage3_38[34]}
   );
   gpc606_5 gpc7530 (
      {stage2_38[66], stage2_38[67], stage2_38[68], stage2_38[69], stage2_38[70], stage2_38[71]},
      {stage2_40[18], stage2_40[19], stage2_40[20], stage2_40[21], stage2_40[22], stage2_40[23]},
      {stage3_42[3],stage3_41[10],stage3_40[17],stage3_39[22],stage3_38[35]}
   );
   gpc606_5 gpc7531 (
      {stage2_38[72], stage2_38[73], stage2_38[74], stage2_38[75], stage2_38[76], stage2_38[77]},
      {stage2_40[24], stage2_40[25], stage2_40[26], stage2_40[27], stage2_40[28], stage2_40[29]},
      {stage3_42[4],stage3_41[11],stage3_40[18],stage3_39[23],stage3_38[36]}
   );
   gpc606_5 gpc7532 (
      {stage2_38[78], stage2_38[79], stage2_38[80], stage2_38[81], stage2_38[82], stage2_38[83]},
      {stage2_40[30], stage2_40[31], stage2_40[32], stage2_40[33], stage2_40[34], stage2_40[35]},
      {stage3_42[5],stage3_41[12],stage3_40[19],stage3_39[24],stage3_38[37]}
   );
   gpc606_5 gpc7533 (
      {stage2_38[84], stage2_38[85], stage2_38[86], stage2_38[87], stage2_38[88], stage2_38[89]},
      {stage2_40[36], stage2_40[37], stage2_40[38], stage2_40[39], stage2_40[40], stage2_40[41]},
      {stage3_42[6],stage3_41[13],stage3_40[20],stage3_39[25],stage3_38[38]}
   );
   gpc606_5 gpc7534 (
      {stage2_38[90], stage2_38[91], stage2_38[92], stage2_38[93], stage2_38[94], stage2_38[95]},
      {stage2_40[42], stage2_40[43], stage2_40[44], stage2_40[45], stage2_40[46], stage2_40[47]},
      {stage3_42[7],stage3_41[14],stage3_40[21],stage3_39[26],stage3_38[39]}
   );
   gpc606_5 gpc7535 (
      {stage2_38[96], stage2_38[97], stage2_38[98], stage2_38[99], stage2_38[100], stage2_38[101]},
      {stage2_40[48], stage2_40[49], stage2_40[50], stage2_40[51], stage2_40[52], stage2_40[53]},
      {stage3_42[8],stage3_41[15],stage3_40[22],stage3_39[27],stage3_38[40]}
   );
   gpc606_5 gpc7536 (
      {stage2_38[102], stage2_38[103], stage2_38[104], stage2_38[105], stage2_38[106], stage2_38[107]},
      {stage2_40[54], stage2_40[55], stage2_40[56], stage2_40[57], stage2_40[58], stage2_40[59]},
      {stage3_42[9],stage3_41[16],stage3_40[23],stage3_39[28],stage3_38[41]}
   );
   gpc606_5 gpc7537 (
      {stage2_38[108], stage2_38[109], stage2_38[110], stage2_38[111], stage2_38[112], stage2_38[113]},
      {stage2_40[60], stage2_40[61], stage2_40[62], stage2_40[63], stage2_40[64], stage2_40[65]},
      {stage3_42[10],stage3_41[17],stage3_40[24],stage3_39[29],stage3_38[42]}
   );
   gpc606_5 gpc7538 (
      {stage2_38[114], stage2_38[115], stage2_38[116], stage2_38[117], stage2_38[118], stage2_38[119]},
      {stage2_40[66], stage2_40[67], stage2_40[68], stage2_40[69], stage2_40[70], stage2_40[71]},
      {stage3_42[11],stage3_41[18],stage3_40[25],stage3_39[30],stage3_38[43]}
   );
   gpc615_5 gpc7539 (
      {stage2_38[120], stage2_38[121], stage2_38[122], stage2_38[123], stage2_38[124]},
      {stage2_39[42]},
      {stage2_40[72], stage2_40[73], stage2_40[74], stage2_40[75], stage2_40[76], stage2_40[77]},
      {stage3_42[12],stage3_41[19],stage3_40[26],stage3_39[31],stage3_38[44]}
   );
   gpc615_5 gpc7540 (
      {stage2_39[43], stage2_39[44], stage2_39[45], stage2_39[46], stage2_39[47]},
      {stage2_40[78]},
      {stage2_41[0], stage2_41[1], stage2_41[2], stage2_41[3], stage2_41[4], stage2_41[5]},
      {stage3_43[0],stage3_42[13],stage3_41[20],stage3_40[27],stage3_39[32]}
   );
   gpc615_5 gpc7541 (
      {stage2_39[48], stage2_39[49], stage2_39[50], stage2_39[51], stage2_39[52]},
      {stage2_40[79]},
      {stage2_41[6], stage2_41[7], stage2_41[8], stage2_41[9], stage2_41[10], stage2_41[11]},
      {stage3_43[1],stage3_42[14],stage3_41[21],stage3_40[28],stage3_39[33]}
   );
   gpc615_5 gpc7542 (
      {stage2_39[53], stage2_39[54], stage2_39[55], stage2_39[56], stage2_39[57]},
      {stage2_40[80]},
      {stage2_41[12], stage2_41[13], stage2_41[14], stage2_41[15], stage2_41[16], stage2_41[17]},
      {stage3_43[2],stage3_42[15],stage3_41[22],stage3_40[29],stage3_39[34]}
   );
   gpc615_5 gpc7543 (
      {stage2_39[58], stage2_39[59], stage2_39[60], stage2_39[61], stage2_39[62]},
      {stage2_40[81]},
      {stage2_41[18], stage2_41[19], stage2_41[20], stage2_41[21], stage2_41[22], stage2_41[23]},
      {stage3_43[3],stage3_42[16],stage3_41[23],stage3_40[30],stage3_39[35]}
   );
   gpc615_5 gpc7544 (
      {stage2_39[63], stage2_39[64], stage2_39[65], stage2_39[66], stage2_39[67]},
      {stage2_40[82]},
      {stage2_41[24], stage2_41[25], stage2_41[26], stage2_41[27], stage2_41[28], stage2_41[29]},
      {stage3_43[4],stage3_42[17],stage3_41[24],stage3_40[31],stage3_39[36]}
   );
   gpc615_5 gpc7545 (
      {stage2_39[68], stage2_39[69], stage2_39[70], stage2_39[71], stage2_39[72]},
      {stage2_40[83]},
      {stage2_41[30], stage2_41[31], stage2_41[32], stage2_41[33], stage2_41[34], stage2_41[35]},
      {stage3_43[5],stage3_42[18],stage3_41[25],stage3_40[32],stage3_39[37]}
   );
   gpc615_5 gpc7546 (
      {stage2_39[73], stage2_39[74], stage2_39[75], stage2_39[76], stage2_39[77]},
      {stage2_40[84]},
      {stage2_41[36], stage2_41[37], stage2_41[38], stage2_41[39], stage2_41[40], stage2_41[41]},
      {stage3_43[6],stage3_42[19],stage3_41[26],stage3_40[33],stage3_39[38]}
   );
   gpc615_5 gpc7547 (
      {stage2_39[78], stage2_39[79], stage2_39[80], stage2_39[81], stage2_39[82]},
      {stage2_40[85]},
      {stage2_41[42], stage2_41[43], stage2_41[44], stage2_41[45], stage2_41[46], stage2_41[47]},
      {stage3_43[7],stage3_42[20],stage3_41[27],stage3_40[34],stage3_39[39]}
   );
   gpc615_5 gpc7548 (
      {stage2_39[83], stage2_39[84], stage2_39[85], stage2_39[86], stage2_39[87]},
      {stage2_40[86]},
      {stage2_41[48], stage2_41[49], stage2_41[50], stage2_41[51], stage2_41[52], stage2_41[53]},
      {stage3_43[8],stage3_42[21],stage3_41[28],stage3_40[35],stage3_39[40]}
   );
   gpc615_5 gpc7549 (
      {stage2_39[88], stage2_39[89], stage2_39[90], stage2_39[91], stage2_39[92]},
      {stage2_40[87]},
      {stage2_41[54], stage2_41[55], stage2_41[56], stage2_41[57], stage2_41[58], stage2_41[59]},
      {stage3_43[9],stage3_42[22],stage3_41[29],stage3_40[36],stage3_39[41]}
   );
   gpc615_5 gpc7550 (
      {stage2_39[93], stage2_39[94], stage2_39[95], stage2_39[96], stage2_39[97]},
      {stage2_40[88]},
      {stage2_41[60], stage2_41[61], stage2_41[62], stage2_41[63], stage2_41[64], stage2_41[65]},
      {stage3_43[10],stage3_42[23],stage3_41[30],stage3_40[37],stage3_39[42]}
   );
   gpc615_5 gpc7551 (
      {stage2_39[98], stage2_39[99], stage2_39[100], stage2_39[101], stage2_39[102]},
      {stage2_40[89]},
      {stage2_41[66], stage2_41[67], stage2_41[68], stage2_41[69], stage2_41[70], stage2_41[71]},
      {stage3_43[11],stage3_42[24],stage3_41[31],stage3_40[38],stage3_39[43]}
   );
   gpc615_5 gpc7552 (
      {stage2_39[103], stage2_39[104], stage2_39[105], stage2_39[106], stage2_39[107]},
      {stage2_40[90]},
      {stage2_41[72], stage2_41[73], stage2_41[74], stage2_41[75], stage2_41[76], stage2_41[77]},
      {stage3_43[12],stage3_42[25],stage3_41[32],stage3_40[39],stage3_39[44]}
   );
   gpc615_5 gpc7553 (
      {stage2_39[108], stage2_39[109], stage2_39[110], stage2_39[111], stage2_39[112]},
      {stage2_40[91]},
      {stage2_41[78], stage2_41[79], stage2_41[80], stage2_41[81], stage2_41[82], stage2_41[83]},
      {stage3_43[13],stage3_42[26],stage3_41[33],stage3_40[40],stage3_39[45]}
   );
   gpc615_5 gpc7554 (
      {stage2_39[113], stage2_39[114], stage2_39[115], stage2_39[116], stage2_39[117]},
      {stage2_40[92]},
      {stage2_41[84], stage2_41[85], stage2_41[86], stage2_41[87], stage2_41[88], stage2_41[89]},
      {stage3_43[14],stage3_42[27],stage3_41[34],stage3_40[41],stage3_39[46]}
   );
   gpc615_5 gpc7555 (
      {stage2_39[118], stage2_39[119], stage2_39[120], stage2_39[121], stage2_39[122]},
      {stage2_40[93]},
      {stage2_41[90], stage2_41[91], stage2_41[92], stage2_41[93], stage2_41[94], stage2_41[95]},
      {stage3_43[15],stage3_42[28],stage3_41[35],stage3_40[42],stage3_39[47]}
   );
   gpc615_5 gpc7556 (
      {stage2_39[123], stage2_39[124], stage2_39[125], stage2_39[126], stage2_39[127]},
      {stage2_40[94]},
      {stage2_41[96], stage2_41[97], stage2_41[98], stage2_41[99], stage2_41[100], stage2_41[101]},
      {stage3_43[16],stage3_42[29],stage3_41[36],stage3_40[43],stage3_39[48]}
   );
   gpc606_5 gpc7557 (
      {stage2_40[95], stage2_40[96], stage2_40[97], stage2_40[98], stage2_40[99], stage2_40[100]},
      {stage2_42[0], stage2_42[1], stage2_42[2], stage2_42[3], stage2_42[4], stage2_42[5]},
      {stage3_44[0],stage3_43[17],stage3_42[30],stage3_41[37],stage3_40[44]}
   );
   gpc606_5 gpc7558 (
      {stage2_40[101], stage2_40[102], stage2_40[103], stage2_40[104], stage2_40[105], stage2_40[106]},
      {stage2_42[6], stage2_42[7], stage2_42[8], stage2_42[9], stage2_42[10], stage2_42[11]},
      {stage3_44[1],stage3_43[18],stage3_42[31],stage3_41[38],stage3_40[45]}
   );
   gpc615_5 gpc7559 (
      {stage2_42[12], stage2_42[13], stage2_42[14], stage2_42[15], stage2_42[16]},
      {stage2_43[0]},
      {stage2_44[0], stage2_44[1], stage2_44[2], stage2_44[3], stage2_44[4], stage2_44[5]},
      {stage3_46[0],stage3_45[0],stage3_44[2],stage3_43[19],stage3_42[32]}
   );
   gpc615_5 gpc7560 (
      {stage2_42[17], stage2_42[18], stage2_42[19], stage2_42[20], stage2_42[21]},
      {stage2_43[1]},
      {stage2_44[6], stage2_44[7], stage2_44[8], stage2_44[9], stage2_44[10], stage2_44[11]},
      {stage3_46[1],stage3_45[1],stage3_44[3],stage3_43[20],stage3_42[33]}
   );
   gpc615_5 gpc7561 (
      {stage2_42[22], stage2_42[23], stage2_42[24], stage2_42[25], stage2_42[26]},
      {stage2_43[2]},
      {stage2_44[12], stage2_44[13], stage2_44[14], stage2_44[15], stage2_44[16], stage2_44[17]},
      {stage3_46[2],stage3_45[2],stage3_44[4],stage3_43[21],stage3_42[34]}
   );
   gpc615_5 gpc7562 (
      {stage2_42[27], stage2_42[28], stage2_42[29], stage2_42[30], stage2_42[31]},
      {stage2_43[3]},
      {stage2_44[18], stage2_44[19], stage2_44[20], stage2_44[21], stage2_44[22], stage2_44[23]},
      {stage3_46[3],stage3_45[3],stage3_44[5],stage3_43[22],stage3_42[35]}
   );
   gpc615_5 gpc7563 (
      {stage2_42[32], stage2_42[33], stage2_42[34], stage2_42[35], stage2_42[36]},
      {stage2_43[4]},
      {stage2_44[24], stage2_44[25], stage2_44[26], stage2_44[27], stage2_44[28], stage2_44[29]},
      {stage3_46[4],stage3_45[4],stage3_44[6],stage3_43[23],stage3_42[36]}
   );
   gpc615_5 gpc7564 (
      {stage2_42[37], stage2_42[38], stage2_42[39], stage2_42[40], stage2_42[41]},
      {stage2_43[5]},
      {stage2_44[30], stage2_44[31], stage2_44[32], stage2_44[33], stage2_44[34], stage2_44[35]},
      {stage3_46[5],stage3_45[5],stage3_44[7],stage3_43[24],stage3_42[37]}
   );
   gpc615_5 gpc7565 (
      {stage2_42[42], stage2_42[43], stage2_42[44], stage2_42[45], stage2_42[46]},
      {stage2_43[6]},
      {stage2_44[36], stage2_44[37], stage2_44[38], stage2_44[39], stage2_44[40], stage2_44[41]},
      {stage3_46[6],stage3_45[6],stage3_44[8],stage3_43[25],stage3_42[38]}
   );
   gpc615_5 gpc7566 (
      {stage2_42[47], stage2_42[48], stage2_42[49], stage2_42[50], stage2_42[51]},
      {stage2_43[7]},
      {stage2_44[42], stage2_44[43], stage2_44[44], stage2_44[45], stage2_44[46], stage2_44[47]},
      {stage3_46[7],stage3_45[7],stage3_44[9],stage3_43[26],stage3_42[39]}
   );
   gpc615_5 gpc7567 (
      {stage2_42[52], stage2_42[53], stage2_42[54], stage2_42[55], stage2_42[56]},
      {stage2_43[8]},
      {stage2_44[48], stage2_44[49], stage2_44[50], stage2_44[51], stage2_44[52], stage2_44[53]},
      {stage3_46[8],stage3_45[8],stage3_44[10],stage3_43[27],stage3_42[40]}
   );
   gpc615_5 gpc7568 (
      {stage2_42[57], stage2_42[58], stage2_42[59], stage2_42[60], stage2_42[61]},
      {stage2_43[9]},
      {stage2_44[54], stage2_44[55], stage2_44[56], stage2_44[57], stage2_44[58], stage2_44[59]},
      {stage3_46[9],stage3_45[9],stage3_44[11],stage3_43[28],stage3_42[41]}
   );
   gpc615_5 gpc7569 (
      {stage2_42[62], stage2_42[63], stage2_42[64], stage2_42[65], stage2_42[66]},
      {stage2_43[10]},
      {stage2_44[60], stage2_44[61], stage2_44[62], stage2_44[63], stage2_44[64], stage2_44[65]},
      {stage3_46[10],stage3_45[10],stage3_44[12],stage3_43[29],stage3_42[42]}
   );
   gpc615_5 gpc7570 (
      {stage2_42[67], stage2_42[68], stage2_42[69], stage2_42[70], stage2_42[71]},
      {stage2_43[11]},
      {stage2_44[66], stage2_44[67], stage2_44[68], stage2_44[69], stage2_44[70], stage2_44[71]},
      {stage3_46[11],stage3_45[11],stage3_44[13],stage3_43[30],stage3_42[43]}
   );
   gpc615_5 gpc7571 (
      {stage2_42[72], stage2_42[73], stage2_42[74], stage2_42[75], stage2_42[76]},
      {stage2_43[12]},
      {stage2_44[72], stage2_44[73], stage2_44[74], stage2_44[75], stage2_44[76], stage2_44[77]},
      {stage3_46[12],stage3_45[12],stage3_44[14],stage3_43[31],stage3_42[44]}
   );
   gpc615_5 gpc7572 (
      {stage2_42[77], stage2_42[78], stage2_42[79], stage2_42[80], stage2_42[81]},
      {stage2_43[13]},
      {stage2_44[78], stage2_44[79], stage2_44[80], stage2_44[81], stage2_44[82], stage2_44[83]},
      {stage3_46[13],stage3_45[13],stage3_44[15],stage3_43[32],stage3_42[45]}
   );
   gpc615_5 gpc7573 (
      {stage2_43[14], stage2_43[15], stage2_43[16], stage2_43[17], stage2_43[18]},
      {stage2_44[84]},
      {stage2_45[0], stage2_45[1], stage2_45[2], stage2_45[3], stage2_45[4], stage2_45[5]},
      {stage3_47[0],stage3_46[14],stage3_45[14],stage3_44[16],stage3_43[33]}
   );
   gpc615_5 gpc7574 (
      {stage2_43[19], stage2_43[20], stage2_43[21], stage2_43[22], stage2_43[23]},
      {stage2_44[85]},
      {stage2_45[6], stage2_45[7], stage2_45[8], stage2_45[9], stage2_45[10], stage2_45[11]},
      {stage3_47[1],stage3_46[15],stage3_45[15],stage3_44[17],stage3_43[34]}
   );
   gpc615_5 gpc7575 (
      {stage2_43[24], stage2_43[25], stage2_43[26], stage2_43[27], stage2_43[28]},
      {stage2_44[86]},
      {stage2_45[12], stage2_45[13], stage2_45[14], stage2_45[15], stage2_45[16], stage2_45[17]},
      {stage3_47[2],stage3_46[16],stage3_45[16],stage3_44[18],stage3_43[35]}
   );
   gpc615_5 gpc7576 (
      {stage2_43[29], stage2_43[30], stage2_43[31], stage2_43[32], stage2_43[33]},
      {stage2_44[87]},
      {stage2_45[18], stage2_45[19], stage2_45[20], stage2_45[21], stage2_45[22], stage2_45[23]},
      {stage3_47[3],stage3_46[17],stage3_45[17],stage3_44[19],stage3_43[36]}
   );
   gpc615_5 gpc7577 (
      {stage2_43[34], stage2_43[35], stage2_43[36], stage2_43[37], stage2_43[38]},
      {stage2_44[88]},
      {stage2_45[24], stage2_45[25], stage2_45[26], stage2_45[27], stage2_45[28], stage2_45[29]},
      {stage3_47[4],stage3_46[18],stage3_45[18],stage3_44[20],stage3_43[37]}
   );
   gpc615_5 gpc7578 (
      {stage2_43[39], stage2_43[40], stage2_43[41], stage2_43[42], stage2_43[43]},
      {stage2_44[89]},
      {stage2_45[30], stage2_45[31], stage2_45[32], stage2_45[33], stage2_45[34], stage2_45[35]},
      {stage3_47[5],stage3_46[19],stage3_45[19],stage3_44[21],stage3_43[38]}
   );
   gpc615_5 gpc7579 (
      {stage2_43[44], stage2_43[45], stage2_43[46], stage2_43[47], stage2_43[48]},
      {stage2_44[90]},
      {stage2_45[36], stage2_45[37], stage2_45[38], stage2_45[39], stage2_45[40], stage2_45[41]},
      {stage3_47[6],stage3_46[20],stage3_45[20],stage3_44[22],stage3_43[39]}
   );
   gpc615_5 gpc7580 (
      {stage2_43[49], stage2_43[50], stage2_43[51], stage2_43[52], stage2_43[53]},
      {stage2_44[91]},
      {stage2_45[42], stage2_45[43], stage2_45[44], stage2_45[45], stage2_45[46], stage2_45[47]},
      {stage3_47[7],stage3_46[21],stage3_45[21],stage3_44[23],stage3_43[40]}
   );
   gpc615_5 gpc7581 (
      {stage2_43[54], stage2_43[55], stage2_43[56], stage2_43[57], stage2_43[58]},
      {stage2_44[92]},
      {stage2_45[48], stage2_45[49], stage2_45[50], stage2_45[51], stage2_45[52], stage2_45[53]},
      {stage3_47[8],stage3_46[22],stage3_45[22],stage3_44[24],stage3_43[41]}
   );
   gpc615_5 gpc7582 (
      {stage2_43[59], stage2_43[60], stage2_43[61], stage2_43[62], stage2_43[63]},
      {stage2_44[93]},
      {stage2_45[54], stage2_45[55], stage2_45[56], stage2_45[57], stage2_45[58], stage2_45[59]},
      {stage3_47[9],stage3_46[23],stage3_45[23],stage3_44[25],stage3_43[42]}
   );
   gpc615_5 gpc7583 (
      {stage2_43[64], stage2_43[65], stage2_43[66], stage2_43[67], stage2_43[68]},
      {stage2_44[94]},
      {stage2_45[60], stage2_45[61], stage2_45[62], stage2_45[63], stage2_45[64], stage2_45[65]},
      {stage3_47[10],stage3_46[24],stage3_45[24],stage3_44[26],stage3_43[43]}
   );
   gpc615_5 gpc7584 (
      {stage2_43[69], stage2_43[70], stage2_43[71], stage2_43[72], stage2_43[73]},
      {stage2_44[95]},
      {stage2_45[66], stage2_45[67], stage2_45[68], stage2_45[69], stage2_45[70], stage2_45[71]},
      {stage3_47[11],stage3_46[25],stage3_45[25],stage3_44[27],stage3_43[44]}
   );
   gpc615_5 gpc7585 (
      {stage2_43[74], stage2_43[75], stage2_43[76], stage2_43[77], stage2_43[78]},
      {stage2_44[96]},
      {stage2_45[72], stage2_45[73], stage2_45[74], stage2_45[75], stage2_45[76], stage2_45[77]},
      {stage3_47[12],stage3_46[26],stage3_45[26],stage3_44[28],stage3_43[45]}
   );
   gpc606_5 gpc7586 (
      {stage2_44[97], stage2_44[98], stage2_44[99], stage2_44[100], stage2_44[101], stage2_44[102]},
      {stage2_46[0], stage2_46[1], stage2_46[2], stage2_46[3], stage2_46[4], stage2_46[5]},
      {stage3_48[0],stage3_47[13],stage3_46[27],stage3_45[27],stage3_44[29]}
   );
   gpc606_5 gpc7587 (
      {stage2_44[103], stage2_44[104], stage2_44[105], stage2_44[106], stage2_44[107], stage2_44[108]},
      {stage2_46[6], stage2_46[7], stage2_46[8], stage2_46[9], stage2_46[10], stage2_46[11]},
      {stage3_48[1],stage3_47[14],stage3_46[28],stage3_45[28],stage3_44[30]}
   );
   gpc606_5 gpc7588 (
      {stage2_45[78], stage2_45[79], stage2_45[80], stage2_45[81], stage2_45[82], stage2_45[83]},
      {stage2_47[0], stage2_47[1], stage2_47[2], stage2_47[3], stage2_47[4], stage2_47[5]},
      {stage3_49[0],stage3_48[2],stage3_47[15],stage3_46[29],stage3_45[29]}
   );
   gpc606_5 gpc7589 (
      {stage2_45[84], stage2_45[85], stage2_45[86], stage2_45[87], stage2_45[88], stage2_45[89]},
      {stage2_47[6], stage2_47[7], stage2_47[8], stage2_47[9], stage2_47[10], stage2_47[11]},
      {stage3_49[1],stage3_48[3],stage3_47[16],stage3_46[30],stage3_45[30]}
   );
   gpc606_5 gpc7590 (
      {stage2_45[90], stage2_45[91], stage2_45[92], stage2_45[93], stage2_45[94], stage2_45[95]},
      {stage2_47[12], stage2_47[13], stage2_47[14], stage2_47[15], stage2_47[16], stage2_47[17]},
      {stage3_49[2],stage3_48[4],stage3_47[17],stage3_46[31],stage3_45[31]}
   );
   gpc606_5 gpc7591 (
      {stage2_45[96], stage2_45[97], stage2_45[98], stage2_45[99], stage2_45[100], stage2_45[101]},
      {stage2_47[18], stage2_47[19], stage2_47[20], stage2_47[21], stage2_47[22], stage2_47[23]},
      {stage3_49[3],stage3_48[5],stage3_47[18],stage3_46[32],stage3_45[32]}
   );
   gpc606_5 gpc7592 (
      {stage2_45[102], stage2_45[103], stage2_45[104], stage2_45[105], stage2_45[106], stage2_45[107]},
      {stage2_47[24], stage2_47[25], stage2_47[26], stage2_47[27], stage2_47[28], stage2_47[29]},
      {stage3_49[4],stage3_48[6],stage3_47[19],stage3_46[33],stage3_45[33]}
   );
   gpc1163_5 gpc7593 (
      {stage2_46[12], stage2_46[13], stage2_46[14]},
      {stage2_47[30], stage2_47[31], stage2_47[32], stage2_47[33], stage2_47[34], stage2_47[35]},
      {stage2_48[0]},
      {stage2_49[0]},
      {stage3_50[0],stage3_49[5],stage3_48[7],stage3_47[20],stage3_46[34]}
   );
   gpc1163_5 gpc7594 (
      {stage2_46[15], stage2_46[16], stage2_46[17]},
      {stage2_47[36], stage2_47[37], stage2_47[38], stage2_47[39], stage2_47[40], stage2_47[41]},
      {stage2_48[1]},
      {stage2_49[1]},
      {stage3_50[1],stage3_49[6],stage3_48[8],stage3_47[21],stage3_46[35]}
   );
   gpc615_5 gpc7595 (
      {stage2_46[18], stage2_46[19], stage2_46[20], stage2_46[21], stage2_46[22]},
      {stage2_47[42]},
      {stage2_48[2], stage2_48[3], stage2_48[4], stage2_48[5], stage2_48[6], stage2_48[7]},
      {stage3_50[2],stage3_49[7],stage3_48[9],stage3_47[22],stage3_46[36]}
   );
   gpc615_5 gpc7596 (
      {stage2_46[23], stage2_46[24], stage2_46[25], stage2_46[26], stage2_46[27]},
      {stage2_47[43]},
      {stage2_48[8], stage2_48[9], stage2_48[10], stage2_48[11], stage2_48[12], stage2_48[13]},
      {stage3_50[3],stage3_49[8],stage3_48[10],stage3_47[23],stage3_46[37]}
   );
   gpc615_5 gpc7597 (
      {stage2_46[28], stage2_46[29], stage2_46[30], stage2_46[31], stage2_46[32]},
      {stage2_47[44]},
      {stage2_48[14], stage2_48[15], stage2_48[16], stage2_48[17], stage2_48[18], stage2_48[19]},
      {stage3_50[4],stage3_49[9],stage3_48[11],stage3_47[24],stage3_46[38]}
   );
   gpc615_5 gpc7598 (
      {stage2_46[33], stage2_46[34], stage2_46[35], stage2_46[36], stage2_46[37]},
      {stage2_47[45]},
      {stage2_48[20], stage2_48[21], stage2_48[22], stage2_48[23], stage2_48[24], stage2_48[25]},
      {stage3_50[5],stage3_49[10],stage3_48[12],stage3_47[25],stage3_46[39]}
   );
   gpc615_5 gpc7599 (
      {stage2_46[38], stage2_46[39], stage2_46[40], stage2_46[41], stage2_46[42]},
      {stage2_47[46]},
      {stage2_48[26], stage2_48[27], stage2_48[28], stage2_48[29], stage2_48[30], stage2_48[31]},
      {stage3_50[6],stage3_49[11],stage3_48[13],stage3_47[26],stage3_46[40]}
   );
   gpc615_5 gpc7600 (
      {stage2_46[43], stage2_46[44], stage2_46[45], stage2_46[46], stage2_46[47]},
      {stage2_47[47]},
      {stage2_48[32], stage2_48[33], stage2_48[34], stage2_48[35], stage2_48[36], stage2_48[37]},
      {stage3_50[7],stage3_49[12],stage3_48[14],stage3_47[27],stage3_46[41]}
   );
   gpc615_5 gpc7601 (
      {stage2_46[48], stage2_46[49], stage2_46[50], stage2_46[51], stage2_46[52]},
      {stage2_47[48]},
      {stage2_48[38], stage2_48[39], stage2_48[40], stage2_48[41], stage2_48[42], stage2_48[43]},
      {stage3_50[8],stage3_49[13],stage3_48[15],stage3_47[28],stage3_46[42]}
   );
   gpc615_5 gpc7602 (
      {stage2_46[53], stage2_46[54], stage2_46[55], stage2_46[56], stage2_46[57]},
      {stage2_47[49]},
      {stage2_48[44], stage2_48[45], stage2_48[46], stage2_48[47], stage2_48[48], stage2_48[49]},
      {stage3_50[9],stage3_49[14],stage3_48[16],stage3_47[29],stage3_46[43]}
   );
   gpc615_5 gpc7603 (
      {stage2_46[58], stage2_46[59], stage2_46[60], stage2_46[61], stage2_46[62]},
      {stage2_47[50]},
      {stage2_48[50], stage2_48[51], stage2_48[52], stage2_48[53], stage2_48[54], stage2_48[55]},
      {stage3_50[10],stage3_49[15],stage3_48[17],stage3_47[30],stage3_46[44]}
   );
   gpc615_5 gpc7604 (
      {stage2_46[63], stage2_46[64], stage2_46[65], stage2_46[66], stage2_46[67]},
      {stage2_47[51]},
      {stage2_48[56], stage2_48[57], stage2_48[58], stage2_48[59], stage2_48[60], stage2_48[61]},
      {stage3_50[11],stage3_49[16],stage3_48[18],stage3_47[31],stage3_46[45]}
   );
   gpc615_5 gpc7605 (
      {stage2_46[68], stage2_46[69], stage2_46[70], stage2_46[71], stage2_46[72]},
      {stage2_47[52]},
      {stage2_48[62], stage2_48[63], stage2_48[64], stage2_48[65], stage2_48[66], stage2_48[67]},
      {stage3_50[12],stage3_49[17],stage3_48[19],stage3_47[32],stage3_46[46]}
   );
   gpc615_5 gpc7606 (
      {stage2_46[73], stage2_46[74], stage2_46[75], stage2_46[76], stage2_46[77]},
      {stage2_47[53]},
      {stage2_48[68], stage2_48[69], stage2_48[70], stage2_48[71], stage2_48[72], stage2_48[73]},
      {stage3_50[13],stage3_49[18],stage3_48[20],stage3_47[33],stage3_46[47]}
   );
   gpc615_5 gpc7607 (
      {stage2_47[54], stage2_47[55], stage2_47[56], stage2_47[57], stage2_47[58]},
      {stage2_48[74]},
      {stage2_49[2], stage2_49[3], stage2_49[4], stage2_49[5], stage2_49[6], stage2_49[7]},
      {stage3_51[0],stage3_50[14],stage3_49[19],stage3_48[21],stage3_47[34]}
   );
   gpc615_5 gpc7608 (
      {stage2_47[59], stage2_47[60], stage2_47[61], stage2_47[62], stage2_47[63]},
      {stage2_48[75]},
      {stage2_49[8], stage2_49[9], stage2_49[10], stage2_49[11], stage2_49[12], stage2_49[13]},
      {stage3_51[1],stage3_50[15],stage3_49[20],stage3_48[22],stage3_47[35]}
   );
   gpc615_5 gpc7609 (
      {stage2_47[64], stage2_47[65], stage2_47[66], stage2_47[67], stage2_47[68]},
      {stage2_48[76]},
      {stage2_49[14], stage2_49[15], stage2_49[16], stage2_49[17], stage2_49[18], stage2_49[19]},
      {stage3_51[2],stage3_50[16],stage3_49[21],stage3_48[23],stage3_47[36]}
   );
   gpc615_5 gpc7610 (
      {stage2_47[69], stage2_47[70], stage2_47[71], stage2_47[72], stage2_47[73]},
      {stage2_48[77]},
      {stage2_49[20], stage2_49[21], stage2_49[22], stage2_49[23], stage2_49[24], stage2_49[25]},
      {stage3_51[3],stage3_50[17],stage3_49[22],stage3_48[24],stage3_47[37]}
   );
   gpc615_5 gpc7611 (
      {stage2_47[74], stage2_47[75], stage2_47[76], stage2_47[77], stage2_47[78]},
      {stage2_48[78]},
      {stage2_49[26], stage2_49[27], stage2_49[28], stage2_49[29], stage2_49[30], stage2_49[31]},
      {stage3_51[4],stage3_50[18],stage3_49[23],stage3_48[25],stage3_47[38]}
   );
   gpc615_5 gpc7612 (
      {stage2_47[79], stage2_47[80], stage2_47[81], stage2_47[82], stage2_47[83]},
      {stage2_48[79]},
      {stage2_49[32], stage2_49[33], stage2_49[34], stage2_49[35], stage2_49[36], stage2_49[37]},
      {stage3_51[5],stage3_50[19],stage3_49[24],stage3_48[26],stage3_47[39]}
   );
   gpc615_5 gpc7613 (
      {stage2_47[84], stage2_47[85], stage2_47[86], stage2_47[87], stage2_47[88]},
      {stage2_48[80]},
      {stage2_49[38], stage2_49[39], stage2_49[40], stage2_49[41], stage2_49[42], stage2_49[43]},
      {stage3_51[6],stage3_50[20],stage3_49[25],stage3_48[27],stage3_47[40]}
   );
   gpc615_5 gpc7614 (
      {stage2_47[89], stage2_47[90], stage2_47[91], stage2_47[92], stage2_47[93]},
      {stage2_48[81]},
      {stage2_49[44], stage2_49[45], stage2_49[46], stage2_49[47], stage2_49[48], stage2_49[49]},
      {stage3_51[7],stage3_50[21],stage3_49[26],stage3_48[28],stage3_47[41]}
   );
   gpc615_5 gpc7615 (
      {stage2_47[94], stage2_47[95], stage2_47[96], stage2_47[97], stage2_47[98]},
      {stage2_48[82]},
      {stage2_49[50], stage2_49[51], stage2_49[52], stage2_49[53], stage2_49[54], stage2_49[55]},
      {stage3_51[8],stage3_50[22],stage3_49[27],stage3_48[29],stage3_47[42]}
   );
   gpc615_5 gpc7616 (
      {stage2_47[99], stage2_47[100], stage2_47[101], stage2_47[102], stage2_47[103]},
      {stage2_48[83]},
      {stage2_49[56], stage2_49[57], stage2_49[58], stage2_49[59], stage2_49[60], stage2_49[61]},
      {stage3_51[9],stage3_50[23],stage3_49[28],stage3_48[30],stage3_47[43]}
   );
   gpc606_5 gpc7617 (
      {stage2_48[84], stage2_48[85], stage2_48[86], stage2_48[87], stage2_48[88], stage2_48[89]},
      {stage2_50[0], stage2_50[1], stage2_50[2], stage2_50[3], stage2_50[4], stage2_50[5]},
      {stage3_52[0],stage3_51[10],stage3_50[24],stage3_49[29],stage3_48[31]}
   );
   gpc606_5 gpc7618 (
      {stage2_48[90], stage2_48[91], stage2_48[92], stage2_48[93], stage2_48[94], stage2_48[95]},
      {stage2_50[6], stage2_50[7], stage2_50[8], stage2_50[9], stage2_50[10], stage2_50[11]},
      {stage3_52[1],stage3_51[11],stage3_50[25],stage3_49[30],stage3_48[32]}
   );
   gpc606_5 gpc7619 (
      {stage2_48[96], stage2_48[97], stage2_48[98], stage2_48[99], stage2_48[100], stage2_48[101]},
      {stage2_50[12], stage2_50[13], stage2_50[14], stage2_50[15], stage2_50[16], stage2_50[17]},
      {stage3_52[2],stage3_51[12],stage3_50[26],stage3_49[31],stage3_48[33]}
   );
   gpc606_5 gpc7620 (
      {stage2_48[102], stage2_48[103], stage2_48[104], stage2_48[105], stage2_48[106], stage2_48[107]},
      {stage2_50[18], stage2_50[19], stage2_50[20], stage2_50[21], stage2_50[22], stage2_50[23]},
      {stage3_52[3],stage3_51[13],stage3_50[27],stage3_49[32],stage3_48[34]}
   );
   gpc606_5 gpc7621 (
      {stage2_48[108], stage2_48[109], stage2_48[110], stage2_48[111], stage2_48[112], stage2_48[113]},
      {stage2_50[24], stage2_50[25], stage2_50[26], stage2_50[27], stage2_50[28], stage2_50[29]},
      {stage3_52[4],stage3_51[14],stage3_50[28],stage3_49[33],stage3_48[35]}
   );
   gpc606_5 gpc7622 (
      {stage2_48[114], stage2_48[115], stage2_48[116], stage2_48[117], stage2_48[118], stage2_48[119]},
      {stage2_50[30], stage2_50[31], stage2_50[32], stage2_50[33], stage2_50[34], stage2_50[35]},
      {stage3_52[5],stage3_51[15],stage3_50[29],stage3_49[34],stage3_48[36]}
   );
   gpc606_5 gpc7623 (
      {stage2_48[120], stage2_48[121], stage2_48[122], stage2_48[123], stage2_48[124], stage2_48[125]},
      {stage2_50[36], stage2_50[37], stage2_50[38], stage2_50[39], stage2_50[40], stage2_50[41]},
      {stage3_52[6],stage3_51[16],stage3_50[30],stage3_49[35],stage3_48[37]}
   );
   gpc606_5 gpc7624 (
      {stage2_49[62], stage2_49[63], stage2_49[64], stage2_49[65], stage2_49[66], stage2_49[67]},
      {stage2_51[0], stage2_51[1], stage2_51[2], stage2_51[3], stage2_51[4], stage2_51[5]},
      {stage3_53[0],stage3_52[7],stage3_51[17],stage3_50[31],stage3_49[36]}
   );
   gpc606_5 gpc7625 (
      {stage2_49[68], stage2_49[69], stage2_49[70], stage2_49[71], stage2_49[72], stage2_49[73]},
      {stage2_51[6], stage2_51[7], stage2_51[8], stage2_51[9], stage2_51[10], stage2_51[11]},
      {stage3_53[1],stage3_52[8],stage3_51[18],stage3_50[32],stage3_49[37]}
   );
   gpc606_5 gpc7626 (
      {stage2_49[74], stage2_49[75], stage2_49[76], stage2_49[77], stage2_49[78], stage2_49[79]},
      {stage2_51[12], stage2_51[13], stage2_51[14], stage2_51[15], stage2_51[16], stage2_51[17]},
      {stage3_53[2],stage3_52[9],stage3_51[19],stage3_50[33],stage3_49[38]}
   );
   gpc606_5 gpc7627 (
      {stage2_49[80], stage2_49[81], stage2_49[82], stage2_49[83], stage2_49[84], stage2_49[85]},
      {stage2_51[18], stage2_51[19], stage2_51[20], stage2_51[21], stage2_51[22], stage2_51[23]},
      {stage3_53[3],stage3_52[10],stage3_51[20],stage3_50[34],stage3_49[39]}
   );
   gpc615_5 gpc7628 (
      {stage2_49[86], stage2_49[87], stage2_49[88], stage2_49[89], stage2_49[90]},
      {stage2_50[42]},
      {stage2_51[24], stage2_51[25], stage2_51[26], stage2_51[27], stage2_51[28], stage2_51[29]},
      {stage3_53[4],stage3_52[11],stage3_51[21],stage3_50[35],stage3_49[40]}
   );
   gpc615_5 gpc7629 (
      {stage2_49[91], stage2_49[92], stage2_49[93], stage2_49[94], stage2_49[95]},
      {stage2_50[43]},
      {stage2_51[30], stage2_51[31], stage2_51[32], stage2_51[33], stage2_51[34], stage2_51[35]},
      {stage3_53[5],stage3_52[12],stage3_51[22],stage3_50[36],stage3_49[41]}
   );
   gpc615_5 gpc7630 (
      {stage2_50[44], stage2_50[45], stage2_50[46], stage2_50[47], stage2_50[48]},
      {stage2_51[36]},
      {stage2_52[0], stage2_52[1], stage2_52[2], stage2_52[3], stage2_52[4], stage2_52[5]},
      {stage3_54[0],stage3_53[6],stage3_52[13],stage3_51[23],stage3_50[37]}
   );
   gpc615_5 gpc7631 (
      {stage2_50[49], stage2_50[50], stage2_50[51], stage2_50[52], stage2_50[53]},
      {stage2_51[37]},
      {stage2_52[6], stage2_52[7], stage2_52[8], stage2_52[9], stage2_52[10], stage2_52[11]},
      {stage3_54[1],stage3_53[7],stage3_52[14],stage3_51[24],stage3_50[38]}
   );
   gpc615_5 gpc7632 (
      {stage2_50[54], stage2_50[55], stage2_50[56], stage2_50[57], stage2_50[58]},
      {stage2_51[38]},
      {stage2_52[12], stage2_52[13], stage2_52[14], stage2_52[15], stage2_52[16], stage2_52[17]},
      {stage3_54[2],stage3_53[8],stage3_52[15],stage3_51[25],stage3_50[39]}
   );
   gpc615_5 gpc7633 (
      {stage2_50[59], stage2_50[60], stage2_50[61], stage2_50[62], stage2_50[63]},
      {stage2_51[39]},
      {stage2_52[18], stage2_52[19], stage2_52[20], stage2_52[21], stage2_52[22], stage2_52[23]},
      {stage3_54[3],stage3_53[9],stage3_52[16],stage3_51[26],stage3_50[40]}
   );
   gpc615_5 gpc7634 (
      {stage2_50[64], stage2_50[65], stage2_50[66], stage2_50[67], stage2_50[68]},
      {stage2_51[40]},
      {stage2_52[24], stage2_52[25], stage2_52[26], stage2_52[27], stage2_52[28], stage2_52[29]},
      {stage3_54[4],stage3_53[10],stage3_52[17],stage3_51[27],stage3_50[41]}
   );
   gpc615_5 gpc7635 (
      {stage2_50[69], stage2_50[70], stage2_50[71], stage2_50[72], stage2_50[73]},
      {stage2_51[41]},
      {stage2_52[30], stage2_52[31], stage2_52[32], stage2_52[33], stage2_52[34], stage2_52[35]},
      {stage3_54[5],stage3_53[11],stage3_52[18],stage3_51[28],stage3_50[42]}
   );
   gpc615_5 gpc7636 (
      {stage2_50[74], stage2_50[75], stage2_50[76], stage2_50[77], stage2_50[78]},
      {stage2_51[42]},
      {stage2_52[36], stage2_52[37], stage2_52[38], stage2_52[39], stage2_52[40], stage2_52[41]},
      {stage3_54[6],stage3_53[12],stage3_52[19],stage3_51[29],stage3_50[43]}
   );
   gpc615_5 gpc7637 (
      {stage2_50[79], stage2_50[80], stage2_50[81], stage2_50[82], stage2_50[83]},
      {stage2_51[43]},
      {stage2_52[42], stage2_52[43], stage2_52[44], stage2_52[45], stage2_52[46], stage2_52[47]},
      {stage3_54[7],stage3_53[13],stage3_52[20],stage3_51[30],stage3_50[44]}
   );
   gpc615_5 gpc7638 (
      {stage2_51[44], stage2_51[45], stage2_51[46], stage2_51[47], stage2_51[48]},
      {stage2_52[48]},
      {stage2_53[0], stage2_53[1], stage2_53[2], stage2_53[3], stage2_53[4], stage2_53[5]},
      {stage3_55[0],stage3_54[8],stage3_53[14],stage3_52[21],stage3_51[31]}
   );
   gpc615_5 gpc7639 (
      {stage2_51[49], stage2_51[50], stage2_51[51], stage2_51[52], stage2_51[53]},
      {stage2_52[49]},
      {stage2_53[6], stage2_53[7], stage2_53[8], stage2_53[9], stage2_53[10], stage2_53[11]},
      {stage3_55[1],stage3_54[9],stage3_53[15],stage3_52[22],stage3_51[32]}
   );
   gpc615_5 gpc7640 (
      {stage2_51[54], stage2_51[55], stage2_51[56], stage2_51[57], stage2_51[58]},
      {stage2_52[50]},
      {stage2_53[12], stage2_53[13], stage2_53[14], stage2_53[15], stage2_53[16], stage2_53[17]},
      {stage3_55[2],stage3_54[10],stage3_53[16],stage3_52[23],stage3_51[33]}
   );
   gpc606_5 gpc7641 (
      {stage2_52[51], stage2_52[52], stage2_52[53], stage2_52[54], stage2_52[55], stage2_52[56]},
      {stage2_54[0], stage2_54[1], stage2_54[2], stage2_54[3], stage2_54[4], stage2_54[5]},
      {stage3_56[0],stage3_55[3],stage3_54[11],stage3_53[17],stage3_52[24]}
   );
   gpc606_5 gpc7642 (
      {stage2_52[57], stage2_52[58], stage2_52[59], stage2_52[60], stage2_52[61], stage2_52[62]},
      {stage2_54[6], stage2_54[7], stage2_54[8], stage2_54[9], stage2_54[10], stage2_54[11]},
      {stage3_56[1],stage3_55[4],stage3_54[12],stage3_53[18],stage3_52[25]}
   );
   gpc606_5 gpc7643 (
      {stage2_52[63], stage2_52[64], stage2_52[65], stage2_52[66], stage2_52[67], stage2_52[68]},
      {stage2_54[12], stage2_54[13], stage2_54[14], stage2_54[15], stage2_54[16], stage2_54[17]},
      {stage3_56[2],stage3_55[5],stage3_54[13],stage3_53[19],stage3_52[26]}
   );
   gpc606_5 gpc7644 (
      {stage2_53[18], stage2_53[19], stage2_53[20], stage2_53[21], stage2_53[22], stage2_53[23]},
      {stage2_55[0], stage2_55[1], stage2_55[2], stage2_55[3], stage2_55[4], stage2_55[5]},
      {stage3_57[0],stage3_56[3],stage3_55[6],stage3_54[14],stage3_53[20]}
   );
   gpc606_5 gpc7645 (
      {stage2_53[24], stage2_53[25], stage2_53[26], stage2_53[27], stage2_53[28], stage2_53[29]},
      {stage2_55[6], stage2_55[7], stage2_55[8], stage2_55[9], stage2_55[10], stage2_55[11]},
      {stage3_57[1],stage3_56[4],stage3_55[7],stage3_54[15],stage3_53[21]}
   );
   gpc606_5 gpc7646 (
      {stage2_53[30], stage2_53[31], stage2_53[32], stage2_53[33], stage2_53[34], stage2_53[35]},
      {stage2_55[12], stage2_55[13], stage2_55[14], stage2_55[15], stage2_55[16], stage2_55[17]},
      {stage3_57[2],stage3_56[5],stage3_55[8],stage3_54[16],stage3_53[22]}
   );
   gpc606_5 gpc7647 (
      {stage2_53[36], stage2_53[37], stage2_53[38], stage2_53[39], stage2_53[40], stage2_53[41]},
      {stage2_55[18], stage2_55[19], stage2_55[20], stage2_55[21], stage2_55[22], stage2_55[23]},
      {stage3_57[3],stage3_56[6],stage3_55[9],stage3_54[17],stage3_53[23]}
   );
   gpc606_5 gpc7648 (
      {stage2_53[42], stage2_53[43], stage2_53[44], stage2_53[45], stage2_53[46], stage2_53[47]},
      {stage2_55[24], stage2_55[25], stage2_55[26], stage2_55[27], stage2_55[28], stage2_55[29]},
      {stage3_57[4],stage3_56[7],stage3_55[10],stage3_54[18],stage3_53[24]}
   );
   gpc606_5 gpc7649 (
      {stage2_53[48], stage2_53[49], stage2_53[50], stage2_53[51], stage2_53[52], stage2_53[53]},
      {stage2_55[30], stage2_55[31], stage2_55[32], stage2_55[33], stage2_55[34], stage2_55[35]},
      {stage3_57[5],stage3_56[8],stage3_55[11],stage3_54[19],stage3_53[25]}
   );
   gpc615_5 gpc7650 (
      {stage2_53[54], stage2_53[55], stage2_53[56], stage2_53[57], stage2_53[58]},
      {stage2_54[18]},
      {stage2_55[36], stage2_55[37], stage2_55[38], stage2_55[39], stage2_55[40], stage2_55[41]},
      {stage3_57[6],stage3_56[9],stage3_55[12],stage3_54[20],stage3_53[26]}
   );
   gpc615_5 gpc7651 (
      {stage2_53[59], stage2_53[60], stage2_53[61], stage2_53[62], stage2_53[63]},
      {stage2_54[19]},
      {stage2_55[42], stage2_55[43], stage2_55[44], stage2_55[45], stage2_55[46], stage2_55[47]},
      {stage3_57[7],stage3_56[10],stage3_55[13],stage3_54[21],stage3_53[27]}
   );
   gpc615_5 gpc7652 (
      {stage2_53[64], stage2_53[65], stage2_53[66], stage2_53[67], stage2_53[68]},
      {stage2_54[20]},
      {stage2_55[48], stage2_55[49], stage2_55[50], stage2_55[51], stage2_55[52], stage2_55[53]},
      {stage3_57[8],stage3_56[11],stage3_55[14],stage3_54[22],stage3_53[28]}
   );
   gpc615_5 gpc7653 (
      {stage2_54[21], stage2_54[22], stage2_54[23], stage2_54[24], stage2_54[25]},
      {stage2_55[54]},
      {stage2_56[0], stage2_56[1], stage2_56[2], stage2_56[3], stage2_56[4], stage2_56[5]},
      {stage3_58[0],stage3_57[9],stage3_56[12],stage3_55[15],stage3_54[23]}
   );
   gpc615_5 gpc7654 (
      {stage2_54[26], stage2_54[27], stage2_54[28], stage2_54[29], stage2_54[30]},
      {stage2_55[55]},
      {stage2_56[6], stage2_56[7], stage2_56[8], stage2_56[9], stage2_56[10], stage2_56[11]},
      {stage3_58[1],stage3_57[10],stage3_56[13],stage3_55[16],stage3_54[24]}
   );
   gpc615_5 gpc7655 (
      {stage2_54[31], stage2_54[32], stage2_54[33], stage2_54[34], stage2_54[35]},
      {stage2_55[56]},
      {stage2_56[12], stage2_56[13], stage2_56[14], stage2_56[15], stage2_56[16], stage2_56[17]},
      {stage3_58[2],stage3_57[11],stage3_56[14],stage3_55[17],stage3_54[25]}
   );
   gpc615_5 gpc7656 (
      {stage2_54[36], stage2_54[37], stage2_54[38], stage2_54[39], stage2_54[40]},
      {stage2_55[57]},
      {stage2_56[18], stage2_56[19], stage2_56[20], stage2_56[21], stage2_56[22], stage2_56[23]},
      {stage3_58[3],stage3_57[12],stage3_56[15],stage3_55[18],stage3_54[26]}
   );
   gpc615_5 gpc7657 (
      {stage2_54[41], stage2_54[42], stage2_54[43], stage2_54[44], stage2_54[45]},
      {stage2_55[58]},
      {stage2_56[24], stage2_56[25], stage2_56[26], stage2_56[27], stage2_56[28], stage2_56[29]},
      {stage3_58[4],stage3_57[13],stage3_56[16],stage3_55[19],stage3_54[27]}
   );
   gpc615_5 gpc7658 (
      {stage2_54[46], stage2_54[47], stage2_54[48], stage2_54[49], stage2_54[50]},
      {stage2_55[59]},
      {stage2_56[30], stage2_56[31], stage2_56[32], stage2_56[33], stage2_56[34], stage2_56[35]},
      {stage3_58[5],stage3_57[14],stage3_56[17],stage3_55[20],stage3_54[28]}
   );
   gpc615_5 gpc7659 (
      {stage2_54[51], stage2_54[52], stage2_54[53], stage2_54[54], stage2_54[55]},
      {stage2_55[60]},
      {stage2_56[36], stage2_56[37], stage2_56[38], stage2_56[39], stage2_56[40], stage2_56[41]},
      {stage3_58[6],stage3_57[15],stage3_56[18],stage3_55[21],stage3_54[29]}
   );
   gpc615_5 gpc7660 (
      {stage2_54[56], stage2_54[57], stage2_54[58], stage2_54[59], stage2_54[60]},
      {stage2_55[61]},
      {stage2_56[42], stage2_56[43], stage2_56[44], stage2_56[45], stage2_56[46], stage2_56[47]},
      {stage3_58[7],stage3_57[16],stage3_56[19],stage3_55[22],stage3_54[30]}
   );
   gpc615_5 gpc7661 (
      {stage2_54[61], stage2_54[62], stage2_54[63], stage2_54[64], stage2_54[65]},
      {stage2_55[62]},
      {stage2_56[48], stage2_56[49], stage2_56[50], stage2_56[51], stage2_56[52], stage2_56[53]},
      {stage3_58[8],stage3_57[17],stage3_56[20],stage3_55[23],stage3_54[31]}
   );
   gpc615_5 gpc7662 (
      {stage2_54[66], stage2_54[67], stage2_54[68], stage2_54[69], stage2_54[70]},
      {stage2_55[63]},
      {stage2_56[54], stage2_56[55], stage2_56[56], stage2_56[57], stage2_56[58], stage2_56[59]},
      {stage3_58[9],stage3_57[18],stage3_56[21],stage3_55[24],stage3_54[32]}
   );
   gpc615_5 gpc7663 (
      {stage2_54[71], stage2_54[72], stage2_54[73], stage2_54[74], stage2_54[75]},
      {stage2_55[64]},
      {stage2_56[60], stage2_56[61], stage2_56[62], stage2_56[63], stage2_56[64], stage2_56[65]},
      {stage3_58[10],stage3_57[19],stage3_56[22],stage3_55[25],stage3_54[33]}
   );
   gpc615_5 gpc7664 (
      {stage2_54[76], stage2_54[77], stage2_54[78], stage2_54[79], stage2_54[80]},
      {stage2_55[65]},
      {stage2_56[66], stage2_56[67], stage2_56[68], stage2_56[69], stage2_56[70], stage2_56[71]},
      {stage3_58[11],stage3_57[20],stage3_56[23],stage3_55[26],stage3_54[34]}
   );
   gpc615_5 gpc7665 (
      {stage2_54[81], stage2_54[82], stage2_54[83], stage2_54[84], stage2_54[85]},
      {stage2_55[66]},
      {stage2_56[72], stage2_56[73], stage2_56[74], stage2_56[75], stage2_56[76], stage2_56[77]},
      {stage3_58[12],stage3_57[21],stage3_56[24],stage3_55[27],stage3_54[35]}
   );
   gpc615_5 gpc7666 (
      {stage2_54[86], stage2_54[87], stage2_54[88], stage2_54[89], stage2_54[90]},
      {stage2_55[67]},
      {stage2_56[78], stage2_56[79], stage2_56[80], stage2_56[81], stage2_56[82], stage2_56[83]},
      {stage3_58[13],stage3_57[22],stage3_56[25],stage3_55[28],stage3_54[36]}
   );
   gpc615_5 gpc7667 (
      {stage2_54[91], stage2_54[92], stage2_54[93], stage2_54[94], stage2_54[95]},
      {stage2_55[68]},
      {stage2_56[84], stage2_56[85], stage2_56[86], stage2_56[87], stage2_56[88], stage2_56[89]},
      {stage3_58[14],stage3_57[23],stage3_56[26],stage3_55[29],stage3_54[37]}
   );
   gpc615_5 gpc7668 (
      {stage2_54[96], stage2_54[97], stage2_54[98], stage2_54[99], 1'b0},
      {stage2_55[69]},
      {stage2_56[90], stage2_56[91], stage2_56[92], stage2_56[93], stage2_56[94], stage2_56[95]},
      {stage3_58[15],stage3_57[24],stage3_56[27],stage3_55[30],stage3_54[38]}
   );
   gpc615_5 gpc7669 (
      {stage2_56[96], stage2_56[97], stage2_56[98], stage2_56[99], stage2_56[100]},
      {stage2_57[0]},
      {stage2_58[0], stage2_58[1], stage2_58[2], stage2_58[3], stage2_58[4], stage2_58[5]},
      {stage3_60[0],stage3_59[0],stage3_58[16],stage3_57[25],stage3_56[28]}
   );
   gpc615_5 gpc7670 (
      {stage2_56[101], stage2_56[102], stage2_56[103], stage2_56[104], stage2_56[105]},
      {stage2_57[1]},
      {stage2_58[6], stage2_58[7], stage2_58[8], stage2_58[9], stage2_58[10], stage2_58[11]},
      {stage3_60[1],stage3_59[1],stage3_58[17],stage3_57[26],stage3_56[29]}
   );
   gpc615_5 gpc7671 (
      {stage2_56[106], stage2_56[107], stage2_56[108], stage2_56[109], stage2_56[110]},
      {stage2_57[2]},
      {stage2_58[12], stage2_58[13], stage2_58[14], stage2_58[15], stage2_58[16], stage2_58[17]},
      {stage3_60[2],stage3_59[2],stage3_58[18],stage3_57[27],stage3_56[30]}
   );
   gpc615_5 gpc7672 (
      {stage2_56[111], stage2_56[112], stage2_56[113], stage2_56[114], 1'b0},
      {stage2_57[3]},
      {stage2_58[18], stage2_58[19], stage2_58[20], stage2_58[21], stage2_58[22], stage2_58[23]},
      {stage3_60[3],stage3_59[3],stage3_58[19],stage3_57[28],stage3_56[31]}
   );
   gpc207_4 gpc7673 (
      {stage2_57[4], stage2_57[5], stage2_57[6], stage2_57[7], stage2_57[8], stage2_57[9], stage2_57[10]},
      {stage2_59[0], stage2_59[1]},
      {stage3_60[4],stage3_59[4],stage3_58[20],stage3_57[29]}
   );
   gpc606_5 gpc7674 (
      {stage2_57[11], stage2_57[12], stage2_57[13], stage2_57[14], stage2_57[15], stage2_57[16]},
      {stage2_59[2], stage2_59[3], stage2_59[4], stage2_59[5], stage2_59[6], stage2_59[7]},
      {stage3_61[0],stage3_60[5],stage3_59[5],stage3_58[21],stage3_57[30]}
   );
   gpc606_5 gpc7675 (
      {stage2_57[17], stage2_57[18], stage2_57[19], stage2_57[20], stage2_57[21], stage2_57[22]},
      {stage2_59[8], stage2_59[9], stage2_59[10], stage2_59[11], stage2_59[12], stage2_59[13]},
      {stage3_61[1],stage3_60[6],stage3_59[6],stage3_58[22],stage3_57[31]}
   );
   gpc606_5 gpc7676 (
      {stage2_57[23], stage2_57[24], stage2_57[25], stage2_57[26], stage2_57[27], stage2_57[28]},
      {stage2_59[14], stage2_59[15], stage2_59[16], stage2_59[17], stage2_59[18], stage2_59[19]},
      {stage3_61[2],stage3_60[7],stage3_59[7],stage3_58[23],stage3_57[32]}
   );
   gpc615_5 gpc7677 (
      {stage2_57[29], stage2_57[30], stage2_57[31], stage2_57[32], stage2_57[33]},
      {stage2_58[24]},
      {stage2_59[20], stage2_59[21], stage2_59[22], stage2_59[23], stage2_59[24], stage2_59[25]},
      {stage3_61[3],stage3_60[8],stage3_59[8],stage3_58[24],stage3_57[33]}
   );
   gpc615_5 gpc7678 (
      {stage2_57[34], stage2_57[35], stage2_57[36], stage2_57[37], stage2_57[38]},
      {stage2_58[25]},
      {stage2_59[26], stage2_59[27], stage2_59[28], stage2_59[29], stage2_59[30], stage2_59[31]},
      {stage3_61[4],stage3_60[9],stage3_59[9],stage3_58[25],stage3_57[34]}
   );
   gpc615_5 gpc7679 (
      {stage2_57[39], stage2_57[40], stage2_57[41], stage2_57[42], stage2_57[43]},
      {stage2_58[26]},
      {stage2_59[32], stage2_59[33], stage2_59[34], stage2_59[35], stage2_59[36], stage2_59[37]},
      {stage3_61[5],stage3_60[10],stage3_59[10],stage3_58[26],stage3_57[35]}
   );
   gpc615_5 gpc7680 (
      {stage2_57[44], stage2_57[45], stage2_57[46], stage2_57[47], stage2_57[48]},
      {stage2_58[27]},
      {stage2_59[38], stage2_59[39], stage2_59[40], stage2_59[41], stage2_59[42], stage2_59[43]},
      {stage3_61[6],stage3_60[11],stage3_59[11],stage3_58[27],stage3_57[36]}
   );
   gpc615_5 gpc7681 (
      {stage2_58[28], stage2_58[29], stage2_58[30], stage2_58[31], stage2_58[32]},
      {stage2_59[44]},
      {stage2_60[0], stage2_60[1], stage2_60[2], stage2_60[3], stage2_60[4], stage2_60[5]},
      {stage3_62[0],stage3_61[7],stage3_60[12],stage3_59[12],stage3_58[28]}
   );
   gpc615_5 gpc7682 (
      {stage2_58[33], stage2_58[34], stage2_58[35], stage2_58[36], stage2_58[37]},
      {stage2_59[45]},
      {stage2_60[6], stage2_60[7], stage2_60[8], stage2_60[9], stage2_60[10], stage2_60[11]},
      {stage3_62[1],stage3_61[8],stage3_60[13],stage3_59[13],stage3_58[29]}
   );
   gpc615_5 gpc7683 (
      {stage2_58[38], stage2_58[39], stage2_58[40], stage2_58[41], stage2_58[42]},
      {stage2_59[46]},
      {stage2_60[12], stage2_60[13], stage2_60[14], stage2_60[15], stage2_60[16], stage2_60[17]},
      {stage3_62[2],stage3_61[9],stage3_60[14],stage3_59[14],stage3_58[30]}
   );
   gpc615_5 gpc7684 (
      {stage2_58[43], stage2_58[44], stage2_58[45], stage2_58[46], stage2_58[47]},
      {stage2_59[47]},
      {stage2_60[18], stage2_60[19], stage2_60[20], stage2_60[21], stage2_60[22], stage2_60[23]},
      {stage3_62[3],stage3_61[10],stage3_60[15],stage3_59[15],stage3_58[31]}
   );
   gpc615_5 gpc7685 (
      {stage2_58[48], stage2_58[49], stage2_58[50], stage2_58[51], stage2_58[52]},
      {stage2_59[48]},
      {stage2_60[24], stage2_60[25], stage2_60[26], stage2_60[27], stage2_60[28], stage2_60[29]},
      {stage3_62[4],stage3_61[11],stage3_60[16],stage3_59[16],stage3_58[32]}
   );
   gpc615_5 gpc7686 (
      {stage2_58[53], stage2_58[54], stage2_58[55], stage2_58[56], stage2_58[57]},
      {stage2_59[49]},
      {stage2_60[30], stage2_60[31], stage2_60[32], stage2_60[33], stage2_60[34], stage2_60[35]},
      {stage3_62[5],stage3_61[12],stage3_60[17],stage3_59[17],stage3_58[33]}
   );
   gpc615_5 gpc7687 (
      {stage2_59[50], stage2_59[51], stage2_59[52], stage2_59[53], stage2_59[54]},
      {stage2_60[36]},
      {stage2_61[0], stage2_61[1], stage2_61[2], stage2_61[3], stage2_61[4], stage2_61[5]},
      {stage3_63[0],stage3_62[6],stage3_61[13],stage3_60[18],stage3_59[18]}
   );
   gpc615_5 gpc7688 (
      {stage2_59[55], stage2_59[56], stage2_59[57], stage2_59[58], stage2_59[59]},
      {stage2_60[37]},
      {stage2_61[6], stage2_61[7], stage2_61[8], stage2_61[9], stage2_61[10], stage2_61[11]},
      {stage3_63[1],stage3_62[7],stage3_61[14],stage3_60[19],stage3_59[19]}
   );
   gpc615_5 gpc7689 (
      {stage2_59[60], stage2_59[61], stage2_59[62], stage2_59[63], stage2_59[64]},
      {stage2_60[38]},
      {stage2_61[12], stage2_61[13], stage2_61[14], stage2_61[15], stage2_61[16], stage2_61[17]},
      {stage3_63[2],stage3_62[8],stage3_61[15],stage3_60[20],stage3_59[20]}
   );
   gpc615_5 gpc7690 (
      {stage2_59[65], stage2_59[66], stage2_59[67], stage2_59[68], stage2_59[69]},
      {stage2_60[39]},
      {stage2_61[18], stage2_61[19], stage2_61[20], stage2_61[21], stage2_61[22], stage2_61[23]},
      {stage3_63[3],stage3_62[9],stage3_61[16],stage3_60[21],stage3_59[21]}
   );
   gpc615_5 gpc7691 (
      {stage2_59[70], stage2_59[71], stage2_59[72], stage2_59[73], stage2_59[74]},
      {stage2_60[40]},
      {stage2_61[24], stage2_61[25], stage2_61[26], stage2_61[27], stage2_61[28], stage2_61[29]},
      {stage3_63[4],stage3_62[10],stage3_61[17],stage3_60[22],stage3_59[22]}
   );
   gpc615_5 gpc7692 (
      {stage2_59[75], stage2_59[76], stage2_59[77], stage2_59[78], stage2_59[79]},
      {stage2_60[41]},
      {stage2_61[30], stage2_61[31], stage2_61[32], stage2_61[33], stage2_61[34], stage2_61[35]},
      {stage3_63[5],stage3_62[11],stage3_61[18],stage3_60[23],stage3_59[23]}
   );
   gpc615_5 gpc7693 (
      {stage2_59[80], stage2_59[81], stage2_59[82], stage2_59[83], stage2_59[84]},
      {stage2_60[42]},
      {stage2_61[36], stage2_61[37], stage2_61[38], stage2_61[39], stage2_61[40], stage2_61[41]},
      {stage3_63[6],stage3_62[12],stage3_61[19],stage3_60[24],stage3_59[24]}
   );
   gpc606_5 gpc7694 (
      {stage2_60[43], stage2_60[44], stage2_60[45], stage2_60[46], stage2_60[47], stage2_60[48]},
      {stage2_62[0], stage2_62[1], stage2_62[2], stage2_62[3], stage2_62[4], stage2_62[5]},
      {stage3_64[0],stage3_63[7],stage3_62[13],stage3_61[20],stage3_60[25]}
   );
   gpc606_5 gpc7695 (
      {stage2_60[49], stage2_60[50], stage2_60[51], stage2_60[52], stage2_60[53], stage2_60[54]},
      {stage2_62[6], stage2_62[7], stage2_62[8], stage2_62[9], stage2_62[10], stage2_62[11]},
      {stage3_64[1],stage3_63[8],stage3_62[14],stage3_61[21],stage3_60[26]}
   );
   gpc606_5 gpc7696 (
      {stage2_60[55], stage2_60[56], stage2_60[57], stage2_60[58], stage2_60[59], stage2_60[60]},
      {stage2_62[12], stage2_62[13], stage2_62[14], stage2_62[15], stage2_62[16], stage2_62[17]},
      {stage3_64[2],stage3_63[9],stage3_62[15],stage3_61[22],stage3_60[27]}
   );
   gpc606_5 gpc7697 (
      {stage2_60[61], stage2_60[62], stage2_60[63], stage2_60[64], stage2_60[65], stage2_60[66]},
      {stage2_62[18], stage2_62[19], stage2_62[20], stage2_62[21], stage2_62[22], stage2_62[23]},
      {stage3_64[3],stage3_63[10],stage3_62[16],stage3_61[23],stage3_60[28]}
   );
   gpc606_5 gpc7698 (
      {stage2_60[67], stage2_60[68], stage2_60[69], stage2_60[70], stage2_60[71], stage2_60[72]},
      {stage2_62[24], stage2_62[25], stage2_62[26], stage2_62[27], stage2_62[28], stage2_62[29]},
      {stage3_64[4],stage3_63[11],stage3_62[17],stage3_61[24],stage3_60[29]}
   );
   gpc606_5 gpc7699 (
      {stage2_61[42], stage2_61[43], stage2_61[44], stage2_61[45], stage2_61[46], stage2_61[47]},
      {stage2_63[0], stage2_63[1], stage2_63[2], stage2_63[3], stage2_63[4], stage2_63[5]},
      {stage3_65[0],stage3_64[5],stage3_63[12],stage3_62[18],stage3_61[25]}
   );
   gpc615_5 gpc7700 (
      {stage2_62[30], stage2_62[31], stage2_62[32], stage2_62[33], stage2_62[34]},
      {stage2_63[6]},
      {stage2_64[0], stage2_64[1], stage2_64[2], stage2_64[3], stage2_64[4], stage2_64[5]},
      {stage3_66[0],stage3_65[1],stage3_64[6],stage3_63[13],stage3_62[19]}
   );
   gpc615_5 gpc7701 (
      {stage2_62[35], stage2_62[36], stage2_62[37], stage2_62[38], stage2_62[39]},
      {stage2_63[7]},
      {stage2_64[6], stage2_64[7], stage2_64[8], stage2_64[9], stage2_64[10], stage2_64[11]},
      {stage3_66[1],stage3_65[2],stage3_64[7],stage3_63[14],stage3_62[20]}
   );
   gpc615_5 gpc7702 (
      {stage2_62[40], stage2_62[41], stage2_62[42], stage2_62[43], stage2_62[44]},
      {stage2_63[8]},
      {stage2_64[12], stage2_64[13], stage2_64[14], stage2_64[15], stage2_64[16], stage2_64[17]},
      {stage3_66[2],stage3_65[3],stage3_64[8],stage3_63[15],stage3_62[21]}
   );
   gpc615_5 gpc7703 (
      {stage2_62[45], stage2_62[46], stage2_62[47], stage2_62[48], stage2_62[49]},
      {stage2_63[9]},
      {stage2_64[18], stage2_64[19], stage2_64[20], stage2_64[21], stage2_64[22], stage2_64[23]},
      {stage3_66[3],stage3_65[4],stage3_64[9],stage3_63[16],stage3_62[22]}
   );
   gpc615_5 gpc7704 (
      {stage2_62[50], stage2_62[51], stage2_62[52], stage2_62[53], stage2_62[54]},
      {stage2_63[10]},
      {stage2_64[24], stage2_64[25], stage2_64[26], stage2_64[27], stage2_64[28], stage2_64[29]},
      {stage3_66[4],stage3_65[5],stage3_64[10],stage3_63[17],stage3_62[23]}
   );
   gpc615_5 gpc7705 (
      {stage2_62[55], stage2_62[56], stage2_62[57], stage2_62[58], stage2_62[59]},
      {stage2_63[11]},
      {stage2_64[30], stage2_64[31], stage2_64[32], stage2_64[33], stage2_64[34], stage2_64[35]},
      {stage3_66[5],stage3_65[6],stage3_64[11],stage3_63[18],stage3_62[24]}
   );
   gpc615_5 gpc7706 (
      {stage2_62[60], stage2_62[61], stage2_62[62], stage2_62[63], stage2_62[64]},
      {stage2_63[12]},
      {stage2_64[36], stage2_64[37], stage2_64[38], stage2_64[39], stage2_64[40], stage2_64[41]},
      {stage3_66[6],stage3_65[7],stage3_64[12],stage3_63[19],stage3_62[25]}
   );
   gpc615_5 gpc7707 (
      {stage2_62[65], stage2_62[66], stage2_62[67], stage2_62[68], stage2_62[69]},
      {stage2_63[13]},
      {stage2_64[42], stage2_64[43], stage2_64[44], stage2_64[45], stage2_64[46], stage2_64[47]},
      {stage3_66[7],stage3_65[8],stage3_64[13],stage3_63[20],stage3_62[26]}
   );
   gpc615_5 gpc7708 (
      {stage2_62[70], stage2_62[71], stage2_62[72], stage2_62[73], stage2_62[74]},
      {stage2_63[14]},
      {stage2_64[48], stage2_64[49], stage2_64[50], stage2_64[51], stage2_64[52], stage2_64[53]},
      {stage3_66[8],stage3_65[9],stage3_64[14],stage3_63[21],stage3_62[27]}
   );
   gpc615_5 gpc7709 (
      {stage2_62[75], stage2_62[76], stage2_62[77], stage2_62[78], stage2_62[79]},
      {stage2_63[15]},
      {stage2_64[54], stage2_64[55], stage2_64[56], stage2_64[57], stage2_64[58], stage2_64[59]},
      {stage3_66[9],stage3_65[10],stage3_64[15],stage3_63[22],stage3_62[28]}
   );
   gpc615_5 gpc7710 (
      {stage2_62[80], stage2_62[81], stage2_62[82], stage2_62[83], stage2_62[84]},
      {stage2_63[16]},
      {stage2_64[60], stage2_64[61], stage2_64[62], stage2_64[63], stage2_64[64], stage2_64[65]},
      {stage3_66[10],stage3_65[11],stage3_64[16],stage3_63[23],stage3_62[29]}
   );
   gpc615_5 gpc7711 (
      {stage2_62[85], stage2_62[86], stage2_62[87], stage2_62[88], stage2_62[89]},
      {stage2_63[17]},
      {stage2_64[66], stage2_64[67], stage2_64[68], stage2_64[69], stage2_64[70], stage2_64[71]},
      {stage3_66[11],stage3_65[12],stage3_64[17],stage3_63[24],stage3_62[30]}
   );
   gpc615_5 gpc7712 (
      {stage2_62[90], stage2_62[91], stage2_62[92], stage2_62[93], stage2_62[94]},
      {stage2_63[18]},
      {stage2_64[72], stage2_64[73], stage2_64[74], stage2_64[75], stage2_64[76], stage2_64[77]},
      {stage3_66[12],stage3_65[13],stage3_64[18],stage3_63[25],stage3_62[31]}
   );
   gpc615_5 gpc7713 (
      {stage2_62[95], stage2_62[96], stage2_62[97], stage2_62[98], stage2_62[99]},
      {stage2_63[19]},
      {stage2_64[78], stage2_64[79], stage2_64[80], stage2_64[81], stage2_64[82], stage2_64[83]},
      {stage3_66[13],stage3_65[14],stage3_64[19],stage3_63[26],stage3_62[32]}
   );
   gpc615_5 gpc7714 (
      {stage2_62[100], stage2_62[101], stage2_62[102], stage2_62[103], stage2_62[104]},
      {stage2_63[20]},
      {stage2_64[84], stage2_64[85], stage2_64[86], stage2_64[87], stage2_64[88], stage2_64[89]},
      {stage3_66[14],stage3_65[15],stage3_64[20],stage3_63[27],stage3_62[33]}
   );
   gpc117_4 gpc7715 (
      {stage2_63[21], stage2_63[22], stage2_63[23], stage2_63[24], stage2_63[25], stage2_63[26], stage2_63[27]},
      {stage2_64[90]},
      {stage2_65[0]},
      {stage3_66[15],stage3_65[16],stage3_64[21],stage3_63[28]}
   );
   gpc117_4 gpc7716 (
      {stage2_63[28], stage2_63[29], stage2_63[30], stage2_63[31], stage2_63[32], stage2_63[33], stage2_63[34]},
      {stage2_64[91]},
      {stage2_65[1]},
      {stage3_66[16],stage3_65[17],stage3_64[22],stage3_63[29]}
   );
   gpc117_4 gpc7717 (
      {stage2_63[35], stage2_63[36], stage2_63[37], stage2_63[38], stage2_63[39], stage2_63[40], stage2_63[41]},
      {stage2_64[92]},
      {stage2_65[2]},
      {stage3_66[17],stage3_65[18],stage3_64[23],stage3_63[30]}
   );
   gpc606_5 gpc7718 (
      {stage2_63[42], stage2_63[43], stage2_63[44], stage2_63[45], stage2_63[46], stage2_63[47]},
      {stage2_65[3], stage2_65[4], stage2_65[5], stage2_65[6], stage2_65[7], stage2_65[8]},
      {stage3_67[0],stage3_66[18],stage3_65[19],stage3_64[24],stage3_63[31]}
   );
   gpc606_5 gpc7719 (
      {stage2_63[48], stage2_63[49], stage2_63[50], stage2_63[51], stage2_63[52], stage2_63[53]},
      {stage2_65[9], stage2_65[10], stage2_65[11], stage2_65[12], stage2_65[13], stage2_65[14]},
      {stage3_67[1],stage3_66[19],stage3_65[20],stage3_64[25],stage3_63[32]}
   );
   gpc606_5 gpc7720 (
      {stage2_63[54], stage2_63[55], stage2_63[56], stage2_63[57], stage2_63[58], stage2_63[59]},
      {stage2_65[15], stage2_65[16], stage2_65[17], stage2_65[18], stage2_65[19], stage2_65[20]},
      {stage3_67[2],stage3_66[20],stage3_65[21],stage3_64[26],stage3_63[33]}
   );
   gpc606_5 gpc7721 (
      {stage2_63[60], stage2_63[61], stage2_63[62], stage2_63[63], stage2_63[64], stage2_63[65]},
      {stage2_65[21], stage2_65[22], stage2_65[23], stage2_65[24], stage2_65[25], stage2_65[26]},
      {stage3_67[3],stage3_66[21],stage3_65[22],stage3_64[27],stage3_63[34]}
   );
   gpc606_5 gpc7722 (
      {stage2_63[66], stage2_63[67], stage2_63[68], stage2_63[69], stage2_63[70], stage2_63[71]},
      {stage2_65[27], stage2_65[28], stage2_65[29], stage2_65[30], stage2_65[31], stage2_65[32]},
      {stage3_67[4],stage3_66[22],stage3_65[23],stage3_64[28],stage3_63[35]}
   );
   gpc606_5 gpc7723 (
      {stage2_63[72], stage2_63[73], stage2_63[74], stage2_63[75], stage2_63[76], stage2_63[77]},
      {stage2_65[33], stage2_65[34], stage2_65[35], stage2_65[36], stage2_65[37], stage2_65[38]},
      {stage3_67[5],stage3_66[23],stage3_65[24],stage3_64[29],stage3_63[36]}
   );
   gpc606_5 gpc7724 (
      {stage2_63[78], stage2_63[79], stage2_63[80], stage2_63[81], stage2_63[82], stage2_63[83]},
      {stage2_65[39], stage2_65[40], stage2_65[41], stage2_65[42], stage2_65[43], stage2_65[44]},
      {stage3_67[6],stage3_66[24],stage3_65[25],stage3_64[30],stage3_63[37]}
   );
   gpc606_5 gpc7725 (
      {stage2_63[84], stage2_63[85], stage2_63[86], stage2_63[87], stage2_63[88], stage2_63[89]},
      {stage2_65[45], stage2_65[46], stage2_65[47], stage2_65[48], stage2_65[49], stage2_65[50]},
      {stage3_67[7],stage3_66[25],stage3_65[26],stage3_64[31],stage3_63[38]}
   );
   gpc606_5 gpc7726 (
      {stage2_64[93], stage2_64[94], stage2_64[95], stage2_64[96], stage2_64[97], stage2_64[98]},
      {stage2_66[0], stage2_66[1], stage2_66[2], stage2_66[3], stage2_66[4], stage2_66[5]},
      {stage3_68[0],stage3_67[8],stage3_66[26],stage3_65[27],stage3_64[32]}
   );
   gpc606_5 gpc7727 (
      {stage2_64[99], stage2_64[100], stage2_64[101], stage2_64[102], stage2_64[103], stage2_64[104]},
      {stage2_66[6], stage2_66[7], stage2_66[8], stage2_66[9], stage2_66[10], stage2_66[11]},
      {stage3_68[1],stage3_67[9],stage3_66[27],stage3_65[28],stage3_64[33]}
   );
   gpc606_5 gpc7728 (
      {stage2_64[105], stage2_64[106], stage2_64[107], stage2_64[108], stage2_64[109], stage2_64[110]},
      {stage2_66[12], stage2_66[13], stage2_66[14], stage2_66[15], stage2_66[16], stage2_66[17]},
      {stage3_68[2],stage3_67[10],stage3_66[28],stage3_65[29],stage3_64[34]}
   );
   gpc606_5 gpc7729 (
      {stage2_64[111], stage2_64[112], stage2_64[113], stage2_64[114], stage2_64[115], stage2_64[116]},
      {stage2_66[18], stage2_66[19], stage2_66[20], stage2_66[21], stage2_66[22], stage2_66[23]},
      {stage3_68[3],stage3_67[11],stage3_66[29],stage3_65[30],stage3_64[35]}
   );
   gpc606_5 gpc7730 (
      {stage2_64[117], stage2_64[118], stage2_64[119], stage2_64[120], stage2_64[121], stage2_64[122]},
      {stage2_66[24], stage2_66[25], stage2_66[26], stage2_66[27], stage2_66[28], stage2_66[29]},
      {stage3_68[4],stage3_67[12],stage3_66[30],stage3_65[31],stage3_64[36]}
   );
   gpc606_5 gpc7731 (
      {stage2_64[123], stage2_64[124], stage2_64[125], stage2_64[126], stage2_64[127], stage2_64[128]},
      {stage2_66[30], stage2_66[31], stage2_66[32], stage2_66[33], stage2_66[34], stage2_66[35]},
      {stage3_68[5],stage3_67[13],stage3_66[31],stage3_65[32],stage3_64[37]}
   );
   gpc1_1 gpc7732 (
      {stage2_0[23]},
      {stage3_0[6]}
   );
   gpc1_1 gpc7733 (
      {stage2_0[24]},
      {stage3_0[7]}
   );
   gpc1_1 gpc7734 (
      {stage2_0[25]},
      {stage3_0[8]}
   );
   gpc1_1 gpc7735 (
      {stage2_0[26]},
      {stage3_0[9]}
   );
   gpc1_1 gpc7736 (
      {stage2_0[27]},
      {stage3_0[10]}
   );
   gpc1_1 gpc7737 (
      {stage2_0[28]},
      {stage3_0[11]}
   );
   gpc1_1 gpc7738 (
      {stage2_0[29]},
      {stage3_0[12]}
   );
   gpc1_1 gpc7739 (
      {stage2_0[30]},
      {stage3_0[13]}
   );
   gpc1_1 gpc7740 (
      {stage2_0[31]},
      {stage3_0[14]}
   );
   gpc1_1 gpc7741 (
      {stage2_0[32]},
      {stage3_0[15]}
   );
   gpc1_1 gpc7742 (
      {stage2_0[33]},
      {stage3_0[16]}
   );
   gpc1_1 gpc7743 (
      {stage2_0[34]},
      {stage3_0[17]}
   );
   gpc1_1 gpc7744 (
      {stage2_0[35]},
      {stage3_0[18]}
   );
   gpc1_1 gpc7745 (
      {stage2_0[36]},
      {stage3_0[19]}
   );
   gpc1_1 gpc7746 (
      {stage2_0[37]},
      {stage3_0[20]}
   );
   gpc1_1 gpc7747 (
      {stage2_1[42]},
      {stage3_1[10]}
   );
   gpc1_1 gpc7748 (
      {stage2_1[43]},
      {stage3_1[11]}
   );
   gpc1_1 gpc7749 (
      {stage2_1[44]},
      {stage3_1[12]}
   );
   gpc1_1 gpc7750 (
      {stage2_1[45]},
      {stage3_1[13]}
   );
   gpc1_1 gpc7751 (
      {stage2_1[46]},
      {stage3_1[14]}
   );
   gpc1_1 gpc7752 (
      {stage2_1[47]},
      {stage3_1[15]}
   );
   gpc1_1 gpc7753 (
      {stage2_1[48]},
      {stage3_1[16]}
   );
   gpc1_1 gpc7754 (
      {stage2_1[49]},
      {stage3_1[17]}
   );
   gpc1_1 gpc7755 (
      {stage2_1[50]},
      {stage3_1[18]}
   );
   gpc1_1 gpc7756 (
      {stage2_1[51]},
      {stage3_1[19]}
   );
   gpc1_1 gpc7757 (
      {stage2_1[52]},
      {stage3_1[20]}
   );
   gpc1_1 gpc7758 (
      {stage2_1[53]},
      {stage3_1[21]}
   );
   gpc1_1 gpc7759 (
      {stage2_2[32]},
      {stage3_2[12]}
   );
   gpc1_1 gpc7760 (
      {stage2_2[33]},
      {stage3_2[13]}
   );
   gpc1_1 gpc7761 (
      {stage2_2[34]},
      {stage3_2[14]}
   );
   gpc1_1 gpc7762 (
      {stage2_2[35]},
      {stage3_2[15]}
   );
   gpc1_1 gpc7763 (
      {stage2_2[36]},
      {stage3_2[16]}
   );
   gpc1_1 gpc7764 (
      {stage2_2[37]},
      {stage3_2[17]}
   );
   gpc1_1 gpc7765 (
      {stage2_2[38]},
      {stage3_2[18]}
   );
   gpc1_1 gpc7766 (
      {stage2_2[39]},
      {stage3_2[19]}
   );
   gpc1_1 gpc7767 (
      {stage2_2[40]},
      {stage3_2[20]}
   );
   gpc1_1 gpc7768 (
      {stage2_2[41]},
      {stage3_2[21]}
   );
   gpc1_1 gpc7769 (
      {stage2_2[42]},
      {stage3_2[22]}
   );
   gpc1_1 gpc7770 (
      {stage2_2[43]},
      {stage3_2[23]}
   );
   gpc1_1 gpc7771 (
      {stage2_2[44]},
      {stage3_2[24]}
   );
   gpc1_1 gpc7772 (
      {stage2_2[45]},
      {stage3_2[25]}
   );
   gpc1_1 gpc7773 (
      {stage2_2[46]},
      {stage3_2[26]}
   );
   gpc1_1 gpc7774 (
      {stage2_2[47]},
      {stage3_2[27]}
   );
   gpc1_1 gpc7775 (
      {stage2_2[48]},
      {stage3_2[28]}
   );
   gpc1_1 gpc7776 (
      {stage2_2[49]},
      {stage3_2[29]}
   );
   gpc1_1 gpc7777 (
      {stage2_2[50]},
      {stage3_2[30]}
   );
   gpc1_1 gpc7778 (
      {stage2_2[51]},
      {stage3_2[31]}
   );
   gpc1_1 gpc7779 (
      {stage2_2[52]},
      {stage3_2[32]}
   );
   gpc1_1 gpc7780 (
      {stage2_2[53]},
      {stage3_2[33]}
   );
   gpc1_1 gpc7781 (
      {stage2_2[54]},
      {stage3_2[34]}
   );
   gpc1_1 gpc7782 (
      {stage2_2[55]},
      {stage3_2[35]}
   );
   gpc1_1 gpc7783 (
      {stage2_2[56]},
      {stage3_2[36]}
   );
   gpc1_1 gpc7784 (
      {stage2_2[57]},
      {stage3_2[37]}
   );
   gpc1_1 gpc7785 (
      {stage2_2[58]},
      {stage3_2[38]}
   );
   gpc1_1 gpc7786 (
      {stage2_2[59]},
      {stage3_2[39]}
   );
   gpc1_1 gpc7787 (
      {stage2_2[60]},
      {stage3_2[40]}
   );
   gpc1_1 gpc7788 (
      {stage2_2[61]},
      {stage3_2[41]}
   );
   gpc1_1 gpc7789 (
      {stage2_2[62]},
      {stage3_2[42]}
   );
   gpc1_1 gpc7790 (
      {stage2_4[29]},
      {stage3_4[29]}
   );
   gpc1_1 gpc7791 (
      {stage2_4[30]},
      {stage3_4[30]}
   );
   gpc1_1 gpc7792 (
      {stage2_4[31]},
      {stage3_4[31]}
   );
   gpc1_1 gpc7793 (
      {stage2_4[32]},
      {stage3_4[32]}
   );
   gpc1_1 gpc7794 (
      {stage2_4[33]},
      {stage3_4[33]}
   );
   gpc1_1 gpc7795 (
      {stage2_4[34]},
      {stage3_4[34]}
   );
   gpc1_1 gpc7796 (
      {stage2_4[35]},
      {stage3_4[35]}
   );
   gpc1_1 gpc7797 (
      {stage2_4[36]},
      {stage3_4[36]}
   );
   gpc1_1 gpc7798 (
      {stage2_4[37]},
      {stage3_4[37]}
   );
   gpc1_1 gpc7799 (
      {stage2_4[38]},
      {stage3_4[38]}
   );
   gpc1_1 gpc7800 (
      {stage2_4[39]},
      {stage3_4[39]}
   );
   gpc1_1 gpc7801 (
      {stage2_4[40]},
      {stage3_4[40]}
   );
   gpc1_1 gpc7802 (
      {stage2_4[41]},
      {stage3_4[41]}
   );
   gpc1_1 gpc7803 (
      {stage2_4[42]},
      {stage3_4[42]}
   );
   gpc1_1 gpc7804 (
      {stage2_4[43]},
      {stage3_4[43]}
   );
   gpc1_1 gpc7805 (
      {stage2_4[44]},
      {stage3_4[44]}
   );
   gpc1_1 gpc7806 (
      {stage2_4[45]},
      {stage3_4[45]}
   );
   gpc1_1 gpc7807 (
      {stage2_4[46]},
      {stage3_4[46]}
   );
   gpc1_1 gpc7808 (
      {stage2_4[47]},
      {stage3_4[47]}
   );
   gpc1_1 gpc7809 (
      {stage2_4[48]},
      {stage3_4[48]}
   );
   gpc1_1 gpc7810 (
      {stage2_4[49]},
      {stage3_4[49]}
   );
   gpc1_1 gpc7811 (
      {stage2_4[50]},
      {stage3_4[50]}
   );
   gpc1_1 gpc7812 (
      {stage2_4[51]},
      {stage3_4[51]}
   );
   gpc1_1 gpc7813 (
      {stage2_4[52]},
      {stage3_4[52]}
   );
   gpc1_1 gpc7814 (
      {stage2_4[53]},
      {stage3_4[53]}
   );
   gpc1_1 gpc7815 (
      {stage2_4[54]},
      {stage3_4[54]}
   );
   gpc1_1 gpc7816 (
      {stage2_4[55]},
      {stage3_4[55]}
   );
   gpc1_1 gpc7817 (
      {stage2_4[56]},
      {stage3_4[56]}
   );
   gpc1_1 gpc7818 (
      {stage2_4[57]},
      {stage3_4[57]}
   );
   gpc1_1 gpc7819 (
      {stage2_4[58]},
      {stage3_4[58]}
   );
   gpc1_1 gpc7820 (
      {stage2_4[59]},
      {stage3_4[59]}
   );
   gpc1_1 gpc7821 (
      {stage2_4[60]},
      {stage3_4[60]}
   );
   gpc1_1 gpc7822 (
      {stage2_4[61]},
      {stage3_4[61]}
   );
   gpc1_1 gpc7823 (
      {stage2_4[62]},
      {stage3_4[62]}
   );
   gpc1_1 gpc7824 (
      {stage2_4[63]},
      {stage3_4[63]}
   );
   gpc1_1 gpc7825 (
      {stage2_4[64]},
      {stage3_4[64]}
   );
   gpc1_1 gpc7826 (
      {stage2_4[65]},
      {stage3_4[65]}
   );
   gpc1_1 gpc7827 (
      {stage2_4[66]},
      {stage3_4[66]}
   );
   gpc1_1 gpc7828 (
      {stage2_4[67]},
      {stage3_4[67]}
   );
   gpc1_1 gpc7829 (
      {stage2_4[68]},
      {stage3_4[68]}
   );
   gpc1_1 gpc7830 (
      {stage2_4[69]},
      {stage3_4[69]}
   );
   gpc1_1 gpc7831 (
      {stage2_4[70]},
      {stage3_4[70]}
   );
   gpc1_1 gpc7832 (
      {stage2_4[71]},
      {stage3_4[71]}
   );
   gpc1_1 gpc7833 (
      {stage2_4[72]},
      {stage3_4[72]}
   );
   gpc1_1 gpc7834 (
      {stage2_4[73]},
      {stage3_4[73]}
   );
   gpc1_1 gpc7835 (
      {stage2_4[74]},
      {stage3_4[74]}
   );
   gpc1_1 gpc7836 (
      {stage2_4[75]},
      {stage3_4[75]}
   );
   gpc1_1 gpc7837 (
      {stage2_4[76]},
      {stage3_4[76]}
   );
   gpc1_1 gpc7838 (
      {stage2_4[77]},
      {stage3_4[77]}
   );
   gpc1_1 gpc7839 (
      {stage2_4[78]},
      {stage3_4[78]}
   );
   gpc1_1 gpc7840 (
      {stage2_4[79]},
      {stage3_4[79]}
   );
   gpc1_1 gpc7841 (
      {stage2_4[80]},
      {stage3_4[80]}
   );
   gpc1_1 gpc7842 (
      {stage2_4[81]},
      {stage3_4[81]}
   );
   gpc1_1 gpc7843 (
      {stage2_4[82]},
      {stage3_4[82]}
   );
   gpc1_1 gpc7844 (
      {stage2_4[83]},
      {stage3_4[83]}
   );
   gpc1_1 gpc7845 (
      {stage2_4[84]},
      {stage3_4[84]}
   );
   gpc1_1 gpc7846 (
      {stage2_4[85]},
      {stage3_4[85]}
   );
   gpc1_1 gpc7847 (
      {stage2_4[86]},
      {stage3_4[86]}
   );
   gpc1_1 gpc7848 (
      {stage2_4[87]},
      {stage3_4[87]}
   );
   gpc1_1 gpc7849 (
      {stage2_4[88]},
      {stage3_4[88]}
   );
   gpc1_1 gpc7850 (
      {stage2_4[89]},
      {stage3_4[89]}
   );
   gpc1_1 gpc7851 (
      {stage2_4[90]},
      {stage3_4[90]}
   );
   gpc1_1 gpc7852 (
      {stage2_4[91]},
      {stage3_4[91]}
   );
   gpc1_1 gpc7853 (
      {stage2_4[92]},
      {stage3_4[92]}
   );
   gpc1_1 gpc7854 (
      {stage2_4[93]},
      {stage3_4[93]}
   );
   gpc1_1 gpc7855 (
      {stage2_4[94]},
      {stage3_4[94]}
   );
   gpc1_1 gpc7856 (
      {stage2_4[95]},
      {stage3_4[95]}
   );
   gpc1_1 gpc7857 (
      {stage2_4[96]},
      {stage3_4[96]}
   );
   gpc1_1 gpc7858 (
      {stage2_4[97]},
      {stage3_4[97]}
   );
   gpc1_1 gpc7859 (
      {stage2_4[98]},
      {stage3_4[98]}
   );
   gpc1_1 gpc7860 (
      {stage2_4[99]},
      {stage3_4[99]}
   );
   gpc1_1 gpc7861 (
      {stage2_4[100]},
      {stage3_4[100]}
   );
   gpc1_1 gpc7862 (
      {stage2_4[101]},
      {stage3_4[101]}
   );
   gpc1_1 gpc7863 (
      {stage2_4[102]},
      {stage3_4[102]}
   );
   gpc1_1 gpc7864 (
      {stage2_4[103]},
      {stage3_4[103]}
   );
   gpc1_1 gpc7865 (
      {stage2_4[104]},
      {stage3_4[104]}
   );
   gpc1_1 gpc7866 (
      {stage2_4[105]},
      {stage3_4[105]}
   );
   gpc1_1 gpc7867 (
      {stage2_4[106]},
      {stage3_4[106]}
   );
   gpc1_1 gpc7868 (
      {stage2_4[107]},
      {stage3_4[107]}
   );
   gpc1_1 gpc7869 (
      {stage2_4[108]},
      {stage3_4[108]}
   );
   gpc1_1 gpc7870 (
      {stage2_4[109]},
      {stage3_4[109]}
   );
   gpc1_1 gpc7871 (
      {stage2_4[110]},
      {stage3_4[110]}
   );
   gpc1_1 gpc7872 (
      {stage2_4[111]},
      {stage3_4[111]}
   );
   gpc1_1 gpc7873 (
      {stage2_5[126]},
      {stage3_5[27]}
   );
   gpc1_1 gpc7874 (
      {stage2_5[127]},
      {stage3_5[28]}
   );
   gpc1_1 gpc7875 (
      {stage2_5[128]},
      {stage3_5[29]}
   );
   gpc1_1 gpc7876 (
      {stage2_5[129]},
      {stage3_5[30]}
   );
   gpc1_1 gpc7877 (
      {stage2_5[130]},
      {stage3_5[31]}
   );
   gpc1_1 gpc7878 (
      {stage2_5[131]},
      {stage3_5[32]}
   );
   gpc1_1 gpc7879 (
      {stage2_5[132]},
      {stage3_5[33]}
   );
   gpc1_1 gpc7880 (
      {stage2_5[133]},
      {stage3_5[34]}
   );
   gpc1_1 gpc7881 (
      {stage2_5[134]},
      {stage3_5[35]}
   );
   gpc1_1 gpc7882 (
      {stage2_5[135]},
      {stage3_5[36]}
   );
   gpc1_1 gpc7883 (
      {stage2_5[136]},
      {stage3_5[37]}
   );
   gpc1_1 gpc7884 (
      {stage2_5[137]},
      {stage3_5[38]}
   );
   gpc1_1 gpc7885 (
      {stage2_5[138]},
      {stage3_5[39]}
   );
   gpc1_1 gpc7886 (
      {stage2_5[139]},
      {stage3_5[40]}
   );
   gpc1_1 gpc7887 (
      {stage2_5[140]},
      {stage3_5[41]}
   );
   gpc1_1 gpc7888 (
      {stage2_5[141]},
      {stage3_5[42]}
   );
   gpc1_1 gpc7889 (
      {stage2_5[142]},
      {stage3_5[43]}
   );
   gpc1_1 gpc7890 (
      {stage2_5[143]},
      {stage3_5[44]}
   );
   gpc1_1 gpc7891 (
      {stage2_5[144]},
      {stage3_5[45]}
   );
   gpc1_1 gpc7892 (
      {stage2_5[145]},
      {stage3_5[46]}
   );
   gpc1_1 gpc7893 (
      {stage2_5[146]},
      {stage3_5[47]}
   );
   gpc1_1 gpc7894 (
      {stage2_5[147]},
      {stage3_5[48]}
   );
   gpc1_1 gpc7895 (
      {stage2_5[148]},
      {stage3_5[49]}
   );
   gpc1_1 gpc7896 (
      {stage2_5[149]},
      {stage3_5[50]}
   );
   gpc1_1 gpc7897 (
      {stage2_5[150]},
      {stage3_5[51]}
   );
   gpc1_1 gpc7898 (
      {stage2_5[151]},
      {stage3_5[52]}
   );
   gpc1_1 gpc7899 (
      {stage2_6[46]},
      {stage3_6[32]}
   );
   gpc1_1 gpc7900 (
      {stage2_6[47]},
      {stage3_6[33]}
   );
   gpc1_1 gpc7901 (
      {stage2_6[48]},
      {stage3_6[34]}
   );
   gpc1_1 gpc7902 (
      {stage2_6[49]},
      {stage3_6[35]}
   );
   gpc1_1 gpc7903 (
      {stage2_6[50]},
      {stage3_6[36]}
   );
   gpc1_1 gpc7904 (
      {stage2_6[51]},
      {stage3_6[37]}
   );
   gpc1_1 gpc7905 (
      {stage2_6[52]},
      {stage3_6[38]}
   );
   gpc1_1 gpc7906 (
      {stage2_6[53]},
      {stage3_6[39]}
   );
   gpc1_1 gpc7907 (
      {stage2_6[54]},
      {stage3_6[40]}
   );
   gpc1_1 gpc7908 (
      {stage2_6[55]},
      {stage3_6[41]}
   );
   gpc1_1 gpc7909 (
      {stage2_6[56]},
      {stage3_6[42]}
   );
   gpc1_1 gpc7910 (
      {stage2_6[57]},
      {stage3_6[43]}
   );
   gpc1_1 gpc7911 (
      {stage2_6[58]},
      {stage3_6[44]}
   );
   gpc1_1 gpc7912 (
      {stage2_6[59]},
      {stage3_6[45]}
   );
   gpc1_1 gpc7913 (
      {stage2_6[60]},
      {stage3_6[46]}
   );
   gpc1_1 gpc7914 (
      {stage2_6[61]},
      {stage3_6[47]}
   );
   gpc1_1 gpc7915 (
      {stage2_6[62]},
      {stage3_6[48]}
   );
   gpc1_1 gpc7916 (
      {stage2_6[63]},
      {stage3_6[49]}
   );
   gpc1_1 gpc7917 (
      {stage2_6[64]},
      {stage3_6[50]}
   );
   gpc1_1 gpc7918 (
      {stage2_6[65]},
      {stage3_6[51]}
   );
   gpc1_1 gpc7919 (
      {stage2_6[66]},
      {stage3_6[52]}
   );
   gpc1_1 gpc7920 (
      {stage2_6[67]},
      {stage3_6[53]}
   );
   gpc1_1 gpc7921 (
      {stage2_6[68]},
      {stage3_6[54]}
   );
   gpc1_1 gpc7922 (
      {stage2_6[69]},
      {stage3_6[55]}
   );
   gpc1_1 gpc7923 (
      {stage2_6[70]},
      {stage3_6[56]}
   );
   gpc1_1 gpc7924 (
      {stage2_6[71]},
      {stage3_6[57]}
   );
   gpc1_1 gpc7925 (
      {stage2_6[72]},
      {stage3_6[58]}
   );
   gpc1_1 gpc7926 (
      {stage2_6[73]},
      {stage3_6[59]}
   );
   gpc1_1 gpc7927 (
      {stage2_6[74]},
      {stage3_6[60]}
   );
   gpc1_1 gpc7928 (
      {stage2_6[75]},
      {stage3_6[61]}
   );
   gpc1_1 gpc7929 (
      {stage2_6[76]},
      {stage3_6[62]}
   );
   gpc1_1 gpc7930 (
      {stage2_6[77]},
      {stage3_6[63]}
   );
   gpc1_1 gpc7931 (
      {stage2_6[78]},
      {stage3_6[64]}
   );
   gpc1_1 gpc7932 (
      {stage2_6[79]},
      {stage3_6[65]}
   );
   gpc1_1 gpc7933 (
      {stage2_6[80]},
      {stage3_6[66]}
   );
   gpc1_1 gpc7934 (
      {stage2_6[81]},
      {stage3_6[67]}
   );
   gpc1_1 gpc7935 (
      {stage2_6[82]},
      {stage3_6[68]}
   );
   gpc1_1 gpc7936 (
      {stage2_6[83]},
      {stage3_6[69]}
   );
   gpc1_1 gpc7937 (
      {stage2_6[84]},
      {stage3_6[70]}
   );
   gpc1_1 gpc7938 (
      {stage2_6[85]},
      {stage3_6[71]}
   );
   gpc1_1 gpc7939 (
      {stage2_6[86]},
      {stage3_6[72]}
   );
   gpc1_1 gpc7940 (
      {stage2_6[87]},
      {stage3_6[73]}
   );
   gpc1_1 gpc7941 (
      {stage2_6[88]},
      {stage3_6[74]}
   );
   gpc1_1 gpc7942 (
      {stage2_6[89]},
      {stage3_6[75]}
   );
   gpc1_1 gpc7943 (
      {stage2_6[90]},
      {stage3_6[76]}
   );
   gpc1_1 gpc7944 (
      {stage2_6[91]},
      {stage3_6[77]}
   );
   gpc1_1 gpc7945 (
      {stage2_7[57]},
      {stage3_7[35]}
   );
   gpc1_1 gpc7946 (
      {stage2_7[58]},
      {stage3_7[36]}
   );
   gpc1_1 gpc7947 (
      {stage2_7[59]},
      {stage3_7[37]}
   );
   gpc1_1 gpc7948 (
      {stage2_7[60]},
      {stage3_7[38]}
   );
   gpc1_1 gpc7949 (
      {stage2_7[61]},
      {stage3_7[39]}
   );
   gpc1_1 gpc7950 (
      {stage2_7[62]},
      {stage3_7[40]}
   );
   gpc1_1 gpc7951 (
      {stage2_7[63]},
      {stage3_7[41]}
   );
   gpc1_1 gpc7952 (
      {stage2_7[64]},
      {stage3_7[42]}
   );
   gpc1_1 gpc7953 (
      {stage2_7[65]},
      {stage3_7[43]}
   );
   gpc1_1 gpc7954 (
      {stage2_7[66]},
      {stage3_7[44]}
   );
   gpc1_1 gpc7955 (
      {stage2_7[67]},
      {stage3_7[45]}
   );
   gpc1_1 gpc7956 (
      {stage2_7[68]},
      {stage3_7[46]}
   );
   gpc1_1 gpc7957 (
      {stage2_7[69]},
      {stage3_7[47]}
   );
   gpc1_1 gpc7958 (
      {stage2_7[70]},
      {stage3_7[48]}
   );
   gpc1_1 gpc7959 (
      {stage2_7[71]},
      {stage3_7[49]}
   );
   gpc1_1 gpc7960 (
      {stage2_7[72]},
      {stage3_7[50]}
   );
   gpc1_1 gpc7961 (
      {stage2_10[117]},
      {stage3_10[53]}
   );
   gpc1_1 gpc7962 (
      {stage2_10[118]},
      {stage3_10[54]}
   );
   gpc1_1 gpc7963 (
      {stage2_10[119]},
      {stage3_10[55]}
   );
   gpc1_1 gpc7964 (
      {stage2_10[120]},
      {stage3_10[56]}
   );
   gpc1_1 gpc7965 (
      {stage2_10[121]},
      {stage3_10[57]}
   );
   gpc1_1 gpc7966 (
      {stage2_10[122]},
      {stage3_10[58]}
   );
   gpc1_1 gpc7967 (
      {stage2_10[123]},
      {stage3_10[59]}
   );
   gpc1_1 gpc7968 (
      {stage2_10[124]},
      {stage3_10[60]}
   );
   gpc1_1 gpc7969 (
      {stage2_10[125]},
      {stage3_10[61]}
   );
   gpc1_1 gpc7970 (
      {stage2_10[126]},
      {stage3_10[62]}
   );
   gpc1_1 gpc7971 (
      {stage2_10[127]},
      {stage3_10[63]}
   );
   gpc1_1 gpc7972 (
      {stage2_10[128]},
      {stage3_10[64]}
   );
   gpc1_1 gpc7973 (
      {stage2_10[129]},
      {stage3_10[65]}
   );
   gpc1_1 gpc7974 (
      {stage2_10[130]},
      {stage3_10[66]}
   );
   gpc1_1 gpc7975 (
      {stage2_10[131]},
      {stage3_10[67]}
   );
   gpc1_1 gpc7976 (
      {stage2_10[132]},
      {stage3_10[68]}
   );
   gpc1_1 gpc7977 (
      {stage2_10[133]},
      {stage3_10[69]}
   );
   gpc1_1 gpc7978 (
      {stage2_10[134]},
      {stage3_10[70]}
   );
   gpc1_1 gpc7979 (
      {stage2_10[135]},
      {stage3_10[71]}
   );
   gpc1_1 gpc7980 (
      {stage2_10[136]},
      {stage3_10[72]}
   );
   gpc1_1 gpc7981 (
      {stage2_10[137]},
      {stage3_10[73]}
   );
   gpc1_1 gpc7982 (
      {stage2_10[138]},
      {stage3_10[74]}
   );
   gpc1_1 gpc7983 (
      {stage2_10[139]},
      {stage3_10[75]}
   );
   gpc1_1 gpc7984 (
      {stage2_10[140]},
      {stage3_10[76]}
   );
   gpc1_1 gpc7985 (
      {stage2_10[141]},
      {stage3_10[77]}
   );
   gpc1_1 gpc7986 (
      {stage2_10[142]},
      {stage3_10[78]}
   );
   gpc1_1 gpc7987 (
      {stage2_10[143]},
      {stage3_10[79]}
   );
   gpc1_1 gpc7988 (
      {stage2_10[144]},
      {stage3_10[80]}
   );
   gpc1_1 gpc7989 (
      {stage2_10[145]},
      {stage3_10[81]}
   );
   gpc1_1 gpc7990 (
      {stage2_10[146]},
      {stage3_10[82]}
   );
   gpc1_1 gpc7991 (
      {stage2_10[147]},
      {stage3_10[83]}
   );
   gpc1_1 gpc7992 (
      {stage2_10[148]},
      {stage3_10[84]}
   );
   gpc1_1 gpc7993 (
      {stage2_10[149]},
      {stage3_10[85]}
   );
   gpc1_1 gpc7994 (
      {stage2_10[150]},
      {stage3_10[86]}
   );
   gpc1_1 gpc7995 (
      {stage2_10[151]},
      {stage3_10[87]}
   );
   gpc1_1 gpc7996 (
      {stage2_10[152]},
      {stage3_10[88]}
   );
   gpc1_1 gpc7997 (
      {stage2_10[153]},
      {stage3_10[89]}
   );
   gpc1_1 gpc7998 (
      {stage2_10[154]},
      {stage3_10[90]}
   );
   gpc1_1 gpc7999 (
      {stage2_10[155]},
      {stage3_10[91]}
   );
   gpc1_1 gpc8000 (
      {stage2_10[156]},
      {stage3_10[92]}
   );
   gpc1_1 gpc8001 (
      {stage2_10[157]},
      {stage3_10[93]}
   );
   gpc1_1 gpc8002 (
      {stage2_10[158]},
      {stage3_10[94]}
   );
   gpc1_1 gpc8003 (
      {stage2_10[159]},
      {stage3_10[95]}
   );
   gpc1_1 gpc8004 (
      {stage2_10[160]},
      {stage3_10[96]}
   );
   gpc1_1 gpc8005 (
      {stage2_10[161]},
      {stage3_10[97]}
   );
   gpc1_1 gpc8006 (
      {stage2_10[162]},
      {stage3_10[98]}
   );
   gpc1_1 gpc8007 (
      {stage2_10[163]},
      {stage3_10[99]}
   );
   gpc1_1 gpc8008 (
      {stage2_11[127]},
      {stage3_11[46]}
   );
   gpc1_1 gpc8009 (
      {stage2_11[128]},
      {stage3_11[47]}
   );
   gpc1_1 gpc8010 (
      {stage2_11[129]},
      {stage3_11[48]}
   );
   gpc1_1 gpc8011 (
      {stage2_11[130]},
      {stage3_11[49]}
   );
   gpc1_1 gpc8012 (
      {stage2_11[131]},
      {stage3_11[50]}
   );
   gpc1_1 gpc8013 (
      {stage2_11[132]},
      {stage3_11[51]}
   );
   gpc1_1 gpc8014 (
      {stage2_11[133]},
      {stage3_11[52]}
   );
   gpc1_1 gpc8015 (
      {stage2_11[134]},
      {stage3_11[53]}
   );
   gpc1_1 gpc8016 (
      {stage2_11[135]},
      {stage3_11[54]}
   );
   gpc1_1 gpc8017 (
      {stage2_11[136]},
      {stage3_11[55]}
   );
   gpc1_1 gpc8018 (
      {stage2_11[137]},
      {stage3_11[56]}
   );
   gpc1_1 gpc8019 (
      {stage2_11[138]},
      {stage3_11[57]}
   );
   gpc1_1 gpc8020 (
      {stage2_12[92]},
      {stage3_12[53]}
   );
   gpc1_1 gpc8021 (
      {stage2_12[93]},
      {stage3_12[54]}
   );
   gpc1_1 gpc8022 (
      {stage2_12[94]},
      {stage3_12[55]}
   );
   gpc1_1 gpc8023 (
      {stage2_12[95]},
      {stage3_12[56]}
   );
   gpc1_1 gpc8024 (
      {stage2_12[96]},
      {stage3_12[57]}
   );
   gpc1_1 gpc8025 (
      {stage2_12[97]},
      {stage3_12[58]}
   );
   gpc1_1 gpc8026 (
      {stage2_12[98]},
      {stage3_12[59]}
   );
   gpc1_1 gpc8027 (
      {stage2_12[99]},
      {stage3_12[60]}
   );
   gpc1_1 gpc8028 (
      {stage2_12[100]},
      {stage3_12[61]}
   );
   gpc1_1 gpc8029 (
      {stage2_12[101]},
      {stage3_12[62]}
   );
   gpc1_1 gpc8030 (
      {stage2_12[102]},
      {stage3_12[63]}
   );
   gpc1_1 gpc8031 (
      {stage2_12[103]},
      {stage3_12[64]}
   );
   gpc1_1 gpc8032 (
      {stage2_12[104]},
      {stage3_12[65]}
   );
   gpc1_1 gpc8033 (
      {stage2_12[105]},
      {stage3_12[66]}
   );
   gpc1_1 gpc8034 (
      {stage2_12[106]},
      {stage3_12[67]}
   );
   gpc1_1 gpc8035 (
      {stage2_13[66]},
      {stage3_13[45]}
   );
   gpc1_1 gpc8036 (
      {stage2_13[67]},
      {stage3_13[46]}
   );
   gpc1_1 gpc8037 (
      {stage2_13[68]},
      {stage3_13[47]}
   );
   gpc1_1 gpc8038 (
      {stage2_13[69]},
      {stage3_13[48]}
   );
   gpc1_1 gpc8039 (
      {stage2_13[70]},
      {stage3_13[49]}
   );
   gpc1_1 gpc8040 (
      {stage2_13[71]},
      {stage3_13[50]}
   );
   gpc1_1 gpc8041 (
      {stage2_13[72]},
      {stage3_13[51]}
   );
   gpc1_1 gpc8042 (
      {stage2_13[73]},
      {stage3_13[52]}
   );
   gpc1_1 gpc8043 (
      {stage2_13[74]},
      {stage3_13[53]}
   );
   gpc1_1 gpc8044 (
      {stage2_13[75]},
      {stage3_13[54]}
   );
   gpc1_1 gpc8045 (
      {stage2_13[76]},
      {stage3_13[55]}
   );
   gpc1_1 gpc8046 (
      {stage2_13[77]},
      {stage3_13[56]}
   );
   gpc1_1 gpc8047 (
      {stage2_15[138]},
      {stage3_15[45]}
   );
   gpc1_1 gpc8048 (
      {stage2_15[139]},
      {stage3_15[46]}
   );
   gpc1_1 gpc8049 (
      {stage2_15[140]},
      {stage3_15[47]}
   );
   gpc1_1 gpc8050 (
      {stage2_16[80]},
      {stage3_16[48]}
   );
   gpc1_1 gpc8051 (
      {stage2_16[81]},
      {stage3_16[49]}
   );
   gpc1_1 gpc8052 (
      {stage2_16[82]},
      {stage3_16[50]}
   );
   gpc1_1 gpc8053 (
      {stage2_18[100]},
      {stage3_18[41]}
   );
   gpc1_1 gpc8054 (
      {stage2_18[101]},
      {stage3_18[42]}
   );
   gpc1_1 gpc8055 (
      {stage2_18[102]},
      {stage3_18[43]}
   );
   gpc1_1 gpc8056 (
      {stage2_18[103]},
      {stage3_18[44]}
   );
   gpc1_1 gpc8057 (
      {stage2_18[104]},
      {stage3_18[45]}
   );
   gpc1_1 gpc8058 (
      {stage2_18[105]},
      {stage3_18[46]}
   );
   gpc1_1 gpc8059 (
      {stage2_18[106]},
      {stage3_18[47]}
   );
   gpc1_1 gpc8060 (
      {stage2_18[107]},
      {stage3_18[48]}
   );
   gpc1_1 gpc8061 (
      {stage2_18[108]},
      {stage3_18[49]}
   );
   gpc1_1 gpc8062 (
      {stage2_18[109]},
      {stage3_18[50]}
   );
   gpc1_1 gpc8063 (
      {stage2_18[110]},
      {stage3_18[51]}
   );
   gpc1_1 gpc8064 (
      {stage2_18[111]},
      {stage3_18[52]}
   );
   gpc1_1 gpc8065 (
      {stage2_18[112]},
      {stage3_18[53]}
   );
   gpc1_1 gpc8066 (
      {stage2_18[113]},
      {stage3_18[54]}
   );
   gpc1_1 gpc8067 (
      {stage2_18[114]},
      {stage3_18[55]}
   );
   gpc1_1 gpc8068 (
      {stage2_18[115]},
      {stage3_18[56]}
   );
   gpc1_1 gpc8069 (
      {stage2_18[116]},
      {stage3_18[57]}
   );
   gpc1_1 gpc8070 (
      {stage2_18[117]},
      {stage3_18[58]}
   );
   gpc1_1 gpc8071 (
      {stage2_18[118]},
      {stage3_18[59]}
   );
   gpc1_1 gpc8072 (
      {stage2_20[45]},
      {stage3_20[35]}
   );
   gpc1_1 gpc8073 (
      {stage2_20[46]},
      {stage3_20[36]}
   );
   gpc1_1 gpc8074 (
      {stage2_20[47]},
      {stage3_20[37]}
   );
   gpc1_1 gpc8075 (
      {stage2_20[48]},
      {stage3_20[38]}
   );
   gpc1_1 gpc8076 (
      {stage2_20[49]},
      {stage3_20[39]}
   );
   gpc1_1 gpc8077 (
      {stage2_20[50]},
      {stage3_20[40]}
   );
   gpc1_1 gpc8078 (
      {stage2_20[51]},
      {stage3_20[41]}
   );
   gpc1_1 gpc8079 (
      {stage2_20[52]},
      {stage3_20[42]}
   );
   gpc1_1 gpc8080 (
      {stage2_20[53]},
      {stage3_20[43]}
   );
   gpc1_1 gpc8081 (
      {stage2_20[54]},
      {stage3_20[44]}
   );
   gpc1_1 gpc8082 (
      {stage2_20[55]},
      {stage3_20[45]}
   );
   gpc1_1 gpc8083 (
      {stage2_20[56]},
      {stage3_20[46]}
   );
   gpc1_1 gpc8084 (
      {stage2_20[57]},
      {stage3_20[47]}
   );
   gpc1_1 gpc8085 (
      {stage2_20[58]},
      {stage3_20[48]}
   );
   gpc1_1 gpc8086 (
      {stage2_20[59]},
      {stage3_20[49]}
   );
   gpc1_1 gpc8087 (
      {stage2_20[60]},
      {stage3_20[50]}
   );
   gpc1_1 gpc8088 (
      {stage2_20[61]},
      {stage3_20[51]}
   );
   gpc1_1 gpc8089 (
      {stage2_20[62]},
      {stage3_20[52]}
   );
   gpc1_1 gpc8090 (
      {stage2_20[63]},
      {stage3_20[53]}
   );
   gpc1_1 gpc8091 (
      {stage2_20[64]},
      {stage3_20[54]}
   );
   gpc1_1 gpc8092 (
      {stage2_20[65]},
      {stage3_20[55]}
   );
   gpc1_1 gpc8093 (
      {stage2_20[66]},
      {stage3_20[56]}
   );
   gpc1_1 gpc8094 (
      {stage2_20[67]},
      {stage3_20[57]}
   );
   gpc1_1 gpc8095 (
      {stage2_20[68]},
      {stage3_20[58]}
   );
   gpc1_1 gpc8096 (
      {stage2_20[69]},
      {stage3_20[59]}
   );
   gpc1_1 gpc8097 (
      {stage2_20[70]},
      {stage3_20[60]}
   );
   gpc1_1 gpc8098 (
      {stage2_20[71]},
      {stage3_20[61]}
   );
   gpc1_1 gpc8099 (
      {stage2_20[72]},
      {stage3_20[62]}
   );
   gpc1_1 gpc8100 (
      {stage2_20[73]},
      {stage3_20[63]}
   );
   gpc1_1 gpc8101 (
      {stage2_20[74]},
      {stage3_20[64]}
   );
   gpc1_1 gpc8102 (
      {stage2_20[75]},
      {stage3_20[65]}
   );
   gpc1_1 gpc8103 (
      {stage2_20[76]},
      {stage3_20[66]}
   );
   gpc1_1 gpc8104 (
      {stage2_20[77]},
      {stage3_20[67]}
   );
   gpc1_1 gpc8105 (
      {stage2_20[78]},
      {stage3_20[68]}
   );
   gpc1_1 gpc8106 (
      {stage2_20[79]},
      {stage3_20[69]}
   );
   gpc1_1 gpc8107 (
      {stage2_20[80]},
      {stage3_20[70]}
   );
   gpc1_1 gpc8108 (
      {stage2_20[81]},
      {stage3_20[71]}
   );
   gpc1_1 gpc8109 (
      {stage2_20[82]},
      {stage3_20[72]}
   );
   gpc1_1 gpc8110 (
      {stage2_20[83]},
      {stage3_20[73]}
   );
   gpc1_1 gpc8111 (
      {stage2_20[84]},
      {stage3_20[74]}
   );
   gpc1_1 gpc8112 (
      {stage2_20[85]},
      {stage3_20[75]}
   );
   gpc1_1 gpc8113 (
      {stage2_20[86]},
      {stage3_20[76]}
   );
   gpc1_1 gpc8114 (
      {stage2_20[87]},
      {stage3_20[77]}
   );
   gpc1_1 gpc8115 (
      {stage2_20[88]},
      {stage3_20[78]}
   );
   gpc1_1 gpc8116 (
      {stage2_20[89]},
      {stage3_20[79]}
   );
   gpc1_1 gpc8117 (
      {stage2_20[90]},
      {stage3_20[80]}
   );
   gpc1_1 gpc8118 (
      {stage2_20[91]},
      {stage3_20[81]}
   );
   gpc1_1 gpc8119 (
      {stage2_20[92]},
      {stage3_20[82]}
   );
   gpc1_1 gpc8120 (
      {stage2_21[120]},
      {stage3_21[31]}
   );
   gpc1_1 gpc8121 (
      {stage2_21[121]},
      {stage3_21[32]}
   );
   gpc1_1 gpc8122 (
      {stage2_21[122]},
      {stage3_21[33]}
   );
   gpc1_1 gpc8123 (
      {stage2_21[123]},
      {stage3_21[34]}
   );
   gpc1_1 gpc8124 (
      {stage2_21[124]},
      {stage3_21[35]}
   );
   gpc1_1 gpc8125 (
      {stage2_21[125]},
      {stage3_21[36]}
   );
   gpc1_1 gpc8126 (
      {stage2_21[126]},
      {stage3_21[37]}
   );
   gpc1_1 gpc8127 (
      {stage2_21[127]},
      {stage3_21[38]}
   );
   gpc1_1 gpc8128 (
      {stage2_22[80]},
      {stage3_22[45]}
   );
   gpc1_1 gpc8129 (
      {stage2_22[81]},
      {stage3_22[46]}
   );
   gpc1_1 gpc8130 (
      {stage2_22[82]},
      {stage3_22[47]}
   );
   gpc1_1 gpc8131 (
      {stage2_22[83]},
      {stage3_22[48]}
   );
   gpc1_1 gpc8132 (
      {stage2_22[84]},
      {stage3_22[49]}
   );
   gpc1_1 gpc8133 (
      {stage2_22[85]},
      {stage3_22[50]}
   );
   gpc1_1 gpc8134 (
      {stage2_22[86]},
      {stage3_22[51]}
   );
   gpc1_1 gpc8135 (
      {stage2_22[87]},
      {stage3_22[52]}
   );
   gpc1_1 gpc8136 (
      {stage2_22[88]},
      {stage3_22[53]}
   );
   gpc1_1 gpc8137 (
      {stage2_22[89]},
      {stage3_22[54]}
   );
   gpc1_1 gpc8138 (
      {stage2_22[90]},
      {stage3_22[55]}
   );
   gpc1_1 gpc8139 (
      {stage2_22[91]},
      {stage3_22[56]}
   );
   gpc1_1 gpc8140 (
      {stage2_22[92]},
      {stage3_22[57]}
   );
   gpc1_1 gpc8141 (
      {stage2_22[93]},
      {stage3_22[58]}
   );
   gpc1_1 gpc8142 (
      {stage2_22[94]},
      {stage3_22[59]}
   );
   gpc1_1 gpc8143 (
      {stage2_22[95]},
      {stage3_22[60]}
   );
   gpc1_1 gpc8144 (
      {stage2_22[96]},
      {stage3_22[61]}
   );
   gpc1_1 gpc8145 (
      {stage2_22[97]},
      {stage3_22[62]}
   );
   gpc1_1 gpc8146 (
      {stage2_22[98]},
      {stage3_22[63]}
   );
   gpc1_1 gpc8147 (
      {stage2_22[99]},
      {stage3_22[64]}
   );
   gpc1_1 gpc8148 (
      {stage2_22[100]},
      {stage3_22[65]}
   );
   gpc1_1 gpc8149 (
      {stage2_22[101]},
      {stage3_22[66]}
   );
   gpc1_1 gpc8150 (
      {stage2_22[102]},
      {stage3_22[67]}
   );
   gpc1_1 gpc8151 (
      {stage2_22[103]},
      {stage3_22[68]}
   );
   gpc1_1 gpc8152 (
      {stage2_22[104]},
      {stage3_22[69]}
   );
   gpc1_1 gpc8153 (
      {stage2_22[105]},
      {stage3_22[70]}
   );
   gpc1_1 gpc8154 (
      {stage2_22[106]},
      {stage3_22[71]}
   );
   gpc1_1 gpc8155 (
      {stage2_22[107]},
      {stage3_22[72]}
   );
   gpc1_1 gpc8156 (
      {stage2_26[83]},
      {stage3_26[47]}
   );
   gpc1_1 gpc8157 (
      {stage2_26[84]},
      {stage3_26[48]}
   );
   gpc1_1 gpc8158 (
      {stage2_27[93]},
      {stage3_27[36]}
   );
   gpc1_1 gpc8159 (
      {stage2_27[94]},
      {stage3_27[37]}
   );
   gpc1_1 gpc8160 (
      {stage2_27[95]},
      {stage3_27[38]}
   );
   gpc1_1 gpc8161 (
      {stage2_27[96]},
      {stage3_27[39]}
   );
   gpc1_1 gpc8162 (
      {stage2_27[97]},
      {stage3_27[40]}
   );
   gpc1_1 gpc8163 (
      {stage2_27[98]},
      {stage3_27[41]}
   );
   gpc1_1 gpc8164 (
      {stage2_27[99]},
      {stage3_27[42]}
   );
   gpc1_1 gpc8165 (
      {stage2_27[100]},
      {stage3_27[43]}
   );
   gpc1_1 gpc8166 (
      {stage2_27[101]},
      {stage3_27[44]}
   );
   gpc1_1 gpc8167 (
      {stage2_27[102]},
      {stage3_27[45]}
   );
   gpc1_1 gpc8168 (
      {stage2_27[103]},
      {stage3_27[46]}
   );
   gpc1_1 gpc8169 (
      {stage2_27[104]},
      {stage3_27[47]}
   );
   gpc1_1 gpc8170 (
      {stage2_27[105]},
      {stage3_27[48]}
   );
   gpc1_1 gpc8171 (
      {stage2_28[69]},
      {stage3_28[34]}
   );
   gpc1_1 gpc8172 (
      {stage2_28[70]},
      {stage3_28[35]}
   );
   gpc1_1 gpc8173 (
      {stage2_28[71]},
      {stage3_28[36]}
   );
   gpc1_1 gpc8174 (
      {stage2_28[72]},
      {stage3_28[37]}
   );
   gpc1_1 gpc8175 (
      {stage2_28[73]},
      {stage3_28[38]}
   );
   gpc1_1 gpc8176 (
      {stage2_28[74]},
      {stage3_28[39]}
   );
   gpc1_1 gpc8177 (
      {stage2_28[75]},
      {stage3_28[40]}
   );
   gpc1_1 gpc8178 (
      {stage2_28[76]},
      {stage3_28[41]}
   );
   gpc1_1 gpc8179 (
      {stage2_28[77]},
      {stage3_28[42]}
   );
   gpc1_1 gpc8180 (
      {stage2_28[78]},
      {stage3_28[43]}
   );
   gpc1_1 gpc8181 (
      {stage2_28[79]},
      {stage3_28[44]}
   );
   gpc1_1 gpc8182 (
      {stage2_28[80]},
      {stage3_28[45]}
   );
   gpc1_1 gpc8183 (
      {stage2_28[81]},
      {stage3_28[46]}
   );
   gpc1_1 gpc8184 (
      {stage2_28[82]},
      {stage3_28[47]}
   );
   gpc1_1 gpc8185 (
      {stage2_28[83]},
      {stage3_28[48]}
   );
   gpc1_1 gpc8186 (
      {stage2_28[84]},
      {stage3_28[49]}
   );
   gpc1_1 gpc8187 (
      {stage2_28[85]},
      {stage3_28[50]}
   );
   gpc1_1 gpc8188 (
      {stage2_28[86]},
      {stage3_28[51]}
   );
   gpc1_1 gpc8189 (
      {stage2_28[87]},
      {stage3_28[52]}
   );
   gpc1_1 gpc8190 (
      {stage2_28[88]},
      {stage3_28[53]}
   );
   gpc1_1 gpc8191 (
      {stage2_28[89]},
      {stage3_28[54]}
   );
   gpc1_1 gpc8192 (
      {stage2_28[90]},
      {stage3_28[55]}
   );
   gpc1_1 gpc8193 (
      {stage2_28[91]},
      {stage3_28[56]}
   );
   gpc1_1 gpc8194 (
      {stage2_30[103]},
      {stage3_30[28]}
   );
   gpc1_1 gpc8195 (
      {stage2_30[104]},
      {stage3_30[29]}
   );
   gpc1_1 gpc8196 (
      {stage2_30[105]},
      {stage3_30[30]}
   );
   gpc1_1 gpc8197 (
      {stage2_30[106]},
      {stage3_30[31]}
   );
   gpc1_1 gpc8198 (
      {stage2_30[107]},
      {stage3_30[32]}
   );
   gpc1_1 gpc8199 (
      {stage2_30[108]},
      {stage3_30[33]}
   );
   gpc1_1 gpc8200 (
      {stage2_30[109]},
      {stage3_30[34]}
   );
   gpc1_1 gpc8201 (
      {stage2_30[110]},
      {stage3_30[35]}
   );
   gpc1_1 gpc8202 (
      {stage2_30[111]},
      {stage3_30[36]}
   );
   gpc1_1 gpc8203 (
      {stage2_30[112]},
      {stage3_30[37]}
   );
   gpc1_1 gpc8204 (
      {stage2_30[113]},
      {stage3_30[38]}
   );
   gpc1_1 gpc8205 (
      {stage2_30[114]},
      {stage3_30[39]}
   );
   gpc1_1 gpc8206 (
      {stage2_30[115]},
      {stage3_30[40]}
   );
   gpc1_1 gpc8207 (
      {stage2_30[116]},
      {stage3_30[41]}
   );
   gpc1_1 gpc8208 (
      {stage2_31[95]},
      {stage3_31[34]}
   );
   gpc1_1 gpc8209 (
      {stage2_31[96]},
      {stage3_31[35]}
   );
   gpc1_1 gpc8210 (
      {stage2_31[97]},
      {stage3_31[36]}
   );
   gpc1_1 gpc8211 (
      {stage2_31[98]},
      {stage3_31[37]}
   );
   gpc1_1 gpc8212 (
      {stage2_32[99]},
      {stage3_32[47]}
   );
   gpc1_1 gpc8213 (
      {stage2_32[100]},
      {stage3_32[48]}
   );
   gpc1_1 gpc8214 (
      {stage2_32[101]},
      {stage3_32[49]}
   );
   gpc1_1 gpc8215 (
      {stage2_32[102]},
      {stage3_32[50]}
   );
   gpc1_1 gpc8216 (
      {stage2_32[103]},
      {stage3_32[51]}
   );
   gpc1_1 gpc8217 (
      {stage2_32[104]},
      {stage3_32[52]}
   );
   gpc1_1 gpc8218 (
      {stage2_32[105]},
      {stage3_32[53]}
   );
   gpc1_1 gpc8219 (
      {stage2_33[72]},
      {stage3_33[42]}
   );
   gpc1_1 gpc8220 (
      {stage2_33[73]},
      {stage3_33[43]}
   );
   gpc1_1 gpc8221 (
      {stage2_33[74]},
      {stage3_33[44]}
   );
   gpc1_1 gpc8222 (
      {stage2_33[75]},
      {stage3_33[45]}
   );
   gpc1_1 gpc8223 (
      {stage2_34[129]},
      {stage3_34[39]}
   );
   gpc1_1 gpc8224 (
      {stage2_34[130]},
      {stage3_34[40]}
   );
   gpc1_1 gpc8225 (
      {stage2_34[131]},
      {stage3_34[41]}
   );
   gpc1_1 gpc8226 (
      {stage2_35[120]},
      {stage3_35[44]}
   );
   gpc1_1 gpc8227 (
      {stage2_35[121]},
      {stage3_35[45]}
   );
   gpc1_1 gpc8228 (
      {stage2_35[122]},
      {stage3_35[46]}
   );
   gpc1_1 gpc8229 (
      {stage2_35[123]},
      {stage3_35[47]}
   );
   gpc1_1 gpc8230 (
      {stage2_35[124]},
      {stage3_35[48]}
   );
   gpc1_1 gpc8231 (
      {stage2_35[125]},
      {stage3_35[49]}
   );
   gpc1_1 gpc8232 (
      {stage2_35[126]},
      {stage3_35[50]}
   );
   gpc1_1 gpc8233 (
      {stage2_35[127]},
      {stage3_35[51]}
   );
   gpc1_1 gpc8234 (
      {stage2_35[128]},
      {stage3_35[52]}
   );
   gpc1_1 gpc8235 (
      {stage2_35[129]},
      {stage3_35[53]}
   );
   gpc1_1 gpc8236 (
      {stage2_35[130]},
      {stage3_35[54]}
   );
   gpc1_1 gpc8237 (
      {stage2_35[131]},
      {stage3_35[55]}
   );
   gpc1_1 gpc8238 (
      {stage2_35[132]},
      {stage3_35[56]}
   );
   gpc1_1 gpc8239 (
      {stage2_36[73]},
      {stage3_36[44]}
   );
   gpc1_1 gpc8240 (
      {stage2_36[74]},
      {stage3_36[45]}
   );
   gpc1_1 gpc8241 (
      {stage2_37[74]},
      {stage3_37[37]}
   );
   gpc1_1 gpc8242 (
      {stage2_37[75]},
      {stage3_37[38]}
   );
   gpc1_1 gpc8243 (
      {stage2_37[76]},
      {stage3_37[39]}
   );
   gpc1_1 gpc8244 (
      {stage2_37[77]},
      {stage3_37[40]}
   );
   gpc1_1 gpc8245 (
      {stage2_37[78]},
      {stage3_37[41]}
   );
   gpc1_1 gpc8246 (
      {stage2_37[79]},
      {stage3_37[42]}
   );
   gpc1_1 gpc8247 (
      {stage2_37[80]},
      {stage3_37[43]}
   );
   gpc1_1 gpc8248 (
      {stage2_37[81]},
      {stage3_37[44]}
   );
   gpc1_1 gpc8249 (
      {stage2_37[82]},
      {stage3_37[45]}
   );
   gpc1_1 gpc8250 (
      {stage2_37[83]},
      {stage3_37[46]}
   );
   gpc1_1 gpc8251 (
      {stage2_37[84]},
      {stage3_37[47]}
   );
   gpc1_1 gpc8252 (
      {stage2_37[85]},
      {stage3_37[48]}
   );
   gpc1_1 gpc8253 (
      {stage2_37[86]},
      {stage3_37[49]}
   );
   gpc1_1 gpc8254 (
      {stage2_37[87]},
      {stage3_37[50]}
   );
   gpc1_1 gpc8255 (
      {stage2_37[88]},
      {stage3_37[51]}
   );
   gpc1_1 gpc8256 (
      {stage2_37[89]},
      {stage3_37[52]}
   );
   gpc1_1 gpc8257 (
      {stage2_38[125]},
      {stage3_38[45]}
   );
   gpc1_1 gpc8258 (
      {stage2_38[126]},
      {stage3_38[46]}
   );
   gpc1_1 gpc8259 (
      {stage2_38[127]},
      {stage3_38[47]}
   );
   gpc1_1 gpc8260 (
      {stage2_38[128]},
      {stage3_38[48]}
   );
   gpc1_1 gpc8261 (
      {stage2_38[129]},
      {stage3_38[49]}
   );
   gpc1_1 gpc8262 (
      {stage2_38[130]},
      {stage3_38[50]}
   );
   gpc1_1 gpc8263 (
      {stage2_38[131]},
      {stage3_38[51]}
   );
   gpc1_1 gpc8264 (
      {stage2_38[132]},
      {stage3_38[52]}
   );
   gpc1_1 gpc8265 (
      {stage2_38[133]},
      {stage3_38[53]}
   );
   gpc1_1 gpc8266 (
      {stage2_38[134]},
      {stage3_38[54]}
   );
   gpc1_1 gpc8267 (
      {stage2_38[135]},
      {stage3_38[55]}
   );
   gpc1_1 gpc8268 (
      {stage2_38[136]},
      {stage3_38[56]}
   );
   gpc1_1 gpc8269 (
      {stage2_38[137]},
      {stage3_38[57]}
   );
   gpc1_1 gpc8270 (
      {stage2_38[138]},
      {stage3_38[58]}
   );
   gpc1_1 gpc8271 (
      {stage2_38[139]},
      {stage3_38[59]}
   );
   gpc1_1 gpc8272 (
      {stage2_39[128]},
      {stage3_39[49]}
   );
   gpc1_1 gpc8273 (
      {stage2_39[129]},
      {stage3_39[50]}
   );
   gpc1_1 gpc8274 (
      {stage2_39[130]},
      {stage3_39[51]}
   );
   gpc1_1 gpc8275 (
      {stage2_39[131]},
      {stage3_39[52]}
   );
   gpc1_1 gpc8276 (
      {stage2_39[132]},
      {stage3_39[53]}
   );
   gpc1_1 gpc8277 (
      {stage2_39[133]},
      {stage3_39[54]}
   );
   gpc1_1 gpc8278 (
      {stage2_39[134]},
      {stage3_39[55]}
   );
   gpc1_1 gpc8279 (
      {stage2_39[135]},
      {stage3_39[56]}
   );
   gpc1_1 gpc8280 (
      {stage2_39[136]},
      {stage3_39[57]}
   );
   gpc1_1 gpc8281 (
      {stage2_40[107]},
      {stage3_40[46]}
   );
   gpc1_1 gpc8282 (
      {stage2_40[108]},
      {stage3_40[47]}
   );
   gpc1_1 gpc8283 (
      {stage2_40[109]},
      {stage3_40[48]}
   );
   gpc1_1 gpc8284 (
      {stage2_40[110]},
      {stage3_40[49]}
   );
   gpc1_1 gpc8285 (
      {stage2_40[111]},
      {stage3_40[50]}
   );
   gpc1_1 gpc8286 (
      {stage2_40[112]},
      {stage3_40[51]}
   );
   gpc1_1 gpc8287 (
      {stage2_41[102]},
      {stage3_41[39]}
   );
   gpc1_1 gpc8288 (
      {stage2_41[103]},
      {stage3_41[40]}
   );
   gpc1_1 gpc8289 (
      {stage2_41[104]},
      {stage3_41[41]}
   );
   gpc1_1 gpc8290 (
      {stage2_41[105]},
      {stage3_41[42]}
   );
   gpc1_1 gpc8291 (
      {stage2_42[82]},
      {stage3_42[46]}
   );
   gpc1_1 gpc8292 (
      {stage2_42[83]},
      {stage3_42[47]}
   );
   gpc1_1 gpc8293 (
      {stage2_42[84]},
      {stage3_42[48]}
   );
   gpc1_1 gpc8294 (
      {stage2_42[85]},
      {stage3_42[49]}
   );
   gpc1_1 gpc8295 (
      {stage2_44[109]},
      {stage3_44[31]}
   );
   gpc1_1 gpc8296 (
      {stage2_44[110]},
      {stage3_44[32]}
   );
   gpc1_1 gpc8297 (
      {stage2_44[111]},
      {stage3_44[33]}
   );
   gpc1_1 gpc8298 (
      {stage2_44[112]},
      {stage3_44[34]}
   );
   gpc1_1 gpc8299 (
      {stage2_44[113]},
      {stage3_44[35]}
   );
   gpc1_1 gpc8300 (
      {stage2_44[114]},
      {stage3_44[36]}
   );
   gpc1_1 gpc8301 (
      {stage2_44[115]},
      {stage3_44[37]}
   );
   gpc1_1 gpc8302 (
      {stage2_44[116]},
      {stage3_44[38]}
   );
   gpc1_1 gpc8303 (
      {stage2_44[117]},
      {stage3_44[39]}
   );
   gpc1_1 gpc8304 (
      {stage2_44[118]},
      {stage3_44[40]}
   );
   gpc1_1 gpc8305 (
      {stage2_45[108]},
      {stage3_45[34]}
   );
   gpc1_1 gpc8306 (
      {stage2_45[109]},
      {stage3_45[35]}
   );
   gpc1_1 gpc8307 (
      {stage2_45[110]},
      {stage3_45[36]}
   );
   gpc1_1 gpc8308 (
      {stage2_45[111]},
      {stage3_45[37]}
   );
   gpc1_1 gpc8309 (
      {stage2_45[112]},
      {stage3_45[38]}
   );
   gpc1_1 gpc8310 (
      {stage2_45[113]},
      {stage3_45[39]}
   );
   gpc1_1 gpc8311 (
      {stage2_45[114]},
      {stage3_45[40]}
   );
   gpc1_1 gpc8312 (
      {stage2_45[115]},
      {stage3_45[41]}
   );
   gpc1_1 gpc8313 (
      {stage2_45[116]},
      {stage3_45[42]}
   );
   gpc1_1 gpc8314 (
      {stage2_45[117]},
      {stage3_45[43]}
   );
   gpc1_1 gpc8315 (
      {stage2_46[78]},
      {stage3_46[48]}
   );
   gpc1_1 gpc8316 (
      {stage2_46[79]},
      {stage3_46[49]}
   );
   gpc1_1 gpc8317 (
      {stage2_46[80]},
      {stage3_46[50]}
   );
   gpc1_1 gpc8318 (
      {stage2_46[81]},
      {stage3_46[51]}
   );
   gpc1_1 gpc8319 (
      {stage2_46[82]},
      {stage3_46[52]}
   );
   gpc1_1 gpc8320 (
      {stage2_46[83]},
      {stage3_46[53]}
   );
   gpc1_1 gpc8321 (
      {stage2_46[84]},
      {stage3_46[54]}
   );
   gpc1_1 gpc8322 (
      {stage2_46[85]},
      {stage3_46[55]}
   );
   gpc1_1 gpc8323 (
      {stage2_46[86]},
      {stage3_46[56]}
   );
   gpc1_1 gpc8324 (
      {stage2_46[87]},
      {stage3_46[57]}
   );
   gpc1_1 gpc8325 (
      {stage2_48[126]},
      {stage3_48[38]}
   );
   gpc1_1 gpc8326 (
      {stage2_48[127]},
      {stage3_48[39]}
   );
   gpc1_1 gpc8327 (
      {stage2_48[128]},
      {stage3_48[40]}
   );
   gpc1_1 gpc8328 (
      {stage2_48[129]},
      {stage3_48[41]}
   );
   gpc1_1 gpc8329 (
      {stage2_50[84]},
      {stage3_50[45]}
   );
   gpc1_1 gpc8330 (
      {stage2_50[85]},
      {stage3_50[46]}
   );
   gpc1_1 gpc8331 (
      {stage2_51[59]},
      {stage3_51[34]}
   );
   gpc1_1 gpc8332 (
      {stage2_51[60]},
      {stage3_51[35]}
   );
   gpc1_1 gpc8333 (
      {stage2_51[61]},
      {stage3_51[36]}
   );
   gpc1_1 gpc8334 (
      {stage2_51[62]},
      {stage3_51[37]}
   );
   gpc1_1 gpc8335 (
      {stage2_51[63]},
      {stage3_51[38]}
   );
   gpc1_1 gpc8336 (
      {stage2_51[64]},
      {stage3_51[39]}
   );
   gpc1_1 gpc8337 (
      {stage2_51[65]},
      {stage3_51[40]}
   );
   gpc1_1 gpc8338 (
      {stage2_51[66]},
      {stage3_51[41]}
   );
   gpc1_1 gpc8339 (
      {stage2_51[67]},
      {stage3_51[42]}
   );
   gpc1_1 gpc8340 (
      {stage2_51[68]},
      {stage3_51[43]}
   );
   gpc1_1 gpc8341 (
      {stage2_51[69]},
      {stage3_51[44]}
   );
   gpc1_1 gpc8342 (
      {stage2_51[70]},
      {stage3_51[45]}
   );
   gpc1_1 gpc8343 (
      {stage2_51[71]},
      {stage3_51[46]}
   );
   gpc1_1 gpc8344 (
      {stage2_51[72]},
      {stage3_51[47]}
   );
   gpc1_1 gpc8345 (
      {stage2_51[73]},
      {stage3_51[48]}
   );
   gpc1_1 gpc8346 (
      {stage2_51[74]},
      {stage3_51[49]}
   );
   gpc1_1 gpc8347 (
      {stage2_51[75]},
      {stage3_51[50]}
   );
   gpc1_1 gpc8348 (
      {stage2_51[76]},
      {stage3_51[51]}
   );
   gpc1_1 gpc8349 (
      {stage2_51[77]},
      {stage3_51[52]}
   );
   gpc1_1 gpc8350 (
      {stage2_51[78]},
      {stage3_51[53]}
   );
   gpc1_1 gpc8351 (
      {stage2_51[79]},
      {stage3_51[54]}
   );
   gpc1_1 gpc8352 (
      {stage2_51[80]},
      {stage3_51[55]}
   );
   gpc1_1 gpc8353 (
      {stage2_51[81]},
      {stage3_51[56]}
   );
   gpc1_1 gpc8354 (
      {stage2_51[82]},
      {stage3_51[57]}
   );
   gpc1_1 gpc8355 (
      {stage2_51[83]},
      {stage3_51[58]}
   );
   gpc1_1 gpc8356 (
      {stage2_51[84]},
      {stage3_51[59]}
   );
   gpc1_1 gpc8357 (
      {stage2_51[85]},
      {stage3_51[60]}
   );
   gpc1_1 gpc8358 (
      {stage2_51[86]},
      {stage3_51[61]}
   );
   gpc1_1 gpc8359 (
      {stage2_51[87]},
      {stage3_51[62]}
   );
   gpc1_1 gpc8360 (
      {stage2_52[69]},
      {stage3_52[27]}
   );
   gpc1_1 gpc8361 (
      {stage2_52[70]},
      {stage3_52[28]}
   );
   gpc1_1 gpc8362 (
      {stage2_52[71]},
      {stage3_52[29]}
   );
   gpc1_1 gpc8363 (
      {stage2_52[72]},
      {stage3_52[30]}
   );
   gpc1_1 gpc8364 (
      {stage2_52[73]},
      {stage3_52[31]}
   );
   gpc1_1 gpc8365 (
      {stage2_52[74]},
      {stage3_52[32]}
   );
   gpc1_1 gpc8366 (
      {stage2_52[75]},
      {stage3_52[33]}
   );
   gpc1_1 gpc8367 (
      {stage2_52[76]},
      {stage3_52[34]}
   );
   gpc1_1 gpc8368 (
      {stage2_52[77]},
      {stage3_52[35]}
   );
   gpc1_1 gpc8369 (
      {stage2_52[78]},
      {stage3_52[36]}
   );
   gpc1_1 gpc8370 (
      {stage2_52[79]},
      {stage3_52[37]}
   );
   gpc1_1 gpc8371 (
      {stage2_52[80]},
      {stage3_52[38]}
   );
   gpc1_1 gpc8372 (
      {stage2_52[81]},
      {stage3_52[39]}
   );
   gpc1_1 gpc8373 (
      {stage2_52[82]},
      {stage3_52[40]}
   );
   gpc1_1 gpc8374 (
      {stage2_52[83]},
      {stage3_52[41]}
   );
   gpc1_1 gpc8375 (
      {stage2_52[84]},
      {stage3_52[42]}
   );
   gpc1_1 gpc8376 (
      {stage2_52[85]},
      {stage3_52[43]}
   );
   gpc1_1 gpc8377 (
      {stage2_52[86]},
      {stage3_52[44]}
   );
   gpc1_1 gpc8378 (
      {stage2_52[87]},
      {stage3_52[45]}
   );
   gpc1_1 gpc8379 (
      {stage2_52[88]},
      {stage3_52[46]}
   );
   gpc1_1 gpc8380 (
      {stage2_52[89]},
      {stage3_52[47]}
   );
   gpc1_1 gpc8381 (
      {stage2_52[90]},
      {stage3_52[48]}
   );
   gpc1_1 gpc8382 (
      {stage2_52[91]},
      {stage3_52[49]}
   );
   gpc1_1 gpc8383 (
      {stage2_52[92]},
      {stage3_52[50]}
   );
   gpc1_1 gpc8384 (
      {stage2_52[93]},
      {stage3_52[51]}
   );
   gpc1_1 gpc8385 (
      {stage2_52[94]},
      {stage3_52[52]}
   );
   gpc1_1 gpc8386 (
      {stage2_52[95]},
      {stage3_52[53]}
   );
   gpc1_1 gpc8387 (
      {stage2_52[96]},
      {stage3_52[54]}
   );
   gpc1_1 gpc8388 (
      {stage2_52[97]},
      {stage3_52[55]}
   );
   gpc1_1 gpc8389 (
      {stage2_52[98]},
      {stage3_52[56]}
   );
   gpc1_1 gpc8390 (
      {stage2_52[99]},
      {stage3_52[57]}
   );
   gpc1_1 gpc8391 (
      {stage2_52[100]},
      {stage3_52[58]}
   );
   gpc1_1 gpc8392 (
      {stage2_52[101]},
      {stage3_52[59]}
   );
   gpc1_1 gpc8393 (
      {stage2_52[102]},
      {stage3_52[60]}
   );
   gpc1_1 gpc8394 (
      {stage2_52[103]},
      {stage3_52[61]}
   );
   gpc1_1 gpc8395 (
      {stage2_52[104]},
      {stage3_52[62]}
   );
   gpc1_1 gpc8396 (
      {stage2_53[69]},
      {stage3_53[29]}
   );
   gpc1_1 gpc8397 (
      {stage2_53[70]},
      {stage3_53[30]}
   );
   gpc1_1 gpc8398 (
      {stage2_53[71]},
      {stage3_53[31]}
   );
   gpc1_1 gpc8399 (
      {stage2_53[72]},
      {stage3_53[32]}
   );
   gpc1_1 gpc8400 (
      {stage2_53[73]},
      {stage3_53[33]}
   );
   gpc1_1 gpc8401 (
      {stage2_53[74]},
      {stage3_53[34]}
   );
   gpc1_1 gpc8402 (
      {stage2_53[75]},
      {stage3_53[35]}
   );
   gpc1_1 gpc8403 (
      {stage2_53[76]},
      {stage3_53[36]}
   );
   gpc1_1 gpc8404 (
      {stage2_53[77]},
      {stage3_53[37]}
   );
   gpc1_1 gpc8405 (
      {stage2_53[78]},
      {stage3_53[38]}
   );
   gpc1_1 gpc8406 (
      {stage2_53[79]},
      {stage3_53[39]}
   );
   gpc1_1 gpc8407 (
      {stage2_53[80]},
      {stage3_53[40]}
   );
   gpc1_1 gpc8408 (
      {stage2_53[81]},
      {stage3_53[41]}
   );
   gpc1_1 gpc8409 (
      {stage2_53[82]},
      {stage3_53[42]}
   );
   gpc1_1 gpc8410 (
      {stage2_53[83]},
      {stage3_53[43]}
   );
   gpc1_1 gpc8411 (
      {stage2_53[84]},
      {stage3_53[44]}
   );
   gpc1_1 gpc8412 (
      {stage2_53[85]},
      {stage3_53[45]}
   );
   gpc1_1 gpc8413 (
      {stage2_53[86]},
      {stage3_53[46]}
   );
   gpc1_1 gpc8414 (
      {stage2_53[87]},
      {stage3_53[47]}
   );
   gpc1_1 gpc8415 (
      {stage2_53[88]},
      {stage3_53[48]}
   );
   gpc1_1 gpc8416 (
      {stage2_53[89]},
      {stage3_53[49]}
   );
   gpc1_1 gpc8417 (
      {stage2_53[90]},
      {stage3_53[50]}
   );
   gpc1_1 gpc8418 (
      {stage2_53[91]},
      {stage3_53[51]}
   );
   gpc1_1 gpc8419 (
      {stage2_53[92]},
      {stage3_53[52]}
   );
   gpc1_1 gpc8420 (
      {stage2_53[93]},
      {stage3_53[53]}
   );
   gpc1_1 gpc8421 (
      {stage2_53[94]},
      {stage3_53[54]}
   );
   gpc1_1 gpc8422 (
      {stage2_53[95]},
      {stage3_53[55]}
   );
   gpc1_1 gpc8423 (
      {stage2_53[96]},
      {stage3_53[56]}
   );
   gpc1_1 gpc8424 (
      {stage2_53[97]},
      {stage3_53[57]}
   );
   gpc1_1 gpc8425 (
      {stage2_53[98]},
      {stage3_53[58]}
   );
   gpc1_1 gpc8426 (
      {stage2_53[99]},
      {stage3_53[59]}
   );
   gpc1_1 gpc8427 (
      {stage2_53[100]},
      {stage3_53[60]}
   );
   gpc1_1 gpc8428 (
      {stage2_53[101]},
      {stage3_53[61]}
   );
   gpc1_1 gpc8429 (
      {stage2_53[102]},
      {stage3_53[62]}
   );
   gpc1_1 gpc8430 (
      {stage2_53[103]},
      {stage3_53[63]}
   );
   gpc1_1 gpc8431 (
      {stage2_53[104]},
      {stage3_53[64]}
   );
   gpc1_1 gpc8432 (
      {stage2_53[105]},
      {stage3_53[65]}
   );
   gpc1_1 gpc8433 (
      {stage2_53[106]},
      {stage3_53[66]}
   );
   gpc1_1 gpc8434 (
      {stage2_53[107]},
      {stage3_53[67]}
   );
   gpc1_1 gpc8435 (
      {stage2_53[108]},
      {stage3_53[68]}
   );
   gpc1_1 gpc8436 (
      {stage2_53[109]},
      {stage3_53[69]}
   );
   gpc1_1 gpc8437 (
      {stage2_53[110]},
      {stage3_53[70]}
   );
   gpc1_1 gpc8438 (
      {stage2_53[111]},
      {stage3_53[71]}
   );
   gpc1_1 gpc8439 (
      {stage2_53[112]},
      {stage3_53[72]}
   );
   gpc1_1 gpc8440 (
      {stage2_53[113]},
      {stage3_53[73]}
   );
   gpc1_1 gpc8441 (
      {stage2_53[114]},
      {stage3_53[74]}
   );
   gpc1_1 gpc8442 (
      {stage2_55[70]},
      {stage3_55[31]}
   );
   gpc1_1 gpc8443 (
      {stage2_55[71]},
      {stage3_55[32]}
   );
   gpc1_1 gpc8444 (
      {stage2_55[72]},
      {stage3_55[33]}
   );
   gpc1_1 gpc8445 (
      {stage2_55[73]},
      {stage3_55[34]}
   );
   gpc1_1 gpc8446 (
      {stage2_55[74]},
      {stage3_55[35]}
   );
   gpc1_1 gpc8447 (
      {stage2_55[75]},
      {stage3_55[36]}
   );
   gpc1_1 gpc8448 (
      {stage2_55[76]},
      {stage3_55[37]}
   );
   gpc1_1 gpc8449 (
      {stage2_55[77]},
      {stage3_55[38]}
   );
   gpc1_1 gpc8450 (
      {stage2_55[78]},
      {stage3_55[39]}
   );
   gpc1_1 gpc8451 (
      {stage2_55[79]},
      {stage3_55[40]}
   );
   gpc1_1 gpc8452 (
      {stage2_55[80]},
      {stage3_55[41]}
   );
   gpc1_1 gpc8453 (
      {stage2_55[81]},
      {stage3_55[42]}
   );
   gpc1_1 gpc8454 (
      {stage2_55[82]},
      {stage3_55[43]}
   );
   gpc1_1 gpc8455 (
      {stage2_55[83]},
      {stage3_55[44]}
   );
   gpc1_1 gpc8456 (
      {stage2_55[84]},
      {stage3_55[45]}
   );
   gpc1_1 gpc8457 (
      {stage2_55[85]},
      {stage3_55[46]}
   );
   gpc1_1 gpc8458 (
      {stage2_55[86]},
      {stage3_55[47]}
   );
   gpc1_1 gpc8459 (
      {stage2_55[87]},
      {stage3_55[48]}
   );
   gpc1_1 gpc8460 (
      {stage2_55[88]},
      {stage3_55[49]}
   );
   gpc1_1 gpc8461 (
      {stage2_55[89]},
      {stage3_55[50]}
   );
   gpc1_1 gpc8462 (
      {stage2_55[90]},
      {stage3_55[51]}
   );
   gpc1_1 gpc8463 (
      {stage2_55[91]},
      {stage3_55[52]}
   );
   gpc1_1 gpc8464 (
      {stage2_55[92]},
      {stage3_55[53]}
   );
   gpc1_1 gpc8465 (
      {stage2_55[93]},
      {stage3_55[54]}
   );
   gpc1_1 gpc8466 (
      {stage2_55[94]},
      {stage3_55[55]}
   );
   gpc1_1 gpc8467 (
      {stage2_55[95]},
      {stage3_55[56]}
   );
   gpc1_1 gpc8468 (
      {stage2_55[96]},
      {stage3_55[57]}
   );
   gpc1_1 gpc8469 (
      {stage2_55[97]},
      {stage3_55[58]}
   );
   gpc1_1 gpc8470 (
      {stage2_55[98]},
      {stage3_55[59]}
   );
   gpc1_1 gpc8471 (
      {stage2_55[99]},
      {stage3_55[60]}
   );
   gpc1_1 gpc8472 (
      {stage2_55[100]},
      {stage3_55[61]}
   );
   gpc1_1 gpc8473 (
      {stage2_55[101]},
      {stage3_55[62]}
   );
   gpc1_1 gpc8474 (
      {stage2_55[102]},
      {stage3_55[63]}
   );
   gpc1_1 gpc8475 (
      {stage2_55[103]},
      {stage3_55[64]}
   );
   gpc1_1 gpc8476 (
      {stage2_55[104]},
      {stage3_55[65]}
   );
   gpc1_1 gpc8477 (
      {stage2_55[105]},
      {stage3_55[66]}
   );
   gpc1_1 gpc8478 (
      {stage2_57[49]},
      {stage3_57[37]}
   );
   gpc1_1 gpc8479 (
      {stage2_57[50]},
      {stage3_57[38]}
   );
   gpc1_1 gpc8480 (
      {stage2_57[51]},
      {stage3_57[39]}
   );
   gpc1_1 gpc8481 (
      {stage2_57[52]},
      {stage3_57[40]}
   );
   gpc1_1 gpc8482 (
      {stage2_57[53]},
      {stage3_57[41]}
   );
   gpc1_1 gpc8483 (
      {stage2_57[54]},
      {stage3_57[42]}
   );
   gpc1_1 gpc8484 (
      {stage2_57[55]},
      {stage3_57[43]}
   );
   gpc1_1 gpc8485 (
      {stage2_57[56]},
      {stage3_57[44]}
   );
   gpc1_1 gpc8486 (
      {stage2_57[57]},
      {stage3_57[45]}
   );
   gpc1_1 gpc8487 (
      {stage2_57[58]},
      {stage3_57[46]}
   );
   gpc1_1 gpc8488 (
      {stage2_57[59]},
      {stage3_57[47]}
   );
   gpc1_1 gpc8489 (
      {stage2_57[60]},
      {stage3_57[48]}
   );
   gpc1_1 gpc8490 (
      {stage2_57[61]},
      {stage3_57[49]}
   );
   gpc1_1 gpc8491 (
      {stage2_57[62]},
      {stage3_57[50]}
   );
   gpc1_1 gpc8492 (
      {stage2_57[63]},
      {stage3_57[51]}
   );
   gpc1_1 gpc8493 (
      {stage2_57[64]},
      {stage3_57[52]}
   );
   gpc1_1 gpc8494 (
      {stage2_57[65]},
      {stage3_57[53]}
   );
   gpc1_1 gpc8495 (
      {stage2_58[58]},
      {stage3_58[34]}
   );
   gpc1_1 gpc8496 (
      {stage2_58[59]},
      {stage3_58[35]}
   );
   gpc1_1 gpc8497 (
      {stage2_58[60]},
      {stage3_58[36]}
   );
   gpc1_1 gpc8498 (
      {stage2_58[61]},
      {stage3_58[37]}
   );
   gpc1_1 gpc8499 (
      {stage2_58[62]},
      {stage3_58[38]}
   );
   gpc1_1 gpc8500 (
      {stage2_58[63]},
      {stage3_58[39]}
   );
   gpc1_1 gpc8501 (
      {stage2_58[64]},
      {stage3_58[40]}
   );
   gpc1_1 gpc8502 (
      {stage2_58[65]},
      {stage3_58[41]}
   );
   gpc1_1 gpc8503 (
      {stage2_58[66]},
      {stage3_58[42]}
   );
   gpc1_1 gpc8504 (
      {stage2_58[67]},
      {stage3_58[43]}
   );
   gpc1_1 gpc8505 (
      {stage2_58[68]},
      {stage3_58[44]}
   );
   gpc1_1 gpc8506 (
      {stage2_58[69]},
      {stage3_58[45]}
   );
   gpc1_1 gpc8507 (
      {stage2_58[70]},
      {stage3_58[46]}
   );
   gpc1_1 gpc8508 (
      {stage2_58[71]},
      {stage3_58[47]}
   );
   gpc1_1 gpc8509 (
      {stage2_58[72]},
      {stage3_58[48]}
   );
   gpc1_1 gpc8510 (
      {stage2_58[73]},
      {stage3_58[49]}
   );
   gpc1_1 gpc8511 (
      {stage2_58[74]},
      {stage3_58[50]}
   );
   gpc1_1 gpc8512 (
      {stage2_58[75]},
      {stage3_58[51]}
   );
   gpc1_1 gpc8513 (
      {stage2_58[76]},
      {stage3_58[52]}
   );
   gpc1_1 gpc8514 (
      {stage2_58[77]},
      {stage3_58[53]}
   );
   gpc1_1 gpc8515 (
      {stage2_58[78]},
      {stage3_58[54]}
   );
   gpc1_1 gpc8516 (
      {stage2_58[79]},
      {stage3_58[55]}
   );
   gpc1_1 gpc8517 (
      {stage2_58[80]},
      {stage3_58[56]}
   );
   gpc1_1 gpc8518 (
      {stage2_58[81]},
      {stage3_58[57]}
   );
   gpc1_1 gpc8519 (
      {stage2_58[82]},
      {stage3_58[58]}
   );
   gpc1_1 gpc8520 (
      {stage2_58[83]},
      {stage3_58[59]}
   );
   gpc1_1 gpc8521 (
      {stage2_58[84]},
      {stage3_58[60]}
   );
   gpc1_1 gpc8522 (
      {stage2_58[85]},
      {stage3_58[61]}
   );
   gpc1_1 gpc8523 (
      {stage2_59[85]},
      {stage3_59[25]}
   );
   gpc1_1 gpc8524 (
      {stage2_59[86]},
      {stage3_59[26]}
   );
   gpc1_1 gpc8525 (
      {stage2_59[87]},
      {stage3_59[27]}
   );
   gpc1_1 gpc8526 (
      {stage2_59[88]},
      {stage3_59[28]}
   );
   gpc1_1 gpc8527 (
      {stage2_59[89]},
      {stage3_59[29]}
   );
   gpc1_1 gpc8528 (
      {stage2_59[90]},
      {stage3_59[30]}
   );
   gpc1_1 gpc8529 (
      {stage2_59[91]},
      {stage3_59[31]}
   );
   gpc1_1 gpc8530 (
      {stage2_59[92]},
      {stage3_59[32]}
   );
   gpc1_1 gpc8531 (
      {stage2_59[93]},
      {stage3_59[33]}
   );
   gpc1_1 gpc8532 (
      {stage2_59[94]},
      {stage3_59[34]}
   );
   gpc1_1 gpc8533 (
      {stage2_59[95]},
      {stage3_59[35]}
   );
   gpc1_1 gpc8534 (
      {stage2_59[96]},
      {stage3_59[36]}
   );
   gpc1_1 gpc8535 (
      {stage2_59[97]},
      {stage3_59[37]}
   );
   gpc1_1 gpc8536 (
      {stage2_59[98]},
      {stage3_59[38]}
   );
   gpc1_1 gpc8537 (
      {stage2_59[99]},
      {stage3_59[39]}
   );
   gpc1_1 gpc8538 (
      {stage2_59[100]},
      {stage3_59[40]}
   );
   gpc1_1 gpc8539 (
      {stage2_59[101]},
      {stage3_59[41]}
   );
   gpc1_1 gpc8540 (
      {stage2_59[102]},
      {stage3_59[42]}
   );
   gpc1_1 gpc8541 (
      {stage2_59[103]},
      {stage3_59[43]}
   );
   gpc1_1 gpc8542 (
      {stage2_59[104]},
      {stage3_59[44]}
   );
   gpc1_1 gpc8543 (
      {stage2_59[105]},
      {stage3_59[45]}
   );
   gpc1_1 gpc8544 (
      {stage2_59[106]},
      {stage3_59[46]}
   );
   gpc1_1 gpc8545 (
      {stage2_59[107]},
      {stage3_59[47]}
   );
   gpc1_1 gpc8546 (
      {stage2_59[108]},
      {stage3_59[48]}
   );
   gpc1_1 gpc8547 (
      {stage2_59[109]},
      {stage3_59[49]}
   );
   gpc1_1 gpc8548 (
      {stage2_60[73]},
      {stage3_60[30]}
   );
   gpc1_1 gpc8549 (
      {stage2_60[74]},
      {stage3_60[31]}
   );
   gpc1_1 gpc8550 (
      {stage2_60[75]},
      {stage3_60[32]}
   );
   gpc1_1 gpc8551 (
      {stage2_60[76]},
      {stage3_60[33]}
   );
   gpc1_1 gpc8552 (
      {stage2_60[77]},
      {stage3_60[34]}
   );
   gpc1_1 gpc8553 (
      {stage2_60[78]},
      {stage3_60[35]}
   );
   gpc1_1 gpc8554 (
      {stage2_60[79]},
      {stage3_60[36]}
   );
   gpc1_1 gpc8555 (
      {stage2_60[80]},
      {stage3_60[37]}
   );
   gpc1_1 gpc8556 (
      {stage2_60[81]},
      {stage3_60[38]}
   );
   gpc1_1 gpc8557 (
      {stage2_60[82]},
      {stage3_60[39]}
   );
   gpc1_1 gpc8558 (
      {stage2_60[83]},
      {stage3_60[40]}
   );
   gpc1_1 gpc8559 (
      {stage2_60[84]},
      {stage3_60[41]}
   );
   gpc1_1 gpc8560 (
      {stage2_61[48]},
      {stage3_61[26]}
   );
   gpc1_1 gpc8561 (
      {stage2_61[49]},
      {stage3_61[27]}
   );
   gpc1_1 gpc8562 (
      {stage2_61[50]},
      {stage3_61[28]}
   );
   gpc1_1 gpc8563 (
      {stage2_61[51]},
      {stage3_61[29]}
   );
   gpc1_1 gpc8564 (
      {stage2_61[52]},
      {stage3_61[30]}
   );
   gpc1_1 gpc8565 (
      {stage2_61[53]},
      {stage3_61[31]}
   );
   gpc1_1 gpc8566 (
      {stage2_61[54]},
      {stage3_61[32]}
   );
   gpc1_1 gpc8567 (
      {stage2_61[55]},
      {stage3_61[33]}
   );
   gpc1_1 gpc8568 (
      {stage2_61[56]},
      {stage3_61[34]}
   );
   gpc1_1 gpc8569 (
      {stage2_61[57]},
      {stage3_61[35]}
   );
   gpc1_1 gpc8570 (
      {stage2_61[58]},
      {stage3_61[36]}
   );
   gpc1_1 gpc8571 (
      {stage2_61[59]},
      {stage3_61[37]}
   );
   gpc1_1 gpc8572 (
      {stage2_61[60]},
      {stage3_61[38]}
   );
   gpc1_1 gpc8573 (
      {stage2_61[61]},
      {stage3_61[39]}
   );
   gpc1_1 gpc8574 (
      {stage2_61[62]},
      {stage3_61[40]}
   );
   gpc1_1 gpc8575 (
      {stage2_61[63]},
      {stage3_61[41]}
   );
   gpc1_1 gpc8576 (
      {stage2_61[64]},
      {stage3_61[42]}
   );
   gpc1_1 gpc8577 (
      {stage2_61[65]},
      {stage3_61[43]}
   );
   gpc1_1 gpc8578 (
      {stage2_61[66]},
      {stage3_61[44]}
   );
   gpc1_1 gpc8579 (
      {stage2_61[67]},
      {stage3_61[45]}
   );
   gpc1_1 gpc8580 (
      {stage2_61[68]},
      {stage3_61[46]}
   );
   gpc1_1 gpc8581 (
      {stage2_61[69]},
      {stage3_61[47]}
   );
   gpc1_1 gpc8582 (
      {stage2_61[70]},
      {stage3_61[48]}
   );
   gpc1_1 gpc8583 (
      {stage2_61[71]},
      {stage3_61[49]}
   );
   gpc1_1 gpc8584 (
      {stage2_61[72]},
      {stage3_61[50]}
   );
   gpc1_1 gpc8585 (
      {stage2_61[73]},
      {stage3_61[51]}
   );
   gpc1_1 gpc8586 (
      {stage2_61[74]},
      {stage3_61[52]}
   );
   gpc1_1 gpc8587 (
      {stage2_63[90]},
      {stage3_63[39]}
   );
   gpc1_1 gpc8588 (
      {stage2_63[91]},
      {stage3_63[40]}
   );
   gpc1_1 gpc8589 (
      {stage2_63[92]},
      {stage3_63[41]}
   );
   gpc1_1 gpc8590 (
      {stage2_63[93]},
      {stage3_63[42]}
   );
   gpc1_1 gpc8591 (
      {stage2_63[94]},
      {stage3_63[43]}
   );
   gpc1_1 gpc8592 (
      {stage2_63[95]},
      {stage3_63[44]}
   );
   gpc1_1 gpc8593 (
      {stage2_63[96]},
      {stage3_63[45]}
   );
   gpc1_1 gpc8594 (
      {stage2_63[97]},
      {stage3_63[46]}
   );
   gpc1_1 gpc8595 (
      {stage2_63[98]},
      {stage3_63[47]}
   );
   gpc1_1 gpc8596 (
      {stage2_64[129]},
      {stage3_64[38]}
   );
   gpc1_1 gpc8597 (
      {stage2_64[130]},
      {stage3_64[39]}
   );
   gpc1_1 gpc8598 (
      {stage2_64[131]},
      {stage3_64[40]}
   );
   gpc1_1 gpc8599 (
      {stage2_64[132]},
      {stage3_64[41]}
   );
   gpc1_1 gpc8600 (
      {stage2_64[133]},
      {stage3_64[42]}
   );
   gpc1_1 gpc8601 (
      {stage2_64[134]},
      {stage3_64[43]}
   );
   gpc1_1 gpc8602 (
      {stage2_64[135]},
      {stage3_64[44]}
   );
   gpc1_1 gpc8603 (
      {stage2_64[136]},
      {stage3_64[45]}
   );
   gpc1_1 gpc8604 (
      {stage2_64[137]},
      {stage3_64[46]}
   );
   gpc1_1 gpc8605 (
      {stage2_64[138]},
      {stage3_64[47]}
   );
   gpc1_1 gpc8606 (
      {stage2_64[139]},
      {stage3_64[48]}
   );
   gpc1_1 gpc8607 (
      {stage2_64[140]},
      {stage3_64[49]}
   );
   gpc1_1 gpc8608 (
      {stage2_64[141]},
      {stage3_64[50]}
   );
   gpc1_1 gpc8609 (
      {stage2_65[51]},
      {stage3_65[33]}
   );
   gpc1_1 gpc8610 (
      {stage2_65[52]},
      {stage3_65[34]}
   );
   gpc1_1 gpc8611 (
      {stage2_65[53]},
      {stage3_65[35]}
   );
   gpc1_1 gpc8612 (
      {stage2_65[54]},
      {stage3_65[36]}
   );
   gpc1_1 gpc8613 (
      {stage2_65[55]},
      {stage3_65[37]}
   );
   gpc1_1 gpc8614 (
      {stage2_66[36]},
      {stage3_66[32]}
   );
   gpc1_1 gpc8615 (
      {stage2_66[37]},
      {stage3_66[33]}
   );
   gpc1_1 gpc8616 (
      {stage2_66[38]},
      {stage3_66[34]}
   );
   gpc1_1 gpc8617 (
      {stage2_66[39]},
      {stage3_66[35]}
   );
   gpc1_1 gpc8618 (
      {stage2_66[40]},
      {stage3_66[36]}
   );
   gpc1_1 gpc8619 (
      {stage2_66[41]},
      {stage3_66[37]}
   );
   gpc615_5 gpc8620 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4]},
      {stage3_1[0]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc615_5 gpc8621 (
      {stage3_0[5], stage3_0[6], stage3_0[7], stage3_0[8], stage3_0[9]},
      {stage3_1[1]},
      {stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9], stage3_2[10], stage3_2[11]},
      {stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1],stage4_0[1]}
   );
   gpc615_5 gpc8622 (
      {stage3_0[10], stage3_0[11], stage3_0[12], stage3_0[13], stage3_0[14]},
      {stage3_1[2]},
      {stage3_2[12], stage3_2[13], stage3_2[14], stage3_2[15], stage3_2[16], stage3_2[17]},
      {stage4_4[2],stage4_3[2],stage4_2[2],stage4_1[2],stage4_0[2]}
   );
   gpc606_5 gpc8623 (
      {stage3_1[3], stage3_1[4], stage3_1[5], stage3_1[6], stage3_1[7], stage3_1[8]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[3],stage4_3[3],stage4_2[3],stage4_1[3]}
   );
   gpc606_5 gpc8624 (
      {stage3_1[9], stage3_1[10], stage3_1[11], stage3_1[12], stage3_1[13], stage3_1[14]},
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage4_5[1],stage4_4[4],stage4_3[4],stage4_2[4],stage4_1[4]}
   );
   gpc606_5 gpc8625 (
      {stage3_1[15], stage3_1[16], stage3_1[17], stage3_1[18], stage3_1[19], stage3_1[20]},
      {stage3_3[12], stage3_3[13], stage3_3[14], stage3_3[15], stage3_3[16], stage3_3[17]},
      {stage4_5[2],stage4_4[5],stage4_3[5],stage4_2[5],stage4_1[5]}
   );
   gpc606_5 gpc8626 (
      {stage3_2[18], stage3_2[19], stage3_2[20], stage3_2[21], stage3_2[22], stage3_2[23]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[3],stage4_4[6],stage4_3[6],stage4_2[6]}
   );
   gpc606_5 gpc8627 (
      {stage3_2[24], stage3_2[25], stage3_2[26], stage3_2[27], stage3_2[28], stage3_2[29]},
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage4_6[1],stage4_5[4],stage4_4[7],stage4_3[7],stage4_2[7]}
   );
   gpc606_5 gpc8628 (
      {stage3_2[30], stage3_2[31], stage3_2[32], stage3_2[33], stage3_2[34], stage3_2[35]},
      {stage3_4[12], stage3_4[13], stage3_4[14], stage3_4[15], stage3_4[16], stage3_4[17]},
      {stage4_6[2],stage4_5[5],stage4_4[8],stage4_3[8],stage4_2[8]}
   );
   gpc606_5 gpc8629 (
      {stage3_2[36], stage3_2[37], stage3_2[38], stage3_2[39], stage3_2[40], stage3_2[41]},
      {stage3_4[18], stage3_4[19], stage3_4[20], stage3_4[21], stage3_4[22], stage3_4[23]},
      {stage4_6[3],stage4_5[6],stage4_4[9],stage4_3[9],stage4_2[9]}
   );
   gpc615_5 gpc8630 (
      {stage3_3[18], stage3_3[19], stage3_3[20], stage3_3[21], stage3_3[22]},
      {stage3_4[24]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[4],stage4_5[7],stage4_4[10],stage4_3[10]}
   );
   gpc1163_5 gpc8631 (
      {stage3_4[25], stage3_4[26], stage3_4[27]},
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage3_6[0]},
      {stage3_7[0]},
      {stage4_8[0],stage4_7[1],stage4_6[5],stage4_5[8],stage4_4[11]}
   );
   gpc1163_5 gpc8632 (
      {stage3_4[28], stage3_4[29], stage3_4[30]},
      {stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17]},
      {stage3_6[1]},
      {stage3_7[1]},
      {stage4_8[1],stage4_7[2],stage4_6[6],stage4_5[9],stage4_4[12]}
   );
   gpc1163_5 gpc8633 (
      {stage3_4[31], stage3_4[32], stage3_4[33]},
      {stage3_5[18], stage3_5[19], stage3_5[20], stage3_5[21], stage3_5[22], stage3_5[23]},
      {stage3_6[2]},
      {stage3_7[2]},
      {stage4_8[2],stage4_7[3],stage4_6[7],stage4_5[10],stage4_4[13]}
   );
   gpc1163_5 gpc8634 (
      {stage3_4[34], stage3_4[35], stage3_4[36]},
      {stage3_5[24], stage3_5[25], stage3_5[26], stage3_5[27], stage3_5[28], stage3_5[29]},
      {stage3_6[3]},
      {stage3_7[3]},
      {stage4_8[3],stage4_7[4],stage4_6[8],stage4_5[11],stage4_4[14]}
   );
   gpc1163_5 gpc8635 (
      {stage3_4[37], stage3_4[38], stage3_4[39]},
      {stage3_5[30], stage3_5[31], stage3_5[32], stage3_5[33], stage3_5[34], stage3_5[35]},
      {stage3_6[4]},
      {stage3_7[4]},
      {stage4_8[4],stage4_7[5],stage4_6[9],stage4_5[12],stage4_4[15]}
   );
   gpc1163_5 gpc8636 (
      {stage3_4[40], stage3_4[41], stage3_4[42]},
      {stage3_5[36], stage3_5[37], stage3_5[38], stage3_5[39], stage3_5[40], stage3_5[41]},
      {stage3_6[5]},
      {stage3_7[5]},
      {stage4_8[5],stage4_7[6],stage4_6[10],stage4_5[13],stage4_4[16]}
   );
   gpc606_5 gpc8637 (
      {stage3_4[43], stage3_4[44], stage3_4[45], stage3_4[46], stage3_4[47], stage3_4[48]},
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10], stage3_6[11]},
      {stage4_8[6],stage4_7[7],stage4_6[11],stage4_5[14],stage4_4[17]}
   );
   gpc606_5 gpc8638 (
      {stage3_4[49], stage3_4[50], stage3_4[51], stage3_4[52], stage3_4[53], stage3_4[54]},
      {stage3_6[12], stage3_6[13], stage3_6[14], stage3_6[15], stage3_6[16], stage3_6[17]},
      {stage4_8[7],stage4_7[8],stage4_6[12],stage4_5[15],stage4_4[18]}
   );
   gpc606_5 gpc8639 (
      {stage3_4[55], stage3_4[56], stage3_4[57], stage3_4[58], stage3_4[59], stage3_4[60]},
      {stage3_6[18], stage3_6[19], stage3_6[20], stage3_6[21], stage3_6[22], stage3_6[23]},
      {stage4_8[8],stage4_7[9],stage4_6[13],stage4_5[16],stage4_4[19]}
   );
   gpc606_5 gpc8640 (
      {stage3_4[61], stage3_4[62], stage3_4[63], stage3_4[64], stage3_4[65], stage3_4[66]},
      {stage3_6[24], stage3_6[25], stage3_6[26], stage3_6[27], stage3_6[28], stage3_6[29]},
      {stage4_8[9],stage4_7[10],stage4_6[14],stage4_5[17],stage4_4[20]}
   );
   gpc606_5 gpc8641 (
      {stage3_4[67], stage3_4[68], stage3_4[69], stage3_4[70], stage3_4[71], stage3_4[72]},
      {stage3_6[30], stage3_6[31], stage3_6[32], stage3_6[33], stage3_6[34], stage3_6[35]},
      {stage4_8[10],stage4_7[11],stage4_6[15],stage4_5[18],stage4_4[21]}
   );
   gpc606_5 gpc8642 (
      {stage3_4[73], stage3_4[74], stage3_4[75], stage3_4[76], stage3_4[77], stage3_4[78]},
      {stage3_6[36], stage3_6[37], stage3_6[38], stage3_6[39], stage3_6[40], stage3_6[41]},
      {stage4_8[11],stage4_7[12],stage4_6[16],stage4_5[19],stage4_4[22]}
   );
   gpc606_5 gpc8643 (
      {stage3_4[79], stage3_4[80], stage3_4[81], stage3_4[82], stage3_4[83], stage3_4[84]},
      {stage3_6[42], stage3_6[43], stage3_6[44], stage3_6[45], stage3_6[46], stage3_6[47]},
      {stage4_8[12],stage4_7[13],stage4_6[17],stage4_5[20],stage4_4[23]}
   );
   gpc606_5 gpc8644 (
      {stage3_4[85], stage3_4[86], stage3_4[87], stage3_4[88], stage3_4[89], stage3_4[90]},
      {stage3_6[48], stage3_6[49], stage3_6[50], stage3_6[51], stage3_6[52], stage3_6[53]},
      {stage4_8[13],stage4_7[14],stage4_6[18],stage4_5[21],stage4_4[24]}
   );
   gpc606_5 gpc8645 (
      {stage3_4[91], stage3_4[92], stage3_4[93], stage3_4[94], stage3_4[95], stage3_4[96]},
      {stage3_6[54], stage3_6[55], stage3_6[56], stage3_6[57], stage3_6[58], stage3_6[59]},
      {stage4_8[14],stage4_7[15],stage4_6[19],stage4_5[22],stage4_4[25]}
   );
   gpc606_5 gpc8646 (
      {stage3_4[97], stage3_4[98], stage3_4[99], stage3_4[100], stage3_4[101], stage3_4[102]},
      {stage3_6[60], stage3_6[61], stage3_6[62], stage3_6[63], stage3_6[64], stage3_6[65]},
      {stage4_8[15],stage4_7[16],stage4_6[20],stage4_5[23],stage4_4[26]}
   );
   gpc606_5 gpc8647 (
      {stage3_4[103], stage3_4[104], stage3_4[105], stage3_4[106], stage3_4[107], stage3_4[108]},
      {stage3_6[66], stage3_6[67], stage3_6[68], stage3_6[69], stage3_6[70], stage3_6[71]},
      {stage4_8[16],stage4_7[17],stage4_6[21],stage4_5[24],stage4_4[27]}
   );
   gpc615_5 gpc8648 (
      {stage3_6[72], stage3_6[73], stage3_6[74], stage3_6[75], stage3_6[76]},
      {stage3_7[6]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[17],stage4_7[18],stage4_6[22]}
   );
   gpc615_5 gpc8649 (
      {stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage3_8[6]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[1],stage4_9[1],stage4_8[18],stage4_7[19]}
   );
   gpc615_5 gpc8650 (
      {stage3_7[12], stage3_7[13], stage3_7[14], stage3_7[15], stage3_7[16]},
      {stage3_8[7]},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage4_11[1],stage4_10[2],stage4_9[2],stage4_8[19],stage4_7[20]}
   );
   gpc615_5 gpc8651 (
      {stage3_7[17], stage3_7[18], stage3_7[19], stage3_7[20], stage3_7[21]},
      {stage3_8[8]},
      {stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15], stage3_9[16], stage3_9[17]},
      {stage4_11[2],stage4_10[3],stage4_9[3],stage4_8[20],stage4_7[21]}
   );
   gpc615_5 gpc8652 (
      {stage3_7[22], stage3_7[23], stage3_7[24], stage3_7[25], stage3_7[26]},
      {stage3_8[9]},
      {stage3_9[18], stage3_9[19], stage3_9[20], stage3_9[21], stage3_9[22], stage3_9[23]},
      {stage4_11[3],stage4_10[4],stage4_9[4],stage4_8[21],stage4_7[22]}
   );
   gpc615_5 gpc8653 (
      {stage3_7[27], stage3_7[28], stage3_7[29], stage3_7[30], stage3_7[31]},
      {stage3_8[10]},
      {stage3_9[24], stage3_9[25], stage3_9[26], stage3_9[27], stage3_9[28], stage3_9[29]},
      {stage4_11[4],stage4_10[5],stage4_9[5],stage4_8[22],stage4_7[23]}
   );
   gpc615_5 gpc8654 (
      {stage3_7[32], stage3_7[33], stage3_7[34], stage3_7[35], stage3_7[36]},
      {stage3_8[11]},
      {stage3_9[30], stage3_9[31], stage3_9[32], stage3_9[33], stage3_9[34], stage3_9[35]},
      {stage4_11[5],stage4_10[6],stage4_9[6],stage4_8[23],stage4_7[24]}
   );
   gpc606_5 gpc8655 (
      {stage3_8[12], stage3_8[13], stage3_8[14], stage3_8[15], stage3_8[16], stage3_8[17]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage4_12[0],stage4_11[6],stage4_10[7],stage4_9[7],stage4_8[24]}
   );
   gpc606_5 gpc8656 (
      {stage3_8[18], stage3_8[19], stage3_8[20], stage3_8[21], stage3_8[22], stage3_8[23]},
      {stage3_10[6], stage3_10[7], stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11]},
      {stage4_12[1],stage4_11[7],stage4_10[8],stage4_9[8],stage4_8[25]}
   );
   gpc606_5 gpc8657 (
      {stage3_8[24], stage3_8[25], stage3_8[26], stage3_8[27], stage3_8[28], stage3_8[29]},
      {stage3_10[12], stage3_10[13], stage3_10[14], stage3_10[15], stage3_10[16], stage3_10[17]},
      {stage4_12[2],stage4_11[8],stage4_10[9],stage4_9[9],stage4_8[26]}
   );
   gpc606_5 gpc8658 (
      {stage3_8[30], stage3_8[31], stage3_8[32], stage3_8[33], stage3_8[34], 1'b0},
      {stage3_10[18], stage3_10[19], stage3_10[20], stage3_10[21], stage3_10[22], stage3_10[23]},
      {stage4_12[3],stage4_11[9],stage4_10[10],stage4_9[10],stage4_8[27]}
   );
   gpc606_5 gpc8659 (
      {stage3_9[36], stage3_9[37], stage3_9[38], stage3_9[39], stage3_9[40], stage3_9[41]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[4],stage4_11[10],stage4_10[11],stage4_9[11]}
   );
   gpc606_5 gpc8660 (
      {stage3_9[42], stage3_9[43], stage3_9[44], stage3_9[45], stage3_9[46], stage3_9[47]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[5],stage4_11[11],stage4_10[12],stage4_9[12]}
   );
   gpc606_5 gpc8661 (
      {stage3_9[48], stage3_9[49], stage3_9[50], stage3_9[51], stage3_9[52], stage3_9[53]},
      {stage3_11[12], stage3_11[13], stage3_11[14], stage3_11[15], stage3_11[16], stage3_11[17]},
      {stage4_13[2],stage4_12[6],stage4_11[12],stage4_10[13],stage4_9[13]}
   );
   gpc615_5 gpc8662 (
      {stage3_10[24], stage3_10[25], stage3_10[26], stage3_10[27], stage3_10[28]},
      {stage3_11[18]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[3],stage4_12[7],stage4_11[13],stage4_10[14]}
   );
   gpc615_5 gpc8663 (
      {stage3_10[29], stage3_10[30], stage3_10[31], stage3_10[32], stage3_10[33]},
      {stage3_11[19]},
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage4_14[1],stage4_13[4],stage4_12[8],stage4_11[14],stage4_10[15]}
   );
   gpc615_5 gpc8664 (
      {stage3_10[34], stage3_10[35], stage3_10[36], stage3_10[37], stage3_10[38]},
      {stage3_11[20]},
      {stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15], stage3_12[16], stage3_12[17]},
      {stage4_14[2],stage4_13[5],stage4_12[9],stage4_11[15],stage4_10[16]}
   );
   gpc615_5 gpc8665 (
      {stage3_10[39], stage3_10[40], stage3_10[41], stage3_10[42], stage3_10[43]},
      {stage3_11[21]},
      {stage3_12[18], stage3_12[19], stage3_12[20], stage3_12[21], stage3_12[22], stage3_12[23]},
      {stage4_14[3],stage4_13[6],stage4_12[10],stage4_11[16],stage4_10[17]}
   );
   gpc615_5 gpc8666 (
      {stage3_10[44], stage3_10[45], stage3_10[46], stage3_10[47], stage3_10[48]},
      {stage3_11[22]},
      {stage3_12[24], stage3_12[25], stage3_12[26], stage3_12[27], stage3_12[28], stage3_12[29]},
      {stage4_14[4],stage4_13[7],stage4_12[11],stage4_11[17],stage4_10[18]}
   );
   gpc615_5 gpc8667 (
      {stage3_10[49], stage3_10[50], stage3_10[51], stage3_10[52], stage3_10[53]},
      {stage3_11[23]},
      {stage3_12[30], stage3_12[31], stage3_12[32], stage3_12[33], stage3_12[34], stage3_12[35]},
      {stage4_14[5],stage4_13[8],stage4_12[12],stage4_11[18],stage4_10[19]}
   );
   gpc615_5 gpc8668 (
      {stage3_10[54], stage3_10[55], stage3_10[56], stage3_10[57], stage3_10[58]},
      {stage3_11[24]},
      {stage3_12[36], stage3_12[37], stage3_12[38], stage3_12[39], stage3_12[40], stage3_12[41]},
      {stage4_14[6],stage4_13[9],stage4_12[13],stage4_11[19],stage4_10[20]}
   );
   gpc615_5 gpc8669 (
      {stage3_10[59], stage3_10[60], stage3_10[61], stage3_10[62], stage3_10[63]},
      {stage3_11[25]},
      {stage3_12[42], stage3_12[43], stage3_12[44], stage3_12[45], stage3_12[46], stage3_12[47]},
      {stage4_14[7],stage4_13[10],stage4_12[14],stage4_11[20],stage4_10[21]}
   );
   gpc615_5 gpc8670 (
      {stage3_10[64], stage3_10[65], stage3_10[66], stage3_10[67], stage3_10[68]},
      {stage3_11[26]},
      {stage3_12[48], stage3_12[49], stage3_12[50], stage3_12[51], stage3_12[52], stage3_12[53]},
      {stage4_14[8],stage4_13[11],stage4_12[15],stage4_11[21],stage4_10[22]}
   );
   gpc615_5 gpc8671 (
      {stage3_10[69], stage3_10[70], stage3_10[71], stage3_10[72], stage3_10[73]},
      {stage3_11[27]},
      {stage3_12[54], stage3_12[55], stage3_12[56], stage3_12[57], stage3_12[58], stage3_12[59]},
      {stage4_14[9],stage4_13[12],stage4_12[16],stage4_11[22],stage4_10[23]}
   );
   gpc1325_5 gpc8672 (
      {stage3_10[74], stage3_10[75], stage3_10[76], stage3_10[77], stage3_10[78]},
      {stage3_11[28], stage3_11[29]},
      {stage3_12[60], stage3_12[61], stage3_12[62]},
      {stage3_13[0]},
      {stage4_14[10],stage4_13[13],stage4_12[17],stage4_11[23],stage4_10[24]}
   );
   gpc1325_5 gpc8673 (
      {stage3_10[79], stage3_10[80], stage3_10[81], stage3_10[82], stage3_10[83]},
      {stage3_11[30], stage3_11[31]},
      {stage3_12[63], stage3_12[64], stage3_12[65]},
      {stage3_13[1]},
      {stage4_14[11],stage4_13[14],stage4_12[18],stage4_11[24],stage4_10[25]}
   );
   gpc207_4 gpc8674 (
      {stage3_11[32], stage3_11[33], stage3_11[34], stage3_11[35], stage3_11[36], stage3_11[37], stage3_11[38]},
      {stage3_13[2], stage3_13[3]},
      {stage4_14[12],stage4_13[15],stage4_12[19],stage4_11[25]}
   );
   gpc207_4 gpc8675 (
      {stage3_11[39], stage3_11[40], stage3_11[41], stage3_11[42], stage3_11[43], stage3_11[44], stage3_11[45]},
      {stage3_13[4], stage3_13[5]},
      {stage4_14[13],stage4_13[16],stage4_12[20],stage4_11[26]}
   );
   gpc207_4 gpc8676 (
      {stage3_11[46], stage3_11[47], stage3_11[48], stage3_11[49], stage3_11[50], stage3_11[51], stage3_11[52]},
      {stage3_13[6], stage3_13[7]},
      {stage4_14[14],stage4_13[17],stage4_12[21],stage4_11[27]}
   );
   gpc615_5 gpc8677 (
      {stage3_11[53], stage3_11[54], stage3_11[55], stage3_11[56], stage3_11[57]},
      {stage3_12[66]},
      {stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11], stage3_13[12], stage3_13[13]},
      {stage4_15[0],stage4_14[15],stage4_13[18],stage4_12[22],stage4_11[28]}
   );
   gpc606_5 gpc8678 (
      {stage3_13[14], stage3_13[15], stage3_13[16], stage3_13[17], stage3_13[18], stage3_13[19]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[0],stage4_15[1],stage4_14[16],stage4_13[19]}
   );
   gpc606_5 gpc8679 (
      {stage3_13[20], stage3_13[21], stage3_13[22], stage3_13[23], stage3_13[24], stage3_13[25]},
      {stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11]},
      {stage4_17[1],stage4_16[1],stage4_15[2],stage4_14[17],stage4_13[20]}
   );
   gpc606_5 gpc8680 (
      {stage3_13[26], stage3_13[27], stage3_13[28], stage3_13[29], stage3_13[30], stage3_13[31]},
      {stage3_15[12], stage3_15[13], stage3_15[14], stage3_15[15], stage3_15[16], stage3_15[17]},
      {stage4_17[2],stage4_16[2],stage4_15[3],stage4_14[18],stage4_13[21]}
   );
   gpc606_5 gpc8681 (
      {stage3_13[32], stage3_13[33], stage3_13[34], stage3_13[35], stage3_13[36], stage3_13[37]},
      {stage3_15[18], stage3_15[19], stage3_15[20], stage3_15[21], stage3_15[22], stage3_15[23]},
      {stage4_17[3],stage4_16[3],stage4_15[4],stage4_14[19],stage4_13[22]}
   );
   gpc606_5 gpc8682 (
      {stage3_13[38], stage3_13[39], stage3_13[40], stage3_13[41], stage3_13[42], stage3_13[43]},
      {stage3_15[24], stage3_15[25], stage3_15[26], stage3_15[27], stage3_15[28], stage3_15[29]},
      {stage4_17[4],stage4_16[4],stage4_15[5],stage4_14[20],stage4_13[23]}
   );
   gpc606_5 gpc8683 (
      {stage3_13[44], stage3_13[45], stage3_13[46], stage3_13[47], stage3_13[48], stage3_13[49]},
      {stage3_15[30], stage3_15[31], stage3_15[32], stage3_15[33], stage3_15[34], stage3_15[35]},
      {stage4_17[5],stage4_16[5],stage4_15[6],stage4_14[21],stage4_13[24]}
   );
   gpc615_5 gpc8684 (
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4]},
      {stage3_15[36]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[6],stage4_16[6],stage4_15[7],stage4_14[22]}
   );
   gpc615_5 gpc8685 (
      {stage3_14[5], stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9]},
      {stage3_15[37]},
      {stage3_16[6], stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11]},
      {stage4_18[1],stage4_17[7],stage4_16[7],stage4_15[8],stage4_14[23]}
   );
   gpc615_5 gpc8686 (
      {stage3_14[10], stage3_14[11], stage3_14[12], stage3_14[13], stage3_14[14]},
      {stage3_15[38]},
      {stage3_16[12], stage3_16[13], stage3_16[14], stage3_16[15], stage3_16[16], stage3_16[17]},
      {stage4_18[2],stage4_17[8],stage4_16[8],stage4_15[9],stage4_14[24]}
   );
   gpc615_5 gpc8687 (
      {stage3_14[15], stage3_14[16], stage3_14[17], stage3_14[18], stage3_14[19]},
      {stage3_15[39]},
      {stage3_16[18], stage3_16[19], stage3_16[20], stage3_16[21], stage3_16[22], stage3_16[23]},
      {stage4_18[3],stage4_17[9],stage4_16[9],stage4_15[10],stage4_14[25]}
   );
   gpc615_5 gpc8688 (
      {stage3_14[20], stage3_14[21], stage3_14[22], stage3_14[23], stage3_14[24]},
      {stage3_15[40]},
      {stage3_16[24], stage3_16[25], stage3_16[26], stage3_16[27], stage3_16[28], stage3_16[29]},
      {stage4_18[4],stage4_17[10],stage4_16[10],stage4_15[11],stage4_14[26]}
   );
   gpc615_5 gpc8689 (
      {stage3_14[25], stage3_14[26], stage3_14[27], stage3_14[28], stage3_14[29]},
      {stage3_15[41]},
      {stage3_16[30], stage3_16[31], stage3_16[32], stage3_16[33], stage3_16[34], stage3_16[35]},
      {stage4_18[5],stage4_17[11],stage4_16[11],stage4_15[12],stage4_14[27]}
   );
   gpc615_5 gpc8690 (
      {stage3_15[42], stage3_15[43], stage3_15[44], stage3_15[45], stage3_15[46]},
      {stage3_16[36]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage4_19[0],stage4_18[6],stage4_17[12],stage4_16[12],stage4_15[13]}
   );
   gpc606_5 gpc8691 (
      {stage3_17[6], stage3_17[7], stage3_17[8], stage3_17[9], stage3_17[10], stage3_17[11]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[0],stage4_19[1],stage4_18[7],stage4_17[13]}
   );
   gpc606_5 gpc8692 (
      {stage3_17[12], stage3_17[13], stage3_17[14], stage3_17[15], stage3_17[16], stage3_17[17]},
      {stage3_19[6], stage3_19[7], stage3_19[8], stage3_19[9], stage3_19[10], stage3_19[11]},
      {stage4_21[1],stage4_20[1],stage4_19[2],stage4_18[8],stage4_17[14]}
   );
   gpc606_5 gpc8693 (
      {stage3_17[18], stage3_17[19], stage3_17[20], stage3_17[21], stage3_17[22], stage3_17[23]},
      {stage3_19[12], stage3_19[13], stage3_19[14], stage3_19[15], stage3_19[16], stage3_19[17]},
      {stage4_21[2],stage4_20[2],stage4_19[3],stage4_18[9],stage4_17[15]}
   );
   gpc606_5 gpc8694 (
      {stage3_17[24], stage3_17[25], stage3_17[26], stage3_17[27], stage3_17[28], stage3_17[29]},
      {stage3_19[18], stage3_19[19], stage3_19[20], stage3_19[21], stage3_19[22], stage3_19[23]},
      {stage4_21[3],stage4_20[3],stage4_19[4],stage4_18[10],stage4_17[16]}
   );
   gpc606_5 gpc8695 (
      {stage3_17[30], stage3_17[31], stage3_17[32], stage3_17[33], stage3_17[34], stage3_17[35]},
      {stage3_19[24], stage3_19[25], stage3_19[26], stage3_19[27], stage3_19[28], stage3_19[29]},
      {stage4_21[4],stage4_20[4],stage4_19[5],stage4_18[11],stage4_17[17]}
   );
   gpc207_4 gpc8696 (
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5], stage3_18[6]},
      {stage3_20[0], stage3_20[1]},
      {stage4_21[5],stage4_20[5],stage4_19[6],stage4_18[12]}
   );
   gpc207_4 gpc8697 (
      {stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11], stage3_18[12], stage3_18[13]},
      {stage3_20[2], stage3_20[3]},
      {stage4_21[6],stage4_20[6],stage4_19[7],stage4_18[13]}
   );
   gpc207_4 gpc8698 (
      {stage3_18[14], stage3_18[15], stage3_18[16], stage3_18[17], stage3_18[18], stage3_18[19], stage3_18[20]},
      {stage3_20[4], stage3_20[5]},
      {stage4_21[7],stage4_20[7],stage4_19[8],stage4_18[14]}
   );
   gpc207_4 gpc8699 (
      {stage3_18[21], stage3_18[22], stage3_18[23], stage3_18[24], stage3_18[25], stage3_18[26], stage3_18[27]},
      {stage3_20[6], stage3_20[7]},
      {stage4_21[8],stage4_20[8],stage4_19[9],stage4_18[15]}
   );
   gpc207_4 gpc8700 (
      {stage3_18[28], stage3_18[29], stage3_18[30], stage3_18[31], stage3_18[32], stage3_18[33], stage3_18[34]},
      {stage3_20[8], stage3_20[9]},
      {stage4_21[9],stage4_20[9],stage4_19[10],stage4_18[16]}
   );
   gpc207_4 gpc8701 (
      {stage3_18[35], stage3_18[36], stage3_18[37], stage3_18[38], stage3_18[39], stage3_18[40], stage3_18[41]},
      {stage3_20[10], stage3_20[11]},
      {stage4_21[10],stage4_20[10],stage4_19[11],stage4_18[17]}
   );
   gpc207_4 gpc8702 (
      {stage3_18[42], stage3_18[43], stage3_18[44], stage3_18[45], stage3_18[46], stage3_18[47], stage3_18[48]},
      {stage3_20[12], stage3_20[13]},
      {stage4_21[11],stage4_20[11],stage4_19[12],stage4_18[18]}
   );
   gpc207_4 gpc8703 (
      {stage3_18[49], stage3_18[50], stage3_18[51], stage3_18[52], stage3_18[53], stage3_18[54], stage3_18[55]},
      {stage3_20[14], stage3_20[15]},
      {stage4_21[12],stage4_20[12],stage4_19[13],stage4_18[19]}
   );
   gpc207_4 gpc8704 (
      {stage3_18[56], stage3_18[57], stage3_18[58], stage3_18[59], 1'b0, 1'b0, 1'b0},
      {stage3_20[16], stage3_20[17]},
      {stage4_21[13],stage4_20[13],stage4_19[14],stage4_18[20]}
   );
   gpc615_5 gpc8705 (
      {stage3_19[30], stage3_19[31], stage3_19[32], stage3_19[33], stage3_19[34]},
      {stage3_20[18]},
      {stage3_21[0], stage3_21[1], stage3_21[2], stage3_21[3], stage3_21[4], stage3_21[5]},
      {stage4_23[0],stage4_22[0],stage4_21[14],stage4_20[14],stage4_19[15]}
   );
   gpc606_5 gpc8706 (
      {stage3_20[19], stage3_20[20], stage3_20[21], stage3_20[22], stage3_20[23], stage3_20[24]},
      {stage3_22[0], stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5]},
      {stage4_24[0],stage4_23[1],stage4_22[1],stage4_21[15],stage4_20[15]}
   );
   gpc606_5 gpc8707 (
      {stage3_20[25], stage3_20[26], stage3_20[27], stage3_20[28], stage3_20[29], stage3_20[30]},
      {stage3_22[6], stage3_22[7], stage3_22[8], stage3_22[9], stage3_22[10], stage3_22[11]},
      {stage4_24[1],stage4_23[2],stage4_22[2],stage4_21[16],stage4_20[16]}
   );
   gpc606_5 gpc8708 (
      {stage3_20[31], stage3_20[32], stage3_20[33], stage3_20[34], stage3_20[35], stage3_20[36]},
      {stage3_22[12], stage3_22[13], stage3_22[14], stage3_22[15], stage3_22[16], stage3_22[17]},
      {stage4_24[2],stage4_23[3],stage4_22[3],stage4_21[17],stage4_20[17]}
   );
   gpc606_5 gpc8709 (
      {stage3_20[37], stage3_20[38], stage3_20[39], stage3_20[40], stage3_20[41], stage3_20[42]},
      {stage3_22[18], stage3_22[19], stage3_22[20], stage3_22[21], stage3_22[22], stage3_22[23]},
      {stage4_24[3],stage4_23[4],stage4_22[4],stage4_21[18],stage4_20[18]}
   );
   gpc606_5 gpc8710 (
      {stage3_20[43], stage3_20[44], stage3_20[45], stage3_20[46], stage3_20[47], stage3_20[48]},
      {stage3_22[24], stage3_22[25], stage3_22[26], stage3_22[27], stage3_22[28], stage3_22[29]},
      {stage4_24[4],stage4_23[5],stage4_22[5],stage4_21[19],stage4_20[19]}
   );
   gpc606_5 gpc8711 (
      {stage3_20[49], stage3_20[50], stage3_20[51], stage3_20[52], stage3_20[53], stage3_20[54]},
      {stage3_22[30], stage3_22[31], stage3_22[32], stage3_22[33], stage3_22[34], stage3_22[35]},
      {stage4_24[5],stage4_23[6],stage4_22[6],stage4_21[20],stage4_20[20]}
   );
   gpc606_5 gpc8712 (
      {stage3_20[55], stage3_20[56], stage3_20[57], stage3_20[58], stage3_20[59], stage3_20[60]},
      {stage3_22[36], stage3_22[37], stage3_22[38], stage3_22[39], stage3_22[40], stage3_22[41]},
      {stage4_24[6],stage4_23[7],stage4_22[7],stage4_21[21],stage4_20[21]}
   );
   gpc606_5 gpc8713 (
      {stage3_20[61], stage3_20[62], stage3_20[63], stage3_20[64], stage3_20[65], stage3_20[66]},
      {stage3_22[42], stage3_22[43], stage3_22[44], stage3_22[45], stage3_22[46], stage3_22[47]},
      {stage4_24[7],stage4_23[8],stage4_22[8],stage4_21[22],stage4_20[22]}
   );
   gpc606_5 gpc8714 (
      {stage3_20[67], stage3_20[68], stage3_20[69], stage3_20[70], stage3_20[71], stage3_20[72]},
      {stage3_22[48], stage3_22[49], stage3_22[50], stage3_22[51], stage3_22[52], stage3_22[53]},
      {stage4_24[8],stage4_23[9],stage4_22[9],stage4_21[23],stage4_20[23]}
   );
   gpc606_5 gpc8715 (
      {stage3_21[6], stage3_21[7], stage3_21[8], stage3_21[9], stage3_21[10], stage3_21[11]},
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5]},
      {stage4_25[0],stage4_24[9],stage4_23[10],stage4_22[10],stage4_21[24]}
   );
   gpc606_5 gpc8716 (
      {stage3_21[12], stage3_21[13], stage3_21[14], stage3_21[15], stage3_21[16], stage3_21[17]},
      {stage3_23[6], stage3_23[7], stage3_23[8], stage3_23[9], stage3_23[10], stage3_23[11]},
      {stage4_25[1],stage4_24[10],stage4_23[11],stage4_22[11],stage4_21[25]}
   );
   gpc606_5 gpc8717 (
      {stage3_21[18], stage3_21[19], stage3_21[20], stage3_21[21], stage3_21[22], stage3_21[23]},
      {stage3_23[12], stage3_23[13], stage3_23[14], stage3_23[15], stage3_23[16], stage3_23[17]},
      {stage4_25[2],stage4_24[11],stage4_23[12],stage4_22[12],stage4_21[26]}
   );
   gpc606_5 gpc8718 (
      {stage3_21[24], stage3_21[25], stage3_21[26], stage3_21[27], stage3_21[28], stage3_21[29]},
      {stage3_23[18], stage3_23[19], stage3_23[20], stage3_23[21], stage3_23[22], stage3_23[23]},
      {stage4_25[3],stage4_24[12],stage4_23[13],stage4_22[13],stage4_21[27]}
   );
   gpc615_5 gpc8719 (
      {stage3_22[54], stage3_22[55], stage3_22[56], stage3_22[57], stage3_22[58]},
      {stage3_23[24]},
      {stage3_24[0], stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5]},
      {stage4_26[0],stage4_25[4],stage4_24[13],stage4_23[14],stage4_22[14]}
   );
   gpc615_5 gpc8720 (
      {stage3_22[59], stage3_22[60], stage3_22[61], stage3_22[62], stage3_22[63]},
      {stage3_23[25]},
      {stage3_24[6], stage3_24[7], stage3_24[8], stage3_24[9], stage3_24[10], stage3_24[11]},
      {stage4_26[1],stage4_25[5],stage4_24[14],stage4_23[15],stage4_22[15]}
   );
   gpc615_5 gpc8721 (
      {stage3_22[64], stage3_22[65], stage3_22[66], stage3_22[67], stage3_22[68]},
      {stage3_23[26]},
      {stage3_24[12], stage3_24[13], stage3_24[14], stage3_24[15], stage3_24[16], stage3_24[17]},
      {stage4_26[2],stage4_25[6],stage4_24[15],stage4_23[16],stage4_22[16]}
   );
   gpc615_5 gpc8722 (
      {stage3_22[69], stage3_22[70], stage3_22[71], stage3_22[72], 1'b0},
      {stage3_23[27]},
      {stage3_24[18], stage3_24[19], stage3_24[20], stage3_24[21], stage3_24[22], stage3_24[23]},
      {stage4_26[3],stage4_25[7],stage4_24[16],stage4_23[17],stage4_22[17]}
   );
   gpc615_5 gpc8723 (
      {stage3_23[28], stage3_23[29], stage3_23[30], stage3_23[31], stage3_23[32]},
      {stage3_24[24]},
      {stage3_25[0], stage3_25[1], stage3_25[2], stage3_25[3], stage3_25[4], stage3_25[5]},
      {stage4_27[0],stage4_26[4],stage4_25[8],stage4_24[17],stage4_23[18]}
   );
   gpc615_5 gpc8724 (
      {stage3_23[33], stage3_23[34], stage3_23[35], stage3_23[36], stage3_23[37]},
      {stage3_24[25]},
      {stage3_25[6], stage3_25[7], stage3_25[8], stage3_25[9], stage3_25[10], stage3_25[11]},
      {stage4_27[1],stage4_26[5],stage4_25[9],stage4_24[18],stage4_23[19]}
   );
   gpc615_5 gpc8725 (
      {stage3_23[38], stage3_23[39], stage3_23[40], stage3_23[41], stage3_23[42]},
      {stage3_24[26]},
      {stage3_25[12], stage3_25[13], stage3_25[14], stage3_25[15], stage3_25[16], stage3_25[17]},
      {stage4_27[2],stage4_26[6],stage4_25[10],stage4_24[19],stage4_23[20]}
   );
   gpc606_5 gpc8726 (
      {stage3_25[18], stage3_25[19], stage3_25[20], stage3_25[21], stage3_25[22], stage3_25[23]},
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4], stage3_27[5]},
      {stage4_29[0],stage4_28[0],stage4_27[3],stage4_26[7],stage4_25[11]}
   );
   gpc1163_5 gpc8727 (
      {stage3_26[0], stage3_26[1], stage3_26[2]},
      {stage3_27[6], stage3_27[7], stage3_27[8], stage3_27[9], stage3_27[10], stage3_27[11]},
      {stage3_28[0]},
      {stage3_29[0]},
      {stage4_30[0],stage4_29[1],stage4_28[1],stage4_27[4],stage4_26[8]}
   );
   gpc1163_5 gpc8728 (
      {stage3_26[3], stage3_26[4], stage3_26[5]},
      {stage3_27[12], stage3_27[13], stage3_27[14], stage3_27[15], stage3_27[16], stage3_27[17]},
      {stage3_28[1]},
      {stage3_29[1]},
      {stage4_30[1],stage4_29[2],stage4_28[2],stage4_27[5],stage4_26[9]}
   );
   gpc1163_5 gpc8729 (
      {stage3_26[6], stage3_26[7], stage3_26[8]},
      {stage3_27[18], stage3_27[19], stage3_27[20], stage3_27[21], stage3_27[22], stage3_27[23]},
      {stage3_28[2]},
      {stage3_29[2]},
      {stage4_30[2],stage4_29[3],stage4_28[3],stage4_27[6],stage4_26[10]}
   );
   gpc615_5 gpc8730 (
      {stage3_26[9], stage3_26[10], stage3_26[11], stage3_26[12], stage3_26[13]},
      {stage3_27[24]},
      {stage3_28[3], stage3_28[4], stage3_28[5], stage3_28[6], stage3_28[7], stage3_28[8]},
      {stage4_30[3],stage4_29[4],stage4_28[4],stage4_27[7],stage4_26[11]}
   );
   gpc615_5 gpc8731 (
      {stage3_26[14], stage3_26[15], stage3_26[16], stage3_26[17], stage3_26[18]},
      {stage3_27[25]},
      {stage3_28[9], stage3_28[10], stage3_28[11], stage3_28[12], stage3_28[13], stage3_28[14]},
      {stage4_30[4],stage4_29[5],stage4_28[5],stage4_27[8],stage4_26[12]}
   );
   gpc615_5 gpc8732 (
      {stage3_26[19], stage3_26[20], stage3_26[21], stage3_26[22], stage3_26[23]},
      {stage3_27[26]},
      {stage3_28[15], stage3_28[16], stage3_28[17], stage3_28[18], stage3_28[19], stage3_28[20]},
      {stage4_30[5],stage4_29[6],stage4_28[6],stage4_27[9],stage4_26[13]}
   );
   gpc615_5 gpc8733 (
      {stage3_26[24], stage3_26[25], stage3_26[26], stage3_26[27], stage3_26[28]},
      {stage3_27[27]},
      {stage3_28[21], stage3_28[22], stage3_28[23], stage3_28[24], stage3_28[25], stage3_28[26]},
      {stage4_30[6],stage4_29[7],stage4_28[7],stage4_27[10],stage4_26[14]}
   );
   gpc615_5 gpc8734 (
      {stage3_26[29], stage3_26[30], stage3_26[31], stage3_26[32], stage3_26[33]},
      {stage3_27[28]},
      {stage3_28[27], stage3_28[28], stage3_28[29], stage3_28[30], stage3_28[31], stage3_28[32]},
      {stage4_30[7],stage4_29[8],stage4_28[8],stage4_27[11],stage4_26[15]}
   );
   gpc615_5 gpc8735 (
      {stage3_26[34], stage3_26[35], stage3_26[36], stage3_26[37], stage3_26[38]},
      {stage3_27[29]},
      {stage3_28[33], stage3_28[34], stage3_28[35], stage3_28[36], stage3_28[37], stage3_28[38]},
      {stage4_30[8],stage4_29[9],stage4_28[9],stage4_27[12],stage4_26[16]}
   );
   gpc615_5 gpc8736 (
      {stage3_26[39], stage3_26[40], stage3_26[41], stage3_26[42], stage3_26[43]},
      {stage3_27[30]},
      {stage3_28[39], stage3_28[40], stage3_28[41], stage3_28[42], stage3_28[43], stage3_28[44]},
      {stage4_30[9],stage4_29[10],stage4_28[10],stage4_27[13],stage4_26[17]}
   );
   gpc615_5 gpc8737 (
      {stage3_26[44], stage3_26[45], stage3_26[46], stage3_26[47], stage3_26[48]},
      {stage3_27[31]},
      {stage3_28[45], stage3_28[46], stage3_28[47], stage3_28[48], stage3_28[49], stage3_28[50]},
      {stage4_30[10],stage4_29[11],stage4_28[11],stage4_27[14],stage4_26[18]}
   );
   gpc606_5 gpc8738 (
      {stage3_27[32], stage3_27[33], stage3_27[34], stage3_27[35], stage3_27[36], stage3_27[37]},
      {stage3_29[3], stage3_29[4], stage3_29[5], stage3_29[6], stage3_29[7], stage3_29[8]},
      {stage4_31[0],stage4_30[11],stage4_29[12],stage4_28[12],stage4_27[15]}
   );
   gpc1163_5 gpc8739 (
      {stage3_29[9], stage3_29[10], stage3_29[11]},
      {stage3_30[0], stage3_30[1], stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5]},
      {stage3_31[0]},
      {stage3_32[0]},
      {stage4_33[0],stage4_32[0],stage4_31[1],stage4_30[12],stage4_29[13]}
   );
   gpc1163_5 gpc8740 (
      {stage3_29[12], stage3_29[13], stage3_29[14]},
      {stage3_30[6], stage3_30[7], stage3_30[8], stage3_30[9], stage3_30[10], stage3_30[11]},
      {stage3_31[1]},
      {stage3_32[1]},
      {stage4_33[1],stage4_32[1],stage4_31[2],stage4_30[13],stage4_29[14]}
   );
   gpc1163_5 gpc8741 (
      {stage3_29[15], stage3_29[16], stage3_29[17]},
      {stage3_30[12], stage3_30[13], stage3_30[14], stage3_30[15], stage3_30[16], stage3_30[17]},
      {stage3_31[2]},
      {stage3_32[2]},
      {stage4_33[2],stage4_32[2],stage4_31[3],stage4_30[14],stage4_29[15]}
   );
   gpc1163_5 gpc8742 (
      {stage3_29[18], stage3_29[19], stage3_29[20]},
      {stage3_30[18], stage3_30[19], stage3_30[20], stage3_30[21], stage3_30[22], stage3_30[23]},
      {stage3_31[3]},
      {stage3_32[3]},
      {stage4_33[3],stage4_32[3],stage4_31[4],stage4_30[15],stage4_29[16]}
   );
   gpc1163_5 gpc8743 (
      {stage3_29[21], stage3_29[22], stage3_29[23]},
      {stage3_30[24], stage3_30[25], stage3_30[26], stage3_30[27], stage3_30[28], stage3_30[29]},
      {stage3_31[4]},
      {stage3_32[4]},
      {stage4_33[4],stage4_32[4],stage4_31[5],stage4_30[16],stage4_29[17]}
   );
   gpc606_5 gpc8744 (
      {stage3_29[24], stage3_29[25], stage3_29[26], stage3_29[27], stage3_29[28], stage3_29[29]},
      {stage3_31[5], stage3_31[6], stage3_31[7], stage3_31[8], stage3_31[9], stage3_31[10]},
      {stage4_33[5],stage4_32[5],stage4_31[6],stage4_30[17],stage4_29[18]}
   );
   gpc606_5 gpc8745 (
      {stage3_29[30], stage3_29[31], stage3_29[32], stage3_29[33], stage3_29[34], stage3_29[35]},
      {stage3_31[11], stage3_31[12], stage3_31[13], stage3_31[14], stage3_31[15], stage3_31[16]},
      {stage4_33[6],stage4_32[6],stage4_31[7],stage4_30[18],stage4_29[19]}
   );
   gpc606_5 gpc8746 (
      {stage3_29[36], stage3_29[37], stage3_29[38], stage3_29[39], stage3_29[40], stage3_29[41]},
      {stage3_31[17], stage3_31[18], stage3_31[19], stage3_31[20], stage3_31[21], stage3_31[22]},
      {stage4_33[7],stage4_32[7],stage4_31[8],stage4_30[19],stage4_29[20]}
   );
   gpc606_5 gpc8747 (
      {stage3_29[42], stage3_29[43], stage3_29[44], stage3_29[45], stage3_29[46], stage3_29[47]},
      {stage3_31[23], stage3_31[24], stage3_31[25], stage3_31[26], stage3_31[27], stage3_31[28]},
      {stage4_33[8],stage4_32[8],stage4_31[9],stage4_30[20],stage4_29[21]}
   );
   gpc615_5 gpc8748 (
      {stage3_31[29], stage3_31[30], stage3_31[31], stage3_31[32], stage3_31[33]},
      {stage3_32[5]},
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4], stage3_33[5]},
      {stage4_35[0],stage4_34[0],stage4_33[9],stage4_32[9],stage4_31[10]}
   );
   gpc2135_5 gpc8749 (
      {stage3_32[6], stage3_32[7], stage3_32[8], stage3_32[9], stage3_32[10]},
      {stage3_33[6], stage3_33[7], stage3_33[8]},
      {stage3_34[0]},
      {stage3_35[0], stage3_35[1]},
      {stage4_36[0],stage4_35[1],stage4_34[1],stage4_33[10],stage4_32[10]}
   );
   gpc2135_5 gpc8750 (
      {stage3_32[11], stage3_32[12], stage3_32[13], stage3_32[14], stage3_32[15]},
      {stage3_33[9], stage3_33[10], stage3_33[11]},
      {stage3_34[1]},
      {stage3_35[2], stage3_35[3]},
      {stage4_36[1],stage4_35[2],stage4_34[2],stage4_33[11],stage4_32[11]}
   );
   gpc615_5 gpc8751 (
      {stage3_32[16], stage3_32[17], stage3_32[18], stage3_32[19], stage3_32[20]},
      {stage3_33[12]},
      {stage3_34[2], stage3_34[3], stage3_34[4], stage3_34[5], stage3_34[6], stage3_34[7]},
      {stage4_36[2],stage4_35[3],stage4_34[3],stage4_33[12],stage4_32[12]}
   );
   gpc615_5 gpc8752 (
      {stage3_32[21], stage3_32[22], stage3_32[23], stage3_32[24], stage3_32[25]},
      {stage3_33[13]},
      {stage3_34[8], stage3_34[9], stage3_34[10], stage3_34[11], stage3_34[12], stage3_34[13]},
      {stage4_36[3],stage4_35[4],stage4_34[4],stage4_33[13],stage4_32[13]}
   );
   gpc615_5 gpc8753 (
      {stage3_32[26], stage3_32[27], stage3_32[28], stage3_32[29], stage3_32[30]},
      {stage3_33[14]},
      {stage3_34[14], stage3_34[15], stage3_34[16], stage3_34[17], stage3_34[18], stage3_34[19]},
      {stage4_36[4],stage4_35[5],stage4_34[5],stage4_33[14],stage4_32[14]}
   );
   gpc615_5 gpc8754 (
      {stage3_32[31], stage3_32[32], stage3_32[33], stage3_32[34], stage3_32[35]},
      {stage3_33[15]},
      {stage3_34[20], stage3_34[21], stage3_34[22], stage3_34[23], stage3_34[24], stage3_34[25]},
      {stage4_36[5],stage4_35[6],stage4_34[6],stage4_33[15],stage4_32[15]}
   );
   gpc615_5 gpc8755 (
      {stage3_32[36], stage3_32[37], stage3_32[38], stage3_32[39], stage3_32[40]},
      {stage3_33[16]},
      {stage3_34[26], stage3_34[27], stage3_34[28], stage3_34[29], stage3_34[30], stage3_34[31]},
      {stage4_36[6],stage4_35[7],stage4_34[7],stage4_33[16],stage4_32[16]}
   );
   gpc117_4 gpc8756 (
      {stage3_33[17], stage3_33[18], stage3_33[19], stage3_33[20], stage3_33[21], stage3_33[22], stage3_33[23]},
      {stage3_34[32]},
      {stage3_35[4]},
      {stage4_36[7],stage4_35[8],stage4_34[8],stage4_33[17]}
   );
   gpc117_4 gpc8757 (
      {stage3_33[24], stage3_33[25], stage3_33[26], stage3_33[27], stage3_33[28], stage3_33[29], stage3_33[30]},
      {stage3_34[33]},
      {stage3_35[5]},
      {stage4_36[8],stage4_35[9],stage4_34[9],stage4_33[18]}
   );
   gpc606_5 gpc8758 (
      {stage3_33[31], stage3_33[32], stage3_33[33], stage3_33[34], stage3_33[35], stage3_33[36]},
      {stage3_35[6], stage3_35[7], stage3_35[8], stage3_35[9], stage3_35[10], stage3_35[11]},
      {stage4_37[0],stage4_36[9],stage4_35[10],stage4_34[10],stage4_33[19]}
   );
   gpc615_5 gpc8759 (
      {stage3_35[12], stage3_35[13], stage3_35[14], stage3_35[15], stage3_35[16]},
      {stage3_36[0]},
      {stage3_37[0], stage3_37[1], stage3_37[2], stage3_37[3], stage3_37[4], stage3_37[5]},
      {stage4_39[0],stage4_38[0],stage4_37[1],stage4_36[10],stage4_35[11]}
   );
   gpc615_5 gpc8760 (
      {stage3_35[17], stage3_35[18], stage3_35[19], stage3_35[20], stage3_35[21]},
      {stage3_36[1]},
      {stage3_37[6], stage3_37[7], stage3_37[8], stage3_37[9], stage3_37[10], stage3_37[11]},
      {stage4_39[1],stage4_38[1],stage4_37[2],stage4_36[11],stage4_35[12]}
   );
   gpc615_5 gpc8761 (
      {stage3_35[22], stage3_35[23], stage3_35[24], stage3_35[25], stage3_35[26]},
      {stage3_36[2]},
      {stage3_37[12], stage3_37[13], stage3_37[14], stage3_37[15], stage3_37[16], stage3_37[17]},
      {stage4_39[2],stage4_38[2],stage4_37[3],stage4_36[12],stage4_35[13]}
   );
   gpc615_5 gpc8762 (
      {stage3_35[27], stage3_35[28], stage3_35[29], stage3_35[30], stage3_35[31]},
      {stage3_36[3]},
      {stage3_37[18], stage3_37[19], stage3_37[20], stage3_37[21], stage3_37[22], stage3_37[23]},
      {stage4_39[3],stage4_38[3],stage4_37[4],stage4_36[13],stage4_35[14]}
   );
   gpc615_5 gpc8763 (
      {stage3_35[32], stage3_35[33], stage3_35[34], stage3_35[35], stage3_35[36]},
      {stage3_36[4]},
      {stage3_37[24], stage3_37[25], stage3_37[26], stage3_37[27], stage3_37[28], stage3_37[29]},
      {stage4_39[4],stage4_38[4],stage4_37[5],stage4_36[14],stage4_35[15]}
   );
   gpc606_5 gpc8764 (
      {stage3_36[5], stage3_36[6], stage3_36[7], stage3_36[8], stage3_36[9], stage3_36[10]},
      {stage3_38[0], stage3_38[1], stage3_38[2], stage3_38[3], stage3_38[4], stage3_38[5]},
      {stage4_40[0],stage4_39[5],stage4_38[5],stage4_37[6],stage4_36[15]}
   );
   gpc606_5 gpc8765 (
      {stage3_36[11], stage3_36[12], stage3_36[13], stage3_36[14], stage3_36[15], stage3_36[16]},
      {stage3_38[6], stage3_38[7], stage3_38[8], stage3_38[9], stage3_38[10], stage3_38[11]},
      {stage4_40[1],stage4_39[6],stage4_38[6],stage4_37[7],stage4_36[16]}
   );
   gpc606_5 gpc8766 (
      {stage3_36[17], stage3_36[18], stage3_36[19], stage3_36[20], stage3_36[21], stage3_36[22]},
      {stage3_38[12], stage3_38[13], stage3_38[14], stage3_38[15], stage3_38[16], stage3_38[17]},
      {stage4_40[2],stage4_39[7],stage4_38[7],stage4_37[8],stage4_36[17]}
   );
   gpc606_5 gpc8767 (
      {stage3_36[23], stage3_36[24], stage3_36[25], stage3_36[26], stage3_36[27], stage3_36[28]},
      {stage3_38[18], stage3_38[19], stage3_38[20], stage3_38[21], stage3_38[22], stage3_38[23]},
      {stage4_40[3],stage4_39[8],stage4_38[8],stage4_37[9],stage4_36[18]}
   );
   gpc606_5 gpc8768 (
      {stage3_37[30], stage3_37[31], stage3_37[32], stage3_37[33], stage3_37[34], stage3_37[35]},
      {stage3_39[0], stage3_39[1], stage3_39[2], stage3_39[3], stage3_39[4], stage3_39[5]},
      {stage4_41[0],stage4_40[4],stage4_39[9],stage4_38[9],stage4_37[10]}
   );
   gpc606_5 gpc8769 (
      {stage3_37[36], stage3_37[37], stage3_37[38], stage3_37[39], stage3_37[40], stage3_37[41]},
      {stage3_39[6], stage3_39[7], stage3_39[8], stage3_39[9], stage3_39[10], stage3_39[11]},
      {stage4_41[1],stage4_40[5],stage4_39[10],stage4_38[10],stage4_37[11]}
   );
   gpc606_5 gpc8770 (
      {stage3_37[42], stage3_37[43], stage3_37[44], stage3_37[45], stage3_37[46], stage3_37[47]},
      {stage3_39[12], stage3_39[13], stage3_39[14], stage3_39[15], stage3_39[16], stage3_39[17]},
      {stage4_41[2],stage4_40[6],stage4_39[11],stage4_38[11],stage4_37[12]}
   );
   gpc615_5 gpc8771 (
      {stage3_38[24], stage3_38[25], stage3_38[26], stage3_38[27], stage3_38[28]},
      {stage3_39[18]},
      {stage3_40[0], stage3_40[1], stage3_40[2], stage3_40[3], stage3_40[4], stage3_40[5]},
      {stage4_42[0],stage4_41[3],stage4_40[7],stage4_39[12],stage4_38[12]}
   );
   gpc615_5 gpc8772 (
      {stage3_38[29], stage3_38[30], stage3_38[31], stage3_38[32], stage3_38[33]},
      {stage3_39[19]},
      {stage3_40[6], stage3_40[7], stage3_40[8], stage3_40[9], stage3_40[10], stage3_40[11]},
      {stage4_42[1],stage4_41[4],stage4_40[8],stage4_39[13],stage4_38[13]}
   );
   gpc615_5 gpc8773 (
      {stage3_38[34], stage3_38[35], stage3_38[36], stage3_38[37], stage3_38[38]},
      {stage3_39[20]},
      {stage3_40[12], stage3_40[13], stage3_40[14], stage3_40[15], stage3_40[16], stage3_40[17]},
      {stage4_42[2],stage4_41[5],stage4_40[9],stage4_39[14],stage4_38[14]}
   );
   gpc615_5 gpc8774 (
      {stage3_38[39], stage3_38[40], stage3_38[41], stage3_38[42], stage3_38[43]},
      {stage3_39[21]},
      {stage3_40[18], stage3_40[19], stage3_40[20], stage3_40[21], stage3_40[22], stage3_40[23]},
      {stage4_42[3],stage4_41[6],stage4_40[10],stage4_39[15],stage4_38[15]}
   );
   gpc615_5 gpc8775 (
      {stage3_38[44], stage3_38[45], stage3_38[46], stage3_38[47], stage3_38[48]},
      {stage3_39[22]},
      {stage3_40[24], stage3_40[25], stage3_40[26], stage3_40[27], stage3_40[28], stage3_40[29]},
      {stage4_42[4],stage4_41[7],stage4_40[11],stage4_39[16],stage4_38[16]}
   );
   gpc615_5 gpc8776 (
      {stage3_38[49], stage3_38[50], stage3_38[51], stage3_38[52], stage3_38[53]},
      {stage3_39[23]},
      {stage3_40[30], stage3_40[31], stage3_40[32], stage3_40[33], stage3_40[34], stage3_40[35]},
      {stage4_42[5],stage4_41[8],stage4_40[12],stage4_39[17],stage4_38[17]}
   );
   gpc615_5 gpc8777 (
      {stage3_38[54], stage3_38[55], stage3_38[56], stage3_38[57], stage3_38[58]},
      {stage3_39[24]},
      {stage3_40[36], stage3_40[37], stage3_40[38], stage3_40[39], stage3_40[40], stage3_40[41]},
      {stage4_42[6],stage4_41[9],stage4_40[13],stage4_39[18],stage4_38[18]}
   );
   gpc207_4 gpc8778 (
      {stage3_39[25], stage3_39[26], stage3_39[27], stage3_39[28], stage3_39[29], stage3_39[30], stage3_39[31]},
      {stage3_41[0], stage3_41[1]},
      {stage4_42[7],stage4_41[10],stage4_40[14],stage4_39[19]}
   );
   gpc207_4 gpc8779 (
      {stage3_39[32], stage3_39[33], stage3_39[34], stage3_39[35], stage3_39[36], stage3_39[37], stage3_39[38]},
      {stage3_41[2], stage3_41[3]},
      {stage4_42[8],stage4_41[11],stage4_40[15],stage4_39[20]}
   );
   gpc207_4 gpc8780 (
      {stage3_39[39], stage3_39[40], stage3_39[41], stage3_39[42], stage3_39[43], stage3_39[44], stage3_39[45]},
      {stage3_41[4], stage3_41[5]},
      {stage4_42[9],stage4_41[12],stage4_40[16],stage4_39[21]}
   );
   gpc207_4 gpc8781 (
      {stage3_39[46], stage3_39[47], stage3_39[48], stage3_39[49], stage3_39[50], stage3_39[51], stage3_39[52]},
      {stage3_41[6], stage3_41[7]},
      {stage4_42[10],stage4_41[13],stage4_40[17],stage4_39[22]}
   );
   gpc615_5 gpc8782 (
      {stage3_39[53], stage3_39[54], stage3_39[55], stage3_39[56], stage3_39[57]},
      {stage3_40[42]},
      {stage3_41[8], stage3_41[9], stage3_41[10], stage3_41[11], stage3_41[12], stage3_41[13]},
      {stage4_43[0],stage4_42[11],stage4_41[14],stage4_40[18],stage4_39[23]}
   );
   gpc606_5 gpc8783 (
      {stage3_41[14], stage3_41[15], stage3_41[16], stage3_41[17], stage3_41[18], stage3_41[19]},
      {stage3_43[0], stage3_43[1], stage3_43[2], stage3_43[3], stage3_43[4], stage3_43[5]},
      {stage4_45[0],stage4_44[0],stage4_43[1],stage4_42[12],stage4_41[15]}
   );
   gpc606_5 gpc8784 (
      {stage3_41[20], stage3_41[21], stage3_41[22], stage3_41[23], stage3_41[24], stage3_41[25]},
      {stage3_43[6], stage3_43[7], stage3_43[8], stage3_43[9], stage3_43[10], stage3_43[11]},
      {stage4_45[1],stage4_44[1],stage4_43[2],stage4_42[13],stage4_41[16]}
   );
   gpc606_5 gpc8785 (
      {stage3_41[26], stage3_41[27], stage3_41[28], stage3_41[29], stage3_41[30], stage3_41[31]},
      {stage3_43[12], stage3_43[13], stage3_43[14], stage3_43[15], stage3_43[16], stage3_43[17]},
      {stage4_45[2],stage4_44[2],stage4_43[3],stage4_42[14],stage4_41[17]}
   );
   gpc606_5 gpc8786 (
      {stage3_41[32], stage3_41[33], stage3_41[34], stage3_41[35], stage3_41[36], stage3_41[37]},
      {stage3_43[18], stage3_43[19], stage3_43[20], stage3_43[21], stage3_43[22], stage3_43[23]},
      {stage4_45[3],stage4_44[3],stage4_43[4],stage4_42[15],stage4_41[18]}
   );
   gpc606_5 gpc8787 (
      {stage3_41[38], stage3_41[39], stage3_41[40], stage3_41[41], stage3_41[42], 1'b0},
      {stage3_43[24], stage3_43[25], stage3_43[26], stage3_43[27], stage3_43[28], stage3_43[29]},
      {stage4_45[4],stage4_44[4],stage4_43[5],stage4_42[16],stage4_41[19]}
   );
   gpc207_4 gpc8788 (
      {stage3_42[0], stage3_42[1], stage3_42[2], stage3_42[3], stage3_42[4], stage3_42[5], stage3_42[6]},
      {stage3_44[0], stage3_44[1]},
      {stage4_45[5],stage4_44[5],stage4_43[6],stage4_42[17]}
   );
   gpc207_4 gpc8789 (
      {stage3_42[7], stage3_42[8], stage3_42[9], stage3_42[10], stage3_42[11], stage3_42[12], stage3_42[13]},
      {stage3_44[2], stage3_44[3]},
      {stage4_45[6],stage4_44[6],stage4_43[7],stage4_42[18]}
   );
   gpc207_4 gpc8790 (
      {stage3_42[14], stage3_42[15], stage3_42[16], stage3_42[17], stage3_42[18], stage3_42[19], stage3_42[20]},
      {stage3_44[4], stage3_44[5]},
      {stage4_45[7],stage4_44[7],stage4_43[8],stage4_42[19]}
   );
   gpc207_4 gpc8791 (
      {stage3_42[21], stage3_42[22], stage3_42[23], stage3_42[24], stage3_42[25], stage3_42[26], stage3_42[27]},
      {stage3_44[6], stage3_44[7]},
      {stage4_45[8],stage4_44[8],stage4_43[9],stage4_42[20]}
   );
   gpc606_5 gpc8792 (
      {stage3_42[28], stage3_42[29], stage3_42[30], stage3_42[31], stage3_42[32], stage3_42[33]},
      {stage3_44[8], stage3_44[9], stage3_44[10], stage3_44[11], stage3_44[12], stage3_44[13]},
      {stage4_46[0],stage4_45[9],stage4_44[9],stage4_43[10],stage4_42[21]}
   );
   gpc606_5 gpc8793 (
      {stage3_43[30], stage3_43[31], stage3_43[32], stage3_43[33], stage3_43[34], stage3_43[35]},
      {stage3_45[0], stage3_45[1], stage3_45[2], stage3_45[3], stage3_45[4], stage3_45[5]},
      {stage4_47[0],stage4_46[1],stage4_45[10],stage4_44[10],stage4_43[11]}
   );
   gpc606_5 gpc8794 (
      {stage3_43[36], stage3_43[37], stage3_43[38], stage3_43[39], stage3_43[40], stage3_43[41]},
      {stage3_45[6], stage3_45[7], stage3_45[8], stage3_45[9], stage3_45[10], stage3_45[11]},
      {stage4_47[1],stage4_46[2],stage4_45[11],stage4_44[11],stage4_43[12]}
   );
   gpc615_5 gpc8795 (
      {stage3_43[42], stage3_43[43], stage3_43[44], stage3_43[45], 1'b0},
      {stage3_44[14]},
      {stage3_45[12], stage3_45[13], stage3_45[14], stage3_45[15], stage3_45[16], stage3_45[17]},
      {stage4_47[2],stage4_46[3],stage4_45[12],stage4_44[12],stage4_43[13]}
   );
   gpc606_5 gpc8796 (
      {stage3_44[15], stage3_44[16], stage3_44[17], stage3_44[18], stage3_44[19], stage3_44[20]},
      {stage3_46[0], stage3_46[1], stage3_46[2], stage3_46[3], stage3_46[4], stage3_46[5]},
      {stage4_48[0],stage4_47[3],stage4_46[4],stage4_45[13],stage4_44[13]}
   );
   gpc606_5 gpc8797 (
      {stage3_44[21], stage3_44[22], stage3_44[23], stage3_44[24], stage3_44[25], stage3_44[26]},
      {stage3_46[6], stage3_46[7], stage3_46[8], stage3_46[9], stage3_46[10], stage3_46[11]},
      {stage4_48[1],stage4_47[4],stage4_46[5],stage4_45[14],stage4_44[14]}
   );
   gpc615_5 gpc8798 (
      {stage3_44[27], stage3_44[28], stage3_44[29], stage3_44[30], stage3_44[31]},
      {stage3_45[18]},
      {stage3_46[12], stage3_46[13], stage3_46[14], stage3_46[15], stage3_46[16], stage3_46[17]},
      {stage4_48[2],stage4_47[5],stage4_46[6],stage4_45[15],stage4_44[15]}
   );
   gpc135_4 gpc8799 (
      {stage3_45[19], stage3_45[20], stage3_45[21], stage3_45[22], stage3_45[23]},
      {stage3_46[18], stage3_46[19], stage3_46[20]},
      {stage3_47[0]},
      {stage4_48[3],stage4_47[6],stage4_46[7],stage4_45[16]}
   );
   gpc135_4 gpc8800 (
      {stage3_45[24], stage3_45[25], stage3_45[26], stage3_45[27], stage3_45[28]},
      {stage3_46[21], stage3_46[22], stage3_46[23]},
      {stage3_47[1]},
      {stage4_48[4],stage4_47[7],stage4_46[8],stage4_45[17]}
   );
   gpc135_4 gpc8801 (
      {stage3_45[29], stage3_45[30], stage3_45[31], stage3_45[32], stage3_45[33]},
      {stage3_46[24], stage3_46[25], stage3_46[26]},
      {stage3_47[2]},
      {stage4_48[5],stage4_47[8],stage4_46[9],stage4_45[18]}
   );
   gpc615_5 gpc8802 (
      {stage3_46[27], stage3_46[28], stage3_46[29], stage3_46[30], stage3_46[31]},
      {stage3_47[3]},
      {stage3_48[0], stage3_48[1], stage3_48[2], stage3_48[3], stage3_48[4], stage3_48[5]},
      {stage4_50[0],stage4_49[0],stage4_48[6],stage4_47[9],stage4_46[10]}
   );
   gpc615_5 gpc8803 (
      {stage3_46[32], stage3_46[33], stage3_46[34], stage3_46[35], stage3_46[36]},
      {stage3_47[4]},
      {stage3_48[6], stage3_48[7], stage3_48[8], stage3_48[9], stage3_48[10], stage3_48[11]},
      {stage4_50[1],stage4_49[1],stage4_48[7],stage4_47[10],stage4_46[11]}
   );
   gpc615_5 gpc8804 (
      {stage3_46[37], stage3_46[38], stage3_46[39], stage3_46[40], stage3_46[41]},
      {stage3_47[5]},
      {stage3_48[12], stage3_48[13], stage3_48[14], stage3_48[15], stage3_48[16], stage3_48[17]},
      {stage4_50[2],stage4_49[2],stage4_48[8],stage4_47[11],stage4_46[12]}
   );
   gpc615_5 gpc8805 (
      {stage3_46[42], stage3_46[43], stage3_46[44], stage3_46[45], stage3_46[46]},
      {stage3_47[6]},
      {stage3_48[18], stage3_48[19], stage3_48[20], stage3_48[21], stage3_48[22], stage3_48[23]},
      {stage4_50[3],stage4_49[3],stage4_48[9],stage4_47[12],stage4_46[13]}
   );
   gpc615_5 gpc8806 (
      {stage3_46[47], stage3_46[48], stage3_46[49], stage3_46[50], stage3_46[51]},
      {stage3_47[7]},
      {stage3_48[24], stage3_48[25], stage3_48[26], stage3_48[27], stage3_48[28], stage3_48[29]},
      {stage4_50[4],stage4_49[4],stage4_48[10],stage4_47[13],stage4_46[14]}
   );
   gpc615_5 gpc8807 (
      {stage3_46[52], stage3_46[53], stage3_46[54], stage3_46[55], stage3_46[56]},
      {stage3_47[8]},
      {stage3_48[30], stage3_48[31], stage3_48[32], stage3_48[33], stage3_48[34], stage3_48[35]},
      {stage4_50[5],stage4_49[5],stage4_48[11],stage4_47[14],stage4_46[15]}
   );
   gpc606_5 gpc8808 (
      {stage3_47[9], stage3_47[10], stage3_47[11], stage3_47[12], stage3_47[13], stage3_47[14]},
      {stage3_49[0], stage3_49[1], stage3_49[2], stage3_49[3], stage3_49[4], stage3_49[5]},
      {stage4_51[0],stage4_50[6],stage4_49[6],stage4_48[12],stage4_47[15]}
   );
   gpc606_5 gpc8809 (
      {stage3_47[15], stage3_47[16], stage3_47[17], stage3_47[18], stage3_47[19], stage3_47[20]},
      {stage3_49[6], stage3_49[7], stage3_49[8], stage3_49[9], stage3_49[10], stage3_49[11]},
      {stage4_51[1],stage4_50[7],stage4_49[7],stage4_48[13],stage4_47[16]}
   );
   gpc606_5 gpc8810 (
      {stage3_47[21], stage3_47[22], stage3_47[23], stage3_47[24], stage3_47[25], stage3_47[26]},
      {stage3_49[12], stage3_49[13], stage3_49[14], stage3_49[15], stage3_49[16], stage3_49[17]},
      {stage4_51[2],stage4_50[8],stage4_49[8],stage4_48[14],stage4_47[17]}
   );
   gpc606_5 gpc8811 (
      {stage3_47[27], stage3_47[28], stage3_47[29], stage3_47[30], stage3_47[31], stage3_47[32]},
      {stage3_49[18], stage3_49[19], stage3_49[20], stage3_49[21], stage3_49[22], stage3_49[23]},
      {stage4_51[3],stage4_50[9],stage4_49[9],stage4_48[15],stage4_47[18]}
   );
   gpc606_5 gpc8812 (
      {stage3_47[33], stage3_47[34], stage3_47[35], stage3_47[36], stage3_47[37], stage3_47[38]},
      {stage3_49[24], stage3_49[25], stage3_49[26], stage3_49[27], stage3_49[28], stage3_49[29]},
      {stage4_51[4],stage4_50[10],stage4_49[10],stage4_48[16],stage4_47[19]}
   );
   gpc615_5 gpc8813 (
      {stage3_47[39], stage3_47[40], stage3_47[41], stage3_47[42], stage3_47[43]},
      {stage3_48[36]},
      {stage3_49[30], stage3_49[31], stage3_49[32], stage3_49[33], stage3_49[34], stage3_49[35]},
      {stage4_51[5],stage4_50[11],stage4_49[11],stage4_48[17],stage4_47[20]}
   );
   gpc606_5 gpc8814 (
      {stage3_49[36], stage3_49[37], stage3_49[38], stage3_49[39], stage3_49[40], stage3_49[41]},
      {stage3_51[0], stage3_51[1], stage3_51[2], stage3_51[3], stage3_51[4], stage3_51[5]},
      {stage4_53[0],stage4_52[0],stage4_51[6],stage4_50[12],stage4_49[12]}
   );
   gpc117_4 gpc8815 (
      {stage3_50[0], stage3_50[1], stage3_50[2], stage3_50[3], stage3_50[4], stage3_50[5], stage3_50[6]},
      {stage3_51[6]},
      {stage3_52[0]},
      {stage4_53[1],stage4_52[1],stage4_51[7],stage4_50[13]}
   );
   gpc117_4 gpc8816 (
      {stage3_50[7], stage3_50[8], stage3_50[9], stage3_50[10], stage3_50[11], stage3_50[12], stage3_50[13]},
      {stage3_51[7]},
      {stage3_52[1]},
      {stage4_53[2],stage4_52[2],stage4_51[8],stage4_50[14]}
   );
   gpc615_5 gpc8817 (
      {stage3_50[14], stage3_50[15], stage3_50[16], stage3_50[17], stage3_50[18]},
      {stage3_51[8]},
      {stage3_52[2], stage3_52[3], stage3_52[4], stage3_52[5], stage3_52[6], stage3_52[7]},
      {stage4_54[0],stage4_53[3],stage4_52[3],stage4_51[9],stage4_50[15]}
   );
   gpc615_5 gpc8818 (
      {stage3_50[19], stage3_50[20], stage3_50[21], stage3_50[22], stage3_50[23]},
      {stage3_51[9]},
      {stage3_52[8], stage3_52[9], stage3_52[10], stage3_52[11], stage3_52[12], stage3_52[13]},
      {stage4_54[1],stage4_53[4],stage4_52[4],stage4_51[10],stage4_50[16]}
   );
   gpc615_5 gpc8819 (
      {stage3_50[24], stage3_50[25], stage3_50[26], stage3_50[27], stage3_50[28]},
      {stage3_51[10]},
      {stage3_52[14], stage3_52[15], stage3_52[16], stage3_52[17], stage3_52[18], stage3_52[19]},
      {stage4_54[2],stage4_53[5],stage4_52[5],stage4_51[11],stage4_50[17]}
   );
   gpc615_5 gpc8820 (
      {stage3_50[29], stage3_50[30], stage3_50[31], stage3_50[32], stage3_50[33]},
      {stage3_51[11]},
      {stage3_52[20], stage3_52[21], stage3_52[22], stage3_52[23], stage3_52[24], stage3_52[25]},
      {stage4_54[3],stage4_53[6],stage4_52[6],stage4_51[12],stage4_50[18]}
   );
   gpc615_5 gpc8821 (
      {stage3_50[34], stage3_50[35], stage3_50[36], stage3_50[37], stage3_50[38]},
      {stage3_51[12]},
      {stage3_52[26], stage3_52[27], stage3_52[28], stage3_52[29], stage3_52[30], stage3_52[31]},
      {stage4_54[4],stage4_53[7],stage4_52[7],stage4_51[13],stage4_50[19]}
   );
   gpc615_5 gpc8822 (
      {stage3_50[39], stage3_50[40], stage3_50[41], stage3_50[42], stage3_50[43]},
      {stage3_51[13]},
      {stage3_52[32], stage3_52[33], stage3_52[34], stage3_52[35], stage3_52[36], stage3_52[37]},
      {stage4_54[5],stage4_53[8],stage4_52[8],stage4_51[14],stage4_50[20]}
   );
   gpc615_5 gpc8823 (
      {stage3_50[44], stage3_50[45], stage3_50[46], 1'b0, 1'b0},
      {stage3_51[14]},
      {stage3_52[38], stage3_52[39], stage3_52[40], stage3_52[41], stage3_52[42], stage3_52[43]},
      {stage4_54[6],stage4_53[9],stage4_52[9],stage4_51[15],stage4_50[21]}
   );
   gpc2135_5 gpc8824 (
      {stage3_51[15], stage3_51[16], stage3_51[17], stage3_51[18], stage3_51[19]},
      {stage3_52[44], stage3_52[45], stage3_52[46]},
      {stage3_53[0]},
      {stage3_54[0], stage3_54[1]},
      {stage4_55[0],stage4_54[7],stage4_53[10],stage4_52[10],stage4_51[16]}
   );
   gpc2135_5 gpc8825 (
      {stage3_51[20], stage3_51[21], stage3_51[22], stage3_51[23], stage3_51[24]},
      {stage3_52[47], stage3_52[48], stage3_52[49]},
      {stage3_53[1]},
      {stage3_54[2], stage3_54[3]},
      {stage4_55[1],stage4_54[8],stage4_53[11],stage4_52[11],stage4_51[17]}
   );
   gpc2135_5 gpc8826 (
      {stage3_51[25], stage3_51[26], stage3_51[27], stage3_51[28], stage3_51[29]},
      {stage3_52[50], stage3_52[51], stage3_52[52]},
      {stage3_53[2]},
      {stage3_54[4], stage3_54[5]},
      {stage4_55[2],stage4_54[9],stage4_53[12],stage4_52[12],stage4_51[18]}
   );
   gpc2135_5 gpc8827 (
      {stage3_51[30], stage3_51[31], stage3_51[32], stage3_51[33], stage3_51[34]},
      {stage3_52[53], stage3_52[54], stage3_52[55]},
      {stage3_53[3]},
      {stage3_54[6], stage3_54[7]},
      {stage4_55[3],stage4_54[10],stage4_53[13],stage4_52[13],stage4_51[19]}
   );
   gpc2135_5 gpc8828 (
      {stage3_51[35], stage3_51[36], stage3_51[37], stage3_51[38], stage3_51[39]},
      {stage3_52[56], stage3_52[57], stage3_52[58]},
      {stage3_53[4]},
      {stage3_54[8], stage3_54[9]},
      {stage4_55[4],stage4_54[11],stage4_53[14],stage4_52[14],stage4_51[20]}
   );
   gpc615_5 gpc8829 (
      {stage3_51[40], stage3_51[41], stage3_51[42], stage3_51[43], stage3_51[44]},
      {stage3_52[59]},
      {stage3_53[5], stage3_53[6], stage3_53[7], stage3_53[8], stage3_53[9], stage3_53[10]},
      {stage4_55[5],stage4_54[12],stage4_53[15],stage4_52[15],stage4_51[21]}
   );
   gpc615_5 gpc8830 (
      {stage3_51[45], stage3_51[46], stage3_51[47], stage3_51[48], stage3_51[49]},
      {stage3_52[60]},
      {stage3_53[11], stage3_53[12], stage3_53[13], stage3_53[14], stage3_53[15], stage3_53[16]},
      {stage4_55[6],stage4_54[13],stage4_53[16],stage4_52[16],stage4_51[22]}
   );
   gpc606_5 gpc8831 (
      {stage3_53[17], stage3_53[18], stage3_53[19], stage3_53[20], stage3_53[21], stage3_53[22]},
      {stage3_55[0], stage3_55[1], stage3_55[2], stage3_55[3], stage3_55[4], stage3_55[5]},
      {stage4_57[0],stage4_56[0],stage4_55[7],stage4_54[14],stage4_53[17]}
   );
   gpc606_5 gpc8832 (
      {stage3_53[23], stage3_53[24], stage3_53[25], stage3_53[26], stage3_53[27], stage3_53[28]},
      {stage3_55[6], stage3_55[7], stage3_55[8], stage3_55[9], stage3_55[10], stage3_55[11]},
      {stage4_57[1],stage4_56[1],stage4_55[8],stage4_54[15],stage4_53[18]}
   );
   gpc606_5 gpc8833 (
      {stage3_53[29], stage3_53[30], stage3_53[31], stage3_53[32], stage3_53[33], stage3_53[34]},
      {stage3_55[12], stage3_55[13], stage3_55[14], stage3_55[15], stage3_55[16], stage3_55[17]},
      {stage4_57[2],stage4_56[2],stage4_55[9],stage4_54[16],stage4_53[19]}
   );
   gpc615_5 gpc8834 (
      {stage3_53[35], stage3_53[36], stage3_53[37], stage3_53[38], stage3_53[39]},
      {stage3_54[10]},
      {stage3_55[18], stage3_55[19], stage3_55[20], stage3_55[21], stage3_55[22], stage3_55[23]},
      {stage4_57[3],stage4_56[3],stage4_55[10],stage4_54[17],stage4_53[20]}
   );
   gpc615_5 gpc8835 (
      {stage3_53[40], stage3_53[41], stage3_53[42], stage3_53[43], stage3_53[44]},
      {stage3_54[11]},
      {stage3_55[24], stage3_55[25], stage3_55[26], stage3_55[27], stage3_55[28], stage3_55[29]},
      {stage4_57[4],stage4_56[4],stage4_55[11],stage4_54[18],stage4_53[21]}
   );
   gpc615_5 gpc8836 (
      {stage3_53[45], stage3_53[46], stage3_53[47], stage3_53[48], stage3_53[49]},
      {stage3_54[12]},
      {stage3_55[30], stage3_55[31], stage3_55[32], stage3_55[33], stage3_55[34], stage3_55[35]},
      {stage4_57[5],stage4_56[5],stage4_55[12],stage4_54[19],stage4_53[22]}
   );
   gpc615_5 gpc8837 (
      {stage3_53[50], stage3_53[51], stage3_53[52], stage3_53[53], stage3_53[54]},
      {stage3_54[13]},
      {stage3_55[36], stage3_55[37], stage3_55[38], stage3_55[39], stage3_55[40], stage3_55[41]},
      {stage4_57[6],stage4_56[6],stage4_55[13],stage4_54[20],stage4_53[23]}
   );
   gpc615_5 gpc8838 (
      {stage3_54[14], stage3_54[15], stage3_54[16], stage3_54[17], stage3_54[18]},
      {stage3_55[42]},
      {stage3_56[0], stage3_56[1], stage3_56[2], stage3_56[3], stage3_56[4], stage3_56[5]},
      {stage4_58[0],stage4_57[7],stage4_56[7],stage4_55[14],stage4_54[21]}
   );
   gpc615_5 gpc8839 (
      {stage3_54[19], stage3_54[20], stage3_54[21], stage3_54[22], stage3_54[23]},
      {stage3_55[43]},
      {stage3_56[6], stage3_56[7], stage3_56[8], stage3_56[9], stage3_56[10], stage3_56[11]},
      {stage4_58[1],stage4_57[8],stage4_56[8],stage4_55[15],stage4_54[22]}
   );
   gpc615_5 gpc8840 (
      {stage3_54[24], stage3_54[25], stage3_54[26], stage3_54[27], stage3_54[28]},
      {stage3_55[44]},
      {stage3_56[12], stage3_56[13], stage3_56[14], stage3_56[15], stage3_56[16], stage3_56[17]},
      {stage4_58[2],stage4_57[9],stage4_56[9],stage4_55[16],stage4_54[23]}
   );
   gpc615_5 gpc8841 (
      {stage3_54[29], stage3_54[30], stage3_54[31], stage3_54[32], stage3_54[33]},
      {stage3_55[45]},
      {stage3_56[18], stage3_56[19], stage3_56[20], stage3_56[21], stage3_56[22], stage3_56[23]},
      {stage4_58[3],stage4_57[10],stage4_56[10],stage4_55[17],stage4_54[24]}
   );
   gpc615_5 gpc8842 (
      {stage3_54[34], stage3_54[35], stage3_54[36], stage3_54[37], stage3_54[38]},
      {stage3_55[46]},
      {stage3_56[24], stage3_56[25], stage3_56[26], stage3_56[27], stage3_56[28], stage3_56[29]},
      {stage4_58[4],stage4_57[11],stage4_56[11],stage4_55[18],stage4_54[25]}
   );
   gpc1163_5 gpc8843 (
      {stage3_57[0], stage3_57[1], stage3_57[2]},
      {stage3_58[0], stage3_58[1], stage3_58[2], stage3_58[3], stage3_58[4], stage3_58[5]},
      {stage3_59[0]},
      {stage3_60[0]},
      {stage4_61[0],stage4_60[0],stage4_59[0],stage4_58[5],stage4_57[12]}
   );
   gpc1163_5 gpc8844 (
      {stage3_57[3], stage3_57[4], stage3_57[5]},
      {stage3_58[6], stage3_58[7], stage3_58[8], stage3_58[9], stage3_58[10], stage3_58[11]},
      {stage3_59[1]},
      {stage3_60[1]},
      {stage4_61[1],stage4_60[1],stage4_59[1],stage4_58[6],stage4_57[13]}
   );
   gpc1163_5 gpc8845 (
      {stage3_57[6], stage3_57[7], stage3_57[8]},
      {stage3_58[12], stage3_58[13], stage3_58[14], stage3_58[15], stage3_58[16], stage3_58[17]},
      {stage3_59[2]},
      {stage3_60[2]},
      {stage4_61[2],stage4_60[2],stage4_59[2],stage4_58[7],stage4_57[14]}
   );
   gpc1163_5 gpc8846 (
      {stage3_57[9], stage3_57[10], stage3_57[11]},
      {stage3_58[18], stage3_58[19], stage3_58[20], stage3_58[21], stage3_58[22], stage3_58[23]},
      {stage3_59[3]},
      {stage3_60[3]},
      {stage4_61[3],stage4_60[3],stage4_59[3],stage4_58[8],stage4_57[15]}
   );
   gpc1163_5 gpc8847 (
      {stage3_57[12], stage3_57[13], stage3_57[14]},
      {stage3_58[24], stage3_58[25], stage3_58[26], stage3_58[27], stage3_58[28], stage3_58[29]},
      {stage3_59[4]},
      {stage3_60[4]},
      {stage4_61[4],stage4_60[4],stage4_59[4],stage4_58[9],stage4_57[16]}
   );
   gpc1163_5 gpc8848 (
      {stage3_57[15], stage3_57[16], stage3_57[17]},
      {stage3_58[30], stage3_58[31], stage3_58[32], stage3_58[33], stage3_58[34], stage3_58[35]},
      {stage3_59[5]},
      {stage3_60[5]},
      {stage4_61[5],stage4_60[5],stage4_59[5],stage4_58[10],stage4_57[17]}
   );
   gpc1163_5 gpc8849 (
      {stage3_57[18], stage3_57[19], stage3_57[20]},
      {stage3_58[36], stage3_58[37], stage3_58[38], stage3_58[39], stage3_58[40], stage3_58[41]},
      {stage3_59[6]},
      {stage3_60[6]},
      {stage4_61[6],stage4_60[6],stage4_59[6],stage4_58[11],stage4_57[18]}
   );
   gpc1163_5 gpc8850 (
      {stage3_57[21], stage3_57[22], stage3_57[23]},
      {stage3_58[42], stage3_58[43], stage3_58[44], stage3_58[45], stage3_58[46], stage3_58[47]},
      {stage3_59[7]},
      {stage3_60[7]},
      {stage4_61[7],stage4_60[7],stage4_59[7],stage4_58[12],stage4_57[19]}
   );
   gpc1163_5 gpc8851 (
      {stage3_57[24], stage3_57[25], stage3_57[26]},
      {stage3_58[48], stage3_58[49], stage3_58[50], stage3_58[51], stage3_58[52], stage3_58[53]},
      {stage3_59[8]},
      {stage3_60[8]},
      {stage4_61[8],stage4_60[8],stage4_59[8],stage4_58[13],stage4_57[20]}
   );
   gpc606_5 gpc8852 (
      {stage3_57[27], stage3_57[28], stage3_57[29], stage3_57[30], stage3_57[31], stage3_57[32]},
      {stage3_59[9], stage3_59[10], stage3_59[11], stage3_59[12], stage3_59[13], stage3_59[14]},
      {stage4_61[9],stage4_60[9],stage4_59[9],stage4_58[14],stage4_57[21]}
   );
   gpc606_5 gpc8853 (
      {stage3_57[33], stage3_57[34], stage3_57[35], stage3_57[36], stage3_57[37], stage3_57[38]},
      {stage3_59[15], stage3_59[16], stage3_59[17], stage3_59[18], stage3_59[19], stage3_59[20]},
      {stage4_61[10],stage4_60[10],stage4_59[10],stage4_58[15],stage4_57[22]}
   );
   gpc615_5 gpc8854 (
      {stage3_57[39], stage3_57[40], stage3_57[41], stage3_57[42], stage3_57[43]},
      {stage3_58[54]},
      {stage3_59[21], stage3_59[22], stage3_59[23], stage3_59[24], stage3_59[25], stage3_59[26]},
      {stage4_61[11],stage4_60[11],stage4_59[11],stage4_58[16],stage4_57[23]}
   );
   gpc615_5 gpc8855 (
      {stage3_57[44], stage3_57[45], stage3_57[46], stage3_57[47], stage3_57[48]},
      {stage3_58[55]},
      {stage3_59[27], stage3_59[28], stage3_59[29], stage3_59[30], stage3_59[31], stage3_59[32]},
      {stage4_61[12],stage4_60[12],stage4_59[12],stage4_58[17],stage4_57[24]}
   );
   gpc615_5 gpc8856 (
      {stage3_57[49], stage3_57[50], stage3_57[51], stage3_57[52], stage3_57[53]},
      {stage3_58[56]},
      {stage3_59[33], stage3_59[34], stage3_59[35], stage3_59[36], stage3_59[37], stage3_59[38]},
      {stage4_61[13],stage4_60[13],stage4_59[13],stage4_58[18],stage4_57[25]}
   );
   gpc615_5 gpc8857 (
      {stage3_59[39], stage3_59[40], stage3_59[41], stage3_59[42], stage3_59[43]},
      {stage3_60[9]},
      {stage3_61[0], stage3_61[1], stage3_61[2], stage3_61[3], stage3_61[4], stage3_61[5]},
      {stage4_63[0],stage4_62[0],stage4_61[14],stage4_60[14],stage4_59[14]}
   );
   gpc606_5 gpc8858 (
      {stage3_60[10], stage3_60[11], stage3_60[12], stage3_60[13], stage3_60[14], stage3_60[15]},
      {stage3_62[0], stage3_62[1], stage3_62[2], stage3_62[3], stage3_62[4], stage3_62[5]},
      {stage4_64[0],stage4_63[1],stage4_62[1],stage4_61[15],stage4_60[15]}
   );
   gpc606_5 gpc8859 (
      {stage3_60[16], stage3_60[17], stage3_60[18], stage3_60[19], stage3_60[20], stage3_60[21]},
      {stage3_62[6], stage3_62[7], stage3_62[8], stage3_62[9], stage3_62[10], stage3_62[11]},
      {stage4_64[1],stage4_63[2],stage4_62[2],stage4_61[16],stage4_60[16]}
   );
   gpc606_5 gpc8860 (
      {stage3_60[22], stage3_60[23], stage3_60[24], stage3_60[25], stage3_60[26], stage3_60[27]},
      {stage3_62[12], stage3_62[13], stage3_62[14], stage3_62[15], stage3_62[16], stage3_62[17]},
      {stage4_64[2],stage4_63[3],stage4_62[3],stage4_61[17],stage4_60[17]}
   );
   gpc606_5 gpc8861 (
      {stage3_60[28], stage3_60[29], stage3_60[30], stage3_60[31], stage3_60[32], stage3_60[33]},
      {stage3_62[18], stage3_62[19], stage3_62[20], stage3_62[21], stage3_62[22], stage3_62[23]},
      {stage4_64[3],stage4_63[4],stage4_62[4],stage4_61[18],stage4_60[18]}
   );
   gpc606_5 gpc8862 (
      {stage3_60[34], stage3_60[35], stage3_60[36], stage3_60[37], stage3_60[38], stage3_60[39]},
      {stage3_62[24], stage3_62[25], stage3_62[26], stage3_62[27], stage3_62[28], stage3_62[29]},
      {stage4_64[4],stage4_63[5],stage4_62[5],stage4_61[19],stage4_60[19]}
   );
   gpc606_5 gpc8863 (
      {stage3_61[6], stage3_61[7], stage3_61[8], stage3_61[9], stage3_61[10], stage3_61[11]},
      {stage3_63[0], stage3_63[1], stage3_63[2], stage3_63[3], stage3_63[4], stage3_63[5]},
      {stage4_65[0],stage4_64[5],stage4_63[6],stage4_62[6],stage4_61[20]}
   );
   gpc606_5 gpc8864 (
      {stage3_61[12], stage3_61[13], stage3_61[14], stage3_61[15], stage3_61[16], stage3_61[17]},
      {stage3_63[6], stage3_63[7], stage3_63[8], stage3_63[9], stage3_63[10], stage3_63[11]},
      {stage4_65[1],stage4_64[6],stage4_63[7],stage4_62[7],stage4_61[21]}
   );
   gpc606_5 gpc8865 (
      {stage3_61[18], stage3_61[19], stage3_61[20], stage3_61[21], stage3_61[22], stage3_61[23]},
      {stage3_63[12], stage3_63[13], stage3_63[14], stage3_63[15], stage3_63[16], stage3_63[17]},
      {stage4_65[2],stage4_64[7],stage4_63[8],stage4_62[8],stage4_61[22]}
   );
   gpc606_5 gpc8866 (
      {stage3_61[24], stage3_61[25], stage3_61[26], stage3_61[27], stage3_61[28], stage3_61[29]},
      {stage3_63[18], stage3_63[19], stage3_63[20], stage3_63[21], stage3_63[22], stage3_63[23]},
      {stage4_65[3],stage4_64[8],stage4_63[9],stage4_62[9],stage4_61[23]}
   );
   gpc606_5 gpc8867 (
      {stage3_61[30], stage3_61[31], stage3_61[32], stage3_61[33], stage3_61[34], stage3_61[35]},
      {stage3_63[24], stage3_63[25], stage3_63[26], stage3_63[27], stage3_63[28], stage3_63[29]},
      {stage4_65[4],stage4_64[9],stage4_63[10],stage4_62[10],stage4_61[24]}
   );
   gpc606_5 gpc8868 (
      {stage3_61[36], stage3_61[37], stage3_61[38], stage3_61[39], stage3_61[40], stage3_61[41]},
      {stage3_63[30], stage3_63[31], stage3_63[32], stage3_63[33], stage3_63[34], stage3_63[35]},
      {stage4_65[5],stage4_64[10],stage4_63[11],stage4_62[11],stage4_61[25]}
   );
   gpc606_5 gpc8869 (
      {stage3_61[42], stage3_61[43], stage3_61[44], stage3_61[45], stage3_61[46], stage3_61[47]},
      {stage3_63[36], stage3_63[37], stage3_63[38], stage3_63[39], stage3_63[40], stage3_63[41]},
      {stage4_65[6],stage4_64[11],stage4_63[12],stage4_62[12],stage4_61[26]}
   );
   gpc606_5 gpc8870 (
      {stage3_63[42], stage3_63[43], stage3_63[44], stage3_63[45], stage3_63[46], stage3_63[47]},
      {stage3_65[0], stage3_65[1], stage3_65[2], stage3_65[3], stage3_65[4], stage3_65[5]},
      {stage4_67[0],stage4_66[0],stage4_65[7],stage4_64[12],stage4_63[13]}
   );
   gpc606_5 gpc8871 (
      {stage3_64[0], stage3_64[1], stage3_64[2], stage3_64[3], stage3_64[4], stage3_64[5]},
      {stage3_66[0], stage3_66[1], stage3_66[2], stage3_66[3], stage3_66[4], stage3_66[5]},
      {stage4_68[0],stage4_67[1],stage4_66[1],stage4_65[8],stage4_64[13]}
   );
   gpc606_5 gpc8872 (
      {stage3_64[6], stage3_64[7], stage3_64[8], stage3_64[9], stage3_64[10], stage3_64[11]},
      {stage3_66[6], stage3_66[7], stage3_66[8], stage3_66[9], stage3_66[10], stage3_66[11]},
      {stage4_68[1],stage4_67[2],stage4_66[2],stage4_65[9],stage4_64[14]}
   );
   gpc606_5 gpc8873 (
      {stage3_64[12], stage3_64[13], stage3_64[14], stage3_64[15], stage3_64[16], stage3_64[17]},
      {stage3_66[12], stage3_66[13], stage3_66[14], stage3_66[15], stage3_66[16], stage3_66[17]},
      {stage4_68[2],stage4_67[3],stage4_66[3],stage4_65[10],stage4_64[15]}
   );
   gpc606_5 gpc8874 (
      {stage3_64[18], stage3_64[19], stage3_64[20], stage3_64[21], stage3_64[22], stage3_64[23]},
      {stage3_66[18], stage3_66[19], stage3_66[20], stage3_66[21], stage3_66[22], stage3_66[23]},
      {stage4_68[3],stage4_67[4],stage4_66[4],stage4_65[11],stage4_64[16]}
   );
   gpc606_5 gpc8875 (
      {stage3_64[24], stage3_64[25], stage3_64[26], stage3_64[27], stage3_64[28], stage3_64[29]},
      {stage3_66[24], stage3_66[25], stage3_66[26], stage3_66[27], stage3_66[28], stage3_66[29]},
      {stage4_68[4],stage4_67[5],stage4_66[5],stage4_65[12],stage4_64[17]}
   );
   gpc606_5 gpc8876 (
      {stage3_64[30], stage3_64[31], stage3_64[32], stage3_64[33], stage3_64[34], stage3_64[35]},
      {stage3_66[30], stage3_66[31], stage3_66[32], stage3_66[33], stage3_66[34], stage3_66[35]},
      {stage4_68[5],stage4_67[6],stage4_66[6],stage4_65[13],stage4_64[18]}
   );
   gpc606_5 gpc8877 (
      {stage3_65[6], stage3_65[7], stage3_65[8], stage3_65[9], stage3_65[10], stage3_65[11]},
      {stage3_67[0], stage3_67[1], stage3_67[2], stage3_67[3], stage3_67[4], stage3_67[5]},
      {stage4_69[0],stage4_68[6],stage4_67[7],stage4_66[7],stage4_65[14]}
   );
   gpc606_5 gpc8878 (
      {stage3_65[12], stage3_65[13], stage3_65[14], stage3_65[15], stage3_65[16], stage3_65[17]},
      {stage3_67[6], stage3_67[7], stage3_67[8], stage3_67[9], stage3_67[10], stage3_67[11]},
      {stage4_69[1],stage4_68[7],stage4_67[8],stage4_66[8],stage4_65[15]}
   );
   gpc1_1 gpc8879 (
      {stage3_0[15]},
      {stage4_0[3]}
   );
   gpc1_1 gpc8880 (
      {stage3_0[16]},
      {stage4_0[4]}
   );
   gpc1_1 gpc8881 (
      {stage3_0[17]},
      {stage4_0[5]}
   );
   gpc1_1 gpc8882 (
      {stage3_0[18]},
      {stage4_0[6]}
   );
   gpc1_1 gpc8883 (
      {stage3_0[19]},
      {stage4_0[7]}
   );
   gpc1_1 gpc8884 (
      {stage3_0[20]},
      {stage4_0[8]}
   );
   gpc1_1 gpc8885 (
      {stage3_1[21]},
      {stage4_1[6]}
   );
   gpc1_1 gpc8886 (
      {stage3_2[42]},
      {stage4_2[10]}
   );
   gpc1_1 gpc8887 (
      {stage3_3[23]},
      {stage4_3[11]}
   );
   gpc1_1 gpc8888 (
      {stage3_3[24]},
      {stage4_3[12]}
   );
   gpc1_1 gpc8889 (
      {stage3_3[25]},
      {stage4_3[13]}
   );
   gpc1_1 gpc8890 (
      {stage3_3[26]},
      {stage4_3[14]}
   );
   gpc1_1 gpc8891 (
      {stage3_3[27]},
      {stage4_3[15]}
   );
   gpc1_1 gpc8892 (
      {stage3_3[28]},
      {stage4_3[16]}
   );
   gpc1_1 gpc8893 (
      {stage3_4[109]},
      {stage4_4[28]}
   );
   gpc1_1 gpc8894 (
      {stage3_4[110]},
      {stage4_4[29]}
   );
   gpc1_1 gpc8895 (
      {stage3_4[111]},
      {stage4_4[30]}
   );
   gpc1_1 gpc8896 (
      {stage3_5[42]},
      {stage4_5[25]}
   );
   gpc1_1 gpc8897 (
      {stage3_5[43]},
      {stage4_5[26]}
   );
   gpc1_1 gpc8898 (
      {stage3_5[44]},
      {stage4_5[27]}
   );
   gpc1_1 gpc8899 (
      {stage3_5[45]},
      {stage4_5[28]}
   );
   gpc1_1 gpc8900 (
      {stage3_5[46]},
      {stage4_5[29]}
   );
   gpc1_1 gpc8901 (
      {stage3_5[47]},
      {stage4_5[30]}
   );
   gpc1_1 gpc8902 (
      {stage3_5[48]},
      {stage4_5[31]}
   );
   gpc1_1 gpc8903 (
      {stage3_5[49]},
      {stage4_5[32]}
   );
   gpc1_1 gpc8904 (
      {stage3_5[50]},
      {stage4_5[33]}
   );
   gpc1_1 gpc8905 (
      {stage3_5[51]},
      {stage4_5[34]}
   );
   gpc1_1 gpc8906 (
      {stage3_5[52]},
      {stage4_5[35]}
   );
   gpc1_1 gpc8907 (
      {stage3_6[77]},
      {stage4_6[23]}
   );
   gpc1_1 gpc8908 (
      {stage3_7[37]},
      {stage4_7[25]}
   );
   gpc1_1 gpc8909 (
      {stage3_7[38]},
      {stage4_7[26]}
   );
   gpc1_1 gpc8910 (
      {stage3_7[39]},
      {stage4_7[27]}
   );
   gpc1_1 gpc8911 (
      {stage3_7[40]},
      {stage4_7[28]}
   );
   gpc1_1 gpc8912 (
      {stage3_7[41]},
      {stage4_7[29]}
   );
   gpc1_1 gpc8913 (
      {stage3_7[42]},
      {stage4_7[30]}
   );
   gpc1_1 gpc8914 (
      {stage3_7[43]},
      {stage4_7[31]}
   );
   gpc1_1 gpc8915 (
      {stage3_7[44]},
      {stage4_7[32]}
   );
   gpc1_1 gpc8916 (
      {stage3_7[45]},
      {stage4_7[33]}
   );
   gpc1_1 gpc8917 (
      {stage3_7[46]},
      {stage4_7[34]}
   );
   gpc1_1 gpc8918 (
      {stage3_7[47]},
      {stage4_7[35]}
   );
   gpc1_1 gpc8919 (
      {stage3_7[48]},
      {stage4_7[36]}
   );
   gpc1_1 gpc8920 (
      {stage3_7[49]},
      {stage4_7[37]}
   );
   gpc1_1 gpc8921 (
      {stage3_7[50]},
      {stage4_7[38]}
   );
   gpc1_1 gpc8922 (
      {stage3_10[84]},
      {stage4_10[26]}
   );
   gpc1_1 gpc8923 (
      {stage3_10[85]},
      {stage4_10[27]}
   );
   gpc1_1 gpc8924 (
      {stage3_10[86]},
      {stage4_10[28]}
   );
   gpc1_1 gpc8925 (
      {stage3_10[87]},
      {stage4_10[29]}
   );
   gpc1_1 gpc8926 (
      {stage3_10[88]},
      {stage4_10[30]}
   );
   gpc1_1 gpc8927 (
      {stage3_10[89]},
      {stage4_10[31]}
   );
   gpc1_1 gpc8928 (
      {stage3_10[90]},
      {stage4_10[32]}
   );
   gpc1_1 gpc8929 (
      {stage3_10[91]},
      {stage4_10[33]}
   );
   gpc1_1 gpc8930 (
      {stage3_10[92]},
      {stage4_10[34]}
   );
   gpc1_1 gpc8931 (
      {stage3_10[93]},
      {stage4_10[35]}
   );
   gpc1_1 gpc8932 (
      {stage3_10[94]},
      {stage4_10[36]}
   );
   gpc1_1 gpc8933 (
      {stage3_10[95]},
      {stage4_10[37]}
   );
   gpc1_1 gpc8934 (
      {stage3_10[96]},
      {stage4_10[38]}
   );
   gpc1_1 gpc8935 (
      {stage3_10[97]},
      {stage4_10[39]}
   );
   gpc1_1 gpc8936 (
      {stage3_10[98]},
      {stage4_10[40]}
   );
   gpc1_1 gpc8937 (
      {stage3_10[99]},
      {stage4_10[41]}
   );
   gpc1_1 gpc8938 (
      {stage3_12[67]},
      {stage4_12[23]}
   );
   gpc1_1 gpc8939 (
      {stage3_13[50]},
      {stage4_13[25]}
   );
   gpc1_1 gpc8940 (
      {stage3_13[51]},
      {stage4_13[26]}
   );
   gpc1_1 gpc8941 (
      {stage3_13[52]},
      {stage4_13[27]}
   );
   gpc1_1 gpc8942 (
      {stage3_13[53]},
      {stage4_13[28]}
   );
   gpc1_1 gpc8943 (
      {stage3_13[54]},
      {stage4_13[29]}
   );
   gpc1_1 gpc8944 (
      {stage3_13[55]},
      {stage4_13[30]}
   );
   gpc1_1 gpc8945 (
      {stage3_13[56]},
      {stage4_13[31]}
   );
   gpc1_1 gpc8946 (
      {stage3_14[30]},
      {stage4_14[28]}
   );
   gpc1_1 gpc8947 (
      {stage3_14[31]},
      {stage4_14[29]}
   );
   gpc1_1 gpc8948 (
      {stage3_15[47]},
      {stage4_15[14]}
   );
   gpc1_1 gpc8949 (
      {stage3_16[37]},
      {stage4_16[13]}
   );
   gpc1_1 gpc8950 (
      {stage3_16[38]},
      {stage4_16[14]}
   );
   gpc1_1 gpc8951 (
      {stage3_16[39]},
      {stage4_16[15]}
   );
   gpc1_1 gpc8952 (
      {stage3_16[40]},
      {stage4_16[16]}
   );
   gpc1_1 gpc8953 (
      {stage3_16[41]},
      {stage4_16[17]}
   );
   gpc1_1 gpc8954 (
      {stage3_16[42]},
      {stage4_16[18]}
   );
   gpc1_1 gpc8955 (
      {stage3_16[43]},
      {stage4_16[19]}
   );
   gpc1_1 gpc8956 (
      {stage3_16[44]},
      {stage4_16[20]}
   );
   gpc1_1 gpc8957 (
      {stage3_16[45]},
      {stage4_16[21]}
   );
   gpc1_1 gpc8958 (
      {stage3_16[46]},
      {stage4_16[22]}
   );
   gpc1_1 gpc8959 (
      {stage3_16[47]},
      {stage4_16[23]}
   );
   gpc1_1 gpc8960 (
      {stage3_16[48]},
      {stage4_16[24]}
   );
   gpc1_1 gpc8961 (
      {stage3_16[49]},
      {stage4_16[25]}
   );
   gpc1_1 gpc8962 (
      {stage3_16[50]},
      {stage4_16[26]}
   );
   gpc1_1 gpc8963 (
      {stage3_19[35]},
      {stage4_19[16]}
   );
   gpc1_1 gpc8964 (
      {stage3_19[36]},
      {stage4_19[17]}
   );
   gpc1_1 gpc8965 (
      {stage3_19[37]},
      {stage4_19[18]}
   );
   gpc1_1 gpc8966 (
      {stage3_19[38]},
      {stage4_19[19]}
   );
   gpc1_1 gpc8967 (
      {stage3_19[39]},
      {stage4_19[20]}
   );
   gpc1_1 gpc8968 (
      {stage3_19[40]},
      {stage4_19[21]}
   );
   gpc1_1 gpc8969 (
      {stage3_19[41]},
      {stage4_19[22]}
   );
   gpc1_1 gpc8970 (
      {stage3_19[42]},
      {stage4_19[23]}
   );
   gpc1_1 gpc8971 (
      {stage3_19[43]},
      {stage4_19[24]}
   );
   gpc1_1 gpc8972 (
      {stage3_19[44]},
      {stage4_19[25]}
   );
   gpc1_1 gpc8973 (
      {stage3_19[45]},
      {stage4_19[26]}
   );
   gpc1_1 gpc8974 (
      {stage3_19[46]},
      {stage4_19[27]}
   );
   gpc1_1 gpc8975 (
      {stage3_19[47]},
      {stage4_19[28]}
   );
   gpc1_1 gpc8976 (
      {stage3_20[73]},
      {stage4_20[24]}
   );
   gpc1_1 gpc8977 (
      {stage3_20[74]},
      {stage4_20[25]}
   );
   gpc1_1 gpc8978 (
      {stage3_20[75]},
      {stage4_20[26]}
   );
   gpc1_1 gpc8979 (
      {stage3_20[76]},
      {stage4_20[27]}
   );
   gpc1_1 gpc8980 (
      {stage3_20[77]},
      {stage4_20[28]}
   );
   gpc1_1 gpc8981 (
      {stage3_20[78]},
      {stage4_20[29]}
   );
   gpc1_1 gpc8982 (
      {stage3_20[79]},
      {stage4_20[30]}
   );
   gpc1_1 gpc8983 (
      {stage3_20[80]},
      {stage4_20[31]}
   );
   gpc1_1 gpc8984 (
      {stage3_20[81]},
      {stage4_20[32]}
   );
   gpc1_1 gpc8985 (
      {stage3_20[82]},
      {stage4_20[33]}
   );
   gpc1_1 gpc8986 (
      {stage3_21[30]},
      {stage4_21[28]}
   );
   gpc1_1 gpc8987 (
      {stage3_21[31]},
      {stage4_21[29]}
   );
   gpc1_1 gpc8988 (
      {stage3_21[32]},
      {stage4_21[30]}
   );
   gpc1_1 gpc8989 (
      {stage3_21[33]},
      {stage4_21[31]}
   );
   gpc1_1 gpc8990 (
      {stage3_21[34]},
      {stage4_21[32]}
   );
   gpc1_1 gpc8991 (
      {stage3_21[35]},
      {stage4_21[33]}
   );
   gpc1_1 gpc8992 (
      {stage3_21[36]},
      {stage4_21[34]}
   );
   gpc1_1 gpc8993 (
      {stage3_21[37]},
      {stage4_21[35]}
   );
   gpc1_1 gpc8994 (
      {stage3_21[38]},
      {stage4_21[36]}
   );
   gpc1_1 gpc8995 (
      {stage3_24[27]},
      {stage4_24[20]}
   );
   gpc1_1 gpc8996 (
      {stage3_24[28]},
      {stage4_24[21]}
   );
   gpc1_1 gpc8997 (
      {stage3_25[24]},
      {stage4_25[12]}
   );
   gpc1_1 gpc8998 (
      {stage3_25[25]},
      {stage4_25[13]}
   );
   gpc1_1 gpc8999 (
      {stage3_25[26]},
      {stage4_25[14]}
   );
   gpc1_1 gpc9000 (
      {stage3_25[27]},
      {stage4_25[15]}
   );
   gpc1_1 gpc9001 (
      {stage3_25[28]},
      {stage4_25[16]}
   );
   gpc1_1 gpc9002 (
      {stage3_25[29]},
      {stage4_25[17]}
   );
   gpc1_1 gpc9003 (
      {stage3_25[30]},
      {stage4_25[18]}
   );
   gpc1_1 gpc9004 (
      {stage3_25[31]},
      {stage4_25[19]}
   );
   gpc1_1 gpc9005 (
      {stage3_25[32]},
      {stage4_25[20]}
   );
   gpc1_1 gpc9006 (
      {stage3_27[38]},
      {stage4_27[16]}
   );
   gpc1_1 gpc9007 (
      {stage3_27[39]},
      {stage4_27[17]}
   );
   gpc1_1 gpc9008 (
      {stage3_27[40]},
      {stage4_27[18]}
   );
   gpc1_1 gpc9009 (
      {stage3_27[41]},
      {stage4_27[19]}
   );
   gpc1_1 gpc9010 (
      {stage3_27[42]},
      {stage4_27[20]}
   );
   gpc1_1 gpc9011 (
      {stage3_27[43]},
      {stage4_27[21]}
   );
   gpc1_1 gpc9012 (
      {stage3_27[44]},
      {stage4_27[22]}
   );
   gpc1_1 gpc9013 (
      {stage3_27[45]},
      {stage4_27[23]}
   );
   gpc1_1 gpc9014 (
      {stage3_27[46]},
      {stage4_27[24]}
   );
   gpc1_1 gpc9015 (
      {stage3_27[47]},
      {stage4_27[25]}
   );
   gpc1_1 gpc9016 (
      {stage3_27[48]},
      {stage4_27[26]}
   );
   gpc1_1 gpc9017 (
      {stage3_28[51]},
      {stage4_28[13]}
   );
   gpc1_1 gpc9018 (
      {stage3_28[52]},
      {stage4_28[14]}
   );
   gpc1_1 gpc9019 (
      {stage3_28[53]},
      {stage4_28[15]}
   );
   gpc1_1 gpc9020 (
      {stage3_28[54]},
      {stage4_28[16]}
   );
   gpc1_1 gpc9021 (
      {stage3_28[55]},
      {stage4_28[17]}
   );
   gpc1_1 gpc9022 (
      {stage3_28[56]},
      {stage4_28[18]}
   );
   gpc1_1 gpc9023 (
      {stage3_30[30]},
      {stage4_30[21]}
   );
   gpc1_1 gpc9024 (
      {stage3_30[31]},
      {stage4_30[22]}
   );
   gpc1_1 gpc9025 (
      {stage3_30[32]},
      {stage4_30[23]}
   );
   gpc1_1 gpc9026 (
      {stage3_30[33]},
      {stage4_30[24]}
   );
   gpc1_1 gpc9027 (
      {stage3_30[34]},
      {stage4_30[25]}
   );
   gpc1_1 gpc9028 (
      {stage3_30[35]},
      {stage4_30[26]}
   );
   gpc1_1 gpc9029 (
      {stage3_30[36]},
      {stage4_30[27]}
   );
   gpc1_1 gpc9030 (
      {stage3_30[37]},
      {stage4_30[28]}
   );
   gpc1_1 gpc9031 (
      {stage3_30[38]},
      {stage4_30[29]}
   );
   gpc1_1 gpc9032 (
      {stage3_30[39]},
      {stage4_30[30]}
   );
   gpc1_1 gpc9033 (
      {stage3_30[40]},
      {stage4_30[31]}
   );
   gpc1_1 gpc9034 (
      {stage3_30[41]},
      {stage4_30[32]}
   );
   gpc1_1 gpc9035 (
      {stage3_31[34]},
      {stage4_31[11]}
   );
   gpc1_1 gpc9036 (
      {stage3_31[35]},
      {stage4_31[12]}
   );
   gpc1_1 gpc9037 (
      {stage3_31[36]},
      {stage4_31[13]}
   );
   gpc1_1 gpc9038 (
      {stage3_31[37]},
      {stage4_31[14]}
   );
   gpc1_1 gpc9039 (
      {stage3_32[41]},
      {stage4_32[17]}
   );
   gpc1_1 gpc9040 (
      {stage3_32[42]},
      {stage4_32[18]}
   );
   gpc1_1 gpc9041 (
      {stage3_32[43]},
      {stage4_32[19]}
   );
   gpc1_1 gpc9042 (
      {stage3_32[44]},
      {stage4_32[20]}
   );
   gpc1_1 gpc9043 (
      {stage3_32[45]},
      {stage4_32[21]}
   );
   gpc1_1 gpc9044 (
      {stage3_32[46]},
      {stage4_32[22]}
   );
   gpc1_1 gpc9045 (
      {stage3_32[47]},
      {stage4_32[23]}
   );
   gpc1_1 gpc9046 (
      {stage3_32[48]},
      {stage4_32[24]}
   );
   gpc1_1 gpc9047 (
      {stage3_32[49]},
      {stage4_32[25]}
   );
   gpc1_1 gpc9048 (
      {stage3_32[50]},
      {stage4_32[26]}
   );
   gpc1_1 gpc9049 (
      {stage3_32[51]},
      {stage4_32[27]}
   );
   gpc1_1 gpc9050 (
      {stage3_32[52]},
      {stage4_32[28]}
   );
   gpc1_1 gpc9051 (
      {stage3_32[53]},
      {stage4_32[29]}
   );
   gpc1_1 gpc9052 (
      {stage3_33[37]},
      {stage4_33[20]}
   );
   gpc1_1 gpc9053 (
      {stage3_33[38]},
      {stage4_33[21]}
   );
   gpc1_1 gpc9054 (
      {stage3_33[39]},
      {stage4_33[22]}
   );
   gpc1_1 gpc9055 (
      {stage3_33[40]},
      {stage4_33[23]}
   );
   gpc1_1 gpc9056 (
      {stage3_33[41]},
      {stage4_33[24]}
   );
   gpc1_1 gpc9057 (
      {stage3_33[42]},
      {stage4_33[25]}
   );
   gpc1_1 gpc9058 (
      {stage3_33[43]},
      {stage4_33[26]}
   );
   gpc1_1 gpc9059 (
      {stage3_33[44]},
      {stage4_33[27]}
   );
   gpc1_1 gpc9060 (
      {stage3_33[45]},
      {stage4_33[28]}
   );
   gpc1_1 gpc9061 (
      {stage3_34[34]},
      {stage4_34[11]}
   );
   gpc1_1 gpc9062 (
      {stage3_34[35]},
      {stage4_34[12]}
   );
   gpc1_1 gpc9063 (
      {stage3_34[36]},
      {stage4_34[13]}
   );
   gpc1_1 gpc9064 (
      {stage3_34[37]},
      {stage4_34[14]}
   );
   gpc1_1 gpc9065 (
      {stage3_34[38]},
      {stage4_34[15]}
   );
   gpc1_1 gpc9066 (
      {stage3_34[39]},
      {stage4_34[16]}
   );
   gpc1_1 gpc9067 (
      {stage3_34[40]},
      {stage4_34[17]}
   );
   gpc1_1 gpc9068 (
      {stage3_34[41]},
      {stage4_34[18]}
   );
   gpc1_1 gpc9069 (
      {stage3_35[37]},
      {stage4_35[16]}
   );
   gpc1_1 gpc9070 (
      {stage3_35[38]},
      {stage4_35[17]}
   );
   gpc1_1 gpc9071 (
      {stage3_35[39]},
      {stage4_35[18]}
   );
   gpc1_1 gpc9072 (
      {stage3_35[40]},
      {stage4_35[19]}
   );
   gpc1_1 gpc9073 (
      {stage3_35[41]},
      {stage4_35[20]}
   );
   gpc1_1 gpc9074 (
      {stage3_35[42]},
      {stage4_35[21]}
   );
   gpc1_1 gpc9075 (
      {stage3_35[43]},
      {stage4_35[22]}
   );
   gpc1_1 gpc9076 (
      {stage3_35[44]},
      {stage4_35[23]}
   );
   gpc1_1 gpc9077 (
      {stage3_35[45]},
      {stage4_35[24]}
   );
   gpc1_1 gpc9078 (
      {stage3_35[46]},
      {stage4_35[25]}
   );
   gpc1_1 gpc9079 (
      {stage3_35[47]},
      {stage4_35[26]}
   );
   gpc1_1 gpc9080 (
      {stage3_35[48]},
      {stage4_35[27]}
   );
   gpc1_1 gpc9081 (
      {stage3_35[49]},
      {stage4_35[28]}
   );
   gpc1_1 gpc9082 (
      {stage3_35[50]},
      {stage4_35[29]}
   );
   gpc1_1 gpc9083 (
      {stage3_35[51]},
      {stage4_35[30]}
   );
   gpc1_1 gpc9084 (
      {stage3_35[52]},
      {stage4_35[31]}
   );
   gpc1_1 gpc9085 (
      {stage3_35[53]},
      {stage4_35[32]}
   );
   gpc1_1 gpc9086 (
      {stage3_35[54]},
      {stage4_35[33]}
   );
   gpc1_1 gpc9087 (
      {stage3_35[55]},
      {stage4_35[34]}
   );
   gpc1_1 gpc9088 (
      {stage3_35[56]},
      {stage4_35[35]}
   );
   gpc1_1 gpc9089 (
      {stage3_36[29]},
      {stage4_36[19]}
   );
   gpc1_1 gpc9090 (
      {stage3_36[30]},
      {stage4_36[20]}
   );
   gpc1_1 gpc9091 (
      {stage3_36[31]},
      {stage4_36[21]}
   );
   gpc1_1 gpc9092 (
      {stage3_36[32]},
      {stage4_36[22]}
   );
   gpc1_1 gpc9093 (
      {stage3_36[33]},
      {stage4_36[23]}
   );
   gpc1_1 gpc9094 (
      {stage3_36[34]},
      {stage4_36[24]}
   );
   gpc1_1 gpc9095 (
      {stage3_36[35]},
      {stage4_36[25]}
   );
   gpc1_1 gpc9096 (
      {stage3_36[36]},
      {stage4_36[26]}
   );
   gpc1_1 gpc9097 (
      {stage3_36[37]},
      {stage4_36[27]}
   );
   gpc1_1 gpc9098 (
      {stage3_36[38]},
      {stage4_36[28]}
   );
   gpc1_1 gpc9099 (
      {stage3_36[39]},
      {stage4_36[29]}
   );
   gpc1_1 gpc9100 (
      {stage3_36[40]},
      {stage4_36[30]}
   );
   gpc1_1 gpc9101 (
      {stage3_36[41]},
      {stage4_36[31]}
   );
   gpc1_1 gpc9102 (
      {stage3_36[42]},
      {stage4_36[32]}
   );
   gpc1_1 gpc9103 (
      {stage3_36[43]},
      {stage4_36[33]}
   );
   gpc1_1 gpc9104 (
      {stage3_36[44]},
      {stage4_36[34]}
   );
   gpc1_1 gpc9105 (
      {stage3_36[45]},
      {stage4_36[35]}
   );
   gpc1_1 gpc9106 (
      {stage3_37[48]},
      {stage4_37[13]}
   );
   gpc1_1 gpc9107 (
      {stage3_37[49]},
      {stage4_37[14]}
   );
   gpc1_1 gpc9108 (
      {stage3_37[50]},
      {stage4_37[15]}
   );
   gpc1_1 gpc9109 (
      {stage3_37[51]},
      {stage4_37[16]}
   );
   gpc1_1 gpc9110 (
      {stage3_37[52]},
      {stage4_37[17]}
   );
   gpc1_1 gpc9111 (
      {stage3_38[59]},
      {stage4_38[19]}
   );
   gpc1_1 gpc9112 (
      {stage3_40[43]},
      {stage4_40[19]}
   );
   gpc1_1 gpc9113 (
      {stage3_40[44]},
      {stage4_40[20]}
   );
   gpc1_1 gpc9114 (
      {stage3_40[45]},
      {stage4_40[21]}
   );
   gpc1_1 gpc9115 (
      {stage3_40[46]},
      {stage4_40[22]}
   );
   gpc1_1 gpc9116 (
      {stage3_40[47]},
      {stage4_40[23]}
   );
   gpc1_1 gpc9117 (
      {stage3_40[48]},
      {stage4_40[24]}
   );
   gpc1_1 gpc9118 (
      {stage3_40[49]},
      {stage4_40[25]}
   );
   gpc1_1 gpc9119 (
      {stage3_40[50]},
      {stage4_40[26]}
   );
   gpc1_1 gpc9120 (
      {stage3_40[51]},
      {stage4_40[27]}
   );
   gpc1_1 gpc9121 (
      {stage3_42[34]},
      {stage4_42[22]}
   );
   gpc1_1 gpc9122 (
      {stage3_42[35]},
      {stage4_42[23]}
   );
   gpc1_1 gpc9123 (
      {stage3_42[36]},
      {stage4_42[24]}
   );
   gpc1_1 gpc9124 (
      {stage3_42[37]},
      {stage4_42[25]}
   );
   gpc1_1 gpc9125 (
      {stage3_42[38]},
      {stage4_42[26]}
   );
   gpc1_1 gpc9126 (
      {stage3_42[39]},
      {stage4_42[27]}
   );
   gpc1_1 gpc9127 (
      {stage3_42[40]},
      {stage4_42[28]}
   );
   gpc1_1 gpc9128 (
      {stage3_42[41]},
      {stage4_42[29]}
   );
   gpc1_1 gpc9129 (
      {stage3_42[42]},
      {stage4_42[30]}
   );
   gpc1_1 gpc9130 (
      {stage3_42[43]},
      {stage4_42[31]}
   );
   gpc1_1 gpc9131 (
      {stage3_42[44]},
      {stage4_42[32]}
   );
   gpc1_1 gpc9132 (
      {stage3_42[45]},
      {stage4_42[33]}
   );
   gpc1_1 gpc9133 (
      {stage3_42[46]},
      {stage4_42[34]}
   );
   gpc1_1 gpc9134 (
      {stage3_42[47]},
      {stage4_42[35]}
   );
   gpc1_1 gpc9135 (
      {stage3_42[48]},
      {stage4_42[36]}
   );
   gpc1_1 gpc9136 (
      {stage3_42[49]},
      {stage4_42[37]}
   );
   gpc1_1 gpc9137 (
      {stage3_44[32]},
      {stage4_44[16]}
   );
   gpc1_1 gpc9138 (
      {stage3_44[33]},
      {stage4_44[17]}
   );
   gpc1_1 gpc9139 (
      {stage3_44[34]},
      {stage4_44[18]}
   );
   gpc1_1 gpc9140 (
      {stage3_44[35]},
      {stage4_44[19]}
   );
   gpc1_1 gpc9141 (
      {stage3_44[36]},
      {stage4_44[20]}
   );
   gpc1_1 gpc9142 (
      {stage3_44[37]},
      {stage4_44[21]}
   );
   gpc1_1 gpc9143 (
      {stage3_44[38]},
      {stage4_44[22]}
   );
   gpc1_1 gpc9144 (
      {stage3_44[39]},
      {stage4_44[23]}
   );
   gpc1_1 gpc9145 (
      {stage3_44[40]},
      {stage4_44[24]}
   );
   gpc1_1 gpc9146 (
      {stage3_45[34]},
      {stage4_45[19]}
   );
   gpc1_1 gpc9147 (
      {stage3_45[35]},
      {stage4_45[20]}
   );
   gpc1_1 gpc9148 (
      {stage3_45[36]},
      {stage4_45[21]}
   );
   gpc1_1 gpc9149 (
      {stage3_45[37]},
      {stage4_45[22]}
   );
   gpc1_1 gpc9150 (
      {stage3_45[38]},
      {stage4_45[23]}
   );
   gpc1_1 gpc9151 (
      {stage3_45[39]},
      {stage4_45[24]}
   );
   gpc1_1 gpc9152 (
      {stage3_45[40]},
      {stage4_45[25]}
   );
   gpc1_1 gpc9153 (
      {stage3_45[41]},
      {stage4_45[26]}
   );
   gpc1_1 gpc9154 (
      {stage3_45[42]},
      {stage4_45[27]}
   );
   gpc1_1 gpc9155 (
      {stage3_45[43]},
      {stage4_45[28]}
   );
   gpc1_1 gpc9156 (
      {stage3_46[57]},
      {stage4_46[16]}
   );
   gpc1_1 gpc9157 (
      {stage3_48[37]},
      {stage4_48[18]}
   );
   gpc1_1 gpc9158 (
      {stage3_48[38]},
      {stage4_48[19]}
   );
   gpc1_1 gpc9159 (
      {stage3_48[39]},
      {stage4_48[20]}
   );
   gpc1_1 gpc9160 (
      {stage3_48[40]},
      {stage4_48[21]}
   );
   gpc1_1 gpc9161 (
      {stage3_48[41]},
      {stage4_48[22]}
   );
   gpc1_1 gpc9162 (
      {stage3_51[50]},
      {stage4_51[23]}
   );
   gpc1_1 gpc9163 (
      {stage3_51[51]},
      {stage4_51[24]}
   );
   gpc1_1 gpc9164 (
      {stage3_51[52]},
      {stage4_51[25]}
   );
   gpc1_1 gpc9165 (
      {stage3_51[53]},
      {stage4_51[26]}
   );
   gpc1_1 gpc9166 (
      {stage3_51[54]},
      {stage4_51[27]}
   );
   gpc1_1 gpc9167 (
      {stage3_51[55]},
      {stage4_51[28]}
   );
   gpc1_1 gpc9168 (
      {stage3_51[56]},
      {stage4_51[29]}
   );
   gpc1_1 gpc9169 (
      {stage3_51[57]},
      {stage4_51[30]}
   );
   gpc1_1 gpc9170 (
      {stage3_51[58]},
      {stage4_51[31]}
   );
   gpc1_1 gpc9171 (
      {stage3_51[59]},
      {stage4_51[32]}
   );
   gpc1_1 gpc9172 (
      {stage3_51[60]},
      {stage4_51[33]}
   );
   gpc1_1 gpc9173 (
      {stage3_51[61]},
      {stage4_51[34]}
   );
   gpc1_1 gpc9174 (
      {stage3_51[62]},
      {stage4_51[35]}
   );
   gpc1_1 gpc9175 (
      {stage3_52[61]},
      {stage4_52[17]}
   );
   gpc1_1 gpc9176 (
      {stage3_52[62]},
      {stage4_52[18]}
   );
   gpc1_1 gpc9177 (
      {stage3_53[55]},
      {stage4_53[24]}
   );
   gpc1_1 gpc9178 (
      {stage3_53[56]},
      {stage4_53[25]}
   );
   gpc1_1 gpc9179 (
      {stage3_53[57]},
      {stage4_53[26]}
   );
   gpc1_1 gpc9180 (
      {stage3_53[58]},
      {stage4_53[27]}
   );
   gpc1_1 gpc9181 (
      {stage3_53[59]},
      {stage4_53[28]}
   );
   gpc1_1 gpc9182 (
      {stage3_53[60]},
      {stage4_53[29]}
   );
   gpc1_1 gpc9183 (
      {stage3_53[61]},
      {stage4_53[30]}
   );
   gpc1_1 gpc9184 (
      {stage3_53[62]},
      {stage4_53[31]}
   );
   gpc1_1 gpc9185 (
      {stage3_53[63]},
      {stage4_53[32]}
   );
   gpc1_1 gpc9186 (
      {stage3_53[64]},
      {stage4_53[33]}
   );
   gpc1_1 gpc9187 (
      {stage3_53[65]},
      {stage4_53[34]}
   );
   gpc1_1 gpc9188 (
      {stage3_53[66]},
      {stage4_53[35]}
   );
   gpc1_1 gpc9189 (
      {stage3_53[67]},
      {stage4_53[36]}
   );
   gpc1_1 gpc9190 (
      {stage3_53[68]},
      {stage4_53[37]}
   );
   gpc1_1 gpc9191 (
      {stage3_53[69]},
      {stage4_53[38]}
   );
   gpc1_1 gpc9192 (
      {stage3_53[70]},
      {stage4_53[39]}
   );
   gpc1_1 gpc9193 (
      {stage3_53[71]},
      {stage4_53[40]}
   );
   gpc1_1 gpc9194 (
      {stage3_53[72]},
      {stage4_53[41]}
   );
   gpc1_1 gpc9195 (
      {stage3_53[73]},
      {stage4_53[42]}
   );
   gpc1_1 gpc9196 (
      {stage3_53[74]},
      {stage4_53[43]}
   );
   gpc1_1 gpc9197 (
      {stage3_55[47]},
      {stage4_55[19]}
   );
   gpc1_1 gpc9198 (
      {stage3_55[48]},
      {stage4_55[20]}
   );
   gpc1_1 gpc9199 (
      {stage3_55[49]},
      {stage4_55[21]}
   );
   gpc1_1 gpc9200 (
      {stage3_55[50]},
      {stage4_55[22]}
   );
   gpc1_1 gpc9201 (
      {stage3_55[51]},
      {stage4_55[23]}
   );
   gpc1_1 gpc9202 (
      {stage3_55[52]},
      {stage4_55[24]}
   );
   gpc1_1 gpc9203 (
      {stage3_55[53]},
      {stage4_55[25]}
   );
   gpc1_1 gpc9204 (
      {stage3_55[54]},
      {stage4_55[26]}
   );
   gpc1_1 gpc9205 (
      {stage3_55[55]},
      {stage4_55[27]}
   );
   gpc1_1 gpc9206 (
      {stage3_55[56]},
      {stage4_55[28]}
   );
   gpc1_1 gpc9207 (
      {stage3_55[57]},
      {stage4_55[29]}
   );
   gpc1_1 gpc9208 (
      {stage3_55[58]},
      {stage4_55[30]}
   );
   gpc1_1 gpc9209 (
      {stage3_55[59]},
      {stage4_55[31]}
   );
   gpc1_1 gpc9210 (
      {stage3_55[60]},
      {stage4_55[32]}
   );
   gpc1_1 gpc9211 (
      {stage3_55[61]},
      {stage4_55[33]}
   );
   gpc1_1 gpc9212 (
      {stage3_55[62]},
      {stage4_55[34]}
   );
   gpc1_1 gpc9213 (
      {stage3_55[63]},
      {stage4_55[35]}
   );
   gpc1_1 gpc9214 (
      {stage3_55[64]},
      {stage4_55[36]}
   );
   gpc1_1 gpc9215 (
      {stage3_55[65]},
      {stage4_55[37]}
   );
   gpc1_1 gpc9216 (
      {stage3_55[66]},
      {stage4_55[38]}
   );
   gpc1_1 gpc9217 (
      {stage3_56[30]},
      {stage4_56[12]}
   );
   gpc1_1 gpc9218 (
      {stage3_56[31]},
      {stage4_56[13]}
   );
   gpc1_1 gpc9219 (
      {stage3_58[57]},
      {stage4_58[19]}
   );
   gpc1_1 gpc9220 (
      {stage3_58[58]},
      {stage4_58[20]}
   );
   gpc1_1 gpc9221 (
      {stage3_58[59]},
      {stage4_58[21]}
   );
   gpc1_1 gpc9222 (
      {stage3_58[60]},
      {stage4_58[22]}
   );
   gpc1_1 gpc9223 (
      {stage3_58[61]},
      {stage4_58[23]}
   );
   gpc1_1 gpc9224 (
      {stage3_59[44]},
      {stage4_59[15]}
   );
   gpc1_1 gpc9225 (
      {stage3_59[45]},
      {stage4_59[16]}
   );
   gpc1_1 gpc9226 (
      {stage3_59[46]},
      {stage4_59[17]}
   );
   gpc1_1 gpc9227 (
      {stage3_59[47]},
      {stage4_59[18]}
   );
   gpc1_1 gpc9228 (
      {stage3_59[48]},
      {stage4_59[19]}
   );
   gpc1_1 gpc9229 (
      {stage3_59[49]},
      {stage4_59[20]}
   );
   gpc1_1 gpc9230 (
      {stage3_60[40]},
      {stage4_60[20]}
   );
   gpc1_1 gpc9231 (
      {stage3_60[41]},
      {stage4_60[21]}
   );
   gpc1_1 gpc9232 (
      {stage3_61[48]},
      {stage4_61[27]}
   );
   gpc1_1 gpc9233 (
      {stage3_61[49]},
      {stage4_61[28]}
   );
   gpc1_1 gpc9234 (
      {stage3_61[50]},
      {stage4_61[29]}
   );
   gpc1_1 gpc9235 (
      {stage3_61[51]},
      {stage4_61[30]}
   );
   gpc1_1 gpc9236 (
      {stage3_61[52]},
      {stage4_61[31]}
   );
   gpc1_1 gpc9237 (
      {stage3_62[30]},
      {stage4_62[13]}
   );
   gpc1_1 gpc9238 (
      {stage3_62[31]},
      {stage4_62[14]}
   );
   gpc1_1 gpc9239 (
      {stage3_62[32]},
      {stage4_62[15]}
   );
   gpc1_1 gpc9240 (
      {stage3_62[33]},
      {stage4_62[16]}
   );
   gpc1_1 gpc9241 (
      {stage3_64[36]},
      {stage4_64[19]}
   );
   gpc1_1 gpc9242 (
      {stage3_64[37]},
      {stage4_64[20]}
   );
   gpc1_1 gpc9243 (
      {stage3_64[38]},
      {stage4_64[21]}
   );
   gpc1_1 gpc9244 (
      {stage3_64[39]},
      {stage4_64[22]}
   );
   gpc1_1 gpc9245 (
      {stage3_64[40]},
      {stage4_64[23]}
   );
   gpc1_1 gpc9246 (
      {stage3_64[41]},
      {stage4_64[24]}
   );
   gpc1_1 gpc9247 (
      {stage3_64[42]},
      {stage4_64[25]}
   );
   gpc1_1 gpc9248 (
      {stage3_64[43]},
      {stage4_64[26]}
   );
   gpc1_1 gpc9249 (
      {stage3_64[44]},
      {stage4_64[27]}
   );
   gpc1_1 gpc9250 (
      {stage3_64[45]},
      {stage4_64[28]}
   );
   gpc1_1 gpc9251 (
      {stage3_64[46]},
      {stage4_64[29]}
   );
   gpc1_1 gpc9252 (
      {stage3_64[47]},
      {stage4_64[30]}
   );
   gpc1_1 gpc9253 (
      {stage3_64[48]},
      {stage4_64[31]}
   );
   gpc1_1 gpc9254 (
      {stage3_64[49]},
      {stage4_64[32]}
   );
   gpc1_1 gpc9255 (
      {stage3_64[50]},
      {stage4_64[33]}
   );
   gpc1_1 gpc9256 (
      {stage3_65[18]},
      {stage4_65[16]}
   );
   gpc1_1 gpc9257 (
      {stage3_65[19]},
      {stage4_65[17]}
   );
   gpc1_1 gpc9258 (
      {stage3_65[20]},
      {stage4_65[18]}
   );
   gpc1_1 gpc9259 (
      {stage3_65[21]},
      {stage4_65[19]}
   );
   gpc1_1 gpc9260 (
      {stage3_65[22]},
      {stage4_65[20]}
   );
   gpc1_1 gpc9261 (
      {stage3_65[23]},
      {stage4_65[21]}
   );
   gpc1_1 gpc9262 (
      {stage3_65[24]},
      {stage4_65[22]}
   );
   gpc1_1 gpc9263 (
      {stage3_65[25]},
      {stage4_65[23]}
   );
   gpc1_1 gpc9264 (
      {stage3_65[26]},
      {stage4_65[24]}
   );
   gpc1_1 gpc9265 (
      {stage3_65[27]},
      {stage4_65[25]}
   );
   gpc1_1 gpc9266 (
      {stage3_65[28]},
      {stage4_65[26]}
   );
   gpc1_1 gpc9267 (
      {stage3_65[29]},
      {stage4_65[27]}
   );
   gpc1_1 gpc9268 (
      {stage3_65[30]},
      {stage4_65[28]}
   );
   gpc1_1 gpc9269 (
      {stage3_65[31]},
      {stage4_65[29]}
   );
   gpc1_1 gpc9270 (
      {stage3_65[32]},
      {stage4_65[30]}
   );
   gpc1_1 gpc9271 (
      {stage3_65[33]},
      {stage4_65[31]}
   );
   gpc1_1 gpc9272 (
      {stage3_65[34]},
      {stage4_65[32]}
   );
   gpc1_1 gpc9273 (
      {stage3_65[35]},
      {stage4_65[33]}
   );
   gpc1_1 gpc9274 (
      {stage3_65[36]},
      {stage4_65[34]}
   );
   gpc1_1 gpc9275 (
      {stage3_65[37]},
      {stage4_65[35]}
   );
   gpc1_1 gpc9276 (
      {stage3_66[36]},
      {stage4_66[9]}
   );
   gpc1_1 gpc9277 (
      {stage3_66[37]},
      {stage4_66[10]}
   );
   gpc1_1 gpc9278 (
      {stage3_67[12]},
      {stage4_67[9]}
   );
   gpc1_1 gpc9279 (
      {stage3_67[13]},
      {stage4_67[10]}
   );
   gpc1_1 gpc9280 (
      {stage3_68[0]},
      {stage4_68[8]}
   );
   gpc1_1 gpc9281 (
      {stage3_68[1]},
      {stage4_68[9]}
   );
   gpc1_1 gpc9282 (
      {stage3_68[2]},
      {stage4_68[10]}
   );
   gpc1_1 gpc9283 (
      {stage3_68[3]},
      {stage4_68[11]}
   );
   gpc1_1 gpc9284 (
      {stage3_68[4]},
      {stage4_68[12]}
   );
   gpc1_1 gpc9285 (
      {stage3_68[5]},
      {stage4_68[13]}
   );
   gpc615_5 gpc9286 (
      {stage4_0[0], stage4_0[1], stage4_0[2], stage4_0[3], stage4_0[4]},
      {stage4_1[0]},
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4], stage4_2[5]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc606_5 gpc9287 (
      {stage4_1[1], stage4_1[2], stage4_1[3], stage4_1[4], stage4_1[5], stage4_1[6]},
      {stage4_3[0], stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5]},
      {stage5_5[0],stage5_4[1],stage5_3[1],stage5_2[1],stage5_1[1]}
   );
   gpc1163_5 gpc9288 (
      {stage4_2[6], stage4_2[7], stage4_2[8]},
      {stage4_3[6], stage4_3[7], stage4_3[8], stage4_3[9], stage4_3[10], stage4_3[11]},
      {stage4_4[0]},
      {stage4_5[0]},
      {stage5_6[0],stage5_5[1],stage5_4[2],stage5_3[2],stage5_2[2]}
   );
   gpc1163_5 gpc9289 (
      {stage4_4[1], stage4_4[2], stage4_4[3]},
      {stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5], stage4_5[6]},
      {stage4_6[0]},
      {stage4_7[0]},
      {stage5_8[0],stage5_7[0],stage5_6[1],stage5_5[2],stage5_4[3]}
   );
   gpc606_5 gpc9290 (
      {stage4_4[4], stage4_4[5], stage4_4[6], stage4_4[7], stage4_4[8], stage4_4[9]},
      {stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5], stage4_6[6]},
      {stage5_8[1],stage5_7[1],stage5_6[2],stage5_5[3],stage5_4[4]}
   );
   gpc606_5 gpc9291 (
      {stage4_4[10], stage4_4[11], stage4_4[12], stage4_4[13], stage4_4[14], stage4_4[15]},
      {stage4_6[7], stage4_6[8], stage4_6[9], stage4_6[10], stage4_6[11], stage4_6[12]},
      {stage5_8[2],stage5_7[2],stage5_6[3],stage5_5[4],stage5_4[5]}
   );
   gpc606_5 gpc9292 (
      {stage4_4[16], stage4_4[17], stage4_4[18], stage4_4[19], stage4_4[20], stage4_4[21]},
      {stage4_6[13], stage4_6[14], stage4_6[15], stage4_6[16], stage4_6[17], stage4_6[18]},
      {stage5_8[3],stage5_7[3],stage5_6[4],stage5_5[5],stage5_4[6]}
   );
   gpc606_5 gpc9293 (
      {stage4_4[22], stage4_4[23], stage4_4[24], stage4_4[25], stage4_4[26], stage4_4[27]},
      {stage4_6[19], stage4_6[20], stage4_6[21], stage4_6[22], stage4_6[23], 1'b0},
      {stage5_8[4],stage5_7[4],stage5_6[5],stage5_5[6],stage5_4[7]}
   );
   gpc606_5 gpc9294 (
      {stage4_5[7], stage4_5[8], stage4_5[9], stage4_5[10], stage4_5[11], stage4_5[12]},
      {stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5], stage4_7[6]},
      {stage5_9[0],stage5_8[5],stage5_7[5],stage5_6[6],stage5_5[7]}
   );
   gpc606_5 gpc9295 (
      {stage4_5[13], stage4_5[14], stage4_5[15], stage4_5[16], stage4_5[17], stage4_5[18]},
      {stage4_7[7], stage4_7[8], stage4_7[9], stage4_7[10], stage4_7[11], stage4_7[12]},
      {stage5_9[1],stage5_8[6],stage5_7[6],stage5_6[7],stage5_5[8]}
   );
   gpc606_5 gpc9296 (
      {stage4_5[19], stage4_5[20], stage4_5[21], stage4_5[22], stage4_5[23], stage4_5[24]},
      {stage4_7[13], stage4_7[14], stage4_7[15], stage4_7[16], stage4_7[17], stage4_7[18]},
      {stage5_9[2],stage5_8[7],stage5_7[7],stage5_6[8],stage5_5[9]}
   );
   gpc606_5 gpc9297 (
      {stage4_5[25], stage4_5[26], stage4_5[27], stage4_5[28], stage4_5[29], stage4_5[30]},
      {stage4_7[19], stage4_7[20], stage4_7[21], stage4_7[22], stage4_7[23], stage4_7[24]},
      {stage5_9[3],stage5_8[8],stage5_7[8],stage5_6[9],stage5_5[10]}
   );
   gpc207_4 gpc9298 (
      {stage4_7[25], stage4_7[26], stage4_7[27], stage4_7[28], stage4_7[29], stage4_7[30], stage4_7[31]},
      {stage4_9[0], stage4_9[1]},
      {stage5_10[0],stage5_9[4],stage5_8[9],stage5_7[9]}
   );
   gpc207_4 gpc9299 (
      {stage4_7[32], stage4_7[33], stage4_7[34], stage4_7[35], stage4_7[36], stage4_7[37], stage4_7[38]},
      {stage4_9[2], stage4_9[3]},
      {stage5_10[1],stage5_9[5],stage5_8[10],stage5_7[10]}
   );
   gpc135_4 gpc9300 (
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4]},
      {stage4_9[4], stage4_9[5], stage4_9[6]},
      {stage4_10[0]},
      {stage5_11[0],stage5_10[2],stage5_9[6],stage5_8[11]}
   );
   gpc117_4 gpc9301 (
      {stage4_8[5], stage4_8[6], stage4_8[7], stage4_8[8], stage4_8[9], stage4_8[10], stage4_8[11]},
      {stage4_9[7]},
      {stage4_10[1]},
      {stage5_11[1],stage5_10[3],stage5_9[7],stage5_8[12]}
   );
   gpc606_5 gpc9302 (
      {stage4_8[12], stage4_8[13], stage4_8[14], stage4_8[15], stage4_8[16], stage4_8[17]},
      {stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5], stage4_10[6], stage4_10[7]},
      {stage5_12[0],stage5_11[2],stage5_10[4],stage5_9[8],stage5_8[13]}
   );
   gpc606_5 gpc9303 (
      {stage4_8[18], stage4_8[19], stage4_8[20], stage4_8[21], stage4_8[22], stage4_8[23]},
      {stage4_10[8], stage4_10[9], stage4_10[10], stage4_10[11], stage4_10[12], stage4_10[13]},
      {stage5_12[1],stage5_11[3],stage5_10[5],stage5_9[9],stage5_8[14]}
   );
   gpc606_5 gpc9304 (
      {stage4_9[8], stage4_9[9], stage4_9[10], stage4_9[11], stage4_9[12], stage4_9[13]},
      {stage4_11[0], stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5]},
      {stage5_13[0],stage5_12[2],stage5_11[4],stage5_10[6],stage5_9[10]}
   );
   gpc2135_5 gpc9305 (
      {stage4_10[14], stage4_10[15], stage4_10[16], stage4_10[17], stage4_10[18]},
      {stage4_11[6], stage4_11[7], stage4_11[8]},
      {stage4_12[0]},
      {stage4_13[0], stage4_13[1]},
      {stage5_14[0],stage5_13[1],stage5_12[3],stage5_11[5],stage5_10[7]}
   );
   gpc606_5 gpc9306 (
      {stage4_10[19], stage4_10[20], stage4_10[21], stage4_10[22], stage4_10[23], stage4_10[24]},
      {stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5], stage4_12[6]},
      {stage5_14[1],stage5_13[2],stage5_12[4],stage5_11[6],stage5_10[8]}
   );
   gpc606_5 gpc9307 (
      {stage4_10[25], stage4_10[26], stage4_10[27], stage4_10[28], stage4_10[29], stage4_10[30]},
      {stage4_12[7], stage4_12[8], stage4_12[9], stage4_12[10], stage4_12[11], stage4_12[12]},
      {stage5_14[2],stage5_13[3],stage5_12[5],stage5_11[7],stage5_10[9]}
   );
   gpc615_5 gpc9308 (
      {stage4_11[9], stage4_11[10], stage4_11[11], stage4_11[12], stage4_11[13]},
      {stage4_12[13]},
      {stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5], stage4_13[6], stage4_13[7]},
      {stage5_15[0],stage5_14[3],stage5_13[4],stage5_12[6],stage5_11[8]}
   );
   gpc615_5 gpc9309 (
      {stage4_11[14], stage4_11[15], stage4_11[16], stage4_11[17], stage4_11[18]},
      {stage4_12[14]},
      {stage4_13[8], stage4_13[9], stage4_13[10], stage4_13[11], stage4_13[12], stage4_13[13]},
      {stage5_15[1],stage5_14[4],stage5_13[5],stage5_12[7],stage5_11[9]}
   );
   gpc615_5 gpc9310 (
      {stage4_11[19], stage4_11[20], stage4_11[21], stage4_11[22], stage4_11[23]},
      {stage4_12[15]},
      {stage4_13[14], stage4_13[15], stage4_13[16], stage4_13[17], stage4_13[18], stage4_13[19]},
      {stage5_15[2],stage5_14[5],stage5_13[6],stage5_12[8],stage5_11[10]}
   );
   gpc623_5 gpc9311 (
      {stage4_11[24], stage4_11[25], stage4_11[26]},
      {stage4_12[16], stage4_12[17]},
      {stage4_13[20], stage4_13[21], stage4_13[22], stage4_13[23], stage4_13[24], stage4_13[25]},
      {stage5_15[3],stage5_14[6],stage5_13[7],stage5_12[9],stage5_11[11]}
   );
   gpc606_5 gpc9312 (
      {stage4_12[18], stage4_12[19], stage4_12[20], stage4_12[21], stage4_12[22], stage4_12[23]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[4],stage5_14[7],stage5_13[8],stage5_12[10]}
   );
   gpc615_5 gpc9313 (
      {stage4_14[6], stage4_14[7], stage4_14[8], stage4_14[9], stage4_14[10]},
      {stage4_15[0]},
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage5_18[0],stage5_17[0],stage5_16[1],stage5_15[5],stage5_14[8]}
   );
   gpc615_5 gpc9314 (
      {stage4_14[11], stage4_14[12], stage4_14[13], stage4_14[14], stage4_14[15]},
      {stage4_15[1]},
      {stage4_16[6], stage4_16[7], stage4_16[8], stage4_16[9], stage4_16[10], stage4_16[11]},
      {stage5_18[1],stage5_17[1],stage5_16[2],stage5_15[6],stage5_14[9]}
   );
   gpc615_5 gpc9315 (
      {stage4_14[16], stage4_14[17], stage4_14[18], stage4_14[19], stage4_14[20]},
      {stage4_15[2]},
      {stage4_16[12], stage4_16[13], stage4_16[14], stage4_16[15], stage4_16[16], stage4_16[17]},
      {stage5_18[2],stage5_17[2],stage5_16[3],stage5_15[7],stage5_14[10]}
   );
   gpc615_5 gpc9316 (
      {stage4_14[21], stage4_14[22], stage4_14[23], stage4_14[24], stage4_14[25]},
      {stage4_15[3]},
      {stage4_16[18], stage4_16[19], stage4_16[20], stage4_16[21], stage4_16[22], stage4_16[23]},
      {stage5_18[3],stage5_17[3],stage5_16[4],stage5_15[8],stage5_14[11]}
   );
   gpc615_5 gpc9317 (
      {stage4_15[4], stage4_15[5], stage4_15[6], stage4_15[7], stage4_15[8]},
      {stage4_16[24]},
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage5_19[0],stage5_18[4],stage5_17[4],stage5_16[5],stage5_15[9]}
   );
   gpc615_5 gpc9318 (
      {stage4_15[9], stage4_15[10], stage4_15[11], stage4_15[12], stage4_15[13]},
      {stage4_16[25]},
      {stage4_17[6], stage4_17[7], stage4_17[8], stage4_17[9], stage4_17[10], stage4_17[11]},
      {stage5_19[1],stage5_18[5],stage5_17[5],stage5_16[6],stage5_15[10]}
   );
   gpc615_5 gpc9319 (
      {stage4_15[14], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage4_16[26]},
      {stage4_17[12], stage4_17[13], stage4_17[14], stage4_17[15], stage4_17[16], stage4_17[17]},
      {stage5_19[2],stage5_18[6],stage5_17[6],stage5_16[7],stage5_15[11]}
   );
   gpc615_5 gpc9320 (
      {stage4_18[0], stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4]},
      {stage4_19[0]},
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], stage4_20[4], stage4_20[5]},
      {stage5_22[0],stage5_21[0],stage5_20[0],stage5_19[3],stage5_18[7]}
   );
   gpc615_5 gpc9321 (
      {stage4_18[5], stage4_18[6], stage4_18[7], stage4_18[8], stage4_18[9]},
      {stage4_19[1]},
      {stage4_20[6], stage4_20[7], stage4_20[8], stage4_20[9], stage4_20[10], stage4_20[11]},
      {stage5_22[1],stage5_21[1],stage5_20[1],stage5_19[4],stage5_18[8]}
   );
   gpc615_5 gpc9322 (
      {stage4_18[10], stage4_18[11], stage4_18[12], stage4_18[13], stage4_18[14]},
      {stage4_19[2]},
      {stage4_20[12], stage4_20[13], stage4_20[14], stage4_20[15], stage4_20[16], stage4_20[17]},
      {stage5_22[2],stage5_21[2],stage5_20[2],stage5_19[5],stage5_18[9]}
   );
   gpc615_5 gpc9323 (
      {stage4_18[15], stage4_18[16], stage4_18[17], stage4_18[18], stage4_18[19]},
      {stage4_19[3]},
      {stage4_20[18], stage4_20[19], stage4_20[20], stage4_20[21], stage4_20[22], stage4_20[23]},
      {stage5_22[3],stage5_21[3],stage5_20[3],stage5_19[6],stage5_18[10]}
   );
   gpc615_5 gpc9324 (
      {stage4_19[4], stage4_19[5], stage4_19[6], stage4_19[7], stage4_19[8]},
      {stage4_20[24]},
      {stage4_21[0], stage4_21[1], stage4_21[2], stage4_21[3], stage4_21[4], stage4_21[5]},
      {stage5_23[0],stage5_22[4],stage5_21[4],stage5_20[4],stage5_19[7]}
   );
   gpc615_5 gpc9325 (
      {stage4_19[9], stage4_19[10], stage4_19[11], stage4_19[12], stage4_19[13]},
      {stage4_20[25]},
      {stage4_21[6], stage4_21[7], stage4_21[8], stage4_21[9], stage4_21[10], stage4_21[11]},
      {stage5_23[1],stage5_22[5],stage5_21[5],stage5_20[5],stage5_19[8]}
   );
   gpc615_5 gpc9326 (
      {stage4_19[14], stage4_19[15], stage4_19[16], stage4_19[17], stage4_19[18]},
      {stage4_20[26]},
      {stage4_21[12], stage4_21[13], stage4_21[14], stage4_21[15], stage4_21[16], stage4_21[17]},
      {stage5_23[2],stage5_22[6],stage5_21[6],stage5_20[6],stage5_19[9]}
   );
   gpc615_5 gpc9327 (
      {stage4_19[19], stage4_19[20], stage4_19[21], stage4_19[22], stage4_19[23]},
      {stage4_20[27]},
      {stage4_21[18], stage4_21[19], stage4_21[20], stage4_21[21], stage4_21[22], stage4_21[23]},
      {stage5_23[3],stage5_22[7],stage5_21[7],stage5_20[7],stage5_19[10]}
   );
   gpc606_5 gpc9328 (
      {stage4_21[24], stage4_21[25], stage4_21[26], stage4_21[27], stage4_21[28], stage4_21[29]},
      {stage4_23[0], stage4_23[1], stage4_23[2], stage4_23[3], stage4_23[4], stage4_23[5]},
      {stage5_25[0],stage5_24[0],stage5_23[4],stage5_22[8],stage5_21[8]}
   );
   gpc606_5 gpc9329 (
      {stage4_21[30], stage4_21[31], stage4_21[32], stage4_21[33], stage4_21[34], stage4_21[35]},
      {stage4_23[6], stage4_23[7], stage4_23[8], stage4_23[9], stage4_23[10], stage4_23[11]},
      {stage5_25[1],stage5_24[1],stage5_23[5],stage5_22[9],stage5_21[9]}
   );
   gpc1163_5 gpc9330 (
      {stage4_22[0], stage4_22[1], stage4_22[2]},
      {stage4_23[12], stage4_23[13], stage4_23[14], stage4_23[15], stage4_23[16], stage4_23[17]},
      {stage4_24[0]},
      {stage4_25[0]},
      {stage5_26[0],stage5_25[2],stage5_24[2],stage5_23[6],stage5_22[10]}
   );
   gpc615_5 gpc9331 (
      {stage4_22[3], stage4_22[4], stage4_22[5], stage4_22[6], stage4_22[7]},
      {stage4_23[18]},
      {stage4_24[1], stage4_24[2], stage4_24[3], stage4_24[4], stage4_24[5], stage4_24[6]},
      {stage5_26[1],stage5_25[3],stage5_24[3],stage5_23[7],stage5_22[11]}
   );
   gpc615_5 gpc9332 (
      {stage4_22[8], stage4_22[9], stage4_22[10], stage4_22[11], stage4_22[12]},
      {stage4_23[19]},
      {stage4_24[7], stage4_24[8], stage4_24[9], stage4_24[10], stage4_24[11], stage4_24[12]},
      {stage5_26[2],stage5_25[4],stage5_24[4],stage5_23[8],stage5_22[12]}
   );
   gpc615_5 gpc9333 (
      {stage4_22[13], stage4_22[14], stage4_22[15], stage4_22[16], stage4_22[17]},
      {stage4_23[20]},
      {stage4_24[13], stage4_24[14], stage4_24[15], stage4_24[16], stage4_24[17], stage4_24[18]},
      {stage5_26[3],stage5_25[5],stage5_24[5],stage5_23[9],stage5_22[13]}
   );
   gpc606_5 gpc9334 (
      {stage4_25[1], stage4_25[2], stage4_25[3], stage4_25[4], stage4_25[5], stage4_25[6]},
      {stage4_27[0], stage4_27[1], stage4_27[2], stage4_27[3], stage4_27[4], stage4_27[5]},
      {stage5_29[0],stage5_28[0],stage5_27[0],stage5_26[4],stage5_25[6]}
   );
   gpc606_5 gpc9335 (
      {stage4_25[7], stage4_25[8], stage4_25[9], stage4_25[10], stage4_25[11], stage4_25[12]},
      {stage4_27[6], stage4_27[7], stage4_27[8], stage4_27[9], stage4_27[10], stage4_27[11]},
      {stage5_29[1],stage5_28[1],stage5_27[1],stage5_26[5],stage5_25[7]}
   );
   gpc606_5 gpc9336 (
      {stage4_25[13], stage4_25[14], stage4_25[15], stage4_25[16], stage4_25[17], stage4_25[18]},
      {stage4_27[12], stage4_27[13], stage4_27[14], stage4_27[15], stage4_27[16], stage4_27[17]},
      {stage5_29[2],stage5_28[2],stage5_27[2],stage5_26[6],stage5_25[8]}
   );
   gpc623_5 gpc9337 (
      {stage4_25[19], stage4_25[20], 1'b0},
      {stage4_26[0], stage4_26[1]},
      {stage4_27[18], stage4_27[19], stage4_27[20], stage4_27[21], stage4_27[22], stage4_27[23]},
      {stage5_29[3],stage5_28[3],stage5_27[3],stage5_26[7],stage5_25[9]}
   );
   gpc2135_5 gpc9338 (
      {stage4_26[2], stage4_26[3], stage4_26[4], stage4_26[5], stage4_26[6]},
      {stage4_27[24], stage4_27[25], stage4_27[26]},
      {stage4_28[0]},
      {stage4_29[0], stage4_29[1]},
      {stage5_30[0],stage5_29[4],stage5_28[4],stage5_27[4],stage5_26[8]}
   );
   gpc117_4 gpc9339 (
      {stage4_26[7], stage4_26[8], stage4_26[9], stage4_26[10], stage4_26[11], stage4_26[12], stage4_26[13]},
      {1'b0},
      {stage4_28[1]},
      {stage5_29[5],stage5_28[5],stage5_27[5],stage5_26[9]}
   );
   gpc606_5 gpc9340 (
      {stage4_28[2], stage4_28[3], stage4_28[4], stage4_28[5], stage4_28[6], stage4_28[7]},
      {stage4_30[0], stage4_30[1], stage4_30[2], stage4_30[3], stage4_30[4], stage4_30[5]},
      {stage5_32[0],stage5_31[0],stage5_30[1],stage5_29[6],stage5_28[6]}
   );
   gpc615_5 gpc9341 (
      {stage4_28[8], stage4_28[9], stage4_28[10], stage4_28[11], stage4_28[12]},
      {stage4_29[2]},
      {stage4_30[6], stage4_30[7], stage4_30[8], stage4_30[9], stage4_30[10], stage4_30[11]},
      {stage5_32[1],stage5_31[1],stage5_30[2],stage5_29[7],stage5_28[7]}
   );
   gpc615_5 gpc9342 (
      {stage4_28[13], stage4_28[14], stage4_28[15], stage4_28[16], stage4_28[17]},
      {stage4_29[3]},
      {stage4_30[12], stage4_30[13], stage4_30[14], stage4_30[15], stage4_30[16], stage4_30[17]},
      {stage5_32[2],stage5_31[2],stage5_30[3],stage5_29[8],stage5_28[8]}
   );
   gpc117_4 gpc9343 (
      {stage4_29[4], stage4_29[5], stage4_29[6], stage4_29[7], stage4_29[8], stage4_29[9], stage4_29[10]},
      {stage4_30[18]},
      {stage4_31[0]},
      {stage5_32[3],stage5_31[3],stage5_30[4],stage5_29[9]}
   );
   gpc117_4 gpc9344 (
      {stage4_29[11], stage4_29[12], stage4_29[13], stage4_29[14], stage4_29[15], stage4_29[16], stage4_29[17]},
      {stage4_30[19]},
      {stage4_31[1]},
      {stage5_32[4],stage5_31[4],stage5_30[5],stage5_29[10]}
   );
   gpc615_5 gpc9345 (
      {stage4_30[20], stage4_30[21], stage4_30[22], stage4_30[23], stage4_30[24]},
      {stage4_31[2]},
      {stage4_32[0], stage4_32[1], stage4_32[2], stage4_32[3], stage4_32[4], stage4_32[5]},
      {stage5_34[0],stage5_33[0],stage5_32[5],stage5_31[5],stage5_30[6]}
   );
   gpc615_5 gpc9346 (
      {stage4_30[25], stage4_30[26], stage4_30[27], stage4_30[28], stage4_30[29]},
      {stage4_31[3]},
      {stage4_32[6], stage4_32[7], stage4_32[8], stage4_32[9], stage4_32[10], stage4_32[11]},
      {stage5_34[1],stage5_33[1],stage5_32[6],stage5_31[6],stage5_30[7]}
   );
   gpc615_5 gpc9347 (
      {stage4_30[30], stage4_30[31], stage4_30[32], 1'b0, 1'b0},
      {stage4_31[4]},
      {stage4_32[12], stage4_32[13], stage4_32[14], stage4_32[15], stage4_32[16], stage4_32[17]},
      {stage5_34[2],stage5_33[2],stage5_32[7],stage5_31[7],stage5_30[8]}
   );
   gpc615_5 gpc9348 (
      {stage4_31[5], stage4_31[6], stage4_31[7], stage4_31[8], stage4_31[9]},
      {stage4_32[18]},
      {stage4_33[0], stage4_33[1], stage4_33[2], stage4_33[3], stage4_33[4], stage4_33[5]},
      {stage5_35[0],stage5_34[3],stage5_33[3],stage5_32[8],stage5_31[8]}
   );
   gpc615_5 gpc9349 (
      {stage4_31[10], stage4_31[11], stage4_31[12], stage4_31[13], stage4_31[14]},
      {stage4_32[19]},
      {stage4_33[6], stage4_33[7], stage4_33[8], stage4_33[9], stage4_33[10], stage4_33[11]},
      {stage5_35[1],stage5_34[4],stage5_33[4],stage5_32[9],stage5_31[9]}
   );
   gpc606_5 gpc9350 (
      {stage4_33[12], stage4_33[13], stage4_33[14], stage4_33[15], stage4_33[16], stage4_33[17]},
      {stage4_35[0], stage4_35[1], stage4_35[2], stage4_35[3], stage4_35[4], stage4_35[5]},
      {stage5_37[0],stage5_36[0],stage5_35[2],stage5_34[5],stage5_33[5]}
   );
   gpc606_5 gpc9351 (
      {stage4_33[18], stage4_33[19], stage4_33[20], stage4_33[21], stage4_33[22], stage4_33[23]},
      {stage4_35[6], stage4_35[7], stage4_35[8], stage4_35[9], stage4_35[10], stage4_35[11]},
      {stage5_37[1],stage5_36[1],stage5_35[3],stage5_34[6],stage5_33[6]}
   );
   gpc135_4 gpc9352 (
      {stage4_34[0], stage4_34[1], stage4_34[2], stage4_34[3], stage4_34[4]},
      {stage4_35[12], stage4_35[13], stage4_35[14]},
      {stage4_36[0]},
      {stage5_37[2],stage5_36[2],stage5_35[4],stage5_34[7]}
   );
   gpc615_5 gpc9353 (
      {stage4_34[5], stage4_34[6], stage4_34[7], stage4_34[8], stage4_34[9]},
      {stage4_35[15]},
      {stage4_36[1], stage4_36[2], stage4_36[3], stage4_36[4], stage4_36[5], stage4_36[6]},
      {stage5_38[0],stage5_37[3],stage5_36[3],stage5_35[5],stage5_34[8]}
   );
   gpc615_5 gpc9354 (
      {stage4_34[10], stage4_34[11], stage4_34[12], stage4_34[13], stage4_34[14]},
      {stage4_35[16]},
      {stage4_36[7], stage4_36[8], stage4_36[9], stage4_36[10], stage4_36[11], stage4_36[12]},
      {stage5_38[1],stage5_37[4],stage5_36[4],stage5_35[6],stage5_34[9]}
   );
   gpc615_5 gpc9355 (
      {stage4_35[17], stage4_35[18], stage4_35[19], stage4_35[20], stage4_35[21]},
      {stage4_36[13]},
      {stage4_37[0], stage4_37[1], stage4_37[2], stage4_37[3], stage4_37[4], stage4_37[5]},
      {stage5_39[0],stage5_38[2],stage5_37[5],stage5_36[5],stage5_35[7]}
   );
   gpc615_5 gpc9356 (
      {stage4_35[22], stage4_35[23], stage4_35[24], stage4_35[25], stage4_35[26]},
      {stage4_36[14]},
      {stage4_37[6], stage4_37[7], stage4_37[8], stage4_37[9], stage4_37[10], stage4_37[11]},
      {stage5_39[1],stage5_38[3],stage5_37[6],stage5_36[6],stage5_35[8]}
   );
   gpc615_5 gpc9357 (
      {stage4_35[27], stage4_35[28], stage4_35[29], stage4_35[30], stage4_35[31]},
      {stage4_36[15]},
      {stage4_37[12], stage4_37[13], stage4_37[14], stage4_37[15], stage4_37[16], stage4_37[17]},
      {stage5_39[2],stage5_38[4],stage5_37[7],stage5_36[7],stage5_35[9]}
   );
   gpc606_5 gpc9358 (
      {stage4_36[16], stage4_36[17], stage4_36[18], stage4_36[19], stage4_36[20], stage4_36[21]},
      {stage4_38[0], stage4_38[1], stage4_38[2], stage4_38[3], stage4_38[4], stage4_38[5]},
      {stage5_40[0],stage5_39[3],stage5_38[5],stage5_37[8],stage5_36[8]}
   );
   gpc606_5 gpc9359 (
      {stage4_36[22], stage4_36[23], stage4_36[24], stage4_36[25], stage4_36[26], stage4_36[27]},
      {stage4_38[6], stage4_38[7], stage4_38[8], stage4_38[9], stage4_38[10], stage4_38[11]},
      {stage5_40[1],stage5_39[4],stage5_38[6],stage5_37[9],stage5_36[9]}
   );
   gpc606_5 gpc9360 (
      {stage4_36[28], stage4_36[29], stage4_36[30], stage4_36[31], stage4_36[32], stage4_36[33]},
      {stage4_38[12], stage4_38[13], stage4_38[14], stage4_38[15], stage4_38[16], stage4_38[17]},
      {stage5_40[2],stage5_39[5],stage5_38[7],stage5_37[10],stage5_36[10]}
   );
   gpc117_4 gpc9361 (
      {stage4_39[0], stage4_39[1], stage4_39[2], stage4_39[3], stage4_39[4], stage4_39[5], stage4_39[6]},
      {stage4_40[0]},
      {stage4_41[0]},
      {stage5_42[0],stage5_41[0],stage5_40[3],stage5_39[6]}
   );
   gpc117_4 gpc9362 (
      {stage4_39[7], stage4_39[8], stage4_39[9], stage4_39[10], stage4_39[11], stage4_39[12], stage4_39[13]},
      {stage4_40[1]},
      {stage4_41[1]},
      {stage5_42[1],stage5_41[1],stage5_40[4],stage5_39[7]}
   );
   gpc615_5 gpc9363 (
      {stage4_39[14], stage4_39[15], stage4_39[16], stage4_39[17], stage4_39[18]},
      {stage4_40[2]},
      {stage4_41[2], stage4_41[3], stage4_41[4], stage4_41[5], stage4_41[6], stage4_41[7]},
      {stage5_43[0],stage5_42[2],stage5_41[2],stage5_40[5],stage5_39[8]}
   );
   gpc615_5 gpc9364 (
      {stage4_39[19], stage4_39[20], stage4_39[21], stage4_39[22], stage4_39[23]},
      {stage4_40[3]},
      {stage4_41[8], stage4_41[9], stage4_41[10], stage4_41[11], stage4_41[12], stage4_41[13]},
      {stage5_43[1],stage5_42[3],stage5_41[3],stage5_40[6],stage5_39[9]}
   );
   gpc606_5 gpc9365 (
      {stage4_40[4], stage4_40[5], stage4_40[6], stage4_40[7], stage4_40[8], stage4_40[9]},
      {stage4_42[0], stage4_42[1], stage4_42[2], stage4_42[3], stage4_42[4], stage4_42[5]},
      {stage5_44[0],stage5_43[2],stage5_42[4],stage5_41[4],stage5_40[7]}
   );
   gpc606_5 gpc9366 (
      {stage4_40[10], stage4_40[11], stage4_40[12], stage4_40[13], stage4_40[14], stage4_40[15]},
      {stage4_42[6], stage4_42[7], stage4_42[8], stage4_42[9], stage4_42[10], stage4_42[11]},
      {stage5_44[1],stage5_43[3],stage5_42[5],stage5_41[5],stage5_40[8]}
   );
   gpc606_5 gpc9367 (
      {stage4_40[16], stage4_40[17], stage4_40[18], stage4_40[19], stage4_40[20], stage4_40[21]},
      {stage4_42[12], stage4_42[13], stage4_42[14], stage4_42[15], stage4_42[16], stage4_42[17]},
      {stage5_44[2],stage5_43[4],stage5_42[6],stage5_41[6],stage5_40[9]}
   );
   gpc606_5 gpc9368 (
      {stage4_40[22], stage4_40[23], stage4_40[24], stage4_40[25], stage4_40[26], stage4_40[27]},
      {stage4_42[18], stage4_42[19], stage4_42[20], stage4_42[21], stage4_42[22], stage4_42[23]},
      {stage5_44[3],stage5_43[5],stage5_42[7],stage5_41[7],stage5_40[10]}
   );
   gpc606_5 gpc9369 (
      {stage4_41[14], stage4_41[15], stage4_41[16], stage4_41[17], stage4_41[18], stage4_41[19]},
      {stage4_43[0], stage4_43[1], stage4_43[2], stage4_43[3], stage4_43[4], stage4_43[5]},
      {stage5_45[0],stage5_44[4],stage5_43[6],stage5_42[8],stage5_41[8]}
   );
   gpc615_5 gpc9370 (
      {stage4_42[24], stage4_42[25], stage4_42[26], stage4_42[27], stage4_42[28]},
      {stage4_43[6]},
      {stage4_44[0], stage4_44[1], stage4_44[2], stage4_44[3], stage4_44[4], stage4_44[5]},
      {stage5_46[0],stage5_45[1],stage5_44[5],stage5_43[7],stage5_42[9]}
   );
   gpc615_5 gpc9371 (
      {stage4_43[7], stage4_43[8], stage4_43[9], stage4_43[10], stage4_43[11]},
      {stage4_44[6]},
      {stage4_45[0], stage4_45[1], stage4_45[2], stage4_45[3], stage4_45[4], stage4_45[5]},
      {stage5_47[0],stage5_46[1],stage5_45[2],stage5_44[6],stage5_43[8]}
   );
   gpc135_4 gpc9372 (
      {stage4_44[7], stage4_44[8], stage4_44[9], stage4_44[10], stage4_44[11]},
      {stage4_45[6], stage4_45[7], stage4_45[8]},
      {stage4_46[0]},
      {stage5_47[1],stage5_46[2],stage5_45[3],stage5_44[7]}
   );
   gpc135_4 gpc9373 (
      {stage4_44[12], stage4_44[13], stage4_44[14], stage4_44[15], stage4_44[16]},
      {stage4_45[9], stage4_45[10], stage4_45[11]},
      {stage4_46[1]},
      {stage5_47[2],stage5_46[3],stage5_45[4],stage5_44[8]}
   );
   gpc135_4 gpc9374 (
      {stage4_44[17], stage4_44[18], stage4_44[19], stage4_44[20], stage4_44[21]},
      {stage4_45[12], stage4_45[13], stage4_45[14]},
      {stage4_46[2]},
      {stage5_47[3],stage5_46[4],stage5_45[5],stage5_44[9]}
   );
   gpc606_5 gpc9375 (
      {stage4_45[15], stage4_45[16], stage4_45[17], stage4_45[18], stage4_45[19], stage4_45[20]},
      {stage4_47[0], stage4_47[1], stage4_47[2], stage4_47[3], stage4_47[4], stage4_47[5]},
      {stage5_49[0],stage5_48[0],stage5_47[4],stage5_46[5],stage5_45[6]}
   );
   gpc615_5 gpc9376 (
      {stage4_46[3], stage4_46[4], stage4_46[5], stage4_46[6], stage4_46[7]},
      {stage4_47[6]},
      {stage4_48[0], stage4_48[1], stage4_48[2], stage4_48[3], stage4_48[4], stage4_48[5]},
      {stage5_50[0],stage5_49[1],stage5_48[1],stage5_47[5],stage5_46[6]}
   );
   gpc615_5 gpc9377 (
      {stage4_46[8], stage4_46[9], stage4_46[10], stage4_46[11], stage4_46[12]},
      {stage4_47[7]},
      {stage4_48[6], stage4_48[7], stage4_48[8], stage4_48[9], stage4_48[10], stage4_48[11]},
      {stage5_50[1],stage5_49[2],stage5_48[2],stage5_47[6],stage5_46[7]}
   );
   gpc615_5 gpc9378 (
      {stage4_47[8], stage4_47[9], stage4_47[10], stage4_47[11], stage4_47[12]},
      {stage4_48[12]},
      {stage4_49[0], stage4_49[1], stage4_49[2], stage4_49[3], stage4_49[4], stage4_49[5]},
      {stage5_51[0],stage5_50[2],stage5_49[3],stage5_48[3],stage5_47[7]}
   );
   gpc615_5 gpc9379 (
      {stage4_47[13], stage4_47[14], stage4_47[15], stage4_47[16], stage4_47[17]},
      {stage4_48[13]},
      {stage4_49[6], stage4_49[7], stage4_49[8], stage4_49[9], stage4_49[10], stage4_49[11]},
      {stage5_51[1],stage5_50[3],stage5_49[4],stage5_48[4],stage5_47[8]}
   );
   gpc7_3 gpc9380 (
      {stage4_50[0], stage4_50[1], stage4_50[2], stage4_50[3], stage4_50[4], stage4_50[5], stage4_50[6]},
      {stage5_52[0],stage5_51[2],stage5_50[4]}
   );
   gpc615_5 gpc9381 (
      {stage4_50[7], stage4_50[8], stage4_50[9], stage4_50[10], stage4_50[11]},
      {stage4_51[0]},
      {stage4_52[0], stage4_52[1], stage4_52[2], stage4_52[3], stage4_52[4], stage4_52[5]},
      {stage5_54[0],stage5_53[0],stage5_52[1],stage5_51[3],stage5_50[5]}
   );
   gpc615_5 gpc9382 (
      {stage4_50[12], stage4_50[13], stage4_50[14], stage4_50[15], stage4_50[16]},
      {stage4_51[1]},
      {stage4_52[6], stage4_52[7], stage4_52[8], stage4_52[9], stage4_52[10], stage4_52[11]},
      {stage5_54[1],stage5_53[1],stage5_52[2],stage5_51[4],stage5_50[6]}
   );
   gpc615_5 gpc9383 (
      {stage4_51[2], stage4_51[3], stage4_51[4], stage4_51[5], stage4_51[6]},
      {stage4_52[12]},
      {stage4_53[0], stage4_53[1], stage4_53[2], stage4_53[3], stage4_53[4], stage4_53[5]},
      {stage5_55[0],stage5_54[2],stage5_53[2],stage5_52[3],stage5_51[5]}
   );
   gpc615_5 gpc9384 (
      {stage4_51[7], stage4_51[8], stage4_51[9], stage4_51[10], stage4_51[11]},
      {stage4_52[13]},
      {stage4_53[6], stage4_53[7], stage4_53[8], stage4_53[9], stage4_53[10], stage4_53[11]},
      {stage5_55[1],stage5_54[3],stage5_53[3],stage5_52[4],stage5_51[6]}
   );
   gpc615_5 gpc9385 (
      {stage4_51[12], stage4_51[13], stage4_51[14], stage4_51[15], stage4_51[16]},
      {stage4_52[14]},
      {stage4_53[12], stage4_53[13], stage4_53[14], stage4_53[15], stage4_53[16], stage4_53[17]},
      {stage5_55[2],stage5_54[4],stage5_53[4],stage5_52[5],stage5_51[7]}
   );
   gpc615_5 gpc9386 (
      {stage4_51[17], stage4_51[18], stage4_51[19], stage4_51[20], stage4_51[21]},
      {stage4_52[15]},
      {stage4_53[18], stage4_53[19], stage4_53[20], stage4_53[21], stage4_53[22], stage4_53[23]},
      {stage5_55[3],stage5_54[5],stage5_53[5],stage5_52[6],stage5_51[8]}
   );
   gpc615_5 gpc9387 (
      {stage4_51[22], stage4_51[23], stage4_51[24], stage4_51[25], stage4_51[26]},
      {stage4_52[16]},
      {stage4_53[24], stage4_53[25], stage4_53[26], stage4_53[27], stage4_53[28], stage4_53[29]},
      {stage5_55[4],stage5_54[6],stage5_53[6],stage5_52[7],stage5_51[9]}
   );
   gpc615_5 gpc9388 (
      {stage4_53[30], stage4_53[31], stage4_53[32], stage4_53[33], stage4_53[34]},
      {stage4_54[0]},
      {stage4_55[0], stage4_55[1], stage4_55[2], stage4_55[3], stage4_55[4], stage4_55[5]},
      {stage5_57[0],stage5_56[0],stage5_55[5],stage5_54[7],stage5_53[7]}
   );
   gpc615_5 gpc9389 (
      {stage4_53[35], stage4_53[36], stage4_53[37], stage4_53[38], stage4_53[39]},
      {stage4_54[1]},
      {stage4_55[6], stage4_55[7], stage4_55[8], stage4_55[9], stage4_55[10], stage4_55[11]},
      {stage5_57[1],stage5_56[1],stage5_55[6],stage5_54[8],stage5_53[8]}
   );
   gpc2135_5 gpc9390 (
      {stage4_54[2], stage4_54[3], stage4_54[4], stage4_54[5], stage4_54[6]},
      {stage4_55[12], stage4_55[13], stage4_55[14]},
      {stage4_56[0]},
      {stage4_57[0], stage4_57[1]},
      {stage5_58[0],stage5_57[2],stage5_56[2],stage5_55[7],stage5_54[9]}
   );
   gpc2135_5 gpc9391 (
      {stage4_54[7], stage4_54[8], stage4_54[9], stage4_54[10], stage4_54[11]},
      {stage4_55[15], stage4_55[16], stage4_55[17]},
      {stage4_56[1]},
      {stage4_57[2], stage4_57[3]},
      {stage5_58[1],stage5_57[3],stage5_56[3],stage5_55[8],stage5_54[10]}
   );
   gpc2135_5 gpc9392 (
      {stage4_54[12], stage4_54[13], stage4_54[14], stage4_54[15], stage4_54[16]},
      {stage4_55[18], stage4_55[19], stage4_55[20]},
      {stage4_56[2]},
      {stage4_57[4], stage4_57[5]},
      {stage5_58[2],stage5_57[4],stage5_56[4],stage5_55[9],stage5_54[11]}
   );
   gpc2135_5 gpc9393 (
      {stage4_54[17], stage4_54[18], stage4_54[19], stage4_54[20], stage4_54[21]},
      {stage4_55[21], stage4_55[22], stage4_55[23]},
      {stage4_56[3]},
      {stage4_57[6], stage4_57[7]},
      {stage5_58[3],stage5_57[5],stage5_56[5],stage5_55[10],stage5_54[12]}
   );
   gpc615_5 gpc9394 (
      {stage4_55[24], stage4_55[25], stage4_55[26], stage4_55[27], stage4_55[28]},
      {stage4_56[4]},
      {stage4_57[8], stage4_57[9], stage4_57[10], stage4_57[11], stage4_57[12], stage4_57[13]},
      {stage5_59[0],stage5_58[4],stage5_57[6],stage5_56[6],stage5_55[11]}
   );
   gpc606_5 gpc9395 (
      {stage4_56[5], stage4_56[6], stage4_56[7], stage4_56[8], stage4_56[9], stage4_56[10]},
      {stage4_58[0], stage4_58[1], stage4_58[2], stage4_58[3], stage4_58[4], stage4_58[5]},
      {stage5_60[0],stage5_59[1],stage5_58[5],stage5_57[7],stage5_56[7]}
   );
   gpc623_5 gpc9396 (
      {stage4_56[11], stage4_56[12], stage4_56[13]},
      {stage4_57[14], stage4_57[15]},
      {stage4_58[6], stage4_58[7], stage4_58[8], stage4_58[9], stage4_58[10], stage4_58[11]},
      {stage5_60[1],stage5_59[2],stage5_58[6],stage5_57[8],stage5_56[8]}
   );
   gpc606_5 gpc9397 (
      {stage4_57[16], stage4_57[17], stage4_57[18], stage4_57[19], stage4_57[20], stage4_57[21]},
      {stage4_59[0], stage4_59[1], stage4_59[2], stage4_59[3], stage4_59[4], stage4_59[5]},
      {stage5_61[0],stage5_60[2],stage5_59[3],stage5_58[7],stage5_57[9]}
   );
   gpc615_5 gpc9398 (
      {stage4_58[12], stage4_58[13], stage4_58[14], stage4_58[15], stage4_58[16]},
      {stage4_59[6]},
      {stage4_60[0], stage4_60[1], stage4_60[2], stage4_60[3], stage4_60[4], stage4_60[5]},
      {stage5_62[0],stage5_61[1],stage5_60[3],stage5_59[4],stage5_58[8]}
   );
   gpc615_5 gpc9399 (
      {stage4_59[7], stage4_59[8], stage4_59[9], stage4_59[10], stage4_59[11]},
      {stage4_60[6]},
      {stage4_61[0], stage4_61[1], stage4_61[2], stage4_61[3], stage4_61[4], stage4_61[5]},
      {stage5_63[0],stage5_62[1],stage5_61[2],stage5_60[4],stage5_59[5]}
   );
   gpc615_5 gpc9400 (
      {stage4_59[12], stage4_59[13], stage4_59[14], stage4_59[15], stage4_59[16]},
      {stage4_60[7]},
      {stage4_61[6], stage4_61[7], stage4_61[8], stage4_61[9], stage4_61[10], stage4_61[11]},
      {stage5_63[1],stage5_62[2],stage5_61[3],stage5_60[5],stage5_59[6]}
   );
   gpc615_5 gpc9401 (
      {stage4_59[17], stage4_59[18], stage4_59[19], stage4_59[20], 1'b0},
      {stage4_60[8]},
      {stage4_61[12], stage4_61[13], stage4_61[14], stage4_61[15], stage4_61[16], stage4_61[17]},
      {stage5_63[2],stage5_62[3],stage5_61[4],stage5_60[6],stage5_59[7]}
   );
   gpc606_5 gpc9402 (
      {stage4_60[9], stage4_60[10], stage4_60[11], stage4_60[12], stage4_60[13], stage4_60[14]},
      {stage4_62[0], stage4_62[1], stage4_62[2], stage4_62[3], stage4_62[4], stage4_62[5]},
      {stage5_64[0],stage5_63[3],stage5_62[4],stage5_61[5],stage5_60[7]}
   );
   gpc615_5 gpc9403 (
      {stage4_61[18], stage4_61[19], stage4_61[20], stage4_61[21], stage4_61[22]},
      {stage4_62[6]},
      {stage4_63[0], stage4_63[1], stage4_63[2], stage4_63[3], stage4_63[4], stage4_63[5]},
      {stage5_65[0],stage5_64[1],stage5_63[4],stage5_62[5],stage5_61[6]}
   );
   gpc615_5 gpc9404 (
      {stage4_62[7], stage4_62[8], stage4_62[9], stage4_62[10], stage4_62[11]},
      {stage4_63[6]},
      {stage4_64[0], stage4_64[1], stage4_64[2], stage4_64[3], stage4_64[4], stage4_64[5]},
      {stage5_66[0],stage5_65[1],stage5_64[2],stage5_63[5],stage5_62[6]}
   );
   gpc615_5 gpc9405 (
      {stage4_63[7], stage4_63[8], stage4_63[9], stage4_63[10], stage4_63[11]},
      {stage4_64[6]},
      {stage4_65[0], stage4_65[1], stage4_65[2], stage4_65[3], stage4_65[4], stage4_65[5]},
      {stage5_67[0],stage5_66[1],stage5_65[2],stage5_64[3],stage5_63[6]}
   );
   gpc2135_5 gpc9406 (
      {stage4_64[7], stage4_64[8], stage4_64[9], stage4_64[10], stage4_64[11]},
      {stage4_65[6], stage4_65[7], stage4_65[8]},
      {stage4_66[0]},
      {stage4_67[0], stage4_67[1]},
      {stage5_68[0],stage5_67[1],stage5_66[2],stage5_65[3],stage5_64[4]}
   );
   gpc2135_5 gpc9407 (
      {stage4_64[12], stage4_64[13], stage4_64[14], stage4_64[15], stage4_64[16]},
      {stage4_65[9], stage4_65[10], stage4_65[11]},
      {stage4_66[1]},
      {stage4_67[2], stage4_67[3]},
      {stage5_68[1],stage5_67[2],stage5_66[3],stage5_65[4],stage5_64[5]}
   );
   gpc1163_5 gpc9408 (
      {stage4_64[17], stage4_64[18], stage4_64[19]},
      {stage4_65[12], stage4_65[13], stage4_65[14], stage4_65[15], stage4_65[16], stage4_65[17]},
      {stage4_66[2]},
      {stage4_67[4]},
      {stage5_68[2],stage5_67[3],stage5_66[4],stage5_65[5],stage5_64[6]}
   );
   gpc1163_5 gpc9409 (
      {stage4_64[20], stage4_64[21], stage4_64[22]},
      {stage4_65[18], stage4_65[19], stage4_65[20], stage4_65[21], stage4_65[22], stage4_65[23]},
      {stage4_66[3]},
      {stage4_67[5]},
      {stage5_68[3],stage5_67[4],stage5_66[5],stage5_65[6],stage5_64[7]}
   );
   gpc1325_5 gpc9410 (
      {stage4_64[23], stage4_64[24], stage4_64[25], stage4_64[26], stage4_64[27]},
      {stage4_65[24], stage4_65[25]},
      {stage4_66[4], stage4_66[5], stage4_66[6]},
      {stage4_67[6]},
      {stage5_68[4],stage5_67[5],stage5_66[6],stage5_65[7],stage5_64[8]}
   );
   gpc606_5 gpc9411 (
      {stage4_66[7], stage4_66[8], stage4_66[9], stage4_66[10], 1'b0, 1'b0},
      {stage4_68[0], stage4_68[1], stage4_68[2], stage4_68[3], stage4_68[4], stage4_68[5]},
      {stage5_70[0],stage5_69[0],stage5_68[5],stage5_67[6],stage5_66[7]}
   );
   gpc1_1 gpc9412 (
      {stage4_0[5]},
      {stage5_0[1]}
   );
   gpc1_1 gpc9413 (
      {stage4_0[6]},
      {stage5_0[2]}
   );
   gpc1_1 gpc9414 (
      {stage4_0[7]},
      {stage5_0[3]}
   );
   gpc1_1 gpc9415 (
      {stage4_0[8]},
      {stage5_0[4]}
   );
   gpc1_1 gpc9416 (
      {stage4_2[9]},
      {stage5_2[3]}
   );
   gpc1_1 gpc9417 (
      {stage4_2[10]},
      {stage5_2[4]}
   );
   gpc1_1 gpc9418 (
      {stage4_3[12]},
      {stage5_3[3]}
   );
   gpc1_1 gpc9419 (
      {stage4_3[13]},
      {stage5_3[4]}
   );
   gpc1_1 gpc9420 (
      {stage4_3[14]},
      {stage5_3[5]}
   );
   gpc1_1 gpc9421 (
      {stage4_3[15]},
      {stage5_3[6]}
   );
   gpc1_1 gpc9422 (
      {stage4_3[16]},
      {stage5_3[7]}
   );
   gpc1_1 gpc9423 (
      {stage4_4[28]},
      {stage5_4[8]}
   );
   gpc1_1 gpc9424 (
      {stage4_4[29]},
      {stage5_4[9]}
   );
   gpc1_1 gpc9425 (
      {stage4_4[30]},
      {stage5_4[10]}
   );
   gpc1_1 gpc9426 (
      {stage4_5[31]},
      {stage5_5[11]}
   );
   gpc1_1 gpc9427 (
      {stage4_5[32]},
      {stage5_5[12]}
   );
   gpc1_1 gpc9428 (
      {stage4_5[33]},
      {stage5_5[13]}
   );
   gpc1_1 gpc9429 (
      {stage4_5[34]},
      {stage5_5[14]}
   );
   gpc1_1 gpc9430 (
      {stage4_5[35]},
      {stage5_5[15]}
   );
   gpc1_1 gpc9431 (
      {stage4_8[24]},
      {stage5_8[15]}
   );
   gpc1_1 gpc9432 (
      {stage4_8[25]},
      {stage5_8[16]}
   );
   gpc1_1 gpc9433 (
      {stage4_8[26]},
      {stage5_8[17]}
   );
   gpc1_1 gpc9434 (
      {stage4_8[27]},
      {stage5_8[18]}
   );
   gpc1_1 gpc9435 (
      {stage4_10[31]},
      {stage5_10[10]}
   );
   gpc1_1 gpc9436 (
      {stage4_10[32]},
      {stage5_10[11]}
   );
   gpc1_1 gpc9437 (
      {stage4_10[33]},
      {stage5_10[12]}
   );
   gpc1_1 gpc9438 (
      {stage4_10[34]},
      {stage5_10[13]}
   );
   gpc1_1 gpc9439 (
      {stage4_10[35]},
      {stage5_10[14]}
   );
   gpc1_1 gpc9440 (
      {stage4_10[36]},
      {stage5_10[15]}
   );
   gpc1_1 gpc9441 (
      {stage4_10[37]},
      {stage5_10[16]}
   );
   gpc1_1 gpc9442 (
      {stage4_10[38]},
      {stage5_10[17]}
   );
   gpc1_1 gpc9443 (
      {stage4_10[39]},
      {stage5_10[18]}
   );
   gpc1_1 gpc9444 (
      {stage4_10[40]},
      {stage5_10[19]}
   );
   gpc1_1 gpc9445 (
      {stage4_10[41]},
      {stage5_10[20]}
   );
   gpc1_1 gpc9446 (
      {stage4_11[27]},
      {stage5_11[12]}
   );
   gpc1_1 gpc9447 (
      {stage4_11[28]},
      {stage5_11[13]}
   );
   gpc1_1 gpc9448 (
      {stage4_13[26]},
      {stage5_13[9]}
   );
   gpc1_1 gpc9449 (
      {stage4_13[27]},
      {stage5_13[10]}
   );
   gpc1_1 gpc9450 (
      {stage4_13[28]},
      {stage5_13[11]}
   );
   gpc1_1 gpc9451 (
      {stage4_13[29]},
      {stage5_13[12]}
   );
   gpc1_1 gpc9452 (
      {stage4_13[30]},
      {stage5_13[13]}
   );
   gpc1_1 gpc9453 (
      {stage4_13[31]},
      {stage5_13[14]}
   );
   gpc1_1 gpc9454 (
      {stage4_14[26]},
      {stage5_14[12]}
   );
   gpc1_1 gpc9455 (
      {stage4_14[27]},
      {stage5_14[13]}
   );
   gpc1_1 gpc9456 (
      {stage4_14[28]},
      {stage5_14[14]}
   );
   gpc1_1 gpc9457 (
      {stage4_14[29]},
      {stage5_14[15]}
   );
   gpc1_1 gpc9458 (
      {stage4_18[20]},
      {stage5_18[11]}
   );
   gpc1_1 gpc9459 (
      {stage4_19[24]},
      {stage5_19[11]}
   );
   gpc1_1 gpc9460 (
      {stage4_19[25]},
      {stage5_19[12]}
   );
   gpc1_1 gpc9461 (
      {stage4_19[26]},
      {stage5_19[13]}
   );
   gpc1_1 gpc9462 (
      {stage4_19[27]},
      {stage5_19[14]}
   );
   gpc1_1 gpc9463 (
      {stage4_19[28]},
      {stage5_19[15]}
   );
   gpc1_1 gpc9464 (
      {stage4_20[28]},
      {stage5_20[8]}
   );
   gpc1_1 gpc9465 (
      {stage4_20[29]},
      {stage5_20[9]}
   );
   gpc1_1 gpc9466 (
      {stage4_20[30]},
      {stage5_20[10]}
   );
   gpc1_1 gpc9467 (
      {stage4_20[31]},
      {stage5_20[11]}
   );
   gpc1_1 gpc9468 (
      {stage4_20[32]},
      {stage5_20[12]}
   );
   gpc1_1 gpc9469 (
      {stage4_20[33]},
      {stage5_20[13]}
   );
   gpc1_1 gpc9470 (
      {stage4_21[36]},
      {stage5_21[10]}
   );
   gpc1_1 gpc9471 (
      {stage4_24[19]},
      {stage5_24[6]}
   );
   gpc1_1 gpc9472 (
      {stage4_24[20]},
      {stage5_24[7]}
   );
   gpc1_1 gpc9473 (
      {stage4_24[21]},
      {stage5_24[8]}
   );
   gpc1_1 gpc9474 (
      {stage4_26[14]},
      {stage5_26[10]}
   );
   gpc1_1 gpc9475 (
      {stage4_26[15]},
      {stage5_26[11]}
   );
   gpc1_1 gpc9476 (
      {stage4_26[16]},
      {stage5_26[12]}
   );
   gpc1_1 gpc9477 (
      {stage4_26[17]},
      {stage5_26[13]}
   );
   gpc1_1 gpc9478 (
      {stage4_26[18]},
      {stage5_26[14]}
   );
   gpc1_1 gpc9479 (
      {stage4_28[18]},
      {stage5_28[9]}
   );
   gpc1_1 gpc9480 (
      {stage4_29[18]},
      {stage5_29[11]}
   );
   gpc1_1 gpc9481 (
      {stage4_29[19]},
      {stage5_29[12]}
   );
   gpc1_1 gpc9482 (
      {stage4_29[20]},
      {stage5_29[13]}
   );
   gpc1_1 gpc9483 (
      {stage4_29[21]},
      {stage5_29[14]}
   );
   gpc1_1 gpc9484 (
      {stage4_32[20]},
      {stage5_32[10]}
   );
   gpc1_1 gpc9485 (
      {stage4_32[21]},
      {stage5_32[11]}
   );
   gpc1_1 gpc9486 (
      {stage4_32[22]},
      {stage5_32[12]}
   );
   gpc1_1 gpc9487 (
      {stage4_32[23]},
      {stage5_32[13]}
   );
   gpc1_1 gpc9488 (
      {stage4_32[24]},
      {stage5_32[14]}
   );
   gpc1_1 gpc9489 (
      {stage4_32[25]},
      {stage5_32[15]}
   );
   gpc1_1 gpc9490 (
      {stage4_32[26]},
      {stage5_32[16]}
   );
   gpc1_1 gpc9491 (
      {stage4_32[27]},
      {stage5_32[17]}
   );
   gpc1_1 gpc9492 (
      {stage4_32[28]},
      {stage5_32[18]}
   );
   gpc1_1 gpc9493 (
      {stage4_32[29]},
      {stage5_32[19]}
   );
   gpc1_1 gpc9494 (
      {stage4_33[24]},
      {stage5_33[7]}
   );
   gpc1_1 gpc9495 (
      {stage4_33[25]},
      {stage5_33[8]}
   );
   gpc1_1 gpc9496 (
      {stage4_33[26]},
      {stage5_33[9]}
   );
   gpc1_1 gpc9497 (
      {stage4_33[27]},
      {stage5_33[10]}
   );
   gpc1_1 gpc9498 (
      {stage4_33[28]},
      {stage5_33[11]}
   );
   gpc1_1 gpc9499 (
      {stage4_34[15]},
      {stage5_34[10]}
   );
   gpc1_1 gpc9500 (
      {stage4_34[16]},
      {stage5_34[11]}
   );
   gpc1_1 gpc9501 (
      {stage4_34[17]},
      {stage5_34[12]}
   );
   gpc1_1 gpc9502 (
      {stage4_34[18]},
      {stage5_34[13]}
   );
   gpc1_1 gpc9503 (
      {stage4_35[32]},
      {stage5_35[10]}
   );
   gpc1_1 gpc9504 (
      {stage4_35[33]},
      {stage5_35[11]}
   );
   gpc1_1 gpc9505 (
      {stage4_35[34]},
      {stage5_35[12]}
   );
   gpc1_1 gpc9506 (
      {stage4_35[35]},
      {stage5_35[13]}
   );
   gpc1_1 gpc9507 (
      {stage4_36[34]},
      {stage5_36[11]}
   );
   gpc1_1 gpc9508 (
      {stage4_36[35]},
      {stage5_36[12]}
   );
   gpc1_1 gpc9509 (
      {stage4_38[18]},
      {stage5_38[8]}
   );
   gpc1_1 gpc9510 (
      {stage4_38[19]},
      {stage5_38[9]}
   );
   gpc1_1 gpc9511 (
      {stage4_42[29]},
      {stage5_42[10]}
   );
   gpc1_1 gpc9512 (
      {stage4_42[30]},
      {stage5_42[11]}
   );
   gpc1_1 gpc9513 (
      {stage4_42[31]},
      {stage5_42[12]}
   );
   gpc1_1 gpc9514 (
      {stage4_42[32]},
      {stage5_42[13]}
   );
   gpc1_1 gpc9515 (
      {stage4_42[33]},
      {stage5_42[14]}
   );
   gpc1_1 gpc9516 (
      {stage4_42[34]},
      {stage5_42[15]}
   );
   gpc1_1 gpc9517 (
      {stage4_42[35]},
      {stage5_42[16]}
   );
   gpc1_1 gpc9518 (
      {stage4_42[36]},
      {stage5_42[17]}
   );
   gpc1_1 gpc9519 (
      {stage4_42[37]},
      {stage5_42[18]}
   );
   gpc1_1 gpc9520 (
      {stage4_43[12]},
      {stage5_43[9]}
   );
   gpc1_1 gpc9521 (
      {stage4_43[13]},
      {stage5_43[10]}
   );
   gpc1_1 gpc9522 (
      {stage4_44[22]},
      {stage5_44[10]}
   );
   gpc1_1 gpc9523 (
      {stage4_44[23]},
      {stage5_44[11]}
   );
   gpc1_1 gpc9524 (
      {stage4_44[24]},
      {stage5_44[12]}
   );
   gpc1_1 gpc9525 (
      {stage4_45[21]},
      {stage5_45[7]}
   );
   gpc1_1 gpc9526 (
      {stage4_45[22]},
      {stage5_45[8]}
   );
   gpc1_1 gpc9527 (
      {stage4_45[23]},
      {stage5_45[9]}
   );
   gpc1_1 gpc9528 (
      {stage4_45[24]},
      {stage5_45[10]}
   );
   gpc1_1 gpc9529 (
      {stage4_45[25]},
      {stage5_45[11]}
   );
   gpc1_1 gpc9530 (
      {stage4_45[26]},
      {stage5_45[12]}
   );
   gpc1_1 gpc9531 (
      {stage4_45[27]},
      {stage5_45[13]}
   );
   gpc1_1 gpc9532 (
      {stage4_45[28]},
      {stage5_45[14]}
   );
   gpc1_1 gpc9533 (
      {stage4_46[13]},
      {stage5_46[8]}
   );
   gpc1_1 gpc9534 (
      {stage4_46[14]},
      {stage5_46[9]}
   );
   gpc1_1 gpc9535 (
      {stage4_46[15]},
      {stage5_46[10]}
   );
   gpc1_1 gpc9536 (
      {stage4_46[16]},
      {stage5_46[11]}
   );
   gpc1_1 gpc9537 (
      {stage4_47[18]},
      {stage5_47[9]}
   );
   gpc1_1 gpc9538 (
      {stage4_47[19]},
      {stage5_47[10]}
   );
   gpc1_1 gpc9539 (
      {stage4_47[20]},
      {stage5_47[11]}
   );
   gpc1_1 gpc9540 (
      {stage4_48[14]},
      {stage5_48[5]}
   );
   gpc1_1 gpc9541 (
      {stage4_48[15]},
      {stage5_48[6]}
   );
   gpc1_1 gpc9542 (
      {stage4_48[16]},
      {stage5_48[7]}
   );
   gpc1_1 gpc9543 (
      {stage4_48[17]},
      {stage5_48[8]}
   );
   gpc1_1 gpc9544 (
      {stage4_48[18]},
      {stage5_48[9]}
   );
   gpc1_1 gpc9545 (
      {stage4_48[19]},
      {stage5_48[10]}
   );
   gpc1_1 gpc9546 (
      {stage4_48[20]},
      {stage5_48[11]}
   );
   gpc1_1 gpc9547 (
      {stage4_48[21]},
      {stage5_48[12]}
   );
   gpc1_1 gpc9548 (
      {stage4_48[22]},
      {stage5_48[13]}
   );
   gpc1_1 gpc9549 (
      {stage4_49[12]},
      {stage5_49[5]}
   );
   gpc1_1 gpc9550 (
      {stage4_50[17]},
      {stage5_50[7]}
   );
   gpc1_1 gpc9551 (
      {stage4_50[18]},
      {stage5_50[8]}
   );
   gpc1_1 gpc9552 (
      {stage4_50[19]},
      {stage5_50[9]}
   );
   gpc1_1 gpc9553 (
      {stage4_50[20]},
      {stage5_50[10]}
   );
   gpc1_1 gpc9554 (
      {stage4_50[21]},
      {stage5_50[11]}
   );
   gpc1_1 gpc9555 (
      {stage4_51[27]},
      {stage5_51[10]}
   );
   gpc1_1 gpc9556 (
      {stage4_51[28]},
      {stage5_51[11]}
   );
   gpc1_1 gpc9557 (
      {stage4_51[29]},
      {stage5_51[12]}
   );
   gpc1_1 gpc9558 (
      {stage4_51[30]},
      {stage5_51[13]}
   );
   gpc1_1 gpc9559 (
      {stage4_51[31]},
      {stage5_51[14]}
   );
   gpc1_1 gpc9560 (
      {stage4_51[32]},
      {stage5_51[15]}
   );
   gpc1_1 gpc9561 (
      {stage4_51[33]},
      {stage5_51[16]}
   );
   gpc1_1 gpc9562 (
      {stage4_51[34]},
      {stage5_51[17]}
   );
   gpc1_1 gpc9563 (
      {stage4_51[35]},
      {stage5_51[18]}
   );
   gpc1_1 gpc9564 (
      {stage4_52[17]},
      {stage5_52[8]}
   );
   gpc1_1 gpc9565 (
      {stage4_52[18]},
      {stage5_52[9]}
   );
   gpc1_1 gpc9566 (
      {stage4_53[40]},
      {stage5_53[9]}
   );
   gpc1_1 gpc9567 (
      {stage4_53[41]},
      {stage5_53[10]}
   );
   gpc1_1 gpc9568 (
      {stage4_53[42]},
      {stage5_53[11]}
   );
   gpc1_1 gpc9569 (
      {stage4_53[43]},
      {stage5_53[12]}
   );
   gpc1_1 gpc9570 (
      {stage4_54[22]},
      {stage5_54[13]}
   );
   gpc1_1 gpc9571 (
      {stage4_54[23]},
      {stage5_54[14]}
   );
   gpc1_1 gpc9572 (
      {stage4_54[24]},
      {stage5_54[15]}
   );
   gpc1_1 gpc9573 (
      {stage4_54[25]},
      {stage5_54[16]}
   );
   gpc1_1 gpc9574 (
      {stage4_55[29]},
      {stage5_55[12]}
   );
   gpc1_1 gpc9575 (
      {stage4_55[30]},
      {stage5_55[13]}
   );
   gpc1_1 gpc9576 (
      {stage4_55[31]},
      {stage5_55[14]}
   );
   gpc1_1 gpc9577 (
      {stage4_55[32]},
      {stage5_55[15]}
   );
   gpc1_1 gpc9578 (
      {stage4_55[33]},
      {stage5_55[16]}
   );
   gpc1_1 gpc9579 (
      {stage4_55[34]},
      {stage5_55[17]}
   );
   gpc1_1 gpc9580 (
      {stage4_55[35]},
      {stage5_55[18]}
   );
   gpc1_1 gpc9581 (
      {stage4_55[36]},
      {stage5_55[19]}
   );
   gpc1_1 gpc9582 (
      {stage4_55[37]},
      {stage5_55[20]}
   );
   gpc1_1 gpc9583 (
      {stage4_55[38]},
      {stage5_55[21]}
   );
   gpc1_1 gpc9584 (
      {stage4_57[22]},
      {stage5_57[10]}
   );
   gpc1_1 gpc9585 (
      {stage4_57[23]},
      {stage5_57[11]}
   );
   gpc1_1 gpc9586 (
      {stage4_57[24]},
      {stage5_57[12]}
   );
   gpc1_1 gpc9587 (
      {stage4_57[25]},
      {stage5_57[13]}
   );
   gpc1_1 gpc9588 (
      {stage4_58[17]},
      {stage5_58[9]}
   );
   gpc1_1 gpc9589 (
      {stage4_58[18]},
      {stage5_58[10]}
   );
   gpc1_1 gpc9590 (
      {stage4_58[19]},
      {stage5_58[11]}
   );
   gpc1_1 gpc9591 (
      {stage4_58[20]},
      {stage5_58[12]}
   );
   gpc1_1 gpc9592 (
      {stage4_58[21]},
      {stage5_58[13]}
   );
   gpc1_1 gpc9593 (
      {stage4_58[22]},
      {stage5_58[14]}
   );
   gpc1_1 gpc9594 (
      {stage4_58[23]},
      {stage5_58[15]}
   );
   gpc1_1 gpc9595 (
      {stage4_60[15]},
      {stage5_60[8]}
   );
   gpc1_1 gpc9596 (
      {stage4_60[16]},
      {stage5_60[9]}
   );
   gpc1_1 gpc9597 (
      {stage4_60[17]},
      {stage5_60[10]}
   );
   gpc1_1 gpc9598 (
      {stage4_60[18]},
      {stage5_60[11]}
   );
   gpc1_1 gpc9599 (
      {stage4_60[19]},
      {stage5_60[12]}
   );
   gpc1_1 gpc9600 (
      {stage4_60[20]},
      {stage5_60[13]}
   );
   gpc1_1 gpc9601 (
      {stage4_60[21]},
      {stage5_60[14]}
   );
   gpc1_1 gpc9602 (
      {stage4_61[23]},
      {stage5_61[7]}
   );
   gpc1_1 gpc9603 (
      {stage4_61[24]},
      {stage5_61[8]}
   );
   gpc1_1 gpc9604 (
      {stage4_61[25]},
      {stage5_61[9]}
   );
   gpc1_1 gpc9605 (
      {stage4_61[26]},
      {stage5_61[10]}
   );
   gpc1_1 gpc9606 (
      {stage4_61[27]},
      {stage5_61[11]}
   );
   gpc1_1 gpc9607 (
      {stage4_61[28]},
      {stage5_61[12]}
   );
   gpc1_1 gpc9608 (
      {stage4_61[29]},
      {stage5_61[13]}
   );
   gpc1_1 gpc9609 (
      {stage4_61[30]},
      {stage5_61[14]}
   );
   gpc1_1 gpc9610 (
      {stage4_61[31]},
      {stage5_61[15]}
   );
   gpc1_1 gpc9611 (
      {stage4_62[12]},
      {stage5_62[7]}
   );
   gpc1_1 gpc9612 (
      {stage4_62[13]},
      {stage5_62[8]}
   );
   gpc1_1 gpc9613 (
      {stage4_62[14]},
      {stage5_62[9]}
   );
   gpc1_1 gpc9614 (
      {stage4_62[15]},
      {stage5_62[10]}
   );
   gpc1_1 gpc9615 (
      {stage4_62[16]},
      {stage5_62[11]}
   );
   gpc1_1 gpc9616 (
      {stage4_63[12]},
      {stage5_63[7]}
   );
   gpc1_1 gpc9617 (
      {stage4_63[13]},
      {stage5_63[8]}
   );
   gpc1_1 gpc9618 (
      {stage4_64[28]},
      {stage5_64[9]}
   );
   gpc1_1 gpc9619 (
      {stage4_64[29]},
      {stage5_64[10]}
   );
   gpc1_1 gpc9620 (
      {stage4_64[30]},
      {stage5_64[11]}
   );
   gpc1_1 gpc9621 (
      {stage4_64[31]},
      {stage5_64[12]}
   );
   gpc1_1 gpc9622 (
      {stage4_64[32]},
      {stage5_64[13]}
   );
   gpc1_1 gpc9623 (
      {stage4_64[33]},
      {stage5_64[14]}
   );
   gpc1_1 gpc9624 (
      {stage4_65[26]},
      {stage5_65[8]}
   );
   gpc1_1 gpc9625 (
      {stage4_65[27]},
      {stage5_65[9]}
   );
   gpc1_1 gpc9626 (
      {stage4_65[28]},
      {stage5_65[10]}
   );
   gpc1_1 gpc9627 (
      {stage4_65[29]},
      {stage5_65[11]}
   );
   gpc1_1 gpc9628 (
      {stage4_65[30]},
      {stage5_65[12]}
   );
   gpc1_1 gpc9629 (
      {stage4_65[31]},
      {stage5_65[13]}
   );
   gpc1_1 gpc9630 (
      {stage4_65[32]},
      {stage5_65[14]}
   );
   gpc1_1 gpc9631 (
      {stage4_65[33]},
      {stage5_65[15]}
   );
   gpc1_1 gpc9632 (
      {stage4_65[34]},
      {stage5_65[16]}
   );
   gpc1_1 gpc9633 (
      {stage4_65[35]},
      {stage5_65[17]}
   );
   gpc1_1 gpc9634 (
      {stage4_67[7]},
      {stage5_67[7]}
   );
   gpc1_1 gpc9635 (
      {stage4_67[8]},
      {stage5_67[8]}
   );
   gpc1_1 gpc9636 (
      {stage4_67[9]},
      {stage5_67[9]}
   );
   gpc1_1 gpc9637 (
      {stage4_67[10]},
      {stage5_67[10]}
   );
   gpc1_1 gpc9638 (
      {stage4_68[6]},
      {stage5_68[6]}
   );
   gpc1_1 gpc9639 (
      {stage4_68[7]},
      {stage5_68[7]}
   );
   gpc1_1 gpc9640 (
      {stage4_68[8]},
      {stage5_68[8]}
   );
   gpc1_1 gpc9641 (
      {stage4_68[9]},
      {stage5_68[9]}
   );
   gpc1_1 gpc9642 (
      {stage4_68[10]},
      {stage5_68[10]}
   );
   gpc1_1 gpc9643 (
      {stage4_68[11]},
      {stage5_68[11]}
   );
   gpc1_1 gpc9644 (
      {stage4_68[12]},
      {stage5_68[12]}
   );
   gpc1_1 gpc9645 (
      {stage4_68[13]},
      {stage5_68[13]}
   );
   gpc1_1 gpc9646 (
      {stage4_69[0]},
      {stage5_69[1]}
   );
   gpc1_1 gpc9647 (
      {stage4_69[1]},
      {stage5_69[2]}
   );
   gpc615_5 gpc9648 (
      {stage5_3[0], stage5_3[1], stage5_3[2], stage5_3[3], stage5_3[4]},
      {stage5_4[0]},
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4], stage5_5[5]},
      {stage6_7[0],stage6_6[0],stage6_5[0],stage6_4[0],stage6_3[0]}
   );
   gpc615_5 gpc9649 (
      {stage5_3[5], stage5_3[6], stage5_3[7], 1'b0, 1'b0},
      {stage5_4[1]},
      {stage5_5[6], stage5_5[7], stage5_5[8], stage5_5[9], stage5_5[10], stage5_5[11]},
      {stage6_7[1],stage6_6[1],stage6_5[1],stage6_4[1],stage6_3[1]}
   );
   gpc606_5 gpc9650 (
      {stage5_4[2], stage5_4[3], stage5_4[4], stage5_4[5], stage5_4[6], stage5_4[7]},
      {stage5_6[0], stage5_6[1], stage5_6[2], stage5_6[3], stage5_6[4], stage5_6[5]},
      {stage6_8[0],stage6_7[2],stage6_6[2],stage6_5[2],stage6_4[2]}
   );
   gpc606_5 gpc9651 (
      {stage5_5[12], stage5_5[13], stage5_5[14], stage5_5[15], 1'b0, 1'b0},
      {stage5_7[0], stage5_7[1], stage5_7[2], stage5_7[3], stage5_7[4], stage5_7[5]},
      {stage6_9[0],stage6_8[1],stage6_7[3],stage6_6[3],stage6_5[3]}
   );
   gpc615_5 gpc9652 (
      {stage5_7[6], stage5_7[7], stage5_7[8], stage5_7[9], stage5_7[10]},
      {stage5_8[0]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3], stage5_9[4], stage5_9[5]},
      {stage6_11[0],stage6_10[0],stage6_9[1],stage6_8[2],stage6_7[4]}
   );
   gpc606_5 gpc9653 (
      {stage5_8[1], stage5_8[2], stage5_8[3], stage5_8[4], stage5_8[5], stage5_8[6]},
      {stage5_10[0], stage5_10[1], stage5_10[2], stage5_10[3], stage5_10[4], stage5_10[5]},
      {stage6_12[0],stage6_11[1],stage6_10[1],stage6_9[2],stage6_8[3]}
   );
   gpc606_5 gpc9654 (
      {stage5_8[7], stage5_8[8], stage5_8[9], stage5_8[10], stage5_8[11], stage5_8[12]},
      {stage5_10[6], stage5_10[7], stage5_10[8], stage5_10[9], stage5_10[10], stage5_10[11]},
      {stage6_12[1],stage6_11[2],stage6_10[2],stage6_9[3],stage6_8[4]}
   );
   gpc606_5 gpc9655 (
      {stage5_8[13], stage5_8[14], stage5_8[15], stage5_8[16], stage5_8[17], stage5_8[18]},
      {stage5_10[12], stage5_10[13], stage5_10[14], stage5_10[15], stage5_10[16], stage5_10[17]},
      {stage6_12[2],stage6_11[3],stage6_10[3],stage6_9[4],stage6_8[5]}
   );
   gpc615_5 gpc9656 (
      {stage5_10[18], stage5_10[19], stage5_10[20], 1'b0, 1'b0},
      {stage5_11[0]},
      {stage5_12[0], stage5_12[1], stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5]},
      {stage6_14[0],stage6_13[0],stage6_12[3],stage6_11[4],stage6_10[4]}
   );
   gpc1406_5 gpc9657 (
      {stage5_11[1], stage5_11[2], stage5_11[3], stage5_11[4], stage5_11[5], stage5_11[6]},
      {stage5_13[0], stage5_13[1], stage5_13[2], stage5_13[3]},
      {stage5_14[0]},
      {stage6_15[0],stage6_14[1],stage6_13[1],stage6_12[4],stage6_11[5]}
   );
   gpc7_3 gpc9658 (
      {stage5_11[7], stage5_11[8], stage5_11[9], stage5_11[10], stage5_11[11], stage5_11[12], stage5_11[13]},
      {stage6_13[2],stage6_12[5],stage6_11[6]}
   );
   gpc606_5 gpc9659 (
      {stage5_12[6], stage5_12[7], stage5_12[8], stage5_12[9], stage5_12[10], 1'b0},
      {stage5_14[1], stage5_14[2], stage5_14[3], stage5_14[4], stage5_14[5], stage5_14[6]},
      {stage6_16[0],stage6_15[1],stage6_14[2],stage6_13[3],stage6_12[6]}
   );
   gpc606_5 gpc9660 (
      {stage5_13[4], stage5_13[5], stage5_13[6], stage5_13[7], stage5_13[8], stage5_13[9]},
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3], stage5_15[4], stage5_15[5]},
      {stage6_17[0],stage6_16[1],stage6_15[2],stage6_14[3],stage6_13[4]}
   );
   gpc1343_5 gpc9661 (
      {stage5_14[7], stage5_14[8], stage5_14[9]},
      {stage5_15[6], stage5_15[7], stage5_15[8], stage5_15[9]},
      {stage5_16[0], stage5_16[1], stage5_16[2]},
      {stage5_17[0]},
      {stage6_18[0],stage6_17[1],stage6_16[2],stage6_15[3],stage6_14[4]}
   );
   gpc615_5 gpc9662 (
      {stage5_14[10], stage5_14[11], stage5_14[12], stage5_14[13], stage5_14[14]},
      {stage5_15[10]},
      {stage5_16[3], stage5_16[4], stage5_16[5], stage5_16[6], stage5_16[7], 1'b0},
      {stage6_18[1],stage6_17[2],stage6_16[3],stage6_15[4],stage6_14[5]}
   );
   gpc615_5 gpc9663 (
      {stage5_14[15], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage5_15[11]},
      {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
      {stage6_18[2],stage6_17[3],stage6_16[4],stage6_15[5],stage6_14[6]}
   );
   gpc606_5 gpc9664 (
      {stage5_17[1], stage5_17[2], stage5_17[3], stage5_17[4], stage5_17[5], stage5_17[6]},
      {stage5_19[0], stage5_19[1], stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5]},
      {stage6_21[0],stage6_20[0],stage6_19[0],stage6_18[3],stage6_17[4]}
   );
   gpc117_4 gpc9665 (
      {stage5_18[0], stage5_18[1], stage5_18[2], stage5_18[3], stage5_18[4], stage5_18[5], stage5_18[6]},
      {stage5_19[6]},
      {stage5_20[0]},
      {stage6_21[1],stage6_20[1],stage6_19[1],stage6_18[4]}
   );
   gpc615_5 gpc9666 (
      {stage5_18[7], stage5_18[8], stage5_18[9], stage5_18[10], stage5_18[11]},
      {stage5_19[7]},
      {stage5_20[1], stage5_20[2], stage5_20[3], stage5_20[4], stage5_20[5], stage5_20[6]},
      {stage6_22[0],stage6_21[2],stage6_20[2],stage6_19[2],stage6_18[5]}
   );
   gpc615_5 gpc9667 (
      {stage5_19[8], stage5_19[9], stage5_19[10], stage5_19[11], stage5_19[12]},
      {stage5_20[7]},
      {stage5_21[0], stage5_21[1], stage5_21[2], stage5_21[3], stage5_21[4], stage5_21[5]},
      {stage6_23[0],stage6_22[1],stage6_21[3],stage6_20[3],stage6_19[3]}
   );
   gpc615_5 gpc9668 (
      {stage5_19[13], stage5_19[14], stage5_19[15], 1'b0, 1'b0},
      {stage5_20[8]},
      {stage5_21[6], stage5_21[7], stage5_21[8], stage5_21[9], stage5_21[10], 1'b0},
      {stage6_23[1],stage6_22[2],stage6_21[4],stage6_20[4],stage6_19[4]}
   );
   gpc606_5 gpc9669 (
      {stage5_20[9], stage5_20[10], stage5_20[11], stage5_20[12], stage5_20[13], 1'b0},
      {stage5_22[0], stage5_22[1], stage5_22[2], stage5_22[3], stage5_22[4], stage5_22[5]},
      {stage6_24[0],stage6_23[2],stage6_22[3],stage6_21[5],stage6_20[5]}
   );
   gpc15_3 gpc9670 (
      {stage5_22[6], stage5_22[7], stage5_22[8], stage5_22[9], stage5_22[10]},
      {stage5_23[0]},
      {stage6_24[1],stage6_23[3],stage6_22[4]}
   );
   gpc15_3 gpc9671 (
      {stage5_22[11], stage5_22[12], stage5_22[13], 1'b0, 1'b0},
      {stage5_23[1]},
      {stage6_24[2],stage6_23[4],stage6_22[5]}
   );
   gpc615_5 gpc9672 (
      {stage5_23[2], stage5_23[3], stage5_23[4], stage5_23[5], stage5_23[6]},
      {stage5_24[0]},
      {stage5_25[0], stage5_25[1], stage5_25[2], stage5_25[3], stage5_25[4], stage5_25[5]},
      {stage6_27[0],stage6_26[0],stage6_25[0],stage6_24[3],stage6_23[5]}
   );
   gpc615_5 gpc9673 (
      {stage5_23[7], stage5_23[8], stage5_23[9], 1'b0, 1'b0},
      {stage5_24[1]},
      {stage5_25[6], stage5_25[7], stage5_25[8], stage5_25[9], 1'b0, 1'b0},
      {stage6_27[1],stage6_26[1],stage6_25[1],stage6_24[4],stage6_23[6]}
   );
   gpc606_5 gpc9674 (
      {stage5_24[2], stage5_24[3], stage5_24[4], stage5_24[5], stage5_24[6], stage5_24[7]},
      {stage5_26[0], stage5_26[1], stage5_26[2], stage5_26[3], stage5_26[4], stage5_26[5]},
      {stage6_28[0],stage6_27[2],stage6_26[2],stage6_25[2],stage6_24[5]}
   );
   gpc615_5 gpc9675 (
      {stage5_26[6], stage5_26[7], stage5_26[8], stage5_26[9], stage5_26[10]},
      {stage5_27[0]},
      {stage5_28[0], stage5_28[1], stage5_28[2], stage5_28[3], stage5_28[4], stage5_28[5]},
      {stage6_30[0],stage6_29[0],stage6_28[1],stage6_27[3],stage6_26[3]}
   );
   gpc615_5 gpc9676 (
      {stage5_27[1], stage5_27[2], stage5_27[3], stage5_27[4], stage5_27[5]},
      {stage5_28[6]},
      {stage5_29[0], stage5_29[1], stage5_29[2], stage5_29[3], stage5_29[4], stage5_29[5]},
      {stage6_31[0],stage6_30[1],stage6_29[1],stage6_28[2],stage6_27[4]}
   );
   gpc606_5 gpc9677 (
      {stage5_29[6], stage5_29[7], stage5_29[8], stage5_29[9], stage5_29[10], stage5_29[11]},
      {stage5_31[0], stage5_31[1], stage5_31[2], stage5_31[3], stage5_31[4], stage5_31[5]},
      {stage6_33[0],stage6_32[0],stage6_31[1],stage6_30[2],stage6_29[2]}
   );
   gpc615_5 gpc9678 (
      {stage5_30[0], stage5_30[1], stage5_30[2], stage5_30[3], stage5_30[4]},
      {stage5_31[6]},
      {stage5_32[0], stage5_32[1], stage5_32[2], stage5_32[3], stage5_32[4], stage5_32[5]},
      {stage6_34[0],stage6_33[1],stage6_32[1],stage6_31[2],stage6_30[3]}
   );
   gpc615_5 gpc9679 (
      {stage5_30[5], stage5_30[6], stage5_30[7], stage5_30[8], 1'b0},
      {stage5_31[7]},
      {stage5_32[6], stage5_32[7], stage5_32[8], stage5_32[9], stage5_32[10], stage5_32[11]},
      {stage6_34[1],stage6_33[2],stage6_32[2],stage6_31[3],stage6_30[4]}
   );
   gpc606_5 gpc9680 (
      {stage5_32[12], stage5_32[13], stage5_32[14], stage5_32[15], stage5_32[16], stage5_32[17]},
      {stage5_34[0], stage5_34[1], stage5_34[2], stage5_34[3], stage5_34[4], stage5_34[5]},
      {stage6_36[0],stage6_35[0],stage6_34[2],stage6_33[3],stage6_32[3]}
   );
   gpc606_5 gpc9681 (
      {stage5_33[0], stage5_33[1], stage5_33[2], stage5_33[3], stage5_33[4], stage5_33[5]},
      {stage5_35[0], stage5_35[1], stage5_35[2], stage5_35[3], stage5_35[4], stage5_35[5]},
      {stage6_37[0],stage6_36[1],stage6_35[1],stage6_34[3],stage6_33[4]}
   );
   gpc606_5 gpc9682 (
      {stage5_33[6], stage5_33[7], stage5_33[8], stage5_33[9], stage5_33[10], stage5_33[11]},
      {stage5_35[6], stage5_35[7], stage5_35[8], stage5_35[9], stage5_35[10], stage5_35[11]},
      {stage6_37[1],stage6_36[2],stage6_35[2],stage6_34[4],stage6_33[5]}
   );
   gpc615_5 gpc9683 (
      {stage5_34[6], stage5_34[7], stage5_34[8], stage5_34[9], stage5_34[10]},
      {stage5_35[12]},
      {stage5_36[0], stage5_36[1], stage5_36[2], stage5_36[3], stage5_36[4], stage5_36[5]},
      {stage6_38[0],stage6_37[2],stage6_36[3],stage6_35[3],stage6_34[5]}
   );
   gpc606_5 gpc9684 (
      {stage5_36[6], stage5_36[7], stage5_36[8], stage5_36[9], stage5_36[10], stage5_36[11]},
      {stage5_38[0], stage5_38[1], stage5_38[2], stage5_38[3], stage5_38[4], stage5_38[5]},
      {stage6_40[0],stage6_39[0],stage6_38[1],stage6_37[3],stage6_36[4]}
   );
   gpc2135_5 gpc9685 (
      {stage5_37[0], stage5_37[1], stage5_37[2], stage5_37[3], stage5_37[4]},
      {stage5_38[6], stage5_38[7], stage5_38[8]},
      {stage5_39[0]},
      {stage5_40[0], stage5_40[1]},
      {stage6_41[0],stage6_40[1],stage6_39[1],stage6_38[2],stage6_37[4]}
   );
   gpc606_5 gpc9686 (
      {stage5_37[5], stage5_37[6], stage5_37[7], stage5_37[8], stage5_37[9], stage5_37[10]},
      {stage5_39[1], stage5_39[2], stage5_39[3], stage5_39[4], stage5_39[5], stage5_39[6]},
      {stage6_41[1],stage6_40[2],stage6_39[2],stage6_38[3],stage6_37[5]}
   );
   gpc23_3 gpc9687 (
      {stage5_39[7], stage5_39[8], stage5_39[9]},
      {stage5_40[2], stage5_40[3]},
      {stage6_41[2],stage6_40[3],stage6_39[3]}
   );
   gpc606_5 gpc9688 (
      {stage5_40[4], stage5_40[5], stage5_40[6], stage5_40[7], stage5_40[8], stage5_40[9]},
      {stage5_42[0], stage5_42[1], stage5_42[2], stage5_42[3], stage5_42[4], stage5_42[5]},
      {stage6_44[0],stage6_43[0],stage6_42[0],stage6_41[3],stage6_40[4]}
   );
   gpc606_5 gpc9689 (
      {stage5_41[0], stage5_41[1], stage5_41[2], stage5_41[3], stage5_41[4], stage5_41[5]},
      {stage5_43[0], stage5_43[1], stage5_43[2], stage5_43[3], stage5_43[4], stage5_43[5]},
      {stage6_45[0],stage6_44[1],stage6_43[1],stage6_42[1],stage6_41[4]}
   );
   gpc615_5 gpc9690 (
      {stage5_42[6], stage5_42[7], stage5_42[8], stage5_42[9], stage5_42[10]},
      {stage5_43[6]},
      {stage5_44[0], stage5_44[1], stage5_44[2], stage5_44[3], stage5_44[4], stage5_44[5]},
      {stage6_46[0],stage6_45[1],stage6_44[2],stage6_43[2],stage6_42[2]}
   );
   gpc615_5 gpc9691 (
      {stage5_42[11], stage5_42[12], stage5_42[13], stage5_42[14], stage5_42[15]},
      {stage5_43[7]},
      {stage5_44[6], stage5_44[7], stage5_44[8], stage5_44[9], stage5_44[10], stage5_44[11]},
      {stage6_46[1],stage6_45[2],stage6_44[3],stage6_43[3],stage6_42[3]}
   );
   gpc1163_5 gpc9692 (
      {stage5_45[0], stage5_45[1], stage5_45[2]},
      {stage5_46[0], stage5_46[1], stage5_46[2], stage5_46[3], stage5_46[4], stage5_46[5]},
      {stage5_47[0]},
      {stage5_48[0]},
      {stage6_49[0],stage6_48[0],stage6_47[0],stage6_46[2],stage6_45[3]}
   );
   gpc1163_5 gpc9693 (
      {stage5_45[3], stage5_45[4], stage5_45[5]},
      {stage5_46[6], stage5_46[7], stage5_46[8], stage5_46[9], stage5_46[10], stage5_46[11]},
      {stage5_47[1]},
      {stage5_48[1]},
      {stage6_49[1],stage6_48[1],stage6_47[1],stage6_46[3],stage6_45[4]}
   );
   gpc606_5 gpc9694 (
      {stage5_45[6], stage5_45[7], stage5_45[8], stage5_45[9], stage5_45[10], stage5_45[11]},
      {stage5_47[2], stage5_47[3], stage5_47[4], stage5_47[5], stage5_47[6], stage5_47[7]},
      {stage6_49[2],stage6_48[2],stage6_47[2],stage6_46[4],stage6_45[5]}
   );
   gpc606_5 gpc9695 (
      {stage5_48[2], stage5_48[3], stage5_48[4], stage5_48[5], stage5_48[6], stage5_48[7]},
      {stage5_50[0], stage5_50[1], stage5_50[2], stage5_50[3], stage5_50[4], stage5_50[5]},
      {stage6_52[0],stage6_51[0],stage6_50[0],stage6_49[3],stage6_48[3]}
   );
   gpc606_5 gpc9696 (
      {stage5_48[8], stage5_48[9], stage5_48[10], stage5_48[11], stage5_48[12], stage5_48[13]},
      {stage5_50[6], stage5_50[7], stage5_50[8], stage5_50[9], stage5_50[10], stage5_50[11]},
      {stage6_52[1],stage6_51[1],stage6_50[1],stage6_49[4],stage6_48[4]}
   );
   gpc606_5 gpc9697 (
      {stage5_49[0], stage5_49[1], stage5_49[2], stage5_49[3], stage5_49[4], stage5_49[5]},
      {stage5_51[0], stage5_51[1], stage5_51[2], stage5_51[3], stage5_51[4], stage5_51[5]},
      {stage6_53[0],stage6_52[2],stage6_51[2],stage6_50[2],stage6_49[5]}
   );
   gpc7_3 gpc9698 (
      {stage5_51[6], stage5_51[7], stage5_51[8], stage5_51[9], stage5_51[10], stage5_51[11], stage5_51[12]},
      {stage6_53[1],stage6_52[3],stage6_51[3]}
   );
   gpc623_5 gpc9699 (
      {stage5_51[13], stage5_51[14], stage5_51[15]},
      {stage5_52[0], stage5_52[1]},
      {stage5_53[0], stage5_53[1], stage5_53[2], stage5_53[3], stage5_53[4], stage5_53[5]},
      {stage6_55[0],stage6_54[0],stage6_53[2],stage6_52[4],stage6_51[4]}
   );
   gpc117_4 gpc9700 (
      {stage5_52[2], stage5_52[3], stage5_52[4], stage5_52[5], stage5_52[6], stage5_52[7], stage5_52[8]},
      {stage5_53[6]},
      {stage5_54[0]},
      {stage6_55[1],stage6_54[1],stage6_53[3],stage6_52[5]}
   );
   gpc117_4 gpc9701 (
      {stage5_53[7], stage5_53[8], stage5_53[9], stage5_53[10], stage5_53[11], stage5_53[12], 1'b0},
      {stage5_54[1]},
      {stage5_55[0]},
      {stage6_56[0],stage6_55[2],stage6_54[2],stage6_53[4]}
   );
   gpc135_4 gpc9702 (
      {stage5_54[2], stage5_54[3], stage5_54[4], stage5_54[5], stage5_54[6]},
      {stage5_55[1], stage5_55[2], stage5_55[3]},
      {stage5_56[0]},
      {stage6_57[0],stage6_56[1],stage6_55[3],stage6_54[3]}
   );
   gpc135_4 gpc9703 (
      {stage5_54[7], stage5_54[8], stage5_54[9], stage5_54[10], stage5_54[11]},
      {stage5_55[4], stage5_55[5], stage5_55[6]},
      {stage5_56[1]},
      {stage6_57[1],stage6_56[2],stage6_55[4],stage6_54[4]}
   );
   gpc135_4 gpc9704 (
      {stage5_54[12], stage5_54[13], stage5_54[14], stage5_54[15], stage5_54[16]},
      {stage5_55[7], stage5_55[8], stage5_55[9]},
      {stage5_56[2]},
      {stage6_57[2],stage6_56[3],stage6_55[5],stage6_54[5]}
   );
   gpc615_5 gpc9705 (
      {stage5_55[10], stage5_55[11], stage5_55[12], stage5_55[13], stage5_55[14]},
      {stage5_56[3]},
      {stage5_57[0], stage5_57[1], stage5_57[2], stage5_57[3], stage5_57[4], stage5_57[5]},
      {stage6_59[0],stage6_58[0],stage6_57[3],stage6_56[4],stage6_55[6]}
   );
   gpc615_5 gpc9706 (
      {stage5_55[15], stage5_55[16], stage5_55[17], stage5_55[18], stage5_55[19]},
      {stage5_56[4]},
      {stage5_57[6], stage5_57[7], stage5_57[8], stage5_57[9], stage5_57[10], stage5_57[11]},
      {stage6_59[1],stage6_58[1],stage6_57[4],stage6_56[5],stage6_55[7]}
   );
   gpc2135_5 gpc9707 (
      {stage5_58[0], stage5_58[1], stage5_58[2], stage5_58[3], stage5_58[4]},
      {stage5_59[0], stage5_59[1], stage5_59[2]},
      {stage5_60[0]},
      {stage5_61[0], stage5_61[1]},
      {stage6_62[0],stage6_61[0],stage6_60[0],stage6_59[2],stage6_58[2]}
   );
   gpc2135_5 gpc9708 (
      {stage5_58[5], stage5_58[6], stage5_58[7], stage5_58[8], stage5_58[9]},
      {stage5_59[3], stage5_59[4], stage5_59[5]},
      {stage5_60[1]},
      {stage5_61[2], stage5_61[3]},
      {stage6_62[1],stage6_61[1],stage6_60[1],stage6_59[3],stage6_58[3]}
   );
   gpc2135_5 gpc9709 (
      {stage5_58[10], stage5_58[11], stage5_58[12], stage5_58[13], stage5_58[14]},
      {stage5_59[6], stage5_59[7], 1'b0},
      {stage5_60[2]},
      {stage5_61[4], stage5_61[5]},
      {stage6_62[2],stage6_61[2],stage6_60[2],stage6_59[4],stage6_58[4]}
   );
   gpc606_5 gpc9710 (
      {stage5_60[3], stage5_60[4], stage5_60[5], stage5_60[6], stage5_60[7], stage5_60[8]},
      {stage5_62[0], stage5_62[1], stage5_62[2], stage5_62[3], stage5_62[4], stage5_62[5]},
      {stage6_64[0],stage6_63[0],stage6_62[3],stage6_61[3],stage6_60[3]}
   );
   gpc606_5 gpc9711 (
      {stage5_60[9], stage5_60[10], stage5_60[11], stage5_60[12], stage5_60[13], stage5_60[14]},
      {stage5_62[6], stage5_62[7], stage5_62[8], stage5_62[9], stage5_62[10], stage5_62[11]},
      {stage6_64[1],stage6_63[1],stage6_62[4],stage6_61[4],stage6_60[4]}
   );
   gpc207_4 gpc9712 (
      {stage5_61[6], stage5_61[7], stage5_61[8], stage5_61[9], stage5_61[10], stage5_61[11], stage5_61[12]},
      {stage5_63[0], stage5_63[1]},
      {stage6_64[2],stage6_63[2],stage6_62[5],stage6_61[5]}
   );
   gpc606_5 gpc9713 (
      {stage5_63[2], stage5_63[3], stage5_63[4], stage5_63[5], stage5_63[6], stage5_63[7]},
      {stage5_65[0], stage5_65[1], stage5_65[2], stage5_65[3], stage5_65[4], stage5_65[5]},
      {stage6_67[0],stage6_66[0],stage6_65[0],stage6_64[3],stage6_63[3]}
   );
   gpc1406_5 gpc9714 (
      {stage5_64[0], stage5_64[1], stage5_64[2], stage5_64[3], stage5_64[4], stage5_64[5]},
      {stage5_66[0], stage5_66[1], stage5_66[2], stage5_66[3]},
      {stage5_67[0]},
      {stage6_68[0],stage6_67[1],stage6_66[1],stage6_65[1],stage6_64[4]}
   );
   gpc1406_5 gpc9715 (
      {stage5_64[6], stage5_64[7], stage5_64[8], stage5_64[9], stage5_64[10], stage5_64[11]},
      {stage5_66[4], stage5_66[5], stage5_66[6], stage5_66[7]},
      {stage5_67[1]},
      {stage6_68[1],stage6_67[2],stage6_66[2],stage6_65[2],stage6_64[5]}
   );
   gpc1406_5 gpc9716 (
      {stage5_65[6], stage5_65[7], stage5_65[8], stage5_65[9], stage5_65[10], stage5_65[11]},
      {stage5_67[2], stage5_67[3], stage5_67[4], stage5_67[5]},
      {stage5_68[0]},
      {stage6_69[0],stage6_68[2],stage6_67[3],stage6_66[3],stage6_65[3]}
   );
   gpc606_5 gpc9717 (
      {stage5_65[12], stage5_65[13], stage5_65[14], stage5_65[15], stage5_65[16], stage5_65[17]},
      {stage5_67[6], stage5_67[7], stage5_67[8], stage5_67[9], stage5_67[10], 1'b0},
      {stage6_69[1],stage6_68[3],stage6_67[4],stage6_66[4],stage6_65[4]}
   );
   gpc1_1 gpc9718 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc9719 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc9720 (
      {stage5_0[2]},
      {stage6_0[2]}
   );
   gpc1_1 gpc9721 (
      {stage5_0[3]},
      {stage6_0[3]}
   );
   gpc1_1 gpc9722 (
      {stage5_0[4]},
      {stage6_0[4]}
   );
   gpc1_1 gpc9723 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc9724 (
      {stage5_1[1]},
      {stage6_1[1]}
   );
   gpc1_1 gpc9725 (
      {stage5_2[0]},
      {stage6_2[0]}
   );
   gpc1_1 gpc9726 (
      {stage5_2[1]},
      {stage6_2[1]}
   );
   gpc1_1 gpc9727 (
      {stage5_2[2]},
      {stage6_2[2]}
   );
   gpc1_1 gpc9728 (
      {stage5_2[3]},
      {stage6_2[3]}
   );
   gpc1_1 gpc9729 (
      {stage5_2[4]},
      {stage6_2[4]}
   );
   gpc1_1 gpc9730 (
      {stage5_4[8]},
      {stage6_4[3]}
   );
   gpc1_1 gpc9731 (
      {stage5_4[9]},
      {stage6_4[4]}
   );
   gpc1_1 gpc9732 (
      {stage5_4[10]},
      {stage6_4[5]}
   );
   gpc1_1 gpc9733 (
      {stage5_6[6]},
      {stage6_6[4]}
   );
   gpc1_1 gpc9734 (
      {stage5_6[7]},
      {stage6_6[5]}
   );
   gpc1_1 gpc9735 (
      {stage5_6[8]},
      {stage6_6[6]}
   );
   gpc1_1 gpc9736 (
      {stage5_6[9]},
      {stage6_6[7]}
   );
   gpc1_1 gpc9737 (
      {stage5_9[6]},
      {stage6_9[5]}
   );
   gpc1_1 gpc9738 (
      {stage5_9[7]},
      {stage6_9[6]}
   );
   gpc1_1 gpc9739 (
      {stage5_9[8]},
      {stage6_9[7]}
   );
   gpc1_1 gpc9740 (
      {stage5_9[9]},
      {stage6_9[8]}
   );
   gpc1_1 gpc9741 (
      {stage5_9[10]},
      {stage6_9[9]}
   );
   gpc1_1 gpc9742 (
      {stage5_13[10]},
      {stage6_13[5]}
   );
   gpc1_1 gpc9743 (
      {stage5_13[11]},
      {stage6_13[6]}
   );
   gpc1_1 gpc9744 (
      {stage5_13[12]},
      {stage6_13[7]}
   );
   gpc1_1 gpc9745 (
      {stage5_13[13]},
      {stage6_13[8]}
   );
   gpc1_1 gpc9746 (
      {stage5_13[14]},
      {stage6_13[9]}
   );
   gpc1_1 gpc9747 (
      {stage5_24[8]},
      {stage6_24[6]}
   );
   gpc1_1 gpc9748 (
      {stage5_26[11]},
      {stage6_26[4]}
   );
   gpc1_1 gpc9749 (
      {stage5_26[12]},
      {stage6_26[5]}
   );
   gpc1_1 gpc9750 (
      {stage5_26[13]},
      {stage6_26[6]}
   );
   gpc1_1 gpc9751 (
      {stage5_26[14]},
      {stage6_26[7]}
   );
   gpc1_1 gpc9752 (
      {stage5_28[7]},
      {stage6_28[3]}
   );
   gpc1_1 gpc9753 (
      {stage5_28[8]},
      {stage6_28[4]}
   );
   gpc1_1 gpc9754 (
      {stage5_28[9]},
      {stage6_28[5]}
   );
   gpc1_1 gpc9755 (
      {stage5_29[12]},
      {stage6_29[3]}
   );
   gpc1_1 gpc9756 (
      {stage5_29[13]},
      {stage6_29[4]}
   );
   gpc1_1 gpc9757 (
      {stage5_29[14]},
      {stage6_29[5]}
   );
   gpc1_1 gpc9758 (
      {stage5_31[8]},
      {stage6_31[4]}
   );
   gpc1_1 gpc9759 (
      {stage5_31[9]},
      {stage6_31[5]}
   );
   gpc1_1 gpc9760 (
      {stage5_32[18]},
      {stage6_32[4]}
   );
   gpc1_1 gpc9761 (
      {stage5_32[19]},
      {stage6_32[5]}
   );
   gpc1_1 gpc9762 (
      {stage5_34[11]},
      {stage6_34[6]}
   );
   gpc1_1 gpc9763 (
      {stage5_34[12]},
      {stage6_34[7]}
   );
   gpc1_1 gpc9764 (
      {stage5_34[13]},
      {stage6_34[8]}
   );
   gpc1_1 gpc9765 (
      {stage5_35[13]},
      {stage6_35[4]}
   );
   gpc1_1 gpc9766 (
      {stage5_36[12]},
      {stage6_36[5]}
   );
   gpc1_1 gpc9767 (
      {stage5_38[9]},
      {stage6_38[4]}
   );
   gpc1_1 gpc9768 (
      {stage5_40[10]},
      {stage6_40[5]}
   );
   gpc1_1 gpc9769 (
      {stage5_41[6]},
      {stage6_41[5]}
   );
   gpc1_1 gpc9770 (
      {stage5_41[7]},
      {stage6_41[6]}
   );
   gpc1_1 gpc9771 (
      {stage5_41[8]},
      {stage6_41[7]}
   );
   gpc1_1 gpc9772 (
      {stage5_42[16]},
      {stage6_42[4]}
   );
   gpc1_1 gpc9773 (
      {stage5_42[17]},
      {stage6_42[5]}
   );
   gpc1_1 gpc9774 (
      {stage5_42[18]},
      {stage6_42[6]}
   );
   gpc1_1 gpc9775 (
      {stage5_43[8]},
      {stage6_43[4]}
   );
   gpc1_1 gpc9776 (
      {stage5_43[9]},
      {stage6_43[5]}
   );
   gpc1_1 gpc9777 (
      {stage5_43[10]},
      {stage6_43[6]}
   );
   gpc1_1 gpc9778 (
      {stage5_44[12]},
      {stage6_44[4]}
   );
   gpc1_1 gpc9779 (
      {stage5_45[12]},
      {stage6_45[6]}
   );
   gpc1_1 gpc9780 (
      {stage5_45[13]},
      {stage6_45[7]}
   );
   gpc1_1 gpc9781 (
      {stage5_45[14]},
      {stage6_45[8]}
   );
   gpc1_1 gpc9782 (
      {stage5_47[8]},
      {stage6_47[3]}
   );
   gpc1_1 gpc9783 (
      {stage5_47[9]},
      {stage6_47[4]}
   );
   gpc1_1 gpc9784 (
      {stage5_47[10]},
      {stage6_47[5]}
   );
   gpc1_1 gpc9785 (
      {stage5_47[11]},
      {stage6_47[6]}
   );
   gpc1_1 gpc9786 (
      {stage5_51[16]},
      {stage6_51[5]}
   );
   gpc1_1 gpc9787 (
      {stage5_51[17]},
      {stage6_51[6]}
   );
   gpc1_1 gpc9788 (
      {stage5_51[18]},
      {stage6_51[7]}
   );
   gpc1_1 gpc9789 (
      {stage5_52[9]},
      {stage6_52[6]}
   );
   gpc1_1 gpc9790 (
      {stage5_55[20]},
      {stage6_55[8]}
   );
   gpc1_1 gpc9791 (
      {stage5_55[21]},
      {stage6_55[9]}
   );
   gpc1_1 gpc9792 (
      {stage5_56[5]},
      {stage6_56[6]}
   );
   gpc1_1 gpc9793 (
      {stage5_56[6]},
      {stage6_56[7]}
   );
   gpc1_1 gpc9794 (
      {stage5_56[7]},
      {stage6_56[8]}
   );
   gpc1_1 gpc9795 (
      {stage5_56[8]},
      {stage6_56[9]}
   );
   gpc1_1 gpc9796 (
      {stage5_57[12]},
      {stage6_57[5]}
   );
   gpc1_1 gpc9797 (
      {stage5_57[13]},
      {stage6_57[6]}
   );
   gpc1_1 gpc9798 (
      {stage5_58[15]},
      {stage6_58[5]}
   );
   gpc1_1 gpc9799 (
      {stage5_61[13]},
      {stage6_61[6]}
   );
   gpc1_1 gpc9800 (
      {stage5_61[14]},
      {stage6_61[7]}
   );
   gpc1_1 gpc9801 (
      {stage5_61[15]},
      {stage6_61[8]}
   );
   gpc1_1 gpc9802 (
      {stage5_63[8]},
      {stage6_63[4]}
   );
   gpc1_1 gpc9803 (
      {stage5_64[12]},
      {stage6_64[6]}
   );
   gpc1_1 gpc9804 (
      {stage5_64[13]},
      {stage6_64[7]}
   );
   gpc1_1 gpc9805 (
      {stage5_64[14]},
      {stage6_64[8]}
   );
   gpc1_1 gpc9806 (
      {stage5_68[1]},
      {stage6_68[4]}
   );
   gpc1_1 gpc9807 (
      {stage5_68[2]},
      {stage6_68[5]}
   );
   gpc1_1 gpc9808 (
      {stage5_68[3]},
      {stage6_68[6]}
   );
   gpc1_1 gpc9809 (
      {stage5_68[4]},
      {stage6_68[7]}
   );
   gpc1_1 gpc9810 (
      {stage5_68[5]},
      {stage6_68[8]}
   );
   gpc1_1 gpc9811 (
      {stage5_68[6]},
      {stage6_68[9]}
   );
   gpc1_1 gpc9812 (
      {stage5_68[7]},
      {stage6_68[10]}
   );
   gpc1_1 gpc9813 (
      {stage5_68[8]},
      {stage6_68[11]}
   );
   gpc1_1 gpc9814 (
      {stage5_68[9]},
      {stage6_68[12]}
   );
   gpc1_1 gpc9815 (
      {stage5_68[10]},
      {stage6_68[13]}
   );
   gpc1_1 gpc9816 (
      {stage5_68[11]},
      {stage6_68[14]}
   );
   gpc1_1 gpc9817 (
      {stage5_68[12]},
      {stage6_68[15]}
   );
   gpc1_1 gpc9818 (
      {stage5_68[13]},
      {stage6_68[16]}
   );
   gpc1_1 gpc9819 (
      {stage5_69[0]},
      {stage6_69[2]}
   );
   gpc1_1 gpc9820 (
      {stage5_69[1]},
      {stage6_69[3]}
   );
   gpc1_1 gpc9821 (
      {stage5_69[2]},
      {stage6_69[4]}
   );
   gpc1_1 gpc9822 (
      {stage5_70[0]},
      {stage6_70[0]}
   );
   gpc1406_5 gpc9823 (
      {stage6_4[0], stage6_4[1], stage6_4[2], stage6_4[3], stage6_4[4], stage6_4[5]},
      {stage6_6[0], stage6_6[1], stage6_6[2], stage6_6[3]},
      {stage6_7[0]},
      {stage7_8[0],stage7_7[0],stage7_6[0],stage7_5[0],stage7_4[0]}
   );
   gpc2135_5 gpc9824 (
      {stage6_5[0], stage6_5[1], stage6_5[2], stage6_5[3], 1'b0},
      {stage6_6[4], stage6_6[5], stage6_6[6]},
      {stage6_7[1]},
      {stage6_8[0], stage6_8[1]},
      {stage7_9[0],stage7_8[1],stage7_7[1],stage7_6[1],stage7_5[1]}
   );
   gpc623_5 gpc9825 (
      {stage6_7[2], stage6_7[3], stage6_7[4]},
      {stage6_8[2], stage6_8[3]},
      {stage6_9[0], stage6_9[1], stage6_9[2], stage6_9[3], stage6_9[4], stage6_9[5]},
      {stage7_11[0],stage7_10[0],stage7_9[1],stage7_8[2],stage7_7[2]}
   );
   gpc615_5 gpc9826 (
      {stage6_10[0], stage6_10[1], stage6_10[2], stage6_10[3], stage6_10[4]},
      {stage6_11[0]},
      {stage6_12[0], stage6_12[1], stage6_12[2], stage6_12[3], stage6_12[4], stage6_12[5]},
      {stage7_14[0],stage7_13[0],stage7_12[0],stage7_11[1],stage7_10[1]}
   );
   gpc615_5 gpc9827 (
      {stage6_11[1], stage6_11[2], stage6_11[3], stage6_11[4], stage6_11[5]},
      {stage6_12[6]},
      {stage6_13[0], stage6_13[1], stage6_13[2], stage6_13[3], stage6_13[4], stage6_13[5]},
      {stage7_15[0],stage7_14[1],stage7_13[1],stage7_12[1],stage7_11[2]}
   );
   gpc7_3 gpc9828 (
      {stage6_14[0], stage6_14[1], stage6_14[2], stage6_14[3], stage6_14[4], stage6_14[5], stage6_14[6]},
      {stage7_16[0],stage7_15[1],stage7_14[2]}
   );
   gpc623_5 gpc9829 (
      {stage6_15[0], stage6_15[1], stage6_15[2]},
      {stage6_16[0], stage6_16[1]},
      {stage6_17[0], stage6_17[1], stage6_17[2], stage6_17[3], stage6_17[4], 1'b0},
      {stage7_19[0],stage7_18[0],stage7_17[0],stage7_16[1],stage7_15[2]}
   );
   gpc606_5 gpc9830 (
      {stage6_16[2], stage6_16[3], stage6_16[4], 1'b0, 1'b0, 1'b0},
      {stage6_18[0], stage6_18[1], stage6_18[2], stage6_18[3], stage6_18[4], stage6_18[5]},
      {stage7_20[0],stage7_19[1],stage7_18[1],stage7_17[1],stage7_16[2]}
   );
   gpc15_3 gpc9831 (
      {stage6_20[0], stage6_20[1], stage6_20[2], stage6_20[3], stage6_20[4]},
      {stage6_21[0]},
      {stage7_22[0],stage7_21[0],stage7_20[1]}
   );
   gpc207_4 gpc9832 (
      {stage6_23[0], stage6_23[1], stage6_23[2], stage6_23[3], stage6_23[4], stage6_23[5], stage6_23[6]},
      {stage6_25[0], stage6_25[1]},
      {stage7_26[0],stage7_25[0],stage7_24[0],stage7_23[0]}
   );
   gpc15_3 gpc9833 (
      {stage6_24[0], stage6_24[1], stage6_24[2], stage6_24[3], stage6_24[4]},
      {stage6_25[2]},
      {stage7_26[1],stage7_25[1],stage7_24[1]}
   );
   gpc615_5 gpc9834 (
      {stage6_26[0], stage6_26[1], stage6_26[2], stage6_26[3], stage6_26[4]},
      {stage6_27[0]},
      {stage6_28[0], stage6_28[1], stage6_28[2], stage6_28[3], stage6_28[4], stage6_28[5]},
      {stage7_30[0],stage7_29[0],stage7_28[0],stage7_27[0],stage7_26[2]}
   );
   gpc3_2 gpc9835 (
      {stage6_29[0], stage6_29[1], stage6_29[2]},
      {stage7_30[1],stage7_29[1]}
   );
   gpc615_5 gpc9836 (
      {stage6_31[0], stage6_31[1], stage6_31[2], stage6_31[3], stage6_31[4]},
      {stage6_32[0]},
      {stage6_33[0], stage6_33[1], stage6_33[2], stage6_33[3], stage6_33[4], stage6_33[5]},
      {stage7_35[0],stage7_34[0],stage7_33[0],stage7_32[0],stage7_31[0]}
   );
   gpc615_5 gpc9837 (
      {stage6_34[0], stage6_34[1], stage6_34[2], stage6_34[3], stage6_34[4]},
      {stage6_35[0]},
      {stage6_36[0], stage6_36[1], stage6_36[2], stage6_36[3], stage6_36[4], stage6_36[5]},
      {stage7_38[0],stage7_37[0],stage7_36[0],stage7_35[1],stage7_34[1]}
   );
   gpc606_5 gpc9838 (
      {stage6_37[0], stage6_37[1], stage6_37[2], stage6_37[3], stage6_37[4], stage6_37[5]},
      {stage6_39[0], stage6_39[1], stage6_39[2], stage6_39[3], 1'b0, 1'b0},
      {stage7_41[0],stage7_40[0],stage7_39[0],stage7_38[1],stage7_37[1]}
   );
   gpc15_3 gpc9839 (
      {stage6_41[0], stage6_41[1], stage6_41[2], stage6_41[3], stage6_41[4]},
      {stage6_42[0]},
      {stage7_43[0],stage7_42[0],stage7_41[1]}
   );
   gpc615_5 gpc9840 (
      {stage6_42[1], stage6_42[2], stage6_42[3], stage6_42[4], stage6_42[5]},
      {stage6_43[0]},
      {stage6_44[0], stage6_44[1], stage6_44[2], stage6_44[3], stage6_44[4], 1'b0},
      {stage7_46[0],stage7_45[0],stage7_44[0],stage7_43[1],stage7_42[1]}
   );
   gpc615_5 gpc9841 (
      {stage6_43[1], stage6_43[2], stage6_43[3], stage6_43[4], stage6_43[5]},
      {1'b0},
      {stage6_45[0], stage6_45[1], stage6_45[2], stage6_45[3], stage6_45[4], stage6_45[5]},
      {stage7_47[0],stage7_46[1],stage7_45[1],stage7_44[1],stage7_43[2]}
   );
   gpc615_5 gpc9842 (
      {stage6_46[0], stage6_46[1], stage6_46[2], stage6_46[3], stage6_46[4]},
      {stage6_47[0]},
      {stage6_48[0], stage6_48[1], stage6_48[2], stage6_48[3], stage6_48[4], 1'b0},
      {stage7_50[0],stage7_49[0],stage7_48[0],stage7_47[1],stage7_46[2]}
   );
   gpc606_5 gpc9843 (
      {stage6_49[0], stage6_49[1], stage6_49[2], stage6_49[3], stage6_49[4], stage6_49[5]},
      {stage6_51[0], stage6_51[1], stage6_51[2], stage6_51[3], stage6_51[4], stage6_51[5]},
      {stage7_53[0],stage7_52[0],stage7_51[0],stage7_50[1],stage7_49[1]}
   );
   gpc3_2 gpc9844 (
      {stage6_50[0], stage6_50[1], stage6_50[2]},
      {stage7_51[1],stage7_50[2]}
   );
   gpc615_5 gpc9845 (
      {stage6_52[0], stage6_52[1], stage6_52[2], stage6_52[3], stage6_52[4]},
      {stage6_53[0]},
      {stage6_54[0], stage6_54[1], stage6_54[2], stage6_54[3], stage6_54[4], stage6_54[5]},
      {stage7_56[0],stage7_55[0],stage7_54[0],stage7_53[1],stage7_52[1]}
   );
   gpc615_5 gpc9846 (
      {stage6_55[0], stage6_55[1], stage6_55[2], stage6_55[3], stage6_55[4]},
      {stage6_56[0]},
      {stage6_57[0], stage6_57[1], stage6_57[2], stage6_57[3], stage6_57[4], stage6_57[5]},
      {stage7_59[0],stage7_58[0],stage7_57[0],stage7_56[1],stage7_55[1]}
   );
   gpc615_5 gpc9847 (
      {stage6_56[1], stage6_56[2], stage6_56[3], stage6_56[4], stage6_56[5]},
      {stage6_57[6]},
      {stage6_58[0], stage6_58[1], stage6_58[2], stage6_58[3], stage6_58[4], stage6_58[5]},
      {stage7_60[0],stage7_59[1],stage7_58[1],stage7_57[1],stage7_56[2]}
   );
   gpc135_4 gpc9848 (
      {stage6_61[0], stage6_61[1], stage6_61[2], stage6_61[3], stage6_61[4]},
      {stage6_62[0], stage6_62[1], stage6_62[2]},
      {stage6_63[0]},
      {stage7_64[0],stage7_63[0],stage7_62[0],stage7_61[0]}
   );
   gpc135_4 gpc9849 (
      {stage6_61[5], stage6_61[6], stage6_61[7], stage6_61[8], 1'b0},
      {stage6_62[3], stage6_62[4], stage6_62[5]},
      {stage6_63[1]},
      {stage7_64[1],stage7_63[1],stage7_62[1],stage7_61[1]}
   );
   gpc223_4 gpc9850 (
      {stage6_63[2], stage6_63[3], stage6_63[4]},
      {stage6_64[0], stage6_64[1]},
      {stage6_65[0], stage6_65[1]},
      {stage7_66[0],stage7_65[0],stage7_64[2],stage7_63[2]}
   );
   gpc7_3 gpc9851 (
      {stage6_64[2], stage6_64[3], stage6_64[4], stage6_64[5], stage6_64[6], stage6_64[7], stage6_64[8]},
      {stage7_66[1],stage7_65[1],stage7_64[3]}
   );
   gpc3_2 gpc9852 (
      {stage6_65[2], stage6_65[3], stage6_65[4]},
      {stage7_66[2],stage7_65[2]}
   );
   gpc1163_5 gpc9853 (
      {stage6_66[0], stage6_66[1], stage6_66[2]},
      {stage6_67[0], stage6_67[1], stage6_67[2], stage6_67[3], stage6_67[4], 1'b0},
      {stage6_68[0]},
      {stage6_69[0]},
      {stage7_70[0],stage7_69[0],stage7_68[0],stage7_67[0],stage7_66[3]}
   );
   gpc117_4 gpc9854 (
      {stage6_68[1], stage6_68[2], stage6_68[3], stage6_68[4], stage6_68[5], stage6_68[6], stage6_68[7]},
      {stage6_69[1]},
      {stage6_70[0]},
      {stage7_71[0],stage7_70[1],stage7_69[1],stage7_68[1]}
   );
   gpc117_4 gpc9855 (
      {stage6_68[8], stage6_68[9], stage6_68[10], stage6_68[11], stage6_68[12], stage6_68[13], stage6_68[14]},
      {stage6_69[2]},
      {1'b0},
      {stage7_71[1],stage7_70[2],stage7_69[2],stage7_68[2]}
   );
   gpc1_1 gpc9856 (
      {stage6_0[0]},
      {stage7_0[0]}
   );
   gpc1_1 gpc9857 (
      {stage6_0[1]},
      {stage7_0[1]}
   );
   gpc1_1 gpc9858 (
      {stage6_0[2]},
      {stage7_0[2]}
   );
   gpc1_1 gpc9859 (
      {stage6_0[3]},
      {stage7_0[3]}
   );
   gpc1_1 gpc9860 (
      {stage6_0[4]},
      {stage7_0[4]}
   );
   gpc1_1 gpc9861 (
      {stage6_1[0]},
      {stage7_1[0]}
   );
   gpc1_1 gpc9862 (
      {stage6_1[1]},
      {stage7_1[1]}
   );
   gpc1_1 gpc9863 (
      {stage6_2[0]},
      {stage7_2[0]}
   );
   gpc1_1 gpc9864 (
      {stage6_2[1]},
      {stage7_2[1]}
   );
   gpc1_1 gpc9865 (
      {stage6_2[2]},
      {stage7_2[2]}
   );
   gpc1_1 gpc9866 (
      {stage6_2[3]},
      {stage7_2[3]}
   );
   gpc1_1 gpc9867 (
      {stage6_2[4]},
      {stage7_2[4]}
   );
   gpc1_1 gpc9868 (
      {stage6_3[0]},
      {stage7_3[0]}
   );
   gpc1_1 gpc9869 (
      {stage6_3[1]},
      {stage7_3[1]}
   );
   gpc1_1 gpc9870 (
      {stage6_6[7]},
      {stage7_6[2]}
   );
   gpc1_1 gpc9871 (
      {stage6_8[4]},
      {stage7_8[3]}
   );
   gpc1_1 gpc9872 (
      {stage6_8[5]},
      {stage7_8[4]}
   );
   gpc1_1 gpc9873 (
      {stage6_9[6]},
      {stage7_9[2]}
   );
   gpc1_1 gpc9874 (
      {stage6_9[7]},
      {stage7_9[3]}
   );
   gpc1_1 gpc9875 (
      {stage6_9[8]},
      {stage7_9[4]}
   );
   gpc1_1 gpc9876 (
      {stage6_9[9]},
      {stage7_9[5]}
   );
   gpc1_1 gpc9877 (
      {stage6_11[6]},
      {stage7_11[3]}
   );
   gpc1_1 gpc9878 (
      {stage6_13[6]},
      {stage7_13[2]}
   );
   gpc1_1 gpc9879 (
      {stage6_13[7]},
      {stage7_13[3]}
   );
   gpc1_1 gpc9880 (
      {stage6_13[8]},
      {stage7_13[4]}
   );
   gpc1_1 gpc9881 (
      {stage6_13[9]},
      {stage7_13[5]}
   );
   gpc1_1 gpc9882 (
      {stage6_15[3]},
      {stage7_15[3]}
   );
   gpc1_1 gpc9883 (
      {stage6_15[4]},
      {stage7_15[4]}
   );
   gpc1_1 gpc9884 (
      {stage6_15[5]},
      {stage7_15[5]}
   );
   gpc1_1 gpc9885 (
      {stage6_19[0]},
      {stage7_19[2]}
   );
   gpc1_1 gpc9886 (
      {stage6_19[1]},
      {stage7_19[3]}
   );
   gpc1_1 gpc9887 (
      {stage6_19[2]},
      {stage7_19[4]}
   );
   gpc1_1 gpc9888 (
      {stage6_19[3]},
      {stage7_19[5]}
   );
   gpc1_1 gpc9889 (
      {stage6_19[4]},
      {stage7_19[6]}
   );
   gpc1_1 gpc9890 (
      {stage6_20[5]},
      {stage7_20[2]}
   );
   gpc1_1 gpc9891 (
      {stage6_21[1]},
      {stage7_21[1]}
   );
   gpc1_1 gpc9892 (
      {stage6_21[2]},
      {stage7_21[2]}
   );
   gpc1_1 gpc9893 (
      {stage6_21[3]},
      {stage7_21[3]}
   );
   gpc1_1 gpc9894 (
      {stage6_21[4]},
      {stage7_21[4]}
   );
   gpc1_1 gpc9895 (
      {stage6_21[5]},
      {stage7_21[5]}
   );
   gpc1_1 gpc9896 (
      {stage6_22[0]},
      {stage7_22[1]}
   );
   gpc1_1 gpc9897 (
      {stage6_22[1]},
      {stage7_22[2]}
   );
   gpc1_1 gpc9898 (
      {stage6_22[2]},
      {stage7_22[3]}
   );
   gpc1_1 gpc9899 (
      {stage6_22[3]},
      {stage7_22[4]}
   );
   gpc1_1 gpc9900 (
      {stage6_22[4]},
      {stage7_22[5]}
   );
   gpc1_1 gpc9901 (
      {stage6_22[5]},
      {stage7_22[6]}
   );
   gpc1_1 gpc9902 (
      {stage6_24[5]},
      {stage7_24[2]}
   );
   gpc1_1 gpc9903 (
      {stage6_24[6]},
      {stage7_24[3]}
   );
   gpc1_1 gpc9904 (
      {stage6_26[5]},
      {stage7_26[3]}
   );
   gpc1_1 gpc9905 (
      {stage6_26[6]},
      {stage7_26[4]}
   );
   gpc1_1 gpc9906 (
      {stage6_26[7]},
      {stage7_26[5]}
   );
   gpc1_1 gpc9907 (
      {stage6_27[1]},
      {stage7_27[1]}
   );
   gpc1_1 gpc9908 (
      {stage6_27[2]},
      {stage7_27[2]}
   );
   gpc1_1 gpc9909 (
      {stage6_27[3]},
      {stage7_27[3]}
   );
   gpc1_1 gpc9910 (
      {stage6_27[4]},
      {stage7_27[4]}
   );
   gpc1_1 gpc9911 (
      {stage6_29[3]},
      {stage7_29[2]}
   );
   gpc1_1 gpc9912 (
      {stage6_29[4]},
      {stage7_29[3]}
   );
   gpc1_1 gpc9913 (
      {stage6_29[5]},
      {stage7_29[4]}
   );
   gpc1_1 gpc9914 (
      {stage6_30[0]},
      {stage7_30[2]}
   );
   gpc1_1 gpc9915 (
      {stage6_30[1]},
      {stage7_30[3]}
   );
   gpc1_1 gpc9916 (
      {stage6_30[2]},
      {stage7_30[4]}
   );
   gpc1_1 gpc9917 (
      {stage6_30[3]},
      {stage7_30[5]}
   );
   gpc1_1 gpc9918 (
      {stage6_30[4]},
      {stage7_30[6]}
   );
   gpc1_1 gpc9919 (
      {stage6_31[5]},
      {stage7_31[1]}
   );
   gpc1_1 gpc9920 (
      {stage6_32[1]},
      {stage7_32[1]}
   );
   gpc1_1 gpc9921 (
      {stage6_32[2]},
      {stage7_32[2]}
   );
   gpc1_1 gpc9922 (
      {stage6_32[3]},
      {stage7_32[3]}
   );
   gpc1_1 gpc9923 (
      {stage6_32[4]},
      {stage7_32[4]}
   );
   gpc1_1 gpc9924 (
      {stage6_32[5]},
      {stage7_32[5]}
   );
   gpc1_1 gpc9925 (
      {stage6_34[5]},
      {stage7_34[2]}
   );
   gpc1_1 gpc9926 (
      {stage6_34[6]},
      {stage7_34[3]}
   );
   gpc1_1 gpc9927 (
      {stage6_34[7]},
      {stage7_34[4]}
   );
   gpc1_1 gpc9928 (
      {stage6_34[8]},
      {stage7_34[5]}
   );
   gpc1_1 gpc9929 (
      {stage6_35[1]},
      {stage7_35[2]}
   );
   gpc1_1 gpc9930 (
      {stage6_35[2]},
      {stage7_35[3]}
   );
   gpc1_1 gpc9931 (
      {stage6_35[3]},
      {stage7_35[4]}
   );
   gpc1_1 gpc9932 (
      {stage6_35[4]},
      {stage7_35[5]}
   );
   gpc1_1 gpc9933 (
      {stage6_38[0]},
      {stage7_38[2]}
   );
   gpc1_1 gpc9934 (
      {stage6_38[1]},
      {stage7_38[3]}
   );
   gpc1_1 gpc9935 (
      {stage6_38[2]},
      {stage7_38[4]}
   );
   gpc1_1 gpc9936 (
      {stage6_38[3]},
      {stage7_38[5]}
   );
   gpc1_1 gpc9937 (
      {stage6_38[4]},
      {stage7_38[6]}
   );
   gpc1_1 gpc9938 (
      {stage6_40[0]},
      {stage7_40[1]}
   );
   gpc1_1 gpc9939 (
      {stage6_40[1]},
      {stage7_40[2]}
   );
   gpc1_1 gpc9940 (
      {stage6_40[2]},
      {stage7_40[3]}
   );
   gpc1_1 gpc9941 (
      {stage6_40[3]},
      {stage7_40[4]}
   );
   gpc1_1 gpc9942 (
      {stage6_40[4]},
      {stage7_40[5]}
   );
   gpc1_1 gpc9943 (
      {stage6_40[5]},
      {stage7_40[6]}
   );
   gpc1_1 gpc9944 (
      {stage6_41[5]},
      {stage7_41[2]}
   );
   gpc1_1 gpc9945 (
      {stage6_41[6]},
      {stage7_41[3]}
   );
   gpc1_1 gpc9946 (
      {stage6_41[7]},
      {stage7_41[4]}
   );
   gpc1_1 gpc9947 (
      {stage6_42[6]},
      {stage7_42[2]}
   );
   gpc1_1 gpc9948 (
      {stage6_43[6]},
      {stage7_43[3]}
   );
   gpc1_1 gpc9949 (
      {stage6_45[6]},
      {stage7_45[2]}
   );
   gpc1_1 gpc9950 (
      {stage6_45[7]},
      {stage7_45[3]}
   );
   gpc1_1 gpc9951 (
      {stage6_45[8]},
      {stage7_45[4]}
   );
   gpc1_1 gpc9952 (
      {stage6_47[1]},
      {stage7_47[2]}
   );
   gpc1_1 gpc9953 (
      {stage6_47[2]},
      {stage7_47[3]}
   );
   gpc1_1 gpc9954 (
      {stage6_47[3]},
      {stage7_47[4]}
   );
   gpc1_1 gpc9955 (
      {stage6_47[4]},
      {stage7_47[5]}
   );
   gpc1_1 gpc9956 (
      {stage6_47[5]},
      {stage7_47[6]}
   );
   gpc1_1 gpc9957 (
      {stage6_47[6]},
      {stage7_47[7]}
   );
   gpc1_1 gpc9958 (
      {stage6_51[6]},
      {stage7_51[2]}
   );
   gpc1_1 gpc9959 (
      {stage6_51[7]},
      {stage7_51[3]}
   );
   gpc1_1 gpc9960 (
      {stage6_52[5]},
      {stage7_52[2]}
   );
   gpc1_1 gpc9961 (
      {stage6_52[6]},
      {stage7_52[3]}
   );
   gpc1_1 gpc9962 (
      {stage6_53[1]},
      {stage7_53[2]}
   );
   gpc1_1 gpc9963 (
      {stage6_53[2]},
      {stage7_53[3]}
   );
   gpc1_1 gpc9964 (
      {stage6_53[3]},
      {stage7_53[4]}
   );
   gpc1_1 gpc9965 (
      {stage6_53[4]},
      {stage7_53[5]}
   );
   gpc1_1 gpc9966 (
      {stage6_55[5]},
      {stage7_55[2]}
   );
   gpc1_1 gpc9967 (
      {stage6_55[6]},
      {stage7_55[3]}
   );
   gpc1_1 gpc9968 (
      {stage6_55[7]},
      {stage7_55[4]}
   );
   gpc1_1 gpc9969 (
      {stage6_55[8]},
      {stage7_55[5]}
   );
   gpc1_1 gpc9970 (
      {stage6_55[9]},
      {stage7_55[6]}
   );
   gpc1_1 gpc9971 (
      {stage6_56[6]},
      {stage7_56[3]}
   );
   gpc1_1 gpc9972 (
      {stage6_56[7]},
      {stage7_56[4]}
   );
   gpc1_1 gpc9973 (
      {stage6_56[8]},
      {stage7_56[5]}
   );
   gpc1_1 gpc9974 (
      {stage6_56[9]},
      {stage7_56[6]}
   );
   gpc1_1 gpc9975 (
      {stage6_59[0]},
      {stage7_59[2]}
   );
   gpc1_1 gpc9976 (
      {stage6_59[1]},
      {stage7_59[3]}
   );
   gpc1_1 gpc9977 (
      {stage6_59[2]},
      {stage7_59[4]}
   );
   gpc1_1 gpc9978 (
      {stage6_59[3]},
      {stage7_59[5]}
   );
   gpc1_1 gpc9979 (
      {stage6_59[4]},
      {stage7_59[6]}
   );
   gpc1_1 gpc9980 (
      {stage6_60[0]},
      {stage7_60[1]}
   );
   gpc1_1 gpc9981 (
      {stage6_60[1]},
      {stage7_60[2]}
   );
   gpc1_1 gpc9982 (
      {stage6_60[2]},
      {stage7_60[3]}
   );
   gpc1_1 gpc9983 (
      {stage6_60[3]},
      {stage7_60[4]}
   );
   gpc1_1 gpc9984 (
      {stage6_60[4]},
      {stage7_60[5]}
   );
   gpc1_1 gpc9985 (
      {stage6_66[3]},
      {stage7_66[4]}
   );
   gpc1_1 gpc9986 (
      {stage6_66[4]},
      {stage7_66[5]}
   );
   gpc1_1 gpc9987 (
      {stage6_68[15]},
      {stage7_68[3]}
   );
   gpc1_1 gpc9988 (
      {stage6_68[16]},
      {stage7_68[4]}
   );
   gpc1_1 gpc9989 (
      {stage6_69[3]},
      {stage7_69[3]}
   );
   gpc1_1 gpc9990 (
      {stage6_69[4]},
      {stage7_69[4]}
   );
   gpc1415_5 gpc9991 (
      {stage7_0[0], stage7_0[1], stage7_0[2], stage7_0[3], stage7_0[4]},
      {stage7_1[0]},
      {stage7_2[0], stage7_2[1], stage7_2[2], stage7_2[3]},
      {stage7_3[0]},
      {stage8_4[0],stage8_3[0],stage8_2[0],stage8_1[0],stage8_0[0]}
   );
   gpc3_2 gpc9992 (
      {stage7_6[0], stage7_6[1], stage7_6[2]},
      {stage8_7[0],stage8_6[0]}
   );
   gpc3_2 gpc9993 (
      {stage7_7[0], stage7_7[1], stage7_7[2]},
      {stage8_8[0],stage8_7[1]}
   );
   gpc215_4 gpc9994 (
      {stage7_8[0], stage7_8[1], stage7_8[2], stage7_8[3], stage7_8[4]},
      {stage7_9[0]},
      {stage7_10[0], stage7_10[1]},
      {stage8_11[0],stage8_10[0],stage8_9[0],stage8_8[1]}
   );
   gpc1415_5 gpc9995 (
      {stage7_9[1], stage7_9[2], stage7_9[3], stage7_9[4], stage7_9[5]},
      {1'b0},
      {stage7_11[0], stage7_11[1], stage7_11[2], stage7_11[3]},
      {stage7_12[0]},
      {stage8_13[0],stage8_12[0],stage8_11[1],stage8_10[1],stage8_9[1]}
   );
   gpc207_4 gpc9996 (
      {stage7_13[0], stage7_13[1], stage7_13[2], stage7_13[3], stage7_13[4], stage7_13[5], 1'b0},
      {stage7_15[0], stage7_15[1]},
      {stage8_16[0],stage8_15[0],stage8_14[0],stage8_13[1]}
   );
   gpc1343_5 gpc9997 (
      {stage7_14[0], stage7_14[1], stage7_14[2]},
      {stage7_15[2], stage7_15[3], stage7_15[4], stage7_15[5]},
      {stage7_16[0], stage7_16[1], stage7_16[2]},
      {stage7_17[0]},
      {stage8_18[0],stage8_17[0],stage8_16[1],stage8_15[1],stage8_14[1]}
   );
   gpc623_5 gpc9998 (
      {stage7_17[1], 1'b0, 1'b0},
      {stage7_18[0], stage7_18[1]},
      {stage7_19[0], stage7_19[1], stage7_19[2], stage7_19[3], stage7_19[4], stage7_19[5]},
      {stage8_21[0],stage8_20[0],stage8_19[0],stage8_18[1],stage8_17[1]}
   );
   gpc1163_5 gpc9999 (
      {stage7_20[0], stage7_20[1], stage7_20[2]},
      {stage7_21[0], stage7_21[1], stage7_21[2], stage7_21[3], stage7_21[4], stage7_21[5]},
      {stage7_22[0]},
      {stage7_23[0]},
      {stage8_24[0],stage8_23[0],stage8_22[0],stage8_21[1],stage8_20[1]}
   );
   gpc1406_5 gpc10000 (
      {stage7_22[1], stage7_22[2], stage7_22[3], stage7_22[4], stage7_22[5], stage7_22[6]},
      {stage7_24[0], stage7_24[1], stage7_24[2], stage7_24[3]},
      {stage7_25[0]},
      {stage8_26[0],stage8_25[0],stage8_24[1],stage8_23[1],stage8_22[1]}
   );
   gpc7_3 gpc10001 (
      {stage7_26[0], stage7_26[1], stage7_26[2], stage7_26[3], stage7_26[4], stage7_26[5], 1'b0},
      {stage8_28[0],stage8_27[0],stage8_26[1]}
   );
   gpc15_3 gpc10002 (
      {stage7_27[0], stage7_27[1], stage7_27[2], stage7_27[3], stage7_27[4]},
      {stage7_28[0]},
      {stage8_29[0],stage8_28[1],stage8_27[1]}
   );
   gpc135_4 gpc10003 (
      {stage7_29[0], stage7_29[1], stage7_29[2], stage7_29[3], stage7_29[4]},
      {stage7_30[0], stage7_30[1], stage7_30[2]},
      {stage7_31[0]},
      {stage8_32[0],stage8_31[0],stage8_30[0],stage8_29[1]}
   );
   gpc615_5 gpc10004 (
      {stage7_30[3], stage7_30[4], stage7_30[5], stage7_30[6], 1'b0},
      {stage7_31[1]},
      {stage7_32[0], stage7_32[1], stage7_32[2], stage7_32[3], stage7_32[4], stage7_32[5]},
      {stage8_34[0],stage8_33[0],stage8_32[1],stage8_31[1],stage8_30[1]}
   );
   gpc7_3 gpc10005 (
      {stage7_34[0], stage7_34[1], stage7_34[2], stage7_34[3], stage7_34[4], stage7_34[5], 1'b0},
      {stage8_36[0],stage8_35[0],stage8_34[1]}
   );
   gpc117_4 gpc10006 (
      {stage7_35[0], stage7_35[1], stage7_35[2], stage7_35[3], stage7_35[4], stage7_35[5], 1'b0},
      {stage7_36[0]},
      {stage7_37[0]},
      {stage8_38[0],stage8_37[0],stage8_36[1],stage8_35[1]}
   );
   gpc7_3 gpc10007 (
      {stage7_38[0], stage7_38[1], stage7_38[2], stage7_38[3], stage7_38[4], stage7_38[5], stage7_38[6]},
      {stage8_40[0],stage8_39[0],stage8_38[1]}
   );
   gpc207_4 gpc10008 (
      {stage7_40[0], stage7_40[1], stage7_40[2], stage7_40[3], stage7_40[4], stage7_40[5], stage7_40[6]},
      {stage7_42[0], stage7_42[1]},
      {stage8_43[0],stage8_42[0],stage8_41[0],stage8_40[1]}
   );
   gpc1415_5 gpc10009 (
      {stage7_41[0], stage7_41[1], stage7_41[2], stage7_41[3], stage7_41[4]},
      {stage7_42[2]},
      {stage7_43[0], stage7_43[1], stage7_43[2], stage7_43[3]},
      {stage7_44[0]},
      {stage8_45[0],stage8_44[0],stage8_43[1],stage8_42[1],stage8_41[1]}
   );
   gpc2135_5 gpc10010 (
      {stage7_45[0], stage7_45[1], stage7_45[2], stage7_45[3], stage7_45[4]},
      {stage7_46[0], stage7_46[1], stage7_46[2]},
      {stage7_47[0]},
      {stage7_48[0], 1'b0},
      {stage8_49[0],stage8_48[0],stage8_47[0],stage8_46[0],stage8_45[1]}
   );
   gpc207_4 gpc10011 (
      {stage7_47[1], stage7_47[2], stage7_47[3], stage7_47[4], stage7_47[5], stage7_47[6], stage7_47[7]},
      {stage7_49[0], stage7_49[1]},
      {stage8_50[0],stage8_49[1],stage8_48[1],stage8_47[1]}
   );
   gpc3_2 gpc10012 (
      {stage7_50[0], stage7_50[1], stage7_50[2]},
      {stage8_51[0],stage8_50[1]}
   );
   gpc615_5 gpc10013 (
      {stage7_51[0], stage7_51[1], stage7_51[2], stage7_51[3], 1'b0},
      {stage7_52[0]},
      {stage7_53[0], stage7_53[1], stage7_53[2], stage7_53[3], stage7_53[4], stage7_53[5]},
      {stage8_55[0],stage8_54[0],stage8_53[0],stage8_52[0],stage8_51[1]}
   );
   gpc3_2 gpc10014 (
      {stage7_52[1], stage7_52[2], stage7_52[3]},
      {stage8_53[1],stage8_52[1]}
   );
   gpc207_4 gpc10015 (
      {stage7_55[0], stage7_55[1], stage7_55[2], stage7_55[3], stage7_55[4], stage7_55[5], stage7_55[6]},
      {stage7_57[0], stage7_57[1]},
      {stage8_58[0],stage8_57[0],stage8_56[0],stage8_55[1]}
   );
   gpc207_4 gpc10016 (
      {stage7_56[0], stage7_56[1], stage7_56[2], stage7_56[3], stage7_56[4], stage7_56[5], stage7_56[6]},
      {stage7_58[0], stage7_58[1]},
      {stage8_59[0],stage8_58[1],stage8_57[1],stage8_56[1]}
   );
   gpc117_4 gpc10017 (
      {stage7_59[0], stage7_59[1], stage7_59[2], stage7_59[3], stage7_59[4], stage7_59[5], stage7_59[6]},
      {stage7_60[0]},
      {stage7_61[0]},
      {stage8_62[0],stage8_61[0],stage8_60[0],stage8_59[1]}
   );
   gpc215_4 gpc10018 (
      {stage7_60[1], stage7_60[2], stage7_60[3], stage7_60[4], stage7_60[5]},
      {stage7_61[1]},
      {stage7_62[0], stage7_62[1]},
      {stage8_63[0],stage8_62[1],stage8_61[1],stage8_60[1]}
   );
   gpc3_2 gpc10019 (
      {stage7_63[0], stage7_63[1], stage7_63[2]},
      {stage8_64[0],stage8_63[1]}
   );
   gpc606_5 gpc10020 (
      {stage7_64[0], stage7_64[1], stage7_64[2], stage7_64[3], 1'b0, 1'b0},
      {stage7_66[0], stage7_66[1], stage7_66[2], stage7_66[3], stage7_66[4], stage7_66[5]},
      {stage8_68[0],stage8_67[0],stage8_66[0],stage8_65[0],stage8_64[1]}
   );
   gpc3_2 gpc10021 (
      {stage7_65[0], stage7_65[1], stage7_65[2]},
      {stage8_66[1],stage8_65[1]}
   );
   gpc615_5 gpc10022 (
      {stage7_68[0], stage7_68[1], stage7_68[2], stage7_68[3], stage7_68[4]},
      {stage7_69[0]},
      {stage7_70[0], stage7_70[1], stage7_70[2], 1'b0, 1'b0, 1'b0},
      {stage8_72[0],stage8_71[0],stage8_70[0],stage8_69[0],stage8_68[1]}
   );
   gpc606_5 gpc10023 (
      {stage7_69[1], stage7_69[2], stage7_69[3], stage7_69[4], 1'b0, 1'b0},
      {stage7_71[0], stage7_71[1], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage8_72[1],stage8_71[1],stage8_70[1],stage8_69[1]}
   );
   gpc1_1 gpc10024 (
      {stage7_1[1]},
      {stage8_1[1]}
   );
   gpc1_1 gpc10025 (
      {stage7_2[4]},
      {stage8_2[1]}
   );
   gpc1_1 gpc10026 (
      {stage7_3[1]},
      {stage8_3[1]}
   );
   gpc1_1 gpc10027 (
      {stage7_4[0]},
      {stage8_4[1]}
   );
   gpc1_1 gpc10028 (
      {stage7_5[0]},
      {stage8_5[0]}
   );
   gpc1_1 gpc10029 (
      {stage7_5[1]},
      {stage8_5[1]}
   );
   gpc1_1 gpc10030 (
      {stage7_12[1]},
      {stage8_12[1]}
   );
   gpc1_1 gpc10031 (
      {stage7_19[6]},
      {stage8_19[1]}
   );
   gpc1_1 gpc10032 (
      {stage7_25[1]},
      {stage8_25[1]}
   );
   gpc1_1 gpc10033 (
      {stage7_33[0]},
      {stage8_33[1]}
   );
   gpc1_1 gpc10034 (
      {stage7_37[1]},
      {stage8_37[1]}
   );
   gpc1_1 gpc10035 (
      {stage7_39[0]},
      {stage8_39[1]}
   );
   gpc1_1 gpc10036 (
      {stage7_44[1]},
      {stage8_44[1]}
   );
   gpc1_1 gpc10037 (
      {stage7_54[0]},
      {stage8_54[1]}
   );
   gpc1_1 gpc10038 (
      {stage7_67[0]},
      {stage8_67[1]}
   );
endmodule

module testbench();
    reg [485:0] src0;
    reg [485:0] src1;
    reg [485:0] src2;
    reg [485:0] src3;
    reg [485:0] src4;
    reg [485:0] src5;
    reg [485:0] src6;
    reg [485:0] src7;
    reg [485:0] src8;
    reg [485:0] src9;
    reg [485:0] src10;
    reg [485:0] src11;
    reg [485:0] src12;
    reg [485:0] src13;
    reg [485:0] src14;
    reg [485:0] src15;
    reg [485:0] src16;
    reg [485:0] src17;
    reg [485:0] src18;
    reg [485:0] src19;
    reg [485:0] src20;
    reg [485:0] src21;
    reg [485:0] src22;
    reg [485:0] src23;
    reg [485:0] src24;
    reg [485:0] src25;
    reg [485:0] src26;
    reg [485:0] src27;
    reg [485:0] src28;
    reg [485:0] src29;
    reg [485:0] src30;
    reg [485:0] src31;
    reg [485:0] src32;
    reg [485:0] src33;
    reg [485:0] src34;
    reg [485:0] src35;
    reg [485:0] src36;
    reg [485:0] src37;
    reg [485:0] src38;
    reg [485:0] src39;
    reg [485:0] src40;
    reg [485:0] src41;
    reg [485:0] src42;
    reg [485:0] src43;
    reg [485:0] src44;
    reg [485:0] src45;
    reg [485:0] src46;
    reg [485:0] src47;
    reg [485:0] src48;
    reg [485:0] src49;
    reg [485:0] src50;
    reg [485:0] src51;
    reg [485:0] src52;
    reg [485:0] src53;
    reg [485:0] src54;
    reg [485:0] src55;
    reg [485:0] src56;
    reg [485:0] src57;
    reg [485:0] src58;
    reg [485:0] src59;
    reg [485:0] src60;
    reg [485:0] src61;
    reg [485:0] src62;
    reg [485:0] src63;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [0:0] dst63;
    wire [0:0] dst64;
    wire [0:0] dst65;
    wire [0:0] dst66;
    wire [0:0] dst67;
    wire [0:0] dst68;
    wire [0:0] dst69;
    wire [0:0] dst70;
    wire [0:0] dst71;
    wire [0:0] dst72;
    wire [72:0] srcsum;
    wire [72:0] dstsum;
    wire test;
    compressor_CLA486_64 compressor_CLA486_64(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62),
        .dst63(dst63),
        .dst64(dst64),
        .dst65(dst65),
        .dst66(dst66),
        .dst67(dst67),
        .dst68(dst68),
        .dst69(dst69),
        .dst70(dst70),
        .dst71(dst71),
        .dst72(dst72));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255] + src0[256] + src0[257] + src0[258] + src0[259] + src0[260] + src0[261] + src0[262] + src0[263] + src0[264] + src0[265] + src0[266] + src0[267] + src0[268] + src0[269] + src0[270] + src0[271] + src0[272] + src0[273] + src0[274] + src0[275] + src0[276] + src0[277] + src0[278] + src0[279] + src0[280] + src0[281] + src0[282] + src0[283] + src0[284] + src0[285] + src0[286] + src0[287] + src0[288] + src0[289] + src0[290] + src0[291] + src0[292] + src0[293] + src0[294] + src0[295] + src0[296] + src0[297] + src0[298] + src0[299] + src0[300] + src0[301] + src0[302] + src0[303] + src0[304] + src0[305] + src0[306] + src0[307] + src0[308] + src0[309] + src0[310] + src0[311] + src0[312] + src0[313] + src0[314] + src0[315] + src0[316] + src0[317] + src0[318] + src0[319] + src0[320] + src0[321] + src0[322] + src0[323] + src0[324] + src0[325] + src0[326] + src0[327] + src0[328] + src0[329] + src0[330] + src0[331] + src0[332] + src0[333] + src0[334] + src0[335] + src0[336] + src0[337] + src0[338] + src0[339] + src0[340] + src0[341] + src0[342] + src0[343] + src0[344] + src0[345] + src0[346] + src0[347] + src0[348] + src0[349] + src0[350] + src0[351] + src0[352] + src0[353] + src0[354] + src0[355] + src0[356] + src0[357] + src0[358] + src0[359] + src0[360] + src0[361] + src0[362] + src0[363] + src0[364] + src0[365] + src0[366] + src0[367] + src0[368] + src0[369] + src0[370] + src0[371] + src0[372] + src0[373] + src0[374] + src0[375] + src0[376] + src0[377] + src0[378] + src0[379] + src0[380] + src0[381] + src0[382] + src0[383] + src0[384] + src0[385] + src0[386] + src0[387] + src0[388] + src0[389] + src0[390] + src0[391] + src0[392] + src0[393] + src0[394] + src0[395] + src0[396] + src0[397] + src0[398] + src0[399] + src0[400] + src0[401] + src0[402] + src0[403] + src0[404] + src0[405] + src0[406] + src0[407] + src0[408] + src0[409] + src0[410] + src0[411] + src0[412] + src0[413] + src0[414] + src0[415] + src0[416] + src0[417] + src0[418] + src0[419] + src0[420] + src0[421] + src0[422] + src0[423] + src0[424] + src0[425] + src0[426] + src0[427] + src0[428] + src0[429] + src0[430] + src0[431] + src0[432] + src0[433] + src0[434] + src0[435] + src0[436] + src0[437] + src0[438] + src0[439] + src0[440] + src0[441] + src0[442] + src0[443] + src0[444] + src0[445] + src0[446] + src0[447] + src0[448] + src0[449] + src0[450] + src0[451] + src0[452] + src0[453] + src0[454] + src0[455] + src0[456] + src0[457] + src0[458] + src0[459] + src0[460] + src0[461] + src0[462] + src0[463] + src0[464] + src0[465] + src0[466] + src0[467] + src0[468] + src0[469] + src0[470] + src0[471] + src0[472] + src0[473] + src0[474] + src0[475] + src0[476] + src0[477] + src0[478] + src0[479] + src0[480] + src0[481] + src0[482] + src0[483] + src0[484] + src0[485])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255] + src1[256] + src1[257] + src1[258] + src1[259] + src1[260] + src1[261] + src1[262] + src1[263] + src1[264] + src1[265] + src1[266] + src1[267] + src1[268] + src1[269] + src1[270] + src1[271] + src1[272] + src1[273] + src1[274] + src1[275] + src1[276] + src1[277] + src1[278] + src1[279] + src1[280] + src1[281] + src1[282] + src1[283] + src1[284] + src1[285] + src1[286] + src1[287] + src1[288] + src1[289] + src1[290] + src1[291] + src1[292] + src1[293] + src1[294] + src1[295] + src1[296] + src1[297] + src1[298] + src1[299] + src1[300] + src1[301] + src1[302] + src1[303] + src1[304] + src1[305] + src1[306] + src1[307] + src1[308] + src1[309] + src1[310] + src1[311] + src1[312] + src1[313] + src1[314] + src1[315] + src1[316] + src1[317] + src1[318] + src1[319] + src1[320] + src1[321] + src1[322] + src1[323] + src1[324] + src1[325] + src1[326] + src1[327] + src1[328] + src1[329] + src1[330] + src1[331] + src1[332] + src1[333] + src1[334] + src1[335] + src1[336] + src1[337] + src1[338] + src1[339] + src1[340] + src1[341] + src1[342] + src1[343] + src1[344] + src1[345] + src1[346] + src1[347] + src1[348] + src1[349] + src1[350] + src1[351] + src1[352] + src1[353] + src1[354] + src1[355] + src1[356] + src1[357] + src1[358] + src1[359] + src1[360] + src1[361] + src1[362] + src1[363] + src1[364] + src1[365] + src1[366] + src1[367] + src1[368] + src1[369] + src1[370] + src1[371] + src1[372] + src1[373] + src1[374] + src1[375] + src1[376] + src1[377] + src1[378] + src1[379] + src1[380] + src1[381] + src1[382] + src1[383] + src1[384] + src1[385] + src1[386] + src1[387] + src1[388] + src1[389] + src1[390] + src1[391] + src1[392] + src1[393] + src1[394] + src1[395] + src1[396] + src1[397] + src1[398] + src1[399] + src1[400] + src1[401] + src1[402] + src1[403] + src1[404] + src1[405] + src1[406] + src1[407] + src1[408] + src1[409] + src1[410] + src1[411] + src1[412] + src1[413] + src1[414] + src1[415] + src1[416] + src1[417] + src1[418] + src1[419] + src1[420] + src1[421] + src1[422] + src1[423] + src1[424] + src1[425] + src1[426] + src1[427] + src1[428] + src1[429] + src1[430] + src1[431] + src1[432] + src1[433] + src1[434] + src1[435] + src1[436] + src1[437] + src1[438] + src1[439] + src1[440] + src1[441] + src1[442] + src1[443] + src1[444] + src1[445] + src1[446] + src1[447] + src1[448] + src1[449] + src1[450] + src1[451] + src1[452] + src1[453] + src1[454] + src1[455] + src1[456] + src1[457] + src1[458] + src1[459] + src1[460] + src1[461] + src1[462] + src1[463] + src1[464] + src1[465] + src1[466] + src1[467] + src1[468] + src1[469] + src1[470] + src1[471] + src1[472] + src1[473] + src1[474] + src1[475] + src1[476] + src1[477] + src1[478] + src1[479] + src1[480] + src1[481] + src1[482] + src1[483] + src1[484] + src1[485])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255] + src2[256] + src2[257] + src2[258] + src2[259] + src2[260] + src2[261] + src2[262] + src2[263] + src2[264] + src2[265] + src2[266] + src2[267] + src2[268] + src2[269] + src2[270] + src2[271] + src2[272] + src2[273] + src2[274] + src2[275] + src2[276] + src2[277] + src2[278] + src2[279] + src2[280] + src2[281] + src2[282] + src2[283] + src2[284] + src2[285] + src2[286] + src2[287] + src2[288] + src2[289] + src2[290] + src2[291] + src2[292] + src2[293] + src2[294] + src2[295] + src2[296] + src2[297] + src2[298] + src2[299] + src2[300] + src2[301] + src2[302] + src2[303] + src2[304] + src2[305] + src2[306] + src2[307] + src2[308] + src2[309] + src2[310] + src2[311] + src2[312] + src2[313] + src2[314] + src2[315] + src2[316] + src2[317] + src2[318] + src2[319] + src2[320] + src2[321] + src2[322] + src2[323] + src2[324] + src2[325] + src2[326] + src2[327] + src2[328] + src2[329] + src2[330] + src2[331] + src2[332] + src2[333] + src2[334] + src2[335] + src2[336] + src2[337] + src2[338] + src2[339] + src2[340] + src2[341] + src2[342] + src2[343] + src2[344] + src2[345] + src2[346] + src2[347] + src2[348] + src2[349] + src2[350] + src2[351] + src2[352] + src2[353] + src2[354] + src2[355] + src2[356] + src2[357] + src2[358] + src2[359] + src2[360] + src2[361] + src2[362] + src2[363] + src2[364] + src2[365] + src2[366] + src2[367] + src2[368] + src2[369] + src2[370] + src2[371] + src2[372] + src2[373] + src2[374] + src2[375] + src2[376] + src2[377] + src2[378] + src2[379] + src2[380] + src2[381] + src2[382] + src2[383] + src2[384] + src2[385] + src2[386] + src2[387] + src2[388] + src2[389] + src2[390] + src2[391] + src2[392] + src2[393] + src2[394] + src2[395] + src2[396] + src2[397] + src2[398] + src2[399] + src2[400] + src2[401] + src2[402] + src2[403] + src2[404] + src2[405] + src2[406] + src2[407] + src2[408] + src2[409] + src2[410] + src2[411] + src2[412] + src2[413] + src2[414] + src2[415] + src2[416] + src2[417] + src2[418] + src2[419] + src2[420] + src2[421] + src2[422] + src2[423] + src2[424] + src2[425] + src2[426] + src2[427] + src2[428] + src2[429] + src2[430] + src2[431] + src2[432] + src2[433] + src2[434] + src2[435] + src2[436] + src2[437] + src2[438] + src2[439] + src2[440] + src2[441] + src2[442] + src2[443] + src2[444] + src2[445] + src2[446] + src2[447] + src2[448] + src2[449] + src2[450] + src2[451] + src2[452] + src2[453] + src2[454] + src2[455] + src2[456] + src2[457] + src2[458] + src2[459] + src2[460] + src2[461] + src2[462] + src2[463] + src2[464] + src2[465] + src2[466] + src2[467] + src2[468] + src2[469] + src2[470] + src2[471] + src2[472] + src2[473] + src2[474] + src2[475] + src2[476] + src2[477] + src2[478] + src2[479] + src2[480] + src2[481] + src2[482] + src2[483] + src2[484] + src2[485])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255] + src3[256] + src3[257] + src3[258] + src3[259] + src3[260] + src3[261] + src3[262] + src3[263] + src3[264] + src3[265] + src3[266] + src3[267] + src3[268] + src3[269] + src3[270] + src3[271] + src3[272] + src3[273] + src3[274] + src3[275] + src3[276] + src3[277] + src3[278] + src3[279] + src3[280] + src3[281] + src3[282] + src3[283] + src3[284] + src3[285] + src3[286] + src3[287] + src3[288] + src3[289] + src3[290] + src3[291] + src3[292] + src3[293] + src3[294] + src3[295] + src3[296] + src3[297] + src3[298] + src3[299] + src3[300] + src3[301] + src3[302] + src3[303] + src3[304] + src3[305] + src3[306] + src3[307] + src3[308] + src3[309] + src3[310] + src3[311] + src3[312] + src3[313] + src3[314] + src3[315] + src3[316] + src3[317] + src3[318] + src3[319] + src3[320] + src3[321] + src3[322] + src3[323] + src3[324] + src3[325] + src3[326] + src3[327] + src3[328] + src3[329] + src3[330] + src3[331] + src3[332] + src3[333] + src3[334] + src3[335] + src3[336] + src3[337] + src3[338] + src3[339] + src3[340] + src3[341] + src3[342] + src3[343] + src3[344] + src3[345] + src3[346] + src3[347] + src3[348] + src3[349] + src3[350] + src3[351] + src3[352] + src3[353] + src3[354] + src3[355] + src3[356] + src3[357] + src3[358] + src3[359] + src3[360] + src3[361] + src3[362] + src3[363] + src3[364] + src3[365] + src3[366] + src3[367] + src3[368] + src3[369] + src3[370] + src3[371] + src3[372] + src3[373] + src3[374] + src3[375] + src3[376] + src3[377] + src3[378] + src3[379] + src3[380] + src3[381] + src3[382] + src3[383] + src3[384] + src3[385] + src3[386] + src3[387] + src3[388] + src3[389] + src3[390] + src3[391] + src3[392] + src3[393] + src3[394] + src3[395] + src3[396] + src3[397] + src3[398] + src3[399] + src3[400] + src3[401] + src3[402] + src3[403] + src3[404] + src3[405] + src3[406] + src3[407] + src3[408] + src3[409] + src3[410] + src3[411] + src3[412] + src3[413] + src3[414] + src3[415] + src3[416] + src3[417] + src3[418] + src3[419] + src3[420] + src3[421] + src3[422] + src3[423] + src3[424] + src3[425] + src3[426] + src3[427] + src3[428] + src3[429] + src3[430] + src3[431] + src3[432] + src3[433] + src3[434] + src3[435] + src3[436] + src3[437] + src3[438] + src3[439] + src3[440] + src3[441] + src3[442] + src3[443] + src3[444] + src3[445] + src3[446] + src3[447] + src3[448] + src3[449] + src3[450] + src3[451] + src3[452] + src3[453] + src3[454] + src3[455] + src3[456] + src3[457] + src3[458] + src3[459] + src3[460] + src3[461] + src3[462] + src3[463] + src3[464] + src3[465] + src3[466] + src3[467] + src3[468] + src3[469] + src3[470] + src3[471] + src3[472] + src3[473] + src3[474] + src3[475] + src3[476] + src3[477] + src3[478] + src3[479] + src3[480] + src3[481] + src3[482] + src3[483] + src3[484] + src3[485])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255] + src4[256] + src4[257] + src4[258] + src4[259] + src4[260] + src4[261] + src4[262] + src4[263] + src4[264] + src4[265] + src4[266] + src4[267] + src4[268] + src4[269] + src4[270] + src4[271] + src4[272] + src4[273] + src4[274] + src4[275] + src4[276] + src4[277] + src4[278] + src4[279] + src4[280] + src4[281] + src4[282] + src4[283] + src4[284] + src4[285] + src4[286] + src4[287] + src4[288] + src4[289] + src4[290] + src4[291] + src4[292] + src4[293] + src4[294] + src4[295] + src4[296] + src4[297] + src4[298] + src4[299] + src4[300] + src4[301] + src4[302] + src4[303] + src4[304] + src4[305] + src4[306] + src4[307] + src4[308] + src4[309] + src4[310] + src4[311] + src4[312] + src4[313] + src4[314] + src4[315] + src4[316] + src4[317] + src4[318] + src4[319] + src4[320] + src4[321] + src4[322] + src4[323] + src4[324] + src4[325] + src4[326] + src4[327] + src4[328] + src4[329] + src4[330] + src4[331] + src4[332] + src4[333] + src4[334] + src4[335] + src4[336] + src4[337] + src4[338] + src4[339] + src4[340] + src4[341] + src4[342] + src4[343] + src4[344] + src4[345] + src4[346] + src4[347] + src4[348] + src4[349] + src4[350] + src4[351] + src4[352] + src4[353] + src4[354] + src4[355] + src4[356] + src4[357] + src4[358] + src4[359] + src4[360] + src4[361] + src4[362] + src4[363] + src4[364] + src4[365] + src4[366] + src4[367] + src4[368] + src4[369] + src4[370] + src4[371] + src4[372] + src4[373] + src4[374] + src4[375] + src4[376] + src4[377] + src4[378] + src4[379] + src4[380] + src4[381] + src4[382] + src4[383] + src4[384] + src4[385] + src4[386] + src4[387] + src4[388] + src4[389] + src4[390] + src4[391] + src4[392] + src4[393] + src4[394] + src4[395] + src4[396] + src4[397] + src4[398] + src4[399] + src4[400] + src4[401] + src4[402] + src4[403] + src4[404] + src4[405] + src4[406] + src4[407] + src4[408] + src4[409] + src4[410] + src4[411] + src4[412] + src4[413] + src4[414] + src4[415] + src4[416] + src4[417] + src4[418] + src4[419] + src4[420] + src4[421] + src4[422] + src4[423] + src4[424] + src4[425] + src4[426] + src4[427] + src4[428] + src4[429] + src4[430] + src4[431] + src4[432] + src4[433] + src4[434] + src4[435] + src4[436] + src4[437] + src4[438] + src4[439] + src4[440] + src4[441] + src4[442] + src4[443] + src4[444] + src4[445] + src4[446] + src4[447] + src4[448] + src4[449] + src4[450] + src4[451] + src4[452] + src4[453] + src4[454] + src4[455] + src4[456] + src4[457] + src4[458] + src4[459] + src4[460] + src4[461] + src4[462] + src4[463] + src4[464] + src4[465] + src4[466] + src4[467] + src4[468] + src4[469] + src4[470] + src4[471] + src4[472] + src4[473] + src4[474] + src4[475] + src4[476] + src4[477] + src4[478] + src4[479] + src4[480] + src4[481] + src4[482] + src4[483] + src4[484] + src4[485])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255] + src5[256] + src5[257] + src5[258] + src5[259] + src5[260] + src5[261] + src5[262] + src5[263] + src5[264] + src5[265] + src5[266] + src5[267] + src5[268] + src5[269] + src5[270] + src5[271] + src5[272] + src5[273] + src5[274] + src5[275] + src5[276] + src5[277] + src5[278] + src5[279] + src5[280] + src5[281] + src5[282] + src5[283] + src5[284] + src5[285] + src5[286] + src5[287] + src5[288] + src5[289] + src5[290] + src5[291] + src5[292] + src5[293] + src5[294] + src5[295] + src5[296] + src5[297] + src5[298] + src5[299] + src5[300] + src5[301] + src5[302] + src5[303] + src5[304] + src5[305] + src5[306] + src5[307] + src5[308] + src5[309] + src5[310] + src5[311] + src5[312] + src5[313] + src5[314] + src5[315] + src5[316] + src5[317] + src5[318] + src5[319] + src5[320] + src5[321] + src5[322] + src5[323] + src5[324] + src5[325] + src5[326] + src5[327] + src5[328] + src5[329] + src5[330] + src5[331] + src5[332] + src5[333] + src5[334] + src5[335] + src5[336] + src5[337] + src5[338] + src5[339] + src5[340] + src5[341] + src5[342] + src5[343] + src5[344] + src5[345] + src5[346] + src5[347] + src5[348] + src5[349] + src5[350] + src5[351] + src5[352] + src5[353] + src5[354] + src5[355] + src5[356] + src5[357] + src5[358] + src5[359] + src5[360] + src5[361] + src5[362] + src5[363] + src5[364] + src5[365] + src5[366] + src5[367] + src5[368] + src5[369] + src5[370] + src5[371] + src5[372] + src5[373] + src5[374] + src5[375] + src5[376] + src5[377] + src5[378] + src5[379] + src5[380] + src5[381] + src5[382] + src5[383] + src5[384] + src5[385] + src5[386] + src5[387] + src5[388] + src5[389] + src5[390] + src5[391] + src5[392] + src5[393] + src5[394] + src5[395] + src5[396] + src5[397] + src5[398] + src5[399] + src5[400] + src5[401] + src5[402] + src5[403] + src5[404] + src5[405] + src5[406] + src5[407] + src5[408] + src5[409] + src5[410] + src5[411] + src5[412] + src5[413] + src5[414] + src5[415] + src5[416] + src5[417] + src5[418] + src5[419] + src5[420] + src5[421] + src5[422] + src5[423] + src5[424] + src5[425] + src5[426] + src5[427] + src5[428] + src5[429] + src5[430] + src5[431] + src5[432] + src5[433] + src5[434] + src5[435] + src5[436] + src5[437] + src5[438] + src5[439] + src5[440] + src5[441] + src5[442] + src5[443] + src5[444] + src5[445] + src5[446] + src5[447] + src5[448] + src5[449] + src5[450] + src5[451] + src5[452] + src5[453] + src5[454] + src5[455] + src5[456] + src5[457] + src5[458] + src5[459] + src5[460] + src5[461] + src5[462] + src5[463] + src5[464] + src5[465] + src5[466] + src5[467] + src5[468] + src5[469] + src5[470] + src5[471] + src5[472] + src5[473] + src5[474] + src5[475] + src5[476] + src5[477] + src5[478] + src5[479] + src5[480] + src5[481] + src5[482] + src5[483] + src5[484] + src5[485])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255] + src6[256] + src6[257] + src6[258] + src6[259] + src6[260] + src6[261] + src6[262] + src6[263] + src6[264] + src6[265] + src6[266] + src6[267] + src6[268] + src6[269] + src6[270] + src6[271] + src6[272] + src6[273] + src6[274] + src6[275] + src6[276] + src6[277] + src6[278] + src6[279] + src6[280] + src6[281] + src6[282] + src6[283] + src6[284] + src6[285] + src6[286] + src6[287] + src6[288] + src6[289] + src6[290] + src6[291] + src6[292] + src6[293] + src6[294] + src6[295] + src6[296] + src6[297] + src6[298] + src6[299] + src6[300] + src6[301] + src6[302] + src6[303] + src6[304] + src6[305] + src6[306] + src6[307] + src6[308] + src6[309] + src6[310] + src6[311] + src6[312] + src6[313] + src6[314] + src6[315] + src6[316] + src6[317] + src6[318] + src6[319] + src6[320] + src6[321] + src6[322] + src6[323] + src6[324] + src6[325] + src6[326] + src6[327] + src6[328] + src6[329] + src6[330] + src6[331] + src6[332] + src6[333] + src6[334] + src6[335] + src6[336] + src6[337] + src6[338] + src6[339] + src6[340] + src6[341] + src6[342] + src6[343] + src6[344] + src6[345] + src6[346] + src6[347] + src6[348] + src6[349] + src6[350] + src6[351] + src6[352] + src6[353] + src6[354] + src6[355] + src6[356] + src6[357] + src6[358] + src6[359] + src6[360] + src6[361] + src6[362] + src6[363] + src6[364] + src6[365] + src6[366] + src6[367] + src6[368] + src6[369] + src6[370] + src6[371] + src6[372] + src6[373] + src6[374] + src6[375] + src6[376] + src6[377] + src6[378] + src6[379] + src6[380] + src6[381] + src6[382] + src6[383] + src6[384] + src6[385] + src6[386] + src6[387] + src6[388] + src6[389] + src6[390] + src6[391] + src6[392] + src6[393] + src6[394] + src6[395] + src6[396] + src6[397] + src6[398] + src6[399] + src6[400] + src6[401] + src6[402] + src6[403] + src6[404] + src6[405] + src6[406] + src6[407] + src6[408] + src6[409] + src6[410] + src6[411] + src6[412] + src6[413] + src6[414] + src6[415] + src6[416] + src6[417] + src6[418] + src6[419] + src6[420] + src6[421] + src6[422] + src6[423] + src6[424] + src6[425] + src6[426] + src6[427] + src6[428] + src6[429] + src6[430] + src6[431] + src6[432] + src6[433] + src6[434] + src6[435] + src6[436] + src6[437] + src6[438] + src6[439] + src6[440] + src6[441] + src6[442] + src6[443] + src6[444] + src6[445] + src6[446] + src6[447] + src6[448] + src6[449] + src6[450] + src6[451] + src6[452] + src6[453] + src6[454] + src6[455] + src6[456] + src6[457] + src6[458] + src6[459] + src6[460] + src6[461] + src6[462] + src6[463] + src6[464] + src6[465] + src6[466] + src6[467] + src6[468] + src6[469] + src6[470] + src6[471] + src6[472] + src6[473] + src6[474] + src6[475] + src6[476] + src6[477] + src6[478] + src6[479] + src6[480] + src6[481] + src6[482] + src6[483] + src6[484] + src6[485])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255] + src7[256] + src7[257] + src7[258] + src7[259] + src7[260] + src7[261] + src7[262] + src7[263] + src7[264] + src7[265] + src7[266] + src7[267] + src7[268] + src7[269] + src7[270] + src7[271] + src7[272] + src7[273] + src7[274] + src7[275] + src7[276] + src7[277] + src7[278] + src7[279] + src7[280] + src7[281] + src7[282] + src7[283] + src7[284] + src7[285] + src7[286] + src7[287] + src7[288] + src7[289] + src7[290] + src7[291] + src7[292] + src7[293] + src7[294] + src7[295] + src7[296] + src7[297] + src7[298] + src7[299] + src7[300] + src7[301] + src7[302] + src7[303] + src7[304] + src7[305] + src7[306] + src7[307] + src7[308] + src7[309] + src7[310] + src7[311] + src7[312] + src7[313] + src7[314] + src7[315] + src7[316] + src7[317] + src7[318] + src7[319] + src7[320] + src7[321] + src7[322] + src7[323] + src7[324] + src7[325] + src7[326] + src7[327] + src7[328] + src7[329] + src7[330] + src7[331] + src7[332] + src7[333] + src7[334] + src7[335] + src7[336] + src7[337] + src7[338] + src7[339] + src7[340] + src7[341] + src7[342] + src7[343] + src7[344] + src7[345] + src7[346] + src7[347] + src7[348] + src7[349] + src7[350] + src7[351] + src7[352] + src7[353] + src7[354] + src7[355] + src7[356] + src7[357] + src7[358] + src7[359] + src7[360] + src7[361] + src7[362] + src7[363] + src7[364] + src7[365] + src7[366] + src7[367] + src7[368] + src7[369] + src7[370] + src7[371] + src7[372] + src7[373] + src7[374] + src7[375] + src7[376] + src7[377] + src7[378] + src7[379] + src7[380] + src7[381] + src7[382] + src7[383] + src7[384] + src7[385] + src7[386] + src7[387] + src7[388] + src7[389] + src7[390] + src7[391] + src7[392] + src7[393] + src7[394] + src7[395] + src7[396] + src7[397] + src7[398] + src7[399] + src7[400] + src7[401] + src7[402] + src7[403] + src7[404] + src7[405] + src7[406] + src7[407] + src7[408] + src7[409] + src7[410] + src7[411] + src7[412] + src7[413] + src7[414] + src7[415] + src7[416] + src7[417] + src7[418] + src7[419] + src7[420] + src7[421] + src7[422] + src7[423] + src7[424] + src7[425] + src7[426] + src7[427] + src7[428] + src7[429] + src7[430] + src7[431] + src7[432] + src7[433] + src7[434] + src7[435] + src7[436] + src7[437] + src7[438] + src7[439] + src7[440] + src7[441] + src7[442] + src7[443] + src7[444] + src7[445] + src7[446] + src7[447] + src7[448] + src7[449] + src7[450] + src7[451] + src7[452] + src7[453] + src7[454] + src7[455] + src7[456] + src7[457] + src7[458] + src7[459] + src7[460] + src7[461] + src7[462] + src7[463] + src7[464] + src7[465] + src7[466] + src7[467] + src7[468] + src7[469] + src7[470] + src7[471] + src7[472] + src7[473] + src7[474] + src7[475] + src7[476] + src7[477] + src7[478] + src7[479] + src7[480] + src7[481] + src7[482] + src7[483] + src7[484] + src7[485])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255] + src8[256] + src8[257] + src8[258] + src8[259] + src8[260] + src8[261] + src8[262] + src8[263] + src8[264] + src8[265] + src8[266] + src8[267] + src8[268] + src8[269] + src8[270] + src8[271] + src8[272] + src8[273] + src8[274] + src8[275] + src8[276] + src8[277] + src8[278] + src8[279] + src8[280] + src8[281] + src8[282] + src8[283] + src8[284] + src8[285] + src8[286] + src8[287] + src8[288] + src8[289] + src8[290] + src8[291] + src8[292] + src8[293] + src8[294] + src8[295] + src8[296] + src8[297] + src8[298] + src8[299] + src8[300] + src8[301] + src8[302] + src8[303] + src8[304] + src8[305] + src8[306] + src8[307] + src8[308] + src8[309] + src8[310] + src8[311] + src8[312] + src8[313] + src8[314] + src8[315] + src8[316] + src8[317] + src8[318] + src8[319] + src8[320] + src8[321] + src8[322] + src8[323] + src8[324] + src8[325] + src8[326] + src8[327] + src8[328] + src8[329] + src8[330] + src8[331] + src8[332] + src8[333] + src8[334] + src8[335] + src8[336] + src8[337] + src8[338] + src8[339] + src8[340] + src8[341] + src8[342] + src8[343] + src8[344] + src8[345] + src8[346] + src8[347] + src8[348] + src8[349] + src8[350] + src8[351] + src8[352] + src8[353] + src8[354] + src8[355] + src8[356] + src8[357] + src8[358] + src8[359] + src8[360] + src8[361] + src8[362] + src8[363] + src8[364] + src8[365] + src8[366] + src8[367] + src8[368] + src8[369] + src8[370] + src8[371] + src8[372] + src8[373] + src8[374] + src8[375] + src8[376] + src8[377] + src8[378] + src8[379] + src8[380] + src8[381] + src8[382] + src8[383] + src8[384] + src8[385] + src8[386] + src8[387] + src8[388] + src8[389] + src8[390] + src8[391] + src8[392] + src8[393] + src8[394] + src8[395] + src8[396] + src8[397] + src8[398] + src8[399] + src8[400] + src8[401] + src8[402] + src8[403] + src8[404] + src8[405] + src8[406] + src8[407] + src8[408] + src8[409] + src8[410] + src8[411] + src8[412] + src8[413] + src8[414] + src8[415] + src8[416] + src8[417] + src8[418] + src8[419] + src8[420] + src8[421] + src8[422] + src8[423] + src8[424] + src8[425] + src8[426] + src8[427] + src8[428] + src8[429] + src8[430] + src8[431] + src8[432] + src8[433] + src8[434] + src8[435] + src8[436] + src8[437] + src8[438] + src8[439] + src8[440] + src8[441] + src8[442] + src8[443] + src8[444] + src8[445] + src8[446] + src8[447] + src8[448] + src8[449] + src8[450] + src8[451] + src8[452] + src8[453] + src8[454] + src8[455] + src8[456] + src8[457] + src8[458] + src8[459] + src8[460] + src8[461] + src8[462] + src8[463] + src8[464] + src8[465] + src8[466] + src8[467] + src8[468] + src8[469] + src8[470] + src8[471] + src8[472] + src8[473] + src8[474] + src8[475] + src8[476] + src8[477] + src8[478] + src8[479] + src8[480] + src8[481] + src8[482] + src8[483] + src8[484] + src8[485])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255] + src9[256] + src9[257] + src9[258] + src9[259] + src9[260] + src9[261] + src9[262] + src9[263] + src9[264] + src9[265] + src9[266] + src9[267] + src9[268] + src9[269] + src9[270] + src9[271] + src9[272] + src9[273] + src9[274] + src9[275] + src9[276] + src9[277] + src9[278] + src9[279] + src9[280] + src9[281] + src9[282] + src9[283] + src9[284] + src9[285] + src9[286] + src9[287] + src9[288] + src9[289] + src9[290] + src9[291] + src9[292] + src9[293] + src9[294] + src9[295] + src9[296] + src9[297] + src9[298] + src9[299] + src9[300] + src9[301] + src9[302] + src9[303] + src9[304] + src9[305] + src9[306] + src9[307] + src9[308] + src9[309] + src9[310] + src9[311] + src9[312] + src9[313] + src9[314] + src9[315] + src9[316] + src9[317] + src9[318] + src9[319] + src9[320] + src9[321] + src9[322] + src9[323] + src9[324] + src9[325] + src9[326] + src9[327] + src9[328] + src9[329] + src9[330] + src9[331] + src9[332] + src9[333] + src9[334] + src9[335] + src9[336] + src9[337] + src9[338] + src9[339] + src9[340] + src9[341] + src9[342] + src9[343] + src9[344] + src9[345] + src9[346] + src9[347] + src9[348] + src9[349] + src9[350] + src9[351] + src9[352] + src9[353] + src9[354] + src9[355] + src9[356] + src9[357] + src9[358] + src9[359] + src9[360] + src9[361] + src9[362] + src9[363] + src9[364] + src9[365] + src9[366] + src9[367] + src9[368] + src9[369] + src9[370] + src9[371] + src9[372] + src9[373] + src9[374] + src9[375] + src9[376] + src9[377] + src9[378] + src9[379] + src9[380] + src9[381] + src9[382] + src9[383] + src9[384] + src9[385] + src9[386] + src9[387] + src9[388] + src9[389] + src9[390] + src9[391] + src9[392] + src9[393] + src9[394] + src9[395] + src9[396] + src9[397] + src9[398] + src9[399] + src9[400] + src9[401] + src9[402] + src9[403] + src9[404] + src9[405] + src9[406] + src9[407] + src9[408] + src9[409] + src9[410] + src9[411] + src9[412] + src9[413] + src9[414] + src9[415] + src9[416] + src9[417] + src9[418] + src9[419] + src9[420] + src9[421] + src9[422] + src9[423] + src9[424] + src9[425] + src9[426] + src9[427] + src9[428] + src9[429] + src9[430] + src9[431] + src9[432] + src9[433] + src9[434] + src9[435] + src9[436] + src9[437] + src9[438] + src9[439] + src9[440] + src9[441] + src9[442] + src9[443] + src9[444] + src9[445] + src9[446] + src9[447] + src9[448] + src9[449] + src9[450] + src9[451] + src9[452] + src9[453] + src9[454] + src9[455] + src9[456] + src9[457] + src9[458] + src9[459] + src9[460] + src9[461] + src9[462] + src9[463] + src9[464] + src9[465] + src9[466] + src9[467] + src9[468] + src9[469] + src9[470] + src9[471] + src9[472] + src9[473] + src9[474] + src9[475] + src9[476] + src9[477] + src9[478] + src9[479] + src9[480] + src9[481] + src9[482] + src9[483] + src9[484] + src9[485])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255] + src10[256] + src10[257] + src10[258] + src10[259] + src10[260] + src10[261] + src10[262] + src10[263] + src10[264] + src10[265] + src10[266] + src10[267] + src10[268] + src10[269] + src10[270] + src10[271] + src10[272] + src10[273] + src10[274] + src10[275] + src10[276] + src10[277] + src10[278] + src10[279] + src10[280] + src10[281] + src10[282] + src10[283] + src10[284] + src10[285] + src10[286] + src10[287] + src10[288] + src10[289] + src10[290] + src10[291] + src10[292] + src10[293] + src10[294] + src10[295] + src10[296] + src10[297] + src10[298] + src10[299] + src10[300] + src10[301] + src10[302] + src10[303] + src10[304] + src10[305] + src10[306] + src10[307] + src10[308] + src10[309] + src10[310] + src10[311] + src10[312] + src10[313] + src10[314] + src10[315] + src10[316] + src10[317] + src10[318] + src10[319] + src10[320] + src10[321] + src10[322] + src10[323] + src10[324] + src10[325] + src10[326] + src10[327] + src10[328] + src10[329] + src10[330] + src10[331] + src10[332] + src10[333] + src10[334] + src10[335] + src10[336] + src10[337] + src10[338] + src10[339] + src10[340] + src10[341] + src10[342] + src10[343] + src10[344] + src10[345] + src10[346] + src10[347] + src10[348] + src10[349] + src10[350] + src10[351] + src10[352] + src10[353] + src10[354] + src10[355] + src10[356] + src10[357] + src10[358] + src10[359] + src10[360] + src10[361] + src10[362] + src10[363] + src10[364] + src10[365] + src10[366] + src10[367] + src10[368] + src10[369] + src10[370] + src10[371] + src10[372] + src10[373] + src10[374] + src10[375] + src10[376] + src10[377] + src10[378] + src10[379] + src10[380] + src10[381] + src10[382] + src10[383] + src10[384] + src10[385] + src10[386] + src10[387] + src10[388] + src10[389] + src10[390] + src10[391] + src10[392] + src10[393] + src10[394] + src10[395] + src10[396] + src10[397] + src10[398] + src10[399] + src10[400] + src10[401] + src10[402] + src10[403] + src10[404] + src10[405] + src10[406] + src10[407] + src10[408] + src10[409] + src10[410] + src10[411] + src10[412] + src10[413] + src10[414] + src10[415] + src10[416] + src10[417] + src10[418] + src10[419] + src10[420] + src10[421] + src10[422] + src10[423] + src10[424] + src10[425] + src10[426] + src10[427] + src10[428] + src10[429] + src10[430] + src10[431] + src10[432] + src10[433] + src10[434] + src10[435] + src10[436] + src10[437] + src10[438] + src10[439] + src10[440] + src10[441] + src10[442] + src10[443] + src10[444] + src10[445] + src10[446] + src10[447] + src10[448] + src10[449] + src10[450] + src10[451] + src10[452] + src10[453] + src10[454] + src10[455] + src10[456] + src10[457] + src10[458] + src10[459] + src10[460] + src10[461] + src10[462] + src10[463] + src10[464] + src10[465] + src10[466] + src10[467] + src10[468] + src10[469] + src10[470] + src10[471] + src10[472] + src10[473] + src10[474] + src10[475] + src10[476] + src10[477] + src10[478] + src10[479] + src10[480] + src10[481] + src10[482] + src10[483] + src10[484] + src10[485])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255] + src11[256] + src11[257] + src11[258] + src11[259] + src11[260] + src11[261] + src11[262] + src11[263] + src11[264] + src11[265] + src11[266] + src11[267] + src11[268] + src11[269] + src11[270] + src11[271] + src11[272] + src11[273] + src11[274] + src11[275] + src11[276] + src11[277] + src11[278] + src11[279] + src11[280] + src11[281] + src11[282] + src11[283] + src11[284] + src11[285] + src11[286] + src11[287] + src11[288] + src11[289] + src11[290] + src11[291] + src11[292] + src11[293] + src11[294] + src11[295] + src11[296] + src11[297] + src11[298] + src11[299] + src11[300] + src11[301] + src11[302] + src11[303] + src11[304] + src11[305] + src11[306] + src11[307] + src11[308] + src11[309] + src11[310] + src11[311] + src11[312] + src11[313] + src11[314] + src11[315] + src11[316] + src11[317] + src11[318] + src11[319] + src11[320] + src11[321] + src11[322] + src11[323] + src11[324] + src11[325] + src11[326] + src11[327] + src11[328] + src11[329] + src11[330] + src11[331] + src11[332] + src11[333] + src11[334] + src11[335] + src11[336] + src11[337] + src11[338] + src11[339] + src11[340] + src11[341] + src11[342] + src11[343] + src11[344] + src11[345] + src11[346] + src11[347] + src11[348] + src11[349] + src11[350] + src11[351] + src11[352] + src11[353] + src11[354] + src11[355] + src11[356] + src11[357] + src11[358] + src11[359] + src11[360] + src11[361] + src11[362] + src11[363] + src11[364] + src11[365] + src11[366] + src11[367] + src11[368] + src11[369] + src11[370] + src11[371] + src11[372] + src11[373] + src11[374] + src11[375] + src11[376] + src11[377] + src11[378] + src11[379] + src11[380] + src11[381] + src11[382] + src11[383] + src11[384] + src11[385] + src11[386] + src11[387] + src11[388] + src11[389] + src11[390] + src11[391] + src11[392] + src11[393] + src11[394] + src11[395] + src11[396] + src11[397] + src11[398] + src11[399] + src11[400] + src11[401] + src11[402] + src11[403] + src11[404] + src11[405] + src11[406] + src11[407] + src11[408] + src11[409] + src11[410] + src11[411] + src11[412] + src11[413] + src11[414] + src11[415] + src11[416] + src11[417] + src11[418] + src11[419] + src11[420] + src11[421] + src11[422] + src11[423] + src11[424] + src11[425] + src11[426] + src11[427] + src11[428] + src11[429] + src11[430] + src11[431] + src11[432] + src11[433] + src11[434] + src11[435] + src11[436] + src11[437] + src11[438] + src11[439] + src11[440] + src11[441] + src11[442] + src11[443] + src11[444] + src11[445] + src11[446] + src11[447] + src11[448] + src11[449] + src11[450] + src11[451] + src11[452] + src11[453] + src11[454] + src11[455] + src11[456] + src11[457] + src11[458] + src11[459] + src11[460] + src11[461] + src11[462] + src11[463] + src11[464] + src11[465] + src11[466] + src11[467] + src11[468] + src11[469] + src11[470] + src11[471] + src11[472] + src11[473] + src11[474] + src11[475] + src11[476] + src11[477] + src11[478] + src11[479] + src11[480] + src11[481] + src11[482] + src11[483] + src11[484] + src11[485])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161] + src12[162] + src12[163] + src12[164] + src12[165] + src12[166] + src12[167] + src12[168] + src12[169] + src12[170] + src12[171] + src12[172] + src12[173] + src12[174] + src12[175] + src12[176] + src12[177] + src12[178] + src12[179] + src12[180] + src12[181] + src12[182] + src12[183] + src12[184] + src12[185] + src12[186] + src12[187] + src12[188] + src12[189] + src12[190] + src12[191] + src12[192] + src12[193] + src12[194] + src12[195] + src12[196] + src12[197] + src12[198] + src12[199] + src12[200] + src12[201] + src12[202] + src12[203] + src12[204] + src12[205] + src12[206] + src12[207] + src12[208] + src12[209] + src12[210] + src12[211] + src12[212] + src12[213] + src12[214] + src12[215] + src12[216] + src12[217] + src12[218] + src12[219] + src12[220] + src12[221] + src12[222] + src12[223] + src12[224] + src12[225] + src12[226] + src12[227] + src12[228] + src12[229] + src12[230] + src12[231] + src12[232] + src12[233] + src12[234] + src12[235] + src12[236] + src12[237] + src12[238] + src12[239] + src12[240] + src12[241] + src12[242] + src12[243] + src12[244] + src12[245] + src12[246] + src12[247] + src12[248] + src12[249] + src12[250] + src12[251] + src12[252] + src12[253] + src12[254] + src12[255] + src12[256] + src12[257] + src12[258] + src12[259] + src12[260] + src12[261] + src12[262] + src12[263] + src12[264] + src12[265] + src12[266] + src12[267] + src12[268] + src12[269] + src12[270] + src12[271] + src12[272] + src12[273] + src12[274] + src12[275] + src12[276] + src12[277] + src12[278] + src12[279] + src12[280] + src12[281] + src12[282] + src12[283] + src12[284] + src12[285] + src12[286] + src12[287] + src12[288] + src12[289] + src12[290] + src12[291] + src12[292] + src12[293] + src12[294] + src12[295] + src12[296] + src12[297] + src12[298] + src12[299] + src12[300] + src12[301] + src12[302] + src12[303] + src12[304] + src12[305] + src12[306] + src12[307] + src12[308] + src12[309] + src12[310] + src12[311] + src12[312] + src12[313] + src12[314] + src12[315] + src12[316] + src12[317] + src12[318] + src12[319] + src12[320] + src12[321] + src12[322] + src12[323] + src12[324] + src12[325] + src12[326] + src12[327] + src12[328] + src12[329] + src12[330] + src12[331] + src12[332] + src12[333] + src12[334] + src12[335] + src12[336] + src12[337] + src12[338] + src12[339] + src12[340] + src12[341] + src12[342] + src12[343] + src12[344] + src12[345] + src12[346] + src12[347] + src12[348] + src12[349] + src12[350] + src12[351] + src12[352] + src12[353] + src12[354] + src12[355] + src12[356] + src12[357] + src12[358] + src12[359] + src12[360] + src12[361] + src12[362] + src12[363] + src12[364] + src12[365] + src12[366] + src12[367] + src12[368] + src12[369] + src12[370] + src12[371] + src12[372] + src12[373] + src12[374] + src12[375] + src12[376] + src12[377] + src12[378] + src12[379] + src12[380] + src12[381] + src12[382] + src12[383] + src12[384] + src12[385] + src12[386] + src12[387] + src12[388] + src12[389] + src12[390] + src12[391] + src12[392] + src12[393] + src12[394] + src12[395] + src12[396] + src12[397] + src12[398] + src12[399] + src12[400] + src12[401] + src12[402] + src12[403] + src12[404] + src12[405] + src12[406] + src12[407] + src12[408] + src12[409] + src12[410] + src12[411] + src12[412] + src12[413] + src12[414] + src12[415] + src12[416] + src12[417] + src12[418] + src12[419] + src12[420] + src12[421] + src12[422] + src12[423] + src12[424] + src12[425] + src12[426] + src12[427] + src12[428] + src12[429] + src12[430] + src12[431] + src12[432] + src12[433] + src12[434] + src12[435] + src12[436] + src12[437] + src12[438] + src12[439] + src12[440] + src12[441] + src12[442] + src12[443] + src12[444] + src12[445] + src12[446] + src12[447] + src12[448] + src12[449] + src12[450] + src12[451] + src12[452] + src12[453] + src12[454] + src12[455] + src12[456] + src12[457] + src12[458] + src12[459] + src12[460] + src12[461] + src12[462] + src12[463] + src12[464] + src12[465] + src12[466] + src12[467] + src12[468] + src12[469] + src12[470] + src12[471] + src12[472] + src12[473] + src12[474] + src12[475] + src12[476] + src12[477] + src12[478] + src12[479] + src12[480] + src12[481] + src12[482] + src12[483] + src12[484] + src12[485])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161] + src13[162] + src13[163] + src13[164] + src13[165] + src13[166] + src13[167] + src13[168] + src13[169] + src13[170] + src13[171] + src13[172] + src13[173] + src13[174] + src13[175] + src13[176] + src13[177] + src13[178] + src13[179] + src13[180] + src13[181] + src13[182] + src13[183] + src13[184] + src13[185] + src13[186] + src13[187] + src13[188] + src13[189] + src13[190] + src13[191] + src13[192] + src13[193] + src13[194] + src13[195] + src13[196] + src13[197] + src13[198] + src13[199] + src13[200] + src13[201] + src13[202] + src13[203] + src13[204] + src13[205] + src13[206] + src13[207] + src13[208] + src13[209] + src13[210] + src13[211] + src13[212] + src13[213] + src13[214] + src13[215] + src13[216] + src13[217] + src13[218] + src13[219] + src13[220] + src13[221] + src13[222] + src13[223] + src13[224] + src13[225] + src13[226] + src13[227] + src13[228] + src13[229] + src13[230] + src13[231] + src13[232] + src13[233] + src13[234] + src13[235] + src13[236] + src13[237] + src13[238] + src13[239] + src13[240] + src13[241] + src13[242] + src13[243] + src13[244] + src13[245] + src13[246] + src13[247] + src13[248] + src13[249] + src13[250] + src13[251] + src13[252] + src13[253] + src13[254] + src13[255] + src13[256] + src13[257] + src13[258] + src13[259] + src13[260] + src13[261] + src13[262] + src13[263] + src13[264] + src13[265] + src13[266] + src13[267] + src13[268] + src13[269] + src13[270] + src13[271] + src13[272] + src13[273] + src13[274] + src13[275] + src13[276] + src13[277] + src13[278] + src13[279] + src13[280] + src13[281] + src13[282] + src13[283] + src13[284] + src13[285] + src13[286] + src13[287] + src13[288] + src13[289] + src13[290] + src13[291] + src13[292] + src13[293] + src13[294] + src13[295] + src13[296] + src13[297] + src13[298] + src13[299] + src13[300] + src13[301] + src13[302] + src13[303] + src13[304] + src13[305] + src13[306] + src13[307] + src13[308] + src13[309] + src13[310] + src13[311] + src13[312] + src13[313] + src13[314] + src13[315] + src13[316] + src13[317] + src13[318] + src13[319] + src13[320] + src13[321] + src13[322] + src13[323] + src13[324] + src13[325] + src13[326] + src13[327] + src13[328] + src13[329] + src13[330] + src13[331] + src13[332] + src13[333] + src13[334] + src13[335] + src13[336] + src13[337] + src13[338] + src13[339] + src13[340] + src13[341] + src13[342] + src13[343] + src13[344] + src13[345] + src13[346] + src13[347] + src13[348] + src13[349] + src13[350] + src13[351] + src13[352] + src13[353] + src13[354] + src13[355] + src13[356] + src13[357] + src13[358] + src13[359] + src13[360] + src13[361] + src13[362] + src13[363] + src13[364] + src13[365] + src13[366] + src13[367] + src13[368] + src13[369] + src13[370] + src13[371] + src13[372] + src13[373] + src13[374] + src13[375] + src13[376] + src13[377] + src13[378] + src13[379] + src13[380] + src13[381] + src13[382] + src13[383] + src13[384] + src13[385] + src13[386] + src13[387] + src13[388] + src13[389] + src13[390] + src13[391] + src13[392] + src13[393] + src13[394] + src13[395] + src13[396] + src13[397] + src13[398] + src13[399] + src13[400] + src13[401] + src13[402] + src13[403] + src13[404] + src13[405] + src13[406] + src13[407] + src13[408] + src13[409] + src13[410] + src13[411] + src13[412] + src13[413] + src13[414] + src13[415] + src13[416] + src13[417] + src13[418] + src13[419] + src13[420] + src13[421] + src13[422] + src13[423] + src13[424] + src13[425] + src13[426] + src13[427] + src13[428] + src13[429] + src13[430] + src13[431] + src13[432] + src13[433] + src13[434] + src13[435] + src13[436] + src13[437] + src13[438] + src13[439] + src13[440] + src13[441] + src13[442] + src13[443] + src13[444] + src13[445] + src13[446] + src13[447] + src13[448] + src13[449] + src13[450] + src13[451] + src13[452] + src13[453] + src13[454] + src13[455] + src13[456] + src13[457] + src13[458] + src13[459] + src13[460] + src13[461] + src13[462] + src13[463] + src13[464] + src13[465] + src13[466] + src13[467] + src13[468] + src13[469] + src13[470] + src13[471] + src13[472] + src13[473] + src13[474] + src13[475] + src13[476] + src13[477] + src13[478] + src13[479] + src13[480] + src13[481] + src13[482] + src13[483] + src13[484] + src13[485])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161] + src14[162] + src14[163] + src14[164] + src14[165] + src14[166] + src14[167] + src14[168] + src14[169] + src14[170] + src14[171] + src14[172] + src14[173] + src14[174] + src14[175] + src14[176] + src14[177] + src14[178] + src14[179] + src14[180] + src14[181] + src14[182] + src14[183] + src14[184] + src14[185] + src14[186] + src14[187] + src14[188] + src14[189] + src14[190] + src14[191] + src14[192] + src14[193] + src14[194] + src14[195] + src14[196] + src14[197] + src14[198] + src14[199] + src14[200] + src14[201] + src14[202] + src14[203] + src14[204] + src14[205] + src14[206] + src14[207] + src14[208] + src14[209] + src14[210] + src14[211] + src14[212] + src14[213] + src14[214] + src14[215] + src14[216] + src14[217] + src14[218] + src14[219] + src14[220] + src14[221] + src14[222] + src14[223] + src14[224] + src14[225] + src14[226] + src14[227] + src14[228] + src14[229] + src14[230] + src14[231] + src14[232] + src14[233] + src14[234] + src14[235] + src14[236] + src14[237] + src14[238] + src14[239] + src14[240] + src14[241] + src14[242] + src14[243] + src14[244] + src14[245] + src14[246] + src14[247] + src14[248] + src14[249] + src14[250] + src14[251] + src14[252] + src14[253] + src14[254] + src14[255] + src14[256] + src14[257] + src14[258] + src14[259] + src14[260] + src14[261] + src14[262] + src14[263] + src14[264] + src14[265] + src14[266] + src14[267] + src14[268] + src14[269] + src14[270] + src14[271] + src14[272] + src14[273] + src14[274] + src14[275] + src14[276] + src14[277] + src14[278] + src14[279] + src14[280] + src14[281] + src14[282] + src14[283] + src14[284] + src14[285] + src14[286] + src14[287] + src14[288] + src14[289] + src14[290] + src14[291] + src14[292] + src14[293] + src14[294] + src14[295] + src14[296] + src14[297] + src14[298] + src14[299] + src14[300] + src14[301] + src14[302] + src14[303] + src14[304] + src14[305] + src14[306] + src14[307] + src14[308] + src14[309] + src14[310] + src14[311] + src14[312] + src14[313] + src14[314] + src14[315] + src14[316] + src14[317] + src14[318] + src14[319] + src14[320] + src14[321] + src14[322] + src14[323] + src14[324] + src14[325] + src14[326] + src14[327] + src14[328] + src14[329] + src14[330] + src14[331] + src14[332] + src14[333] + src14[334] + src14[335] + src14[336] + src14[337] + src14[338] + src14[339] + src14[340] + src14[341] + src14[342] + src14[343] + src14[344] + src14[345] + src14[346] + src14[347] + src14[348] + src14[349] + src14[350] + src14[351] + src14[352] + src14[353] + src14[354] + src14[355] + src14[356] + src14[357] + src14[358] + src14[359] + src14[360] + src14[361] + src14[362] + src14[363] + src14[364] + src14[365] + src14[366] + src14[367] + src14[368] + src14[369] + src14[370] + src14[371] + src14[372] + src14[373] + src14[374] + src14[375] + src14[376] + src14[377] + src14[378] + src14[379] + src14[380] + src14[381] + src14[382] + src14[383] + src14[384] + src14[385] + src14[386] + src14[387] + src14[388] + src14[389] + src14[390] + src14[391] + src14[392] + src14[393] + src14[394] + src14[395] + src14[396] + src14[397] + src14[398] + src14[399] + src14[400] + src14[401] + src14[402] + src14[403] + src14[404] + src14[405] + src14[406] + src14[407] + src14[408] + src14[409] + src14[410] + src14[411] + src14[412] + src14[413] + src14[414] + src14[415] + src14[416] + src14[417] + src14[418] + src14[419] + src14[420] + src14[421] + src14[422] + src14[423] + src14[424] + src14[425] + src14[426] + src14[427] + src14[428] + src14[429] + src14[430] + src14[431] + src14[432] + src14[433] + src14[434] + src14[435] + src14[436] + src14[437] + src14[438] + src14[439] + src14[440] + src14[441] + src14[442] + src14[443] + src14[444] + src14[445] + src14[446] + src14[447] + src14[448] + src14[449] + src14[450] + src14[451] + src14[452] + src14[453] + src14[454] + src14[455] + src14[456] + src14[457] + src14[458] + src14[459] + src14[460] + src14[461] + src14[462] + src14[463] + src14[464] + src14[465] + src14[466] + src14[467] + src14[468] + src14[469] + src14[470] + src14[471] + src14[472] + src14[473] + src14[474] + src14[475] + src14[476] + src14[477] + src14[478] + src14[479] + src14[480] + src14[481] + src14[482] + src14[483] + src14[484] + src14[485])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161] + src15[162] + src15[163] + src15[164] + src15[165] + src15[166] + src15[167] + src15[168] + src15[169] + src15[170] + src15[171] + src15[172] + src15[173] + src15[174] + src15[175] + src15[176] + src15[177] + src15[178] + src15[179] + src15[180] + src15[181] + src15[182] + src15[183] + src15[184] + src15[185] + src15[186] + src15[187] + src15[188] + src15[189] + src15[190] + src15[191] + src15[192] + src15[193] + src15[194] + src15[195] + src15[196] + src15[197] + src15[198] + src15[199] + src15[200] + src15[201] + src15[202] + src15[203] + src15[204] + src15[205] + src15[206] + src15[207] + src15[208] + src15[209] + src15[210] + src15[211] + src15[212] + src15[213] + src15[214] + src15[215] + src15[216] + src15[217] + src15[218] + src15[219] + src15[220] + src15[221] + src15[222] + src15[223] + src15[224] + src15[225] + src15[226] + src15[227] + src15[228] + src15[229] + src15[230] + src15[231] + src15[232] + src15[233] + src15[234] + src15[235] + src15[236] + src15[237] + src15[238] + src15[239] + src15[240] + src15[241] + src15[242] + src15[243] + src15[244] + src15[245] + src15[246] + src15[247] + src15[248] + src15[249] + src15[250] + src15[251] + src15[252] + src15[253] + src15[254] + src15[255] + src15[256] + src15[257] + src15[258] + src15[259] + src15[260] + src15[261] + src15[262] + src15[263] + src15[264] + src15[265] + src15[266] + src15[267] + src15[268] + src15[269] + src15[270] + src15[271] + src15[272] + src15[273] + src15[274] + src15[275] + src15[276] + src15[277] + src15[278] + src15[279] + src15[280] + src15[281] + src15[282] + src15[283] + src15[284] + src15[285] + src15[286] + src15[287] + src15[288] + src15[289] + src15[290] + src15[291] + src15[292] + src15[293] + src15[294] + src15[295] + src15[296] + src15[297] + src15[298] + src15[299] + src15[300] + src15[301] + src15[302] + src15[303] + src15[304] + src15[305] + src15[306] + src15[307] + src15[308] + src15[309] + src15[310] + src15[311] + src15[312] + src15[313] + src15[314] + src15[315] + src15[316] + src15[317] + src15[318] + src15[319] + src15[320] + src15[321] + src15[322] + src15[323] + src15[324] + src15[325] + src15[326] + src15[327] + src15[328] + src15[329] + src15[330] + src15[331] + src15[332] + src15[333] + src15[334] + src15[335] + src15[336] + src15[337] + src15[338] + src15[339] + src15[340] + src15[341] + src15[342] + src15[343] + src15[344] + src15[345] + src15[346] + src15[347] + src15[348] + src15[349] + src15[350] + src15[351] + src15[352] + src15[353] + src15[354] + src15[355] + src15[356] + src15[357] + src15[358] + src15[359] + src15[360] + src15[361] + src15[362] + src15[363] + src15[364] + src15[365] + src15[366] + src15[367] + src15[368] + src15[369] + src15[370] + src15[371] + src15[372] + src15[373] + src15[374] + src15[375] + src15[376] + src15[377] + src15[378] + src15[379] + src15[380] + src15[381] + src15[382] + src15[383] + src15[384] + src15[385] + src15[386] + src15[387] + src15[388] + src15[389] + src15[390] + src15[391] + src15[392] + src15[393] + src15[394] + src15[395] + src15[396] + src15[397] + src15[398] + src15[399] + src15[400] + src15[401] + src15[402] + src15[403] + src15[404] + src15[405] + src15[406] + src15[407] + src15[408] + src15[409] + src15[410] + src15[411] + src15[412] + src15[413] + src15[414] + src15[415] + src15[416] + src15[417] + src15[418] + src15[419] + src15[420] + src15[421] + src15[422] + src15[423] + src15[424] + src15[425] + src15[426] + src15[427] + src15[428] + src15[429] + src15[430] + src15[431] + src15[432] + src15[433] + src15[434] + src15[435] + src15[436] + src15[437] + src15[438] + src15[439] + src15[440] + src15[441] + src15[442] + src15[443] + src15[444] + src15[445] + src15[446] + src15[447] + src15[448] + src15[449] + src15[450] + src15[451] + src15[452] + src15[453] + src15[454] + src15[455] + src15[456] + src15[457] + src15[458] + src15[459] + src15[460] + src15[461] + src15[462] + src15[463] + src15[464] + src15[465] + src15[466] + src15[467] + src15[468] + src15[469] + src15[470] + src15[471] + src15[472] + src15[473] + src15[474] + src15[475] + src15[476] + src15[477] + src15[478] + src15[479] + src15[480] + src15[481] + src15[482] + src15[483] + src15[484] + src15[485])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63] + src16[64] + src16[65] + src16[66] + src16[67] + src16[68] + src16[69] + src16[70] + src16[71] + src16[72] + src16[73] + src16[74] + src16[75] + src16[76] + src16[77] + src16[78] + src16[79] + src16[80] + src16[81] + src16[82] + src16[83] + src16[84] + src16[85] + src16[86] + src16[87] + src16[88] + src16[89] + src16[90] + src16[91] + src16[92] + src16[93] + src16[94] + src16[95] + src16[96] + src16[97] + src16[98] + src16[99] + src16[100] + src16[101] + src16[102] + src16[103] + src16[104] + src16[105] + src16[106] + src16[107] + src16[108] + src16[109] + src16[110] + src16[111] + src16[112] + src16[113] + src16[114] + src16[115] + src16[116] + src16[117] + src16[118] + src16[119] + src16[120] + src16[121] + src16[122] + src16[123] + src16[124] + src16[125] + src16[126] + src16[127] + src16[128] + src16[129] + src16[130] + src16[131] + src16[132] + src16[133] + src16[134] + src16[135] + src16[136] + src16[137] + src16[138] + src16[139] + src16[140] + src16[141] + src16[142] + src16[143] + src16[144] + src16[145] + src16[146] + src16[147] + src16[148] + src16[149] + src16[150] + src16[151] + src16[152] + src16[153] + src16[154] + src16[155] + src16[156] + src16[157] + src16[158] + src16[159] + src16[160] + src16[161] + src16[162] + src16[163] + src16[164] + src16[165] + src16[166] + src16[167] + src16[168] + src16[169] + src16[170] + src16[171] + src16[172] + src16[173] + src16[174] + src16[175] + src16[176] + src16[177] + src16[178] + src16[179] + src16[180] + src16[181] + src16[182] + src16[183] + src16[184] + src16[185] + src16[186] + src16[187] + src16[188] + src16[189] + src16[190] + src16[191] + src16[192] + src16[193] + src16[194] + src16[195] + src16[196] + src16[197] + src16[198] + src16[199] + src16[200] + src16[201] + src16[202] + src16[203] + src16[204] + src16[205] + src16[206] + src16[207] + src16[208] + src16[209] + src16[210] + src16[211] + src16[212] + src16[213] + src16[214] + src16[215] + src16[216] + src16[217] + src16[218] + src16[219] + src16[220] + src16[221] + src16[222] + src16[223] + src16[224] + src16[225] + src16[226] + src16[227] + src16[228] + src16[229] + src16[230] + src16[231] + src16[232] + src16[233] + src16[234] + src16[235] + src16[236] + src16[237] + src16[238] + src16[239] + src16[240] + src16[241] + src16[242] + src16[243] + src16[244] + src16[245] + src16[246] + src16[247] + src16[248] + src16[249] + src16[250] + src16[251] + src16[252] + src16[253] + src16[254] + src16[255] + src16[256] + src16[257] + src16[258] + src16[259] + src16[260] + src16[261] + src16[262] + src16[263] + src16[264] + src16[265] + src16[266] + src16[267] + src16[268] + src16[269] + src16[270] + src16[271] + src16[272] + src16[273] + src16[274] + src16[275] + src16[276] + src16[277] + src16[278] + src16[279] + src16[280] + src16[281] + src16[282] + src16[283] + src16[284] + src16[285] + src16[286] + src16[287] + src16[288] + src16[289] + src16[290] + src16[291] + src16[292] + src16[293] + src16[294] + src16[295] + src16[296] + src16[297] + src16[298] + src16[299] + src16[300] + src16[301] + src16[302] + src16[303] + src16[304] + src16[305] + src16[306] + src16[307] + src16[308] + src16[309] + src16[310] + src16[311] + src16[312] + src16[313] + src16[314] + src16[315] + src16[316] + src16[317] + src16[318] + src16[319] + src16[320] + src16[321] + src16[322] + src16[323] + src16[324] + src16[325] + src16[326] + src16[327] + src16[328] + src16[329] + src16[330] + src16[331] + src16[332] + src16[333] + src16[334] + src16[335] + src16[336] + src16[337] + src16[338] + src16[339] + src16[340] + src16[341] + src16[342] + src16[343] + src16[344] + src16[345] + src16[346] + src16[347] + src16[348] + src16[349] + src16[350] + src16[351] + src16[352] + src16[353] + src16[354] + src16[355] + src16[356] + src16[357] + src16[358] + src16[359] + src16[360] + src16[361] + src16[362] + src16[363] + src16[364] + src16[365] + src16[366] + src16[367] + src16[368] + src16[369] + src16[370] + src16[371] + src16[372] + src16[373] + src16[374] + src16[375] + src16[376] + src16[377] + src16[378] + src16[379] + src16[380] + src16[381] + src16[382] + src16[383] + src16[384] + src16[385] + src16[386] + src16[387] + src16[388] + src16[389] + src16[390] + src16[391] + src16[392] + src16[393] + src16[394] + src16[395] + src16[396] + src16[397] + src16[398] + src16[399] + src16[400] + src16[401] + src16[402] + src16[403] + src16[404] + src16[405] + src16[406] + src16[407] + src16[408] + src16[409] + src16[410] + src16[411] + src16[412] + src16[413] + src16[414] + src16[415] + src16[416] + src16[417] + src16[418] + src16[419] + src16[420] + src16[421] + src16[422] + src16[423] + src16[424] + src16[425] + src16[426] + src16[427] + src16[428] + src16[429] + src16[430] + src16[431] + src16[432] + src16[433] + src16[434] + src16[435] + src16[436] + src16[437] + src16[438] + src16[439] + src16[440] + src16[441] + src16[442] + src16[443] + src16[444] + src16[445] + src16[446] + src16[447] + src16[448] + src16[449] + src16[450] + src16[451] + src16[452] + src16[453] + src16[454] + src16[455] + src16[456] + src16[457] + src16[458] + src16[459] + src16[460] + src16[461] + src16[462] + src16[463] + src16[464] + src16[465] + src16[466] + src16[467] + src16[468] + src16[469] + src16[470] + src16[471] + src16[472] + src16[473] + src16[474] + src16[475] + src16[476] + src16[477] + src16[478] + src16[479] + src16[480] + src16[481] + src16[482] + src16[483] + src16[484] + src16[485])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63] + src17[64] + src17[65] + src17[66] + src17[67] + src17[68] + src17[69] + src17[70] + src17[71] + src17[72] + src17[73] + src17[74] + src17[75] + src17[76] + src17[77] + src17[78] + src17[79] + src17[80] + src17[81] + src17[82] + src17[83] + src17[84] + src17[85] + src17[86] + src17[87] + src17[88] + src17[89] + src17[90] + src17[91] + src17[92] + src17[93] + src17[94] + src17[95] + src17[96] + src17[97] + src17[98] + src17[99] + src17[100] + src17[101] + src17[102] + src17[103] + src17[104] + src17[105] + src17[106] + src17[107] + src17[108] + src17[109] + src17[110] + src17[111] + src17[112] + src17[113] + src17[114] + src17[115] + src17[116] + src17[117] + src17[118] + src17[119] + src17[120] + src17[121] + src17[122] + src17[123] + src17[124] + src17[125] + src17[126] + src17[127] + src17[128] + src17[129] + src17[130] + src17[131] + src17[132] + src17[133] + src17[134] + src17[135] + src17[136] + src17[137] + src17[138] + src17[139] + src17[140] + src17[141] + src17[142] + src17[143] + src17[144] + src17[145] + src17[146] + src17[147] + src17[148] + src17[149] + src17[150] + src17[151] + src17[152] + src17[153] + src17[154] + src17[155] + src17[156] + src17[157] + src17[158] + src17[159] + src17[160] + src17[161] + src17[162] + src17[163] + src17[164] + src17[165] + src17[166] + src17[167] + src17[168] + src17[169] + src17[170] + src17[171] + src17[172] + src17[173] + src17[174] + src17[175] + src17[176] + src17[177] + src17[178] + src17[179] + src17[180] + src17[181] + src17[182] + src17[183] + src17[184] + src17[185] + src17[186] + src17[187] + src17[188] + src17[189] + src17[190] + src17[191] + src17[192] + src17[193] + src17[194] + src17[195] + src17[196] + src17[197] + src17[198] + src17[199] + src17[200] + src17[201] + src17[202] + src17[203] + src17[204] + src17[205] + src17[206] + src17[207] + src17[208] + src17[209] + src17[210] + src17[211] + src17[212] + src17[213] + src17[214] + src17[215] + src17[216] + src17[217] + src17[218] + src17[219] + src17[220] + src17[221] + src17[222] + src17[223] + src17[224] + src17[225] + src17[226] + src17[227] + src17[228] + src17[229] + src17[230] + src17[231] + src17[232] + src17[233] + src17[234] + src17[235] + src17[236] + src17[237] + src17[238] + src17[239] + src17[240] + src17[241] + src17[242] + src17[243] + src17[244] + src17[245] + src17[246] + src17[247] + src17[248] + src17[249] + src17[250] + src17[251] + src17[252] + src17[253] + src17[254] + src17[255] + src17[256] + src17[257] + src17[258] + src17[259] + src17[260] + src17[261] + src17[262] + src17[263] + src17[264] + src17[265] + src17[266] + src17[267] + src17[268] + src17[269] + src17[270] + src17[271] + src17[272] + src17[273] + src17[274] + src17[275] + src17[276] + src17[277] + src17[278] + src17[279] + src17[280] + src17[281] + src17[282] + src17[283] + src17[284] + src17[285] + src17[286] + src17[287] + src17[288] + src17[289] + src17[290] + src17[291] + src17[292] + src17[293] + src17[294] + src17[295] + src17[296] + src17[297] + src17[298] + src17[299] + src17[300] + src17[301] + src17[302] + src17[303] + src17[304] + src17[305] + src17[306] + src17[307] + src17[308] + src17[309] + src17[310] + src17[311] + src17[312] + src17[313] + src17[314] + src17[315] + src17[316] + src17[317] + src17[318] + src17[319] + src17[320] + src17[321] + src17[322] + src17[323] + src17[324] + src17[325] + src17[326] + src17[327] + src17[328] + src17[329] + src17[330] + src17[331] + src17[332] + src17[333] + src17[334] + src17[335] + src17[336] + src17[337] + src17[338] + src17[339] + src17[340] + src17[341] + src17[342] + src17[343] + src17[344] + src17[345] + src17[346] + src17[347] + src17[348] + src17[349] + src17[350] + src17[351] + src17[352] + src17[353] + src17[354] + src17[355] + src17[356] + src17[357] + src17[358] + src17[359] + src17[360] + src17[361] + src17[362] + src17[363] + src17[364] + src17[365] + src17[366] + src17[367] + src17[368] + src17[369] + src17[370] + src17[371] + src17[372] + src17[373] + src17[374] + src17[375] + src17[376] + src17[377] + src17[378] + src17[379] + src17[380] + src17[381] + src17[382] + src17[383] + src17[384] + src17[385] + src17[386] + src17[387] + src17[388] + src17[389] + src17[390] + src17[391] + src17[392] + src17[393] + src17[394] + src17[395] + src17[396] + src17[397] + src17[398] + src17[399] + src17[400] + src17[401] + src17[402] + src17[403] + src17[404] + src17[405] + src17[406] + src17[407] + src17[408] + src17[409] + src17[410] + src17[411] + src17[412] + src17[413] + src17[414] + src17[415] + src17[416] + src17[417] + src17[418] + src17[419] + src17[420] + src17[421] + src17[422] + src17[423] + src17[424] + src17[425] + src17[426] + src17[427] + src17[428] + src17[429] + src17[430] + src17[431] + src17[432] + src17[433] + src17[434] + src17[435] + src17[436] + src17[437] + src17[438] + src17[439] + src17[440] + src17[441] + src17[442] + src17[443] + src17[444] + src17[445] + src17[446] + src17[447] + src17[448] + src17[449] + src17[450] + src17[451] + src17[452] + src17[453] + src17[454] + src17[455] + src17[456] + src17[457] + src17[458] + src17[459] + src17[460] + src17[461] + src17[462] + src17[463] + src17[464] + src17[465] + src17[466] + src17[467] + src17[468] + src17[469] + src17[470] + src17[471] + src17[472] + src17[473] + src17[474] + src17[475] + src17[476] + src17[477] + src17[478] + src17[479] + src17[480] + src17[481] + src17[482] + src17[483] + src17[484] + src17[485])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63] + src18[64] + src18[65] + src18[66] + src18[67] + src18[68] + src18[69] + src18[70] + src18[71] + src18[72] + src18[73] + src18[74] + src18[75] + src18[76] + src18[77] + src18[78] + src18[79] + src18[80] + src18[81] + src18[82] + src18[83] + src18[84] + src18[85] + src18[86] + src18[87] + src18[88] + src18[89] + src18[90] + src18[91] + src18[92] + src18[93] + src18[94] + src18[95] + src18[96] + src18[97] + src18[98] + src18[99] + src18[100] + src18[101] + src18[102] + src18[103] + src18[104] + src18[105] + src18[106] + src18[107] + src18[108] + src18[109] + src18[110] + src18[111] + src18[112] + src18[113] + src18[114] + src18[115] + src18[116] + src18[117] + src18[118] + src18[119] + src18[120] + src18[121] + src18[122] + src18[123] + src18[124] + src18[125] + src18[126] + src18[127] + src18[128] + src18[129] + src18[130] + src18[131] + src18[132] + src18[133] + src18[134] + src18[135] + src18[136] + src18[137] + src18[138] + src18[139] + src18[140] + src18[141] + src18[142] + src18[143] + src18[144] + src18[145] + src18[146] + src18[147] + src18[148] + src18[149] + src18[150] + src18[151] + src18[152] + src18[153] + src18[154] + src18[155] + src18[156] + src18[157] + src18[158] + src18[159] + src18[160] + src18[161] + src18[162] + src18[163] + src18[164] + src18[165] + src18[166] + src18[167] + src18[168] + src18[169] + src18[170] + src18[171] + src18[172] + src18[173] + src18[174] + src18[175] + src18[176] + src18[177] + src18[178] + src18[179] + src18[180] + src18[181] + src18[182] + src18[183] + src18[184] + src18[185] + src18[186] + src18[187] + src18[188] + src18[189] + src18[190] + src18[191] + src18[192] + src18[193] + src18[194] + src18[195] + src18[196] + src18[197] + src18[198] + src18[199] + src18[200] + src18[201] + src18[202] + src18[203] + src18[204] + src18[205] + src18[206] + src18[207] + src18[208] + src18[209] + src18[210] + src18[211] + src18[212] + src18[213] + src18[214] + src18[215] + src18[216] + src18[217] + src18[218] + src18[219] + src18[220] + src18[221] + src18[222] + src18[223] + src18[224] + src18[225] + src18[226] + src18[227] + src18[228] + src18[229] + src18[230] + src18[231] + src18[232] + src18[233] + src18[234] + src18[235] + src18[236] + src18[237] + src18[238] + src18[239] + src18[240] + src18[241] + src18[242] + src18[243] + src18[244] + src18[245] + src18[246] + src18[247] + src18[248] + src18[249] + src18[250] + src18[251] + src18[252] + src18[253] + src18[254] + src18[255] + src18[256] + src18[257] + src18[258] + src18[259] + src18[260] + src18[261] + src18[262] + src18[263] + src18[264] + src18[265] + src18[266] + src18[267] + src18[268] + src18[269] + src18[270] + src18[271] + src18[272] + src18[273] + src18[274] + src18[275] + src18[276] + src18[277] + src18[278] + src18[279] + src18[280] + src18[281] + src18[282] + src18[283] + src18[284] + src18[285] + src18[286] + src18[287] + src18[288] + src18[289] + src18[290] + src18[291] + src18[292] + src18[293] + src18[294] + src18[295] + src18[296] + src18[297] + src18[298] + src18[299] + src18[300] + src18[301] + src18[302] + src18[303] + src18[304] + src18[305] + src18[306] + src18[307] + src18[308] + src18[309] + src18[310] + src18[311] + src18[312] + src18[313] + src18[314] + src18[315] + src18[316] + src18[317] + src18[318] + src18[319] + src18[320] + src18[321] + src18[322] + src18[323] + src18[324] + src18[325] + src18[326] + src18[327] + src18[328] + src18[329] + src18[330] + src18[331] + src18[332] + src18[333] + src18[334] + src18[335] + src18[336] + src18[337] + src18[338] + src18[339] + src18[340] + src18[341] + src18[342] + src18[343] + src18[344] + src18[345] + src18[346] + src18[347] + src18[348] + src18[349] + src18[350] + src18[351] + src18[352] + src18[353] + src18[354] + src18[355] + src18[356] + src18[357] + src18[358] + src18[359] + src18[360] + src18[361] + src18[362] + src18[363] + src18[364] + src18[365] + src18[366] + src18[367] + src18[368] + src18[369] + src18[370] + src18[371] + src18[372] + src18[373] + src18[374] + src18[375] + src18[376] + src18[377] + src18[378] + src18[379] + src18[380] + src18[381] + src18[382] + src18[383] + src18[384] + src18[385] + src18[386] + src18[387] + src18[388] + src18[389] + src18[390] + src18[391] + src18[392] + src18[393] + src18[394] + src18[395] + src18[396] + src18[397] + src18[398] + src18[399] + src18[400] + src18[401] + src18[402] + src18[403] + src18[404] + src18[405] + src18[406] + src18[407] + src18[408] + src18[409] + src18[410] + src18[411] + src18[412] + src18[413] + src18[414] + src18[415] + src18[416] + src18[417] + src18[418] + src18[419] + src18[420] + src18[421] + src18[422] + src18[423] + src18[424] + src18[425] + src18[426] + src18[427] + src18[428] + src18[429] + src18[430] + src18[431] + src18[432] + src18[433] + src18[434] + src18[435] + src18[436] + src18[437] + src18[438] + src18[439] + src18[440] + src18[441] + src18[442] + src18[443] + src18[444] + src18[445] + src18[446] + src18[447] + src18[448] + src18[449] + src18[450] + src18[451] + src18[452] + src18[453] + src18[454] + src18[455] + src18[456] + src18[457] + src18[458] + src18[459] + src18[460] + src18[461] + src18[462] + src18[463] + src18[464] + src18[465] + src18[466] + src18[467] + src18[468] + src18[469] + src18[470] + src18[471] + src18[472] + src18[473] + src18[474] + src18[475] + src18[476] + src18[477] + src18[478] + src18[479] + src18[480] + src18[481] + src18[482] + src18[483] + src18[484] + src18[485])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63] + src19[64] + src19[65] + src19[66] + src19[67] + src19[68] + src19[69] + src19[70] + src19[71] + src19[72] + src19[73] + src19[74] + src19[75] + src19[76] + src19[77] + src19[78] + src19[79] + src19[80] + src19[81] + src19[82] + src19[83] + src19[84] + src19[85] + src19[86] + src19[87] + src19[88] + src19[89] + src19[90] + src19[91] + src19[92] + src19[93] + src19[94] + src19[95] + src19[96] + src19[97] + src19[98] + src19[99] + src19[100] + src19[101] + src19[102] + src19[103] + src19[104] + src19[105] + src19[106] + src19[107] + src19[108] + src19[109] + src19[110] + src19[111] + src19[112] + src19[113] + src19[114] + src19[115] + src19[116] + src19[117] + src19[118] + src19[119] + src19[120] + src19[121] + src19[122] + src19[123] + src19[124] + src19[125] + src19[126] + src19[127] + src19[128] + src19[129] + src19[130] + src19[131] + src19[132] + src19[133] + src19[134] + src19[135] + src19[136] + src19[137] + src19[138] + src19[139] + src19[140] + src19[141] + src19[142] + src19[143] + src19[144] + src19[145] + src19[146] + src19[147] + src19[148] + src19[149] + src19[150] + src19[151] + src19[152] + src19[153] + src19[154] + src19[155] + src19[156] + src19[157] + src19[158] + src19[159] + src19[160] + src19[161] + src19[162] + src19[163] + src19[164] + src19[165] + src19[166] + src19[167] + src19[168] + src19[169] + src19[170] + src19[171] + src19[172] + src19[173] + src19[174] + src19[175] + src19[176] + src19[177] + src19[178] + src19[179] + src19[180] + src19[181] + src19[182] + src19[183] + src19[184] + src19[185] + src19[186] + src19[187] + src19[188] + src19[189] + src19[190] + src19[191] + src19[192] + src19[193] + src19[194] + src19[195] + src19[196] + src19[197] + src19[198] + src19[199] + src19[200] + src19[201] + src19[202] + src19[203] + src19[204] + src19[205] + src19[206] + src19[207] + src19[208] + src19[209] + src19[210] + src19[211] + src19[212] + src19[213] + src19[214] + src19[215] + src19[216] + src19[217] + src19[218] + src19[219] + src19[220] + src19[221] + src19[222] + src19[223] + src19[224] + src19[225] + src19[226] + src19[227] + src19[228] + src19[229] + src19[230] + src19[231] + src19[232] + src19[233] + src19[234] + src19[235] + src19[236] + src19[237] + src19[238] + src19[239] + src19[240] + src19[241] + src19[242] + src19[243] + src19[244] + src19[245] + src19[246] + src19[247] + src19[248] + src19[249] + src19[250] + src19[251] + src19[252] + src19[253] + src19[254] + src19[255] + src19[256] + src19[257] + src19[258] + src19[259] + src19[260] + src19[261] + src19[262] + src19[263] + src19[264] + src19[265] + src19[266] + src19[267] + src19[268] + src19[269] + src19[270] + src19[271] + src19[272] + src19[273] + src19[274] + src19[275] + src19[276] + src19[277] + src19[278] + src19[279] + src19[280] + src19[281] + src19[282] + src19[283] + src19[284] + src19[285] + src19[286] + src19[287] + src19[288] + src19[289] + src19[290] + src19[291] + src19[292] + src19[293] + src19[294] + src19[295] + src19[296] + src19[297] + src19[298] + src19[299] + src19[300] + src19[301] + src19[302] + src19[303] + src19[304] + src19[305] + src19[306] + src19[307] + src19[308] + src19[309] + src19[310] + src19[311] + src19[312] + src19[313] + src19[314] + src19[315] + src19[316] + src19[317] + src19[318] + src19[319] + src19[320] + src19[321] + src19[322] + src19[323] + src19[324] + src19[325] + src19[326] + src19[327] + src19[328] + src19[329] + src19[330] + src19[331] + src19[332] + src19[333] + src19[334] + src19[335] + src19[336] + src19[337] + src19[338] + src19[339] + src19[340] + src19[341] + src19[342] + src19[343] + src19[344] + src19[345] + src19[346] + src19[347] + src19[348] + src19[349] + src19[350] + src19[351] + src19[352] + src19[353] + src19[354] + src19[355] + src19[356] + src19[357] + src19[358] + src19[359] + src19[360] + src19[361] + src19[362] + src19[363] + src19[364] + src19[365] + src19[366] + src19[367] + src19[368] + src19[369] + src19[370] + src19[371] + src19[372] + src19[373] + src19[374] + src19[375] + src19[376] + src19[377] + src19[378] + src19[379] + src19[380] + src19[381] + src19[382] + src19[383] + src19[384] + src19[385] + src19[386] + src19[387] + src19[388] + src19[389] + src19[390] + src19[391] + src19[392] + src19[393] + src19[394] + src19[395] + src19[396] + src19[397] + src19[398] + src19[399] + src19[400] + src19[401] + src19[402] + src19[403] + src19[404] + src19[405] + src19[406] + src19[407] + src19[408] + src19[409] + src19[410] + src19[411] + src19[412] + src19[413] + src19[414] + src19[415] + src19[416] + src19[417] + src19[418] + src19[419] + src19[420] + src19[421] + src19[422] + src19[423] + src19[424] + src19[425] + src19[426] + src19[427] + src19[428] + src19[429] + src19[430] + src19[431] + src19[432] + src19[433] + src19[434] + src19[435] + src19[436] + src19[437] + src19[438] + src19[439] + src19[440] + src19[441] + src19[442] + src19[443] + src19[444] + src19[445] + src19[446] + src19[447] + src19[448] + src19[449] + src19[450] + src19[451] + src19[452] + src19[453] + src19[454] + src19[455] + src19[456] + src19[457] + src19[458] + src19[459] + src19[460] + src19[461] + src19[462] + src19[463] + src19[464] + src19[465] + src19[466] + src19[467] + src19[468] + src19[469] + src19[470] + src19[471] + src19[472] + src19[473] + src19[474] + src19[475] + src19[476] + src19[477] + src19[478] + src19[479] + src19[480] + src19[481] + src19[482] + src19[483] + src19[484] + src19[485])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63] + src20[64] + src20[65] + src20[66] + src20[67] + src20[68] + src20[69] + src20[70] + src20[71] + src20[72] + src20[73] + src20[74] + src20[75] + src20[76] + src20[77] + src20[78] + src20[79] + src20[80] + src20[81] + src20[82] + src20[83] + src20[84] + src20[85] + src20[86] + src20[87] + src20[88] + src20[89] + src20[90] + src20[91] + src20[92] + src20[93] + src20[94] + src20[95] + src20[96] + src20[97] + src20[98] + src20[99] + src20[100] + src20[101] + src20[102] + src20[103] + src20[104] + src20[105] + src20[106] + src20[107] + src20[108] + src20[109] + src20[110] + src20[111] + src20[112] + src20[113] + src20[114] + src20[115] + src20[116] + src20[117] + src20[118] + src20[119] + src20[120] + src20[121] + src20[122] + src20[123] + src20[124] + src20[125] + src20[126] + src20[127] + src20[128] + src20[129] + src20[130] + src20[131] + src20[132] + src20[133] + src20[134] + src20[135] + src20[136] + src20[137] + src20[138] + src20[139] + src20[140] + src20[141] + src20[142] + src20[143] + src20[144] + src20[145] + src20[146] + src20[147] + src20[148] + src20[149] + src20[150] + src20[151] + src20[152] + src20[153] + src20[154] + src20[155] + src20[156] + src20[157] + src20[158] + src20[159] + src20[160] + src20[161] + src20[162] + src20[163] + src20[164] + src20[165] + src20[166] + src20[167] + src20[168] + src20[169] + src20[170] + src20[171] + src20[172] + src20[173] + src20[174] + src20[175] + src20[176] + src20[177] + src20[178] + src20[179] + src20[180] + src20[181] + src20[182] + src20[183] + src20[184] + src20[185] + src20[186] + src20[187] + src20[188] + src20[189] + src20[190] + src20[191] + src20[192] + src20[193] + src20[194] + src20[195] + src20[196] + src20[197] + src20[198] + src20[199] + src20[200] + src20[201] + src20[202] + src20[203] + src20[204] + src20[205] + src20[206] + src20[207] + src20[208] + src20[209] + src20[210] + src20[211] + src20[212] + src20[213] + src20[214] + src20[215] + src20[216] + src20[217] + src20[218] + src20[219] + src20[220] + src20[221] + src20[222] + src20[223] + src20[224] + src20[225] + src20[226] + src20[227] + src20[228] + src20[229] + src20[230] + src20[231] + src20[232] + src20[233] + src20[234] + src20[235] + src20[236] + src20[237] + src20[238] + src20[239] + src20[240] + src20[241] + src20[242] + src20[243] + src20[244] + src20[245] + src20[246] + src20[247] + src20[248] + src20[249] + src20[250] + src20[251] + src20[252] + src20[253] + src20[254] + src20[255] + src20[256] + src20[257] + src20[258] + src20[259] + src20[260] + src20[261] + src20[262] + src20[263] + src20[264] + src20[265] + src20[266] + src20[267] + src20[268] + src20[269] + src20[270] + src20[271] + src20[272] + src20[273] + src20[274] + src20[275] + src20[276] + src20[277] + src20[278] + src20[279] + src20[280] + src20[281] + src20[282] + src20[283] + src20[284] + src20[285] + src20[286] + src20[287] + src20[288] + src20[289] + src20[290] + src20[291] + src20[292] + src20[293] + src20[294] + src20[295] + src20[296] + src20[297] + src20[298] + src20[299] + src20[300] + src20[301] + src20[302] + src20[303] + src20[304] + src20[305] + src20[306] + src20[307] + src20[308] + src20[309] + src20[310] + src20[311] + src20[312] + src20[313] + src20[314] + src20[315] + src20[316] + src20[317] + src20[318] + src20[319] + src20[320] + src20[321] + src20[322] + src20[323] + src20[324] + src20[325] + src20[326] + src20[327] + src20[328] + src20[329] + src20[330] + src20[331] + src20[332] + src20[333] + src20[334] + src20[335] + src20[336] + src20[337] + src20[338] + src20[339] + src20[340] + src20[341] + src20[342] + src20[343] + src20[344] + src20[345] + src20[346] + src20[347] + src20[348] + src20[349] + src20[350] + src20[351] + src20[352] + src20[353] + src20[354] + src20[355] + src20[356] + src20[357] + src20[358] + src20[359] + src20[360] + src20[361] + src20[362] + src20[363] + src20[364] + src20[365] + src20[366] + src20[367] + src20[368] + src20[369] + src20[370] + src20[371] + src20[372] + src20[373] + src20[374] + src20[375] + src20[376] + src20[377] + src20[378] + src20[379] + src20[380] + src20[381] + src20[382] + src20[383] + src20[384] + src20[385] + src20[386] + src20[387] + src20[388] + src20[389] + src20[390] + src20[391] + src20[392] + src20[393] + src20[394] + src20[395] + src20[396] + src20[397] + src20[398] + src20[399] + src20[400] + src20[401] + src20[402] + src20[403] + src20[404] + src20[405] + src20[406] + src20[407] + src20[408] + src20[409] + src20[410] + src20[411] + src20[412] + src20[413] + src20[414] + src20[415] + src20[416] + src20[417] + src20[418] + src20[419] + src20[420] + src20[421] + src20[422] + src20[423] + src20[424] + src20[425] + src20[426] + src20[427] + src20[428] + src20[429] + src20[430] + src20[431] + src20[432] + src20[433] + src20[434] + src20[435] + src20[436] + src20[437] + src20[438] + src20[439] + src20[440] + src20[441] + src20[442] + src20[443] + src20[444] + src20[445] + src20[446] + src20[447] + src20[448] + src20[449] + src20[450] + src20[451] + src20[452] + src20[453] + src20[454] + src20[455] + src20[456] + src20[457] + src20[458] + src20[459] + src20[460] + src20[461] + src20[462] + src20[463] + src20[464] + src20[465] + src20[466] + src20[467] + src20[468] + src20[469] + src20[470] + src20[471] + src20[472] + src20[473] + src20[474] + src20[475] + src20[476] + src20[477] + src20[478] + src20[479] + src20[480] + src20[481] + src20[482] + src20[483] + src20[484] + src20[485])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63] + src21[64] + src21[65] + src21[66] + src21[67] + src21[68] + src21[69] + src21[70] + src21[71] + src21[72] + src21[73] + src21[74] + src21[75] + src21[76] + src21[77] + src21[78] + src21[79] + src21[80] + src21[81] + src21[82] + src21[83] + src21[84] + src21[85] + src21[86] + src21[87] + src21[88] + src21[89] + src21[90] + src21[91] + src21[92] + src21[93] + src21[94] + src21[95] + src21[96] + src21[97] + src21[98] + src21[99] + src21[100] + src21[101] + src21[102] + src21[103] + src21[104] + src21[105] + src21[106] + src21[107] + src21[108] + src21[109] + src21[110] + src21[111] + src21[112] + src21[113] + src21[114] + src21[115] + src21[116] + src21[117] + src21[118] + src21[119] + src21[120] + src21[121] + src21[122] + src21[123] + src21[124] + src21[125] + src21[126] + src21[127] + src21[128] + src21[129] + src21[130] + src21[131] + src21[132] + src21[133] + src21[134] + src21[135] + src21[136] + src21[137] + src21[138] + src21[139] + src21[140] + src21[141] + src21[142] + src21[143] + src21[144] + src21[145] + src21[146] + src21[147] + src21[148] + src21[149] + src21[150] + src21[151] + src21[152] + src21[153] + src21[154] + src21[155] + src21[156] + src21[157] + src21[158] + src21[159] + src21[160] + src21[161] + src21[162] + src21[163] + src21[164] + src21[165] + src21[166] + src21[167] + src21[168] + src21[169] + src21[170] + src21[171] + src21[172] + src21[173] + src21[174] + src21[175] + src21[176] + src21[177] + src21[178] + src21[179] + src21[180] + src21[181] + src21[182] + src21[183] + src21[184] + src21[185] + src21[186] + src21[187] + src21[188] + src21[189] + src21[190] + src21[191] + src21[192] + src21[193] + src21[194] + src21[195] + src21[196] + src21[197] + src21[198] + src21[199] + src21[200] + src21[201] + src21[202] + src21[203] + src21[204] + src21[205] + src21[206] + src21[207] + src21[208] + src21[209] + src21[210] + src21[211] + src21[212] + src21[213] + src21[214] + src21[215] + src21[216] + src21[217] + src21[218] + src21[219] + src21[220] + src21[221] + src21[222] + src21[223] + src21[224] + src21[225] + src21[226] + src21[227] + src21[228] + src21[229] + src21[230] + src21[231] + src21[232] + src21[233] + src21[234] + src21[235] + src21[236] + src21[237] + src21[238] + src21[239] + src21[240] + src21[241] + src21[242] + src21[243] + src21[244] + src21[245] + src21[246] + src21[247] + src21[248] + src21[249] + src21[250] + src21[251] + src21[252] + src21[253] + src21[254] + src21[255] + src21[256] + src21[257] + src21[258] + src21[259] + src21[260] + src21[261] + src21[262] + src21[263] + src21[264] + src21[265] + src21[266] + src21[267] + src21[268] + src21[269] + src21[270] + src21[271] + src21[272] + src21[273] + src21[274] + src21[275] + src21[276] + src21[277] + src21[278] + src21[279] + src21[280] + src21[281] + src21[282] + src21[283] + src21[284] + src21[285] + src21[286] + src21[287] + src21[288] + src21[289] + src21[290] + src21[291] + src21[292] + src21[293] + src21[294] + src21[295] + src21[296] + src21[297] + src21[298] + src21[299] + src21[300] + src21[301] + src21[302] + src21[303] + src21[304] + src21[305] + src21[306] + src21[307] + src21[308] + src21[309] + src21[310] + src21[311] + src21[312] + src21[313] + src21[314] + src21[315] + src21[316] + src21[317] + src21[318] + src21[319] + src21[320] + src21[321] + src21[322] + src21[323] + src21[324] + src21[325] + src21[326] + src21[327] + src21[328] + src21[329] + src21[330] + src21[331] + src21[332] + src21[333] + src21[334] + src21[335] + src21[336] + src21[337] + src21[338] + src21[339] + src21[340] + src21[341] + src21[342] + src21[343] + src21[344] + src21[345] + src21[346] + src21[347] + src21[348] + src21[349] + src21[350] + src21[351] + src21[352] + src21[353] + src21[354] + src21[355] + src21[356] + src21[357] + src21[358] + src21[359] + src21[360] + src21[361] + src21[362] + src21[363] + src21[364] + src21[365] + src21[366] + src21[367] + src21[368] + src21[369] + src21[370] + src21[371] + src21[372] + src21[373] + src21[374] + src21[375] + src21[376] + src21[377] + src21[378] + src21[379] + src21[380] + src21[381] + src21[382] + src21[383] + src21[384] + src21[385] + src21[386] + src21[387] + src21[388] + src21[389] + src21[390] + src21[391] + src21[392] + src21[393] + src21[394] + src21[395] + src21[396] + src21[397] + src21[398] + src21[399] + src21[400] + src21[401] + src21[402] + src21[403] + src21[404] + src21[405] + src21[406] + src21[407] + src21[408] + src21[409] + src21[410] + src21[411] + src21[412] + src21[413] + src21[414] + src21[415] + src21[416] + src21[417] + src21[418] + src21[419] + src21[420] + src21[421] + src21[422] + src21[423] + src21[424] + src21[425] + src21[426] + src21[427] + src21[428] + src21[429] + src21[430] + src21[431] + src21[432] + src21[433] + src21[434] + src21[435] + src21[436] + src21[437] + src21[438] + src21[439] + src21[440] + src21[441] + src21[442] + src21[443] + src21[444] + src21[445] + src21[446] + src21[447] + src21[448] + src21[449] + src21[450] + src21[451] + src21[452] + src21[453] + src21[454] + src21[455] + src21[456] + src21[457] + src21[458] + src21[459] + src21[460] + src21[461] + src21[462] + src21[463] + src21[464] + src21[465] + src21[466] + src21[467] + src21[468] + src21[469] + src21[470] + src21[471] + src21[472] + src21[473] + src21[474] + src21[475] + src21[476] + src21[477] + src21[478] + src21[479] + src21[480] + src21[481] + src21[482] + src21[483] + src21[484] + src21[485])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63] + src22[64] + src22[65] + src22[66] + src22[67] + src22[68] + src22[69] + src22[70] + src22[71] + src22[72] + src22[73] + src22[74] + src22[75] + src22[76] + src22[77] + src22[78] + src22[79] + src22[80] + src22[81] + src22[82] + src22[83] + src22[84] + src22[85] + src22[86] + src22[87] + src22[88] + src22[89] + src22[90] + src22[91] + src22[92] + src22[93] + src22[94] + src22[95] + src22[96] + src22[97] + src22[98] + src22[99] + src22[100] + src22[101] + src22[102] + src22[103] + src22[104] + src22[105] + src22[106] + src22[107] + src22[108] + src22[109] + src22[110] + src22[111] + src22[112] + src22[113] + src22[114] + src22[115] + src22[116] + src22[117] + src22[118] + src22[119] + src22[120] + src22[121] + src22[122] + src22[123] + src22[124] + src22[125] + src22[126] + src22[127] + src22[128] + src22[129] + src22[130] + src22[131] + src22[132] + src22[133] + src22[134] + src22[135] + src22[136] + src22[137] + src22[138] + src22[139] + src22[140] + src22[141] + src22[142] + src22[143] + src22[144] + src22[145] + src22[146] + src22[147] + src22[148] + src22[149] + src22[150] + src22[151] + src22[152] + src22[153] + src22[154] + src22[155] + src22[156] + src22[157] + src22[158] + src22[159] + src22[160] + src22[161] + src22[162] + src22[163] + src22[164] + src22[165] + src22[166] + src22[167] + src22[168] + src22[169] + src22[170] + src22[171] + src22[172] + src22[173] + src22[174] + src22[175] + src22[176] + src22[177] + src22[178] + src22[179] + src22[180] + src22[181] + src22[182] + src22[183] + src22[184] + src22[185] + src22[186] + src22[187] + src22[188] + src22[189] + src22[190] + src22[191] + src22[192] + src22[193] + src22[194] + src22[195] + src22[196] + src22[197] + src22[198] + src22[199] + src22[200] + src22[201] + src22[202] + src22[203] + src22[204] + src22[205] + src22[206] + src22[207] + src22[208] + src22[209] + src22[210] + src22[211] + src22[212] + src22[213] + src22[214] + src22[215] + src22[216] + src22[217] + src22[218] + src22[219] + src22[220] + src22[221] + src22[222] + src22[223] + src22[224] + src22[225] + src22[226] + src22[227] + src22[228] + src22[229] + src22[230] + src22[231] + src22[232] + src22[233] + src22[234] + src22[235] + src22[236] + src22[237] + src22[238] + src22[239] + src22[240] + src22[241] + src22[242] + src22[243] + src22[244] + src22[245] + src22[246] + src22[247] + src22[248] + src22[249] + src22[250] + src22[251] + src22[252] + src22[253] + src22[254] + src22[255] + src22[256] + src22[257] + src22[258] + src22[259] + src22[260] + src22[261] + src22[262] + src22[263] + src22[264] + src22[265] + src22[266] + src22[267] + src22[268] + src22[269] + src22[270] + src22[271] + src22[272] + src22[273] + src22[274] + src22[275] + src22[276] + src22[277] + src22[278] + src22[279] + src22[280] + src22[281] + src22[282] + src22[283] + src22[284] + src22[285] + src22[286] + src22[287] + src22[288] + src22[289] + src22[290] + src22[291] + src22[292] + src22[293] + src22[294] + src22[295] + src22[296] + src22[297] + src22[298] + src22[299] + src22[300] + src22[301] + src22[302] + src22[303] + src22[304] + src22[305] + src22[306] + src22[307] + src22[308] + src22[309] + src22[310] + src22[311] + src22[312] + src22[313] + src22[314] + src22[315] + src22[316] + src22[317] + src22[318] + src22[319] + src22[320] + src22[321] + src22[322] + src22[323] + src22[324] + src22[325] + src22[326] + src22[327] + src22[328] + src22[329] + src22[330] + src22[331] + src22[332] + src22[333] + src22[334] + src22[335] + src22[336] + src22[337] + src22[338] + src22[339] + src22[340] + src22[341] + src22[342] + src22[343] + src22[344] + src22[345] + src22[346] + src22[347] + src22[348] + src22[349] + src22[350] + src22[351] + src22[352] + src22[353] + src22[354] + src22[355] + src22[356] + src22[357] + src22[358] + src22[359] + src22[360] + src22[361] + src22[362] + src22[363] + src22[364] + src22[365] + src22[366] + src22[367] + src22[368] + src22[369] + src22[370] + src22[371] + src22[372] + src22[373] + src22[374] + src22[375] + src22[376] + src22[377] + src22[378] + src22[379] + src22[380] + src22[381] + src22[382] + src22[383] + src22[384] + src22[385] + src22[386] + src22[387] + src22[388] + src22[389] + src22[390] + src22[391] + src22[392] + src22[393] + src22[394] + src22[395] + src22[396] + src22[397] + src22[398] + src22[399] + src22[400] + src22[401] + src22[402] + src22[403] + src22[404] + src22[405] + src22[406] + src22[407] + src22[408] + src22[409] + src22[410] + src22[411] + src22[412] + src22[413] + src22[414] + src22[415] + src22[416] + src22[417] + src22[418] + src22[419] + src22[420] + src22[421] + src22[422] + src22[423] + src22[424] + src22[425] + src22[426] + src22[427] + src22[428] + src22[429] + src22[430] + src22[431] + src22[432] + src22[433] + src22[434] + src22[435] + src22[436] + src22[437] + src22[438] + src22[439] + src22[440] + src22[441] + src22[442] + src22[443] + src22[444] + src22[445] + src22[446] + src22[447] + src22[448] + src22[449] + src22[450] + src22[451] + src22[452] + src22[453] + src22[454] + src22[455] + src22[456] + src22[457] + src22[458] + src22[459] + src22[460] + src22[461] + src22[462] + src22[463] + src22[464] + src22[465] + src22[466] + src22[467] + src22[468] + src22[469] + src22[470] + src22[471] + src22[472] + src22[473] + src22[474] + src22[475] + src22[476] + src22[477] + src22[478] + src22[479] + src22[480] + src22[481] + src22[482] + src22[483] + src22[484] + src22[485])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63] + src23[64] + src23[65] + src23[66] + src23[67] + src23[68] + src23[69] + src23[70] + src23[71] + src23[72] + src23[73] + src23[74] + src23[75] + src23[76] + src23[77] + src23[78] + src23[79] + src23[80] + src23[81] + src23[82] + src23[83] + src23[84] + src23[85] + src23[86] + src23[87] + src23[88] + src23[89] + src23[90] + src23[91] + src23[92] + src23[93] + src23[94] + src23[95] + src23[96] + src23[97] + src23[98] + src23[99] + src23[100] + src23[101] + src23[102] + src23[103] + src23[104] + src23[105] + src23[106] + src23[107] + src23[108] + src23[109] + src23[110] + src23[111] + src23[112] + src23[113] + src23[114] + src23[115] + src23[116] + src23[117] + src23[118] + src23[119] + src23[120] + src23[121] + src23[122] + src23[123] + src23[124] + src23[125] + src23[126] + src23[127] + src23[128] + src23[129] + src23[130] + src23[131] + src23[132] + src23[133] + src23[134] + src23[135] + src23[136] + src23[137] + src23[138] + src23[139] + src23[140] + src23[141] + src23[142] + src23[143] + src23[144] + src23[145] + src23[146] + src23[147] + src23[148] + src23[149] + src23[150] + src23[151] + src23[152] + src23[153] + src23[154] + src23[155] + src23[156] + src23[157] + src23[158] + src23[159] + src23[160] + src23[161] + src23[162] + src23[163] + src23[164] + src23[165] + src23[166] + src23[167] + src23[168] + src23[169] + src23[170] + src23[171] + src23[172] + src23[173] + src23[174] + src23[175] + src23[176] + src23[177] + src23[178] + src23[179] + src23[180] + src23[181] + src23[182] + src23[183] + src23[184] + src23[185] + src23[186] + src23[187] + src23[188] + src23[189] + src23[190] + src23[191] + src23[192] + src23[193] + src23[194] + src23[195] + src23[196] + src23[197] + src23[198] + src23[199] + src23[200] + src23[201] + src23[202] + src23[203] + src23[204] + src23[205] + src23[206] + src23[207] + src23[208] + src23[209] + src23[210] + src23[211] + src23[212] + src23[213] + src23[214] + src23[215] + src23[216] + src23[217] + src23[218] + src23[219] + src23[220] + src23[221] + src23[222] + src23[223] + src23[224] + src23[225] + src23[226] + src23[227] + src23[228] + src23[229] + src23[230] + src23[231] + src23[232] + src23[233] + src23[234] + src23[235] + src23[236] + src23[237] + src23[238] + src23[239] + src23[240] + src23[241] + src23[242] + src23[243] + src23[244] + src23[245] + src23[246] + src23[247] + src23[248] + src23[249] + src23[250] + src23[251] + src23[252] + src23[253] + src23[254] + src23[255] + src23[256] + src23[257] + src23[258] + src23[259] + src23[260] + src23[261] + src23[262] + src23[263] + src23[264] + src23[265] + src23[266] + src23[267] + src23[268] + src23[269] + src23[270] + src23[271] + src23[272] + src23[273] + src23[274] + src23[275] + src23[276] + src23[277] + src23[278] + src23[279] + src23[280] + src23[281] + src23[282] + src23[283] + src23[284] + src23[285] + src23[286] + src23[287] + src23[288] + src23[289] + src23[290] + src23[291] + src23[292] + src23[293] + src23[294] + src23[295] + src23[296] + src23[297] + src23[298] + src23[299] + src23[300] + src23[301] + src23[302] + src23[303] + src23[304] + src23[305] + src23[306] + src23[307] + src23[308] + src23[309] + src23[310] + src23[311] + src23[312] + src23[313] + src23[314] + src23[315] + src23[316] + src23[317] + src23[318] + src23[319] + src23[320] + src23[321] + src23[322] + src23[323] + src23[324] + src23[325] + src23[326] + src23[327] + src23[328] + src23[329] + src23[330] + src23[331] + src23[332] + src23[333] + src23[334] + src23[335] + src23[336] + src23[337] + src23[338] + src23[339] + src23[340] + src23[341] + src23[342] + src23[343] + src23[344] + src23[345] + src23[346] + src23[347] + src23[348] + src23[349] + src23[350] + src23[351] + src23[352] + src23[353] + src23[354] + src23[355] + src23[356] + src23[357] + src23[358] + src23[359] + src23[360] + src23[361] + src23[362] + src23[363] + src23[364] + src23[365] + src23[366] + src23[367] + src23[368] + src23[369] + src23[370] + src23[371] + src23[372] + src23[373] + src23[374] + src23[375] + src23[376] + src23[377] + src23[378] + src23[379] + src23[380] + src23[381] + src23[382] + src23[383] + src23[384] + src23[385] + src23[386] + src23[387] + src23[388] + src23[389] + src23[390] + src23[391] + src23[392] + src23[393] + src23[394] + src23[395] + src23[396] + src23[397] + src23[398] + src23[399] + src23[400] + src23[401] + src23[402] + src23[403] + src23[404] + src23[405] + src23[406] + src23[407] + src23[408] + src23[409] + src23[410] + src23[411] + src23[412] + src23[413] + src23[414] + src23[415] + src23[416] + src23[417] + src23[418] + src23[419] + src23[420] + src23[421] + src23[422] + src23[423] + src23[424] + src23[425] + src23[426] + src23[427] + src23[428] + src23[429] + src23[430] + src23[431] + src23[432] + src23[433] + src23[434] + src23[435] + src23[436] + src23[437] + src23[438] + src23[439] + src23[440] + src23[441] + src23[442] + src23[443] + src23[444] + src23[445] + src23[446] + src23[447] + src23[448] + src23[449] + src23[450] + src23[451] + src23[452] + src23[453] + src23[454] + src23[455] + src23[456] + src23[457] + src23[458] + src23[459] + src23[460] + src23[461] + src23[462] + src23[463] + src23[464] + src23[465] + src23[466] + src23[467] + src23[468] + src23[469] + src23[470] + src23[471] + src23[472] + src23[473] + src23[474] + src23[475] + src23[476] + src23[477] + src23[478] + src23[479] + src23[480] + src23[481] + src23[482] + src23[483] + src23[484] + src23[485])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63] + src24[64] + src24[65] + src24[66] + src24[67] + src24[68] + src24[69] + src24[70] + src24[71] + src24[72] + src24[73] + src24[74] + src24[75] + src24[76] + src24[77] + src24[78] + src24[79] + src24[80] + src24[81] + src24[82] + src24[83] + src24[84] + src24[85] + src24[86] + src24[87] + src24[88] + src24[89] + src24[90] + src24[91] + src24[92] + src24[93] + src24[94] + src24[95] + src24[96] + src24[97] + src24[98] + src24[99] + src24[100] + src24[101] + src24[102] + src24[103] + src24[104] + src24[105] + src24[106] + src24[107] + src24[108] + src24[109] + src24[110] + src24[111] + src24[112] + src24[113] + src24[114] + src24[115] + src24[116] + src24[117] + src24[118] + src24[119] + src24[120] + src24[121] + src24[122] + src24[123] + src24[124] + src24[125] + src24[126] + src24[127] + src24[128] + src24[129] + src24[130] + src24[131] + src24[132] + src24[133] + src24[134] + src24[135] + src24[136] + src24[137] + src24[138] + src24[139] + src24[140] + src24[141] + src24[142] + src24[143] + src24[144] + src24[145] + src24[146] + src24[147] + src24[148] + src24[149] + src24[150] + src24[151] + src24[152] + src24[153] + src24[154] + src24[155] + src24[156] + src24[157] + src24[158] + src24[159] + src24[160] + src24[161] + src24[162] + src24[163] + src24[164] + src24[165] + src24[166] + src24[167] + src24[168] + src24[169] + src24[170] + src24[171] + src24[172] + src24[173] + src24[174] + src24[175] + src24[176] + src24[177] + src24[178] + src24[179] + src24[180] + src24[181] + src24[182] + src24[183] + src24[184] + src24[185] + src24[186] + src24[187] + src24[188] + src24[189] + src24[190] + src24[191] + src24[192] + src24[193] + src24[194] + src24[195] + src24[196] + src24[197] + src24[198] + src24[199] + src24[200] + src24[201] + src24[202] + src24[203] + src24[204] + src24[205] + src24[206] + src24[207] + src24[208] + src24[209] + src24[210] + src24[211] + src24[212] + src24[213] + src24[214] + src24[215] + src24[216] + src24[217] + src24[218] + src24[219] + src24[220] + src24[221] + src24[222] + src24[223] + src24[224] + src24[225] + src24[226] + src24[227] + src24[228] + src24[229] + src24[230] + src24[231] + src24[232] + src24[233] + src24[234] + src24[235] + src24[236] + src24[237] + src24[238] + src24[239] + src24[240] + src24[241] + src24[242] + src24[243] + src24[244] + src24[245] + src24[246] + src24[247] + src24[248] + src24[249] + src24[250] + src24[251] + src24[252] + src24[253] + src24[254] + src24[255] + src24[256] + src24[257] + src24[258] + src24[259] + src24[260] + src24[261] + src24[262] + src24[263] + src24[264] + src24[265] + src24[266] + src24[267] + src24[268] + src24[269] + src24[270] + src24[271] + src24[272] + src24[273] + src24[274] + src24[275] + src24[276] + src24[277] + src24[278] + src24[279] + src24[280] + src24[281] + src24[282] + src24[283] + src24[284] + src24[285] + src24[286] + src24[287] + src24[288] + src24[289] + src24[290] + src24[291] + src24[292] + src24[293] + src24[294] + src24[295] + src24[296] + src24[297] + src24[298] + src24[299] + src24[300] + src24[301] + src24[302] + src24[303] + src24[304] + src24[305] + src24[306] + src24[307] + src24[308] + src24[309] + src24[310] + src24[311] + src24[312] + src24[313] + src24[314] + src24[315] + src24[316] + src24[317] + src24[318] + src24[319] + src24[320] + src24[321] + src24[322] + src24[323] + src24[324] + src24[325] + src24[326] + src24[327] + src24[328] + src24[329] + src24[330] + src24[331] + src24[332] + src24[333] + src24[334] + src24[335] + src24[336] + src24[337] + src24[338] + src24[339] + src24[340] + src24[341] + src24[342] + src24[343] + src24[344] + src24[345] + src24[346] + src24[347] + src24[348] + src24[349] + src24[350] + src24[351] + src24[352] + src24[353] + src24[354] + src24[355] + src24[356] + src24[357] + src24[358] + src24[359] + src24[360] + src24[361] + src24[362] + src24[363] + src24[364] + src24[365] + src24[366] + src24[367] + src24[368] + src24[369] + src24[370] + src24[371] + src24[372] + src24[373] + src24[374] + src24[375] + src24[376] + src24[377] + src24[378] + src24[379] + src24[380] + src24[381] + src24[382] + src24[383] + src24[384] + src24[385] + src24[386] + src24[387] + src24[388] + src24[389] + src24[390] + src24[391] + src24[392] + src24[393] + src24[394] + src24[395] + src24[396] + src24[397] + src24[398] + src24[399] + src24[400] + src24[401] + src24[402] + src24[403] + src24[404] + src24[405] + src24[406] + src24[407] + src24[408] + src24[409] + src24[410] + src24[411] + src24[412] + src24[413] + src24[414] + src24[415] + src24[416] + src24[417] + src24[418] + src24[419] + src24[420] + src24[421] + src24[422] + src24[423] + src24[424] + src24[425] + src24[426] + src24[427] + src24[428] + src24[429] + src24[430] + src24[431] + src24[432] + src24[433] + src24[434] + src24[435] + src24[436] + src24[437] + src24[438] + src24[439] + src24[440] + src24[441] + src24[442] + src24[443] + src24[444] + src24[445] + src24[446] + src24[447] + src24[448] + src24[449] + src24[450] + src24[451] + src24[452] + src24[453] + src24[454] + src24[455] + src24[456] + src24[457] + src24[458] + src24[459] + src24[460] + src24[461] + src24[462] + src24[463] + src24[464] + src24[465] + src24[466] + src24[467] + src24[468] + src24[469] + src24[470] + src24[471] + src24[472] + src24[473] + src24[474] + src24[475] + src24[476] + src24[477] + src24[478] + src24[479] + src24[480] + src24[481] + src24[482] + src24[483] + src24[484] + src24[485])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63] + src25[64] + src25[65] + src25[66] + src25[67] + src25[68] + src25[69] + src25[70] + src25[71] + src25[72] + src25[73] + src25[74] + src25[75] + src25[76] + src25[77] + src25[78] + src25[79] + src25[80] + src25[81] + src25[82] + src25[83] + src25[84] + src25[85] + src25[86] + src25[87] + src25[88] + src25[89] + src25[90] + src25[91] + src25[92] + src25[93] + src25[94] + src25[95] + src25[96] + src25[97] + src25[98] + src25[99] + src25[100] + src25[101] + src25[102] + src25[103] + src25[104] + src25[105] + src25[106] + src25[107] + src25[108] + src25[109] + src25[110] + src25[111] + src25[112] + src25[113] + src25[114] + src25[115] + src25[116] + src25[117] + src25[118] + src25[119] + src25[120] + src25[121] + src25[122] + src25[123] + src25[124] + src25[125] + src25[126] + src25[127] + src25[128] + src25[129] + src25[130] + src25[131] + src25[132] + src25[133] + src25[134] + src25[135] + src25[136] + src25[137] + src25[138] + src25[139] + src25[140] + src25[141] + src25[142] + src25[143] + src25[144] + src25[145] + src25[146] + src25[147] + src25[148] + src25[149] + src25[150] + src25[151] + src25[152] + src25[153] + src25[154] + src25[155] + src25[156] + src25[157] + src25[158] + src25[159] + src25[160] + src25[161] + src25[162] + src25[163] + src25[164] + src25[165] + src25[166] + src25[167] + src25[168] + src25[169] + src25[170] + src25[171] + src25[172] + src25[173] + src25[174] + src25[175] + src25[176] + src25[177] + src25[178] + src25[179] + src25[180] + src25[181] + src25[182] + src25[183] + src25[184] + src25[185] + src25[186] + src25[187] + src25[188] + src25[189] + src25[190] + src25[191] + src25[192] + src25[193] + src25[194] + src25[195] + src25[196] + src25[197] + src25[198] + src25[199] + src25[200] + src25[201] + src25[202] + src25[203] + src25[204] + src25[205] + src25[206] + src25[207] + src25[208] + src25[209] + src25[210] + src25[211] + src25[212] + src25[213] + src25[214] + src25[215] + src25[216] + src25[217] + src25[218] + src25[219] + src25[220] + src25[221] + src25[222] + src25[223] + src25[224] + src25[225] + src25[226] + src25[227] + src25[228] + src25[229] + src25[230] + src25[231] + src25[232] + src25[233] + src25[234] + src25[235] + src25[236] + src25[237] + src25[238] + src25[239] + src25[240] + src25[241] + src25[242] + src25[243] + src25[244] + src25[245] + src25[246] + src25[247] + src25[248] + src25[249] + src25[250] + src25[251] + src25[252] + src25[253] + src25[254] + src25[255] + src25[256] + src25[257] + src25[258] + src25[259] + src25[260] + src25[261] + src25[262] + src25[263] + src25[264] + src25[265] + src25[266] + src25[267] + src25[268] + src25[269] + src25[270] + src25[271] + src25[272] + src25[273] + src25[274] + src25[275] + src25[276] + src25[277] + src25[278] + src25[279] + src25[280] + src25[281] + src25[282] + src25[283] + src25[284] + src25[285] + src25[286] + src25[287] + src25[288] + src25[289] + src25[290] + src25[291] + src25[292] + src25[293] + src25[294] + src25[295] + src25[296] + src25[297] + src25[298] + src25[299] + src25[300] + src25[301] + src25[302] + src25[303] + src25[304] + src25[305] + src25[306] + src25[307] + src25[308] + src25[309] + src25[310] + src25[311] + src25[312] + src25[313] + src25[314] + src25[315] + src25[316] + src25[317] + src25[318] + src25[319] + src25[320] + src25[321] + src25[322] + src25[323] + src25[324] + src25[325] + src25[326] + src25[327] + src25[328] + src25[329] + src25[330] + src25[331] + src25[332] + src25[333] + src25[334] + src25[335] + src25[336] + src25[337] + src25[338] + src25[339] + src25[340] + src25[341] + src25[342] + src25[343] + src25[344] + src25[345] + src25[346] + src25[347] + src25[348] + src25[349] + src25[350] + src25[351] + src25[352] + src25[353] + src25[354] + src25[355] + src25[356] + src25[357] + src25[358] + src25[359] + src25[360] + src25[361] + src25[362] + src25[363] + src25[364] + src25[365] + src25[366] + src25[367] + src25[368] + src25[369] + src25[370] + src25[371] + src25[372] + src25[373] + src25[374] + src25[375] + src25[376] + src25[377] + src25[378] + src25[379] + src25[380] + src25[381] + src25[382] + src25[383] + src25[384] + src25[385] + src25[386] + src25[387] + src25[388] + src25[389] + src25[390] + src25[391] + src25[392] + src25[393] + src25[394] + src25[395] + src25[396] + src25[397] + src25[398] + src25[399] + src25[400] + src25[401] + src25[402] + src25[403] + src25[404] + src25[405] + src25[406] + src25[407] + src25[408] + src25[409] + src25[410] + src25[411] + src25[412] + src25[413] + src25[414] + src25[415] + src25[416] + src25[417] + src25[418] + src25[419] + src25[420] + src25[421] + src25[422] + src25[423] + src25[424] + src25[425] + src25[426] + src25[427] + src25[428] + src25[429] + src25[430] + src25[431] + src25[432] + src25[433] + src25[434] + src25[435] + src25[436] + src25[437] + src25[438] + src25[439] + src25[440] + src25[441] + src25[442] + src25[443] + src25[444] + src25[445] + src25[446] + src25[447] + src25[448] + src25[449] + src25[450] + src25[451] + src25[452] + src25[453] + src25[454] + src25[455] + src25[456] + src25[457] + src25[458] + src25[459] + src25[460] + src25[461] + src25[462] + src25[463] + src25[464] + src25[465] + src25[466] + src25[467] + src25[468] + src25[469] + src25[470] + src25[471] + src25[472] + src25[473] + src25[474] + src25[475] + src25[476] + src25[477] + src25[478] + src25[479] + src25[480] + src25[481] + src25[482] + src25[483] + src25[484] + src25[485])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63] + src26[64] + src26[65] + src26[66] + src26[67] + src26[68] + src26[69] + src26[70] + src26[71] + src26[72] + src26[73] + src26[74] + src26[75] + src26[76] + src26[77] + src26[78] + src26[79] + src26[80] + src26[81] + src26[82] + src26[83] + src26[84] + src26[85] + src26[86] + src26[87] + src26[88] + src26[89] + src26[90] + src26[91] + src26[92] + src26[93] + src26[94] + src26[95] + src26[96] + src26[97] + src26[98] + src26[99] + src26[100] + src26[101] + src26[102] + src26[103] + src26[104] + src26[105] + src26[106] + src26[107] + src26[108] + src26[109] + src26[110] + src26[111] + src26[112] + src26[113] + src26[114] + src26[115] + src26[116] + src26[117] + src26[118] + src26[119] + src26[120] + src26[121] + src26[122] + src26[123] + src26[124] + src26[125] + src26[126] + src26[127] + src26[128] + src26[129] + src26[130] + src26[131] + src26[132] + src26[133] + src26[134] + src26[135] + src26[136] + src26[137] + src26[138] + src26[139] + src26[140] + src26[141] + src26[142] + src26[143] + src26[144] + src26[145] + src26[146] + src26[147] + src26[148] + src26[149] + src26[150] + src26[151] + src26[152] + src26[153] + src26[154] + src26[155] + src26[156] + src26[157] + src26[158] + src26[159] + src26[160] + src26[161] + src26[162] + src26[163] + src26[164] + src26[165] + src26[166] + src26[167] + src26[168] + src26[169] + src26[170] + src26[171] + src26[172] + src26[173] + src26[174] + src26[175] + src26[176] + src26[177] + src26[178] + src26[179] + src26[180] + src26[181] + src26[182] + src26[183] + src26[184] + src26[185] + src26[186] + src26[187] + src26[188] + src26[189] + src26[190] + src26[191] + src26[192] + src26[193] + src26[194] + src26[195] + src26[196] + src26[197] + src26[198] + src26[199] + src26[200] + src26[201] + src26[202] + src26[203] + src26[204] + src26[205] + src26[206] + src26[207] + src26[208] + src26[209] + src26[210] + src26[211] + src26[212] + src26[213] + src26[214] + src26[215] + src26[216] + src26[217] + src26[218] + src26[219] + src26[220] + src26[221] + src26[222] + src26[223] + src26[224] + src26[225] + src26[226] + src26[227] + src26[228] + src26[229] + src26[230] + src26[231] + src26[232] + src26[233] + src26[234] + src26[235] + src26[236] + src26[237] + src26[238] + src26[239] + src26[240] + src26[241] + src26[242] + src26[243] + src26[244] + src26[245] + src26[246] + src26[247] + src26[248] + src26[249] + src26[250] + src26[251] + src26[252] + src26[253] + src26[254] + src26[255] + src26[256] + src26[257] + src26[258] + src26[259] + src26[260] + src26[261] + src26[262] + src26[263] + src26[264] + src26[265] + src26[266] + src26[267] + src26[268] + src26[269] + src26[270] + src26[271] + src26[272] + src26[273] + src26[274] + src26[275] + src26[276] + src26[277] + src26[278] + src26[279] + src26[280] + src26[281] + src26[282] + src26[283] + src26[284] + src26[285] + src26[286] + src26[287] + src26[288] + src26[289] + src26[290] + src26[291] + src26[292] + src26[293] + src26[294] + src26[295] + src26[296] + src26[297] + src26[298] + src26[299] + src26[300] + src26[301] + src26[302] + src26[303] + src26[304] + src26[305] + src26[306] + src26[307] + src26[308] + src26[309] + src26[310] + src26[311] + src26[312] + src26[313] + src26[314] + src26[315] + src26[316] + src26[317] + src26[318] + src26[319] + src26[320] + src26[321] + src26[322] + src26[323] + src26[324] + src26[325] + src26[326] + src26[327] + src26[328] + src26[329] + src26[330] + src26[331] + src26[332] + src26[333] + src26[334] + src26[335] + src26[336] + src26[337] + src26[338] + src26[339] + src26[340] + src26[341] + src26[342] + src26[343] + src26[344] + src26[345] + src26[346] + src26[347] + src26[348] + src26[349] + src26[350] + src26[351] + src26[352] + src26[353] + src26[354] + src26[355] + src26[356] + src26[357] + src26[358] + src26[359] + src26[360] + src26[361] + src26[362] + src26[363] + src26[364] + src26[365] + src26[366] + src26[367] + src26[368] + src26[369] + src26[370] + src26[371] + src26[372] + src26[373] + src26[374] + src26[375] + src26[376] + src26[377] + src26[378] + src26[379] + src26[380] + src26[381] + src26[382] + src26[383] + src26[384] + src26[385] + src26[386] + src26[387] + src26[388] + src26[389] + src26[390] + src26[391] + src26[392] + src26[393] + src26[394] + src26[395] + src26[396] + src26[397] + src26[398] + src26[399] + src26[400] + src26[401] + src26[402] + src26[403] + src26[404] + src26[405] + src26[406] + src26[407] + src26[408] + src26[409] + src26[410] + src26[411] + src26[412] + src26[413] + src26[414] + src26[415] + src26[416] + src26[417] + src26[418] + src26[419] + src26[420] + src26[421] + src26[422] + src26[423] + src26[424] + src26[425] + src26[426] + src26[427] + src26[428] + src26[429] + src26[430] + src26[431] + src26[432] + src26[433] + src26[434] + src26[435] + src26[436] + src26[437] + src26[438] + src26[439] + src26[440] + src26[441] + src26[442] + src26[443] + src26[444] + src26[445] + src26[446] + src26[447] + src26[448] + src26[449] + src26[450] + src26[451] + src26[452] + src26[453] + src26[454] + src26[455] + src26[456] + src26[457] + src26[458] + src26[459] + src26[460] + src26[461] + src26[462] + src26[463] + src26[464] + src26[465] + src26[466] + src26[467] + src26[468] + src26[469] + src26[470] + src26[471] + src26[472] + src26[473] + src26[474] + src26[475] + src26[476] + src26[477] + src26[478] + src26[479] + src26[480] + src26[481] + src26[482] + src26[483] + src26[484] + src26[485])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63] + src27[64] + src27[65] + src27[66] + src27[67] + src27[68] + src27[69] + src27[70] + src27[71] + src27[72] + src27[73] + src27[74] + src27[75] + src27[76] + src27[77] + src27[78] + src27[79] + src27[80] + src27[81] + src27[82] + src27[83] + src27[84] + src27[85] + src27[86] + src27[87] + src27[88] + src27[89] + src27[90] + src27[91] + src27[92] + src27[93] + src27[94] + src27[95] + src27[96] + src27[97] + src27[98] + src27[99] + src27[100] + src27[101] + src27[102] + src27[103] + src27[104] + src27[105] + src27[106] + src27[107] + src27[108] + src27[109] + src27[110] + src27[111] + src27[112] + src27[113] + src27[114] + src27[115] + src27[116] + src27[117] + src27[118] + src27[119] + src27[120] + src27[121] + src27[122] + src27[123] + src27[124] + src27[125] + src27[126] + src27[127] + src27[128] + src27[129] + src27[130] + src27[131] + src27[132] + src27[133] + src27[134] + src27[135] + src27[136] + src27[137] + src27[138] + src27[139] + src27[140] + src27[141] + src27[142] + src27[143] + src27[144] + src27[145] + src27[146] + src27[147] + src27[148] + src27[149] + src27[150] + src27[151] + src27[152] + src27[153] + src27[154] + src27[155] + src27[156] + src27[157] + src27[158] + src27[159] + src27[160] + src27[161] + src27[162] + src27[163] + src27[164] + src27[165] + src27[166] + src27[167] + src27[168] + src27[169] + src27[170] + src27[171] + src27[172] + src27[173] + src27[174] + src27[175] + src27[176] + src27[177] + src27[178] + src27[179] + src27[180] + src27[181] + src27[182] + src27[183] + src27[184] + src27[185] + src27[186] + src27[187] + src27[188] + src27[189] + src27[190] + src27[191] + src27[192] + src27[193] + src27[194] + src27[195] + src27[196] + src27[197] + src27[198] + src27[199] + src27[200] + src27[201] + src27[202] + src27[203] + src27[204] + src27[205] + src27[206] + src27[207] + src27[208] + src27[209] + src27[210] + src27[211] + src27[212] + src27[213] + src27[214] + src27[215] + src27[216] + src27[217] + src27[218] + src27[219] + src27[220] + src27[221] + src27[222] + src27[223] + src27[224] + src27[225] + src27[226] + src27[227] + src27[228] + src27[229] + src27[230] + src27[231] + src27[232] + src27[233] + src27[234] + src27[235] + src27[236] + src27[237] + src27[238] + src27[239] + src27[240] + src27[241] + src27[242] + src27[243] + src27[244] + src27[245] + src27[246] + src27[247] + src27[248] + src27[249] + src27[250] + src27[251] + src27[252] + src27[253] + src27[254] + src27[255] + src27[256] + src27[257] + src27[258] + src27[259] + src27[260] + src27[261] + src27[262] + src27[263] + src27[264] + src27[265] + src27[266] + src27[267] + src27[268] + src27[269] + src27[270] + src27[271] + src27[272] + src27[273] + src27[274] + src27[275] + src27[276] + src27[277] + src27[278] + src27[279] + src27[280] + src27[281] + src27[282] + src27[283] + src27[284] + src27[285] + src27[286] + src27[287] + src27[288] + src27[289] + src27[290] + src27[291] + src27[292] + src27[293] + src27[294] + src27[295] + src27[296] + src27[297] + src27[298] + src27[299] + src27[300] + src27[301] + src27[302] + src27[303] + src27[304] + src27[305] + src27[306] + src27[307] + src27[308] + src27[309] + src27[310] + src27[311] + src27[312] + src27[313] + src27[314] + src27[315] + src27[316] + src27[317] + src27[318] + src27[319] + src27[320] + src27[321] + src27[322] + src27[323] + src27[324] + src27[325] + src27[326] + src27[327] + src27[328] + src27[329] + src27[330] + src27[331] + src27[332] + src27[333] + src27[334] + src27[335] + src27[336] + src27[337] + src27[338] + src27[339] + src27[340] + src27[341] + src27[342] + src27[343] + src27[344] + src27[345] + src27[346] + src27[347] + src27[348] + src27[349] + src27[350] + src27[351] + src27[352] + src27[353] + src27[354] + src27[355] + src27[356] + src27[357] + src27[358] + src27[359] + src27[360] + src27[361] + src27[362] + src27[363] + src27[364] + src27[365] + src27[366] + src27[367] + src27[368] + src27[369] + src27[370] + src27[371] + src27[372] + src27[373] + src27[374] + src27[375] + src27[376] + src27[377] + src27[378] + src27[379] + src27[380] + src27[381] + src27[382] + src27[383] + src27[384] + src27[385] + src27[386] + src27[387] + src27[388] + src27[389] + src27[390] + src27[391] + src27[392] + src27[393] + src27[394] + src27[395] + src27[396] + src27[397] + src27[398] + src27[399] + src27[400] + src27[401] + src27[402] + src27[403] + src27[404] + src27[405] + src27[406] + src27[407] + src27[408] + src27[409] + src27[410] + src27[411] + src27[412] + src27[413] + src27[414] + src27[415] + src27[416] + src27[417] + src27[418] + src27[419] + src27[420] + src27[421] + src27[422] + src27[423] + src27[424] + src27[425] + src27[426] + src27[427] + src27[428] + src27[429] + src27[430] + src27[431] + src27[432] + src27[433] + src27[434] + src27[435] + src27[436] + src27[437] + src27[438] + src27[439] + src27[440] + src27[441] + src27[442] + src27[443] + src27[444] + src27[445] + src27[446] + src27[447] + src27[448] + src27[449] + src27[450] + src27[451] + src27[452] + src27[453] + src27[454] + src27[455] + src27[456] + src27[457] + src27[458] + src27[459] + src27[460] + src27[461] + src27[462] + src27[463] + src27[464] + src27[465] + src27[466] + src27[467] + src27[468] + src27[469] + src27[470] + src27[471] + src27[472] + src27[473] + src27[474] + src27[475] + src27[476] + src27[477] + src27[478] + src27[479] + src27[480] + src27[481] + src27[482] + src27[483] + src27[484] + src27[485])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63] + src28[64] + src28[65] + src28[66] + src28[67] + src28[68] + src28[69] + src28[70] + src28[71] + src28[72] + src28[73] + src28[74] + src28[75] + src28[76] + src28[77] + src28[78] + src28[79] + src28[80] + src28[81] + src28[82] + src28[83] + src28[84] + src28[85] + src28[86] + src28[87] + src28[88] + src28[89] + src28[90] + src28[91] + src28[92] + src28[93] + src28[94] + src28[95] + src28[96] + src28[97] + src28[98] + src28[99] + src28[100] + src28[101] + src28[102] + src28[103] + src28[104] + src28[105] + src28[106] + src28[107] + src28[108] + src28[109] + src28[110] + src28[111] + src28[112] + src28[113] + src28[114] + src28[115] + src28[116] + src28[117] + src28[118] + src28[119] + src28[120] + src28[121] + src28[122] + src28[123] + src28[124] + src28[125] + src28[126] + src28[127] + src28[128] + src28[129] + src28[130] + src28[131] + src28[132] + src28[133] + src28[134] + src28[135] + src28[136] + src28[137] + src28[138] + src28[139] + src28[140] + src28[141] + src28[142] + src28[143] + src28[144] + src28[145] + src28[146] + src28[147] + src28[148] + src28[149] + src28[150] + src28[151] + src28[152] + src28[153] + src28[154] + src28[155] + src28[156] + src28[157] + src28[158] + src28[159] + src28[160] + src28[161] + src28[162] + src28[163] + src28[164] + src28[165] + src28[166] + src28[167] + src28[168] + src28[169] + src28[170] + src28[171] + src28[172] + src28[173] + src28[174] + src28[175] + src28[176] + src28[177] + src28[178] + src28[179] + src28[180] + src28[181] + src28[182] + src28[183] + src28[184] + src28[185] + src28[186] + src28[187] + src28[188] + src28[189] + src28[190] + src28[191] + src28[192] + src28[193] + src28[194] + src28[195] + src28[196] + src28[197] + src28[198] + src28[199] + src28[200] + src28[201] + src28[202] + src28[203] + src28[204] + src28[205] + src28[206] + src28[207] + src28[208] + src28[209] + src28[210] + src28[211] + src28[212] + src28[213] + src28[214] + src28[215] + src28[216] + src28[217] + src28[218] + src28[219] + src28[220] + src28[221] + src28[222] + src28[223] + src28[224] + src28[225] + src28[226] + src28[227] + src28[228] + src28[229] + src28[230] + src28[231] + src28[232] + src28[233] + src28[234] + src28[235] + src28[236] + src28[237] + src28[238] + src28[239] + src28[240] + src28[241] + src28[242] + src28[243] + src28[244] + src28[245] + src28[246] + src28[247] + src28[248] + src28[249] + src28[250] + src28[251] + src28[252] + src28[253] + src28[254] + src28[255] + src28[256] + src28[257] + src28[258] + src28[259] + src28[260] + src28[261] + src28[262] + src28[263] + src28[264] + src28[265] + src28[266] + src28[267] + src28[268] + src28[269] + src28[270] + src28[271] + src28[272] + src28[273] + src28[274] + src28[275] + src28[276] + src28[277] + src28[278] + src28[279] + src28[280] + src28[281] + src28[282] + src28[283] + src28[284] + src28[285] + src28[286] + src28[287] + src28[288] + src28[289] + src28[290] + src28[291] + src28[292] + src28[293] + src28[294] + src28[295] + src28[296] + src28[297] + src28[298] + src28[299] + src28[300] + src28[301] + src28[302] + src28[303] + src28[304] + src28[305] + src28[306] + src28[307] + src28[308] + src28[309] + src28[310] + src28[311] + src28[312] + src28[313] + src28[314] + src28[315] + src28[316] + src28[317] + src28[318] + src28[319] + src28[320] + src28[321] + src28[322] + src28[323] + src28[324] + src28[325] + src28[326] + src28[327] + src28[328] + src28[329] + src28[330] + src28[331] + src28[332] + src28[333] + src28[334] + src28[335] + src28[336] + src28[337] + src28[338] + src28[339] + src28[340] + src28[341] + src28[342] + src28[343] + src28[344] + src28[345] + src28[346] + src28[347] + src28[348] + src28[349] + src28[350] + src28[351] + src28[352] + src28[353] + src28[354] + src28[355] + src28[356] + src28[357] + src28[358] + src28[359] + src28[360] + src28[361] + src28[362] + src28[363] + src28[364] + src28[365] + src28[366] + src28[367] + src28[368] + src28[369] + src28[370] + src28[371] + src28[372] + src28[373] + src28[374] + src28[375] + src28[376] + src28[377] + src28[378] + src28[379] + src28[380] + src28[381] + src28[382] + src28[383] + src28[384] + src28[385] + src28[386] + src28[387] + src28[388] + src28[389] + src28[390] + src28[391] + src28[392] + src28[393] + src28[394] + src28[395] + src28[396] + src28[397] + src28[398] + src28[399] + src28[400] + src28[401] + src28[402] + src28[403] + src28[404] + src28[405] + src28[406] + src28[407] + src28[408] + src28[409] + src28[410] + src28[411] + src28[412] + src28[413] + src28[414] + src28[415] + src28[416] + src28[417] + src28[418] + src28[419] + src28[420] + src28[421] + src28[422] + src28[423] + src28[424] + src28[425] + src28[426] + src28[427] + src28[428] + src28[429] + src28[430] + src28[431] + src28[432] + src28[433] + src28[434] + src28[435] + src28[436] + src28[437] + src28[438] + src28[439] + src28[440] + src28[441] + src28[442] + src28[443] + src28[444] + src28[445] + src28[446] + src28[447] + src28[448] + src28[449] + src28[450] + src28[451] + src28[452] + src28[453] + src28[454] + src28[455] + src28[456] + src28[457] + src28[458] + src28[459] + src28[460] + src28[461] + src28[462] + src28[463] + src28[464] + src28[465] + src28[466] + src28[467] + src28[468] + src28[469] + src28[470] + src28[471] + src28[472] + src28[473] + src28[474] + src28[475] + src28[476] + src28[477] + src28[478] + src28[479] + src28[480] + src28[481] + src28[482] + src28[483] + src28[484] + src28[485])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63] + src29[64] + src29[65] + src29[66] + src29[67] + src29[68] + src29[69] + src29[70] + src29[71] + src29[72] + src29[73] + src29[74] + src29[75] + src29[76] + src29[77] + src29[78] + src29[79] + src29[80] + src29[81] + src29[82] + src29[83] + src29[84] + src29[85] + src29[86] + src29[87] + src29[88] + src29[89] + src29[90] + src29[91] + src29[92] + src29[93] + src29[94] + src29[95] + src29[96] + src29[97] + src29[98] + src29[99] + src29[100] + src29[101] + src29[102] + src29[103] + src29[104] + src29[105] + src29[106] + src29[107] + src29[108] + src29[109] + src29[110] + src29[111] + src29[112] + src29[113] + src29[114] + src29[115] + src29[116] + src29[117] + src29[118] + src29[119] + src29[120] + src29[121] + src29[122] + src29[123] + src29[124] + src29[125] + src29[126] + src29[127] + src29[128] + src29[129] + src29[130] + src29[131] + src29[132] + src29[133] + src29[134] + src29[135] + src29[136] + src29[137] + src29[138] + src29[139] + src29[140] + src29[141] + src29[142] + src29[143] + src29[144] + src29[145] + src29[146] + src29[147] + src29[148] + src29[149] + src29[150] + src29[151] + src29[152] + src29[153] + src29[154] + src29[155] + src29[156] + src29[157] + src29[158] + src29[159] + src29[160] + src29[161] + src29[162] + src29[163] + src29[164] + src29[165] + src29[166] + src29[167] + src29[168] + src29[169] + src29[170] + src29[171] + src29[172] + src29[173] + src29[174] + src29[175] + src29[176] + src29[177] + src29[178] + src29[179] + src29[180] + src29[181] + src29[182] + src29[183] + src29[184] + src29[185] + src29[186] + src29[187] + src29[188] + src29[189] + src29[190] + src29[191] + src29[192] + src29[193] + src29[194] + src29[195] + src29[196] + src29[197] + src29[198] + src29[199] + src29[200] + src29[201] + src29[202] + src29[203] + src29[204] + src29[205] + src29[206] + src29[207] + src29[208] + src29[209] + src29[210] + src29[211] + src29[212] + src29[213] + src29[214] + src29[215] + src29[216] + src29[217] + src29[218] + src29[219] + src29[220] + src29[221] + src29[222] + src29[223] + src29[224] + src29[225] + src29[226] + src29[227] + src29[228] + src29[229] + src29[230] + src29[231] + src29[232] + src29[233] + src29[234] + src29[235] + src29[236] + src29[237] + src29[238] + src29[239] + src29[240] + src29[241] + src29[242] + src29[243] + src29[244] + src29[245] + src29[246] + src29[247] + src29[248] + src29[249] + src29[250] + src29[251] + src29[252] + src29[253] + src29[254] + src29[255] + src29[256] + src29[257] + src29[258] + src29[259] + src29[260] + src29[261] + src29[262] + src29[263] + src29[264] + src29[265] + src29[266] + src29[267] + src29[268] + src29[269] + src29[270] + src29[271] + src29[272] + src29[273] + src29[274] + src29[275] + src29[276] + src29[277] + src29[278] + src29[279] + src29[280] + src29[281] + src29[282] + src29[283] + src29[284] + src29[285] + src29[286] + src29[287] + src29[288] + src29[289] + src29[290] + src29[291] + src29[292] + src29[293] + src29[294] + src29[295] + src29[296] + src29[297] + src29[298] + src29[299] + src29[300] + src29[301] + src29[302] + src29[303] + src29[304] + src29[305] + src29[306] + src29[307] + src29[308] + src29[309] + src29[310] + src29[311] + src29[312] + src29[313] + src29[314] + src29[315] + src29[316] + src29[317] + src29[318] + src29[319] + src29[320] + src29[321] + src29[322] + src29[323] + src29[324] + src29[325] + src29[326] + src29[327] + src29[328] + src29[329] + src29[330] + src29[331] + src29[332] + src29[333] + src29[334] + src29[335] + src29[336] + src29[337] + src29[338] + src29[339] + src29[340] + src29[341] + src29[342] + src29[343] + src29[344] + src29[345] + src29[346] + src29[347] + src29[348] + src29[349] + src29[350] + src29[351] + src29[352] + src29[353] + src29[354] + src29[355] + src29[356] + src29[357] + src29[358] + src29[359] + src29[360] + src29[361] + src29[362] + src29[363] + src29[364] + src29[365] + src29[366] + src29[367] + src29[368] + src29[369] + src29[370] + src29[371] + src29[372] + src29[373] + src29[374] + src29[375] + src29[376] + src29[377] + src29[378] + src29[379] + src29[380] + src29[381] + src29[382] + src29[383] + src29[384] + src29[385] + src29[386] + src29[387] + src29[388] + src29[389] + src29[390] + src29[391] + src29[392] + src29[393] + src29[394] + src29[395] + src29[396] + src29[397] + src29[398] + src29[399] + src29[400] + src29[401] + src29[402] + src29[403] + src29[404] + src29[405] + src29[406] + src29[407] + src29[408] + src29[409] + src29[410] + src29[411] + src29[412] + src29[413] + src29[414] + src29[415] + src29[416] + src29[417] + src29[418] + src29[419] + src29[420] + src29[421] + src29[422] + src29[423] + src29[424] + src29[425] + src29[426] + src29[427] + src29[428] + src29[429] + src29[430] + src29[431] + src29[432] + src29[433] + src29[434] + src29[435] + src29[436] + src29[437] + src29[438] + src29[439] + src29[440] + src29[441] + src29[442] + src29[443] + src29[444] + src29[445] + src29[446] + src29[447] + src29[448] + src29[449] + src29[450] + src29[451] + src29[452] + src29[453] + src29[454] + src29[455] + src29[456] + src29[457] + src29[458] + src29[459] + src29[460] + src29[461] + src29[462] + src29[463] + src29[464] + src29[465] + src29[466] + src29[467] + src29[468] + src29[469] + src29[470] + src29[471] + src29[472] + src29[473] + src29[474] + src29[475] + src29[476] + src29[477] + src29[478] + src29[479] + src29[480] + src29[481] + src29[482] + src29[483] + src29[484] + src29[485])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63] + src30[64] + src30[65] + src30[66] + src30[67] + src30[68] + src30[69] + src30[70] + src30[71] + src30[72] + src30[73] + src30[74] + src30[75] + src30[76] + src30[77] + src30[78] + src30[79] + src30[80] + src30[81] + src30[82] + src30[83] + src30[84] + src30[85] + src30[86] + src30[87] + src30[88] + src30[89] + src30[90] + src30[91] + src30[92] + src30[93] + src30[94] + src30[95] + src30[96] + src30[97] + src30[98] + src30[99] + src30[100] + src30[101] + src30[102] + src30[103] + src30[104] + src30[105] + src30[106] + src30[107] + src30[108] + src30[109] + src30[110] + src30[111] + src30[112] + src30[113] + src30[114] + src30[115] + src30[116] + src30[117] + src30[118] + src30[119] + src30[120] + src30[121] + src30[122] + src30[123] + src30[124] + src30[125] + src30[126] + src30[127] + src30[128] + src30[129] + src30[130] + src30[131] + src30[132] + src30[133] + src30[134] + src30[135] + src30[136] + src30[137] + src30[138] + src30[139] + src30[140] + src30[141] + src30[142] + src30[143] + src30[144] + src30[145] + src30[146] + src30[147] + src30[148] + src30[149] + src30[150] + src30[151] + src30[152] + src30[153] + src30[154] + src30[155] + src30[156] + src30[157] + src30[158] + src30[159] + src30[160] + src30[161] + src30[162] + src30[163] + src30[164] + src30[165] + src30[166] + src30[167] + src30[168] + src30[169] + src30[170] + src30[171] + src30[172] + src30[173] + src30[174] + src30[175] + src30[176] + src30[177] + src30[178] + src30[179] + src30[180] + src30[181] + src30[182] + src30[183] + src30[184] + src30[185] + src30[186] + src30[187] + src30[188] + src30[189] + src30[190] + src30[191] + src30[192] + src30[193] + src30[194] + src30[195] + src30[196] + src30[197] + src30[198] + src30[199] + src30[200] + src30[201] + src30[202] + src30[203] + src30[204] + src30[205] + src30[206] + src30[207] + src30[208] + src30[209] + src30[210] + src30[211] + src30[212] + src30[213] + src30[214] + src30[215] + src30[216] + src30[217] + src30[218] + src30[219] + src30[220] + src30[221] + src30[222] + src30[223] + src30[224] + src30[225] + src30[226] + src30[227] + src30[228] + src30[229] + src30[230] + src30[231] + src30[232] + src30[233] + src30[234] + src30[235] + src30[236] + src30[237] + src30[238] + src30[239] + src30[240] + src30[241] + src30[242] + src30[243] + src30[244] + src30[245] + src30[246] + src30[247] + src30[248] + src30[249] + src30[250] + src30[251] + src30[252] + src30[253] + src30[254] + src30[255] + src30[256] + src30[257] + src30[258] + src30[259] + src30[260] + src30[261] + src30[262] + src30[263] + src30[264] + src30[265] + src30[266] + src30[267] + src30[268] + src30[269] + src30[270] + src30[271] + src30[272] + src30[273] + src30[274] + src30[275] + src30[276] + src30[277] + src30[278] + src30[279] + src30[280] + src30[281] + src30[282] + src30[283] + src30[284] + src30[285] + src30[286] + src30[287] + src30[288] + src30[289] + src30[290] + src30[291] + src30[292] + src30[293] + src30[294] + src30[295] + src30[296] + src30[297] + src30[298] + src30[299] + src30[300] + src30[301] + src30[302] + src30[303] + src30[304] + src30[305] + src30[306] + src30[307] + src30[308] + src30[309] + src30[310] + src30[311] + src30[312] + src30[313] + src30[314] + src30[315] + src30[316] + src30[317] + src30[318] + src30[319] + src30[320] + src30[321] + src30[322] + src30[323] + src30[324] + src30[325] + src30[326] + src30[327] + src30[328] + src30[329] + src30[330] + src30[331] + src30[332] + src30[333] + src30[334] + src30[335] + src30[336] + src30[337] + src30[338] + src30[339] + src30[340] + src30[341] + src30[342] + src30[343] + src30[344] + src30[345] + src30[346] + src30[347] + src30[348] + src30[349] + src30[350] + src30[351] + src30[352] + src30[353] + src30[354] + src30[355] + src30[356] + src30[357] + src30[358] + src30[359] + src30[360] + src30[361] + src30[362] + src30[363] + src30[364] + src30[365] + src30[366] + src30[367] + src30[368] + src30[369] + src30[370] + src30[371] + src30[372] + src30[373] + src30[374] + src30[375] + src30[376] + src30[377] + src30[378] + src30[379] + src30[380] + src30[381] + src30[382] + src30[383] + src30[384] + src30[385] + src30[386] + src30[387] + src30[388] + src30[389] + src30[390] + src30[391] + src30[392] + src30[393] + src30[394] + src30[395] + src30[396] + src30[397] + src30[398] + src30[399] + src30[400] + src30[401] + src30[402] + src30[403] + src30[404] + src30[405] + src30[406] + src30[407] + src30[408] + src30[409] + src30[410] + src30[411] + src30[412] + src30[413] + src30[414] + src30[415] + src30[416] + src30[417] + src30[418] + src30[419] + src30[420] + src30[421] + src30[422] + src30[423] + src30[424] + src30[425] + src30[426] + src30[427] + src30[428] + src30[429] + src30[430] + src30[431] + src30[432] + src30[433] + src30[434] + src30[435] + src30[436] + src30[437] + src30[438] + src30[439] + src30[440] + src30[441] + src30[442] + src30[443] + src30[444] + src30[445] + src30[446] + src30[447] + src30[448] + src30[449] + src30[450] + src30[451] + src30[452] + src30[453] + src30[454] + src30[455] + src30[456] + src30[457] + src30[458] + src30[459] + src30[460] + src30[461] + src30[462] + src30[463] + src30[464] + src30[465] + src30[466] + src30[467] + src30[468] + src30[469] + src30[470] + src30[471] + src30[472] + src30[473] + src30[474] + src30[475] + src30[476] + src30[477] + src30[478] + src30[479] + src30[480] + src30[481] + src30[482] + src30[483] + src30[484] + src30[485])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63] + src31[64] + src31[65] + src31[66] + src31[67] + src31[68] + src31[69] + src31[70] + src31[71] + src31[72] + src31[73] + src31[74] + src31[75] + src31[76] + src31[77] + src31[78] + src31[79] + src31[80] + src31[81] + src31[82] + src31[83] + src31[84] + src31[85] + src31[86] + src31[87] + src31[88] + src31[89] + src31[90] + src31[91] + src31[92] + src31[93] + src31[94] + src31[95] + src31[96] + src31[97] + src31[98] + src31[99] + src31[100] + src31[101] + src31[102] + src31[103] + src31[104] + src31[105] + src31[106] + src31[107] + src31[108] + src31[109] + src31[110] + src31[111] + src31[112] + src31[113] + src31[114] + src31[115] + src31[116] + src31[117] + src31[118] + src31[119] + src31[120] + src31[121] + src31[122] + src31[123] + src31[124] + src31[125] + src31[126] + src31[127] + src31[128] + src31[129] + src31[130] + src31[131] + src31[132] + src31[133] + src31[134] + src31[135] + src31[136] + src31[137] + src31[138] + src31[139] + src31[140] + src31[141] + src31[142] + src31[143] + src31[144] + src31[145] + src31[146] + src31[147] + src31[148] + src31[149] + src31[150] + src31[151] + src31[152] + src31[153] + src31[154] + src31[155] + src31[156] + src31[157] + src31[158] + src31[159] + src31[160] + src31[161] + src31[162] + src31[163] + src31[164] + src31[165] + src31[166] + src31[167] + src31[168] + src31[169] + src31[170] + src31[171] + src31[172] + src31[173] + src31[174] + src31[175] + src31[176] + src31[177] + src31[178] + src31[179] + src31[180] + src31[181] + src31[182] + src31[183] + src31[184] + src31[185] + src31[186] + src31[187] + src31[188] + src31[189] + src31[190] + src31[191] + src31[192] + src31[193] + src31[194] + src31[195] + src31[196] + src31[197] + src31[198] + src31[199] + src31[200] + src31[201] + src31[202] + src31[203] + src31[204] + src31[205] + src31[206] + src31[207] + src31[208] + src31[209] + src31[210] + src31[211] + src31[212] + src31[213] + src31[214] + src31[215] + src31[216] + src31[217] + src31[218] + src31[219] + src31[220] + src31[221] + src31[222] + src31[223] + src31[224] + src31[225] + src31[226] + src31[227] + src31[228] + src31[229] + src31[230] + src31[231] + src31[232] + src31[233] + src31[234] + src31[235] + src31[236] + src31[237] + src31[238] + src31[239] + src31[240] + src31[241] + src31[242] + src31[243] + src31[244] + src31[245] + src31[246] + src31[247] + src31[248] + src31[249] + src31[250] + src31[251] + src31[252] + src31[253] + src31[254] + src31[255] + src31[256] + src31[257] + src31[258] + src31[259] + src31[260] + src31[261] + src31[262] + src31[263] + src31[264] + src31[265] + src31[266] + src31[267] + src31[268] + src31[269] + src31[270] + src31[271] + src31[272] + src31[273] + src31[274] + src31[275] + src31[276] + src31[277] + src31[278] + src31[279] + src31[280] + src31[281] + src31[282] + src31[283] + src31[284] + src31[285] + src31[286] + src31[287] + src31[288] + src31[289] + src31[290] + src31[291] + src31[292] + src31[293] + src31[294] + src31[295] + src31[296] + src31[297] + src31[298] + src31[299] + src31[300] + src31[301] + src31[302] + src31[303] + src31[304] + src31[305] + src31[306] + src31[307] + src31[308] + src31[309] + src31[310] + src31[311] + src31[312] + src31[313] + src31[314] + src31[315] + src31[316] + src31[317] + src31[318] + src31[319] + src31[320] + src31[321] + src31[322] + src31[323] + src31[324] + src31[325] + src31[326] + src31[327] + src31[328] + src31[329] + src31[330] + src31[331] + src31[332] + src31[333] + src31[334] + src31[335] + src31[336] + src31[337] + src31[338] + src31[339] + src31[340] + src31[341] + src31[342] + src31[343] + src31[344] + src31[345] + src31[346] + src31[347] + src31[348] + src31[349] + src31[350] + src31[351] + src31[352] + src31[353] + src31[354] + src31[355] + src31[356] + src31[357] + src31[358] + src31[359] + src31[360] + src31[361] + src31[362] + src31[363] + src31[364] + src31[365] + src31[366] + src31[367] + src31[368] + src31[369] + src31[370] + src31[371] + src31[372] + src31[373] + src31[374] + src31[375] + src31[376] + src31[377] + src31[378] + src31[379] + src31[380] + src31[381] + src31[382] + src31[383] + src31[384] + src31[385] + src31[386] + src31[387] + src31[388] + src31[389] + src31[390] + src31[391] + src31[392] + src31[393] + src31[394] + src31[395] + src31[396] + src31[397] + src31[398] + src31[399] + src31[400] + src31[401] + src31[402] + src31[403] + src31[404] + src31[405] + src31[406] + src31[407] + src31[408] + src31[409] + src31[410] + src31[411] + src31[412] + src31[413] + src31[414] + src31[415] + src31[416] + src31[417] + src31[418] + src31[419] + src31[420] + src31[421] + src31[422] + src31[423] + src31[424] + src31[425] + src31[426] + src31[427] + src31[428] + src31[429] + src31[430] + src31[431] + src31[432] + src31[433] + src31[434] + src31[435] + src31[436] + src31[437] + src31[438] + src31[439] + src31[440] + src31[441] + src31[442] + src31[443] + src31[444] + src31[445] + src31[446] + src31[447] + src31[448] + src31[449] + src31[450] + src31[451] + src31[452] + src31[453] + src31[454] + src31[455] + src31[456] + src31[457] + src31[458] + src31[459] + src31[460] + src31[461] + src31[462] + src31[463] + src31[464] + src31[465] + src31[466] + src31[467] + src31[468] + src31[469] + src31[470] + src31[471] + src31[472] + src31[473] + src31[474] + src31[475] + src31[476] + src31[477] + src31[478] + src31[479] + src31[480] + src31[481] + src31[482] + src31[483] + src31[484] + src31[485])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28] + src32[29] + src32[30] + src32[31] + src32[32] + src32[33] + src32[34] + src32[35] + src32[36] + src32[37] + src32[38] + src32[39] + src32[40] + src32[41] + src32[42] + src32[43] + src32[44] + src32[45] + src32[46] + src32[47] + src32[48] + src32[49] + src32[50] + src32[51] + src32[52] + src32[53] + src32[54] + src32[55] + src32[56] + src32[57] + src32[58] + src32[59] + src32[60] + src32[61] + src32[62] + src32[63] + src32[64] + src32[65] + src32[66] + src32[67] + src32[68] + src32[69] + src32[70] + src32[71] + src32[72] + src32[73] + src32[74] + src32[75] + src32[76] + src32[77] + src32[78] + src32[79] + src32[80] + src32[81] + src32[82] + src32[83] + src32[84] + src32[85] + src32[86] + src32[87] + src32[88] + src32[89] + src32[90] + src32[91] + src32[92] + src32[93] + src32[94] + src32[95] + src32[96] + src32[97] + src32[98] + src32[99] + src32[100] + src32[101] + src32[102] + src32[103] + src32[104] + src32[105] + src32[106] + src32[107] + src32[108] + src32[109] + src32[110] + src32[111] + src32[112] + src32[113] + src32[114] + src32[115] + src32[116] + src32[117] + src32[118] + src32[119] + src32[120] + src32[121] + src32[122] + src32[123] + src32[124] + src32[125] + src32[126] + src32[127] + src32[128] + src32[129] + src32[130] + src32[131] + src32[132] + src32[133] + src32[134] + src32[135] + src32[136] + src32[137] + src32[138] + src32[139] + src32[140] + src32[141] + src32[142] + src32[143] + src32[144] + src32[145] + src32[146] + src32[147] + src32[148] + src32[149] + src32[150] + src32[151] + src32[152] + src32[153] + src32[154] + src32[155] + src32[156] + src32[157] + src32[158] + src32[159] + src32[160] + src32[161] + src32[162] + src32[163] + src32[164] + src32[165] + src32[166] + src32[167] + src32[168] + src32[169] + src32[170] + src32[171] + src32[172] + src32[173] + src32[174] + src32[175] + src32[176] + src32[177] + src32[178] + src32[179] + src32[180] + src32[181] + src32[182] + src32[183] + src32[184] + src32[185] + src32[186] + src32[187] + src32[188] + src32[189] + src32[190] + src32[191] + src32[192] + src32[193] + src32[194] + src32[195] + src32[196] + src32[197] + src32[198] + src32[199] + src32[200] + src32[201] + src32[202] + src32[203] + src32[204] + src32[205] + src32[206] + src32[207] + src32[208] + src32[209] + src32[210] + src32[211] + src32[212] + src32[213] + src32[214] + src32[215] + src32[216] + src32[217] + src32[218] + src32[219] + src32[220] + src32[221] + src32[222] + src32[223] + src32[224] + src32[225] + src32[226] + src32[227] + src32[228] + src32[229] + src32[230] + src32[231] + src32[232] + src32[233] + src32[234] + src32[235] + src32[236] + src32[237] + src32[238] + src32[239] + src32[240] + src32[241] + src32[242] + src32[243] + src32[244] + src32[245] + src32[246] + src32[247] + src32[248] + src32[249] + src32[250] + src32[251] + src32[252] + src32[253] + src32[254] + src32[255] + src32[256] + src32[257] + src32[258] + src32[259] + src32[260] + src32[261] + src32[262] + src32[263] + src32[264] + src32[265] + src32[266] + src32[267] + src32[268] + src32[269] + src32[270] + src32[271] + src32[272] + src32[273] + src32[274] + src32[275] + src32[276] + src32[277] + src32[278] + src32[279] + src32[280] + src32[281] + src32[282] + src32[283] + src32[284] + src32[285] + src32[286] + src32[287] + src32[288] + src32[289] + src32[290] + src32[291] + src32[292] + src32[293] + src32[294] + src32[295] + src32[296] + src32[297] + src32[298] + src32[299] + src32[300] + src32[301] + src32[302] + src32[303] + src32[304] + src32[305] + src32[306] + src32[307] + src32[308] + src32[309] + src32[310] + src32[311] + src32[312] + src32[313] + src32[314] + src32[315] + src32[316] + src32[317] + src32[318] + src32[319] + src32[320] + src32[321] + src32[322] + src32[323] + src32[324] + src32[325] + src32[326] + src32[327] + src32[328] + src32[329] + src32[330] + src32[331] + src32[332] + src32[333] + src32[334] + src32[335] + src32[336] + src32[337] + src32[338] + src32[339] + src32[340] + src32[341] + src32[342] + src32[343] + src32[344] + src32[345] + src32[346] + src32[347] + src32[348] + src32[349] + src32[350] + src32[351] + src32[352] + src32[353] + src32[354] + src32[355] + src32[356] + src32[357] + src32[358] + src32[359] + src32[360] + src32[361] + src32[362] + src32[363] + src32[364] + src32[365] + src32[366] + src32[367] + src32[368] + src32[369] + src32[370] + src32[371] + src32[372] + src32[373] + src32[374] + src32[375] + src32[376] + src32[377] + src32[378] + src32[379] + src32[380] + src32[381] + src32[382] + src32[383] + src32[384] + src32[385] + src32[386] + src32[387] + src32[388] + src32[389] + src32[390] + src32[391] + src32[392] + src32[393] + src32[394] + src32[395] + src32[396] + src32[397] + src32[398] + src32[399] + src32[400] + src32[401] + src32[402] + src32[403] + src32[404] + src32[405] + src32[406] + src32[407] + src32[408] + src32[409] + src32[410] + src32[411] + src32[412] + src32[413] + src32[414] + src32[415] + src32[416] + src32[417] + src32[418] + src32[419] + src32[420] + src32[421] + src32[422] + src32[423] + src32[424] + src32[425] + src32[426] + src32[427] + src32[428] + src32[429] + src32[430] + src32[431] + src32[432] + src32[433] + src32[434] + src32[435] + src32[436] + src32[437] + src32[438] + src32[439] + src32[440] + src32[441] + src32[442] + src32[443] + src32[444] + src32[445] + src32[446] + src32[447] + src32[448] + src32[449] + src32[450] + src32[451] + src32[452] + src32[453] + src32[454] + src32[455] + src32[456] + src32[457] + src32[458] + src32[459] + src32[460] + src32[461] + src32[462] + src32[463] + src32[464] + src32[465] + src32[466] + src32[467] + src32[468] + src32[469] + src32[470] + src32[471] + src32[472] + src32[473] + src32[474] + src32[475] + src32[476] + src32[477] + src32[478] + src32[479] + src32[480] + src32[481] + src32[482] + src32[483] + src32[484] + src32[485])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27] + src33[28] + src33[29] + src33[30] + src33[31] + src33[32] + src33[33] + src33[34] + src33[35] + src33[36] + src33[37] + src33[38] + src33[39] + src33[40] + src33[41] + src33[42] + src33[43] + src33[44] + src33[45] + src33[46] + src33[47] + src33[48] + src33[49] + src33[50] + src33[51] + src33[52] + src33[53] + src33[54] + src33[55] + src33[56] + src33[57] + src33[58] + src33[59] + src33[60] + src33[61] + src33[62] + src33[63] + src33[64] + src33[65] + src33[66] + src33[67] + src33[68] + src33[69] + src33[70] + src33[71] + src33[72] + src33[73] + src33[74] + src33[75] + src33[76] + src33[77] + src33[78] + src33[79] + src33[80] + src33[81] + src33[82] + src33[83] + src33[84] + src33[85] + src33[86] + src33[87] + src33[88] + src33[89] + src33[90] + src33[91] + src33[92] + src33[93] + src33[94] + src33[95] + src33[96] + src33[97] + src33[98] + src33[99] + src33[100] + src33[101] + src33[102] + src33[103] + src33[104] + src33[105] + src33[106] + src33[107] + src33[108] + src33[109] + src33[110] + src33[111] + src33[112] + src33[113] + src33[114] + src33[115] + src33[116] + src33[117] + src33[118] + src33[119] + src33[120] + src33[121] + src33[122] + src33[123] + src33[124] + src33[125] + src33[126] + src33[127] + src33[128] + src33[129] + src33[130] + src33[131] + src33[132] + src33[133] + src33[134] + src33[135] + src33[136] + src33[137] + src33[138] + src33[139] + src33[140] + src33[141] + src33[142] + src33[143] + src33[144] + src33[145] + src33[146] + src33[147] + src33[148] + src33[149] + src33[150] + src33[151] + src33[152] + src33[153] + src33[154] + src33[155] + src33[156] + src33[157] + src33[158] + src33[159] + src33[160] + src33[161] + src33[162] + src33[163] + src33[164] + src33[165] + src33[166] + src33[167] + src33[168] + src33[169] + src33[170] + src33[171] + src33[172] + src33[173] + src33[174] + src33[175] + src33[176] + src33[177] + src33[178] + src33[179] + src33[180] + src33[181] + src33[182] + src33[183] + src33[184] + src33[185] + src33[186] + src33[187] + src33[188] + src33[189] + src33[190] + src33[191] + src33[192] + src33[193] + src33[194] + src33[195] + src33[196] + src33[197] + src33[198] + src33[199] + src33[200] + src33[201] + src33[202] + src33[203] + src33[204] + src33[205] + src33[206] + src33[207] + src33[208] + src33[209] + src33[210] + src33[211] + src33[212] + src33[213] + src33[214] + src33[215] + src33[216] + src33[217] + src33[218] + src33[219] + src33[220] + src33[221] + src33[222] + src33[223] + src33[224] + src33[225] + src33[226] + src33[227] + src33[228] + src33[229] + src33[230] + src33[231] + src33[232] + src33[233] + src33[234] + src33[235] + src33[236] + src33[237] + src33[238] + src33[239] + src33[240] + src33[241] + src33[242] + src33[243] + src33[244] + src33[245] + src33[246] + src33[247] + src33[248] + src33[249] + src33[250] + src33[251] + src33[252] + src33[253] + src33[254] + src33[255] + src33[256] + src33[257] + src33[258] + src33[259] + src33[260] + src33[261] + src33[262] + src33[263] + src33[264] + src33[265] + src33[266] + src33[267] + src33[268] + src33[269] + src33[270] + src33[271] + src33[272] + src33[273] + src33[274] + src33[275] + src33[276] + src33[277] + src33[278] + src33[279] + src33[280] + src33[281] + src33[282] + src33[283] + src33[284] + src33[285] + src33[286] + src33[287] + src33[288] + src33[289] + src33[290] + src33[291] + src33[292] + src33[293] + src33[294] + src33[295] + src33[296] + src33[297] + src33[298] + src33[299] + src33[300] + src33[301] + src33[302] + src33[303] + src33[304] + src33[305] + src33[306] + src33[307] + src33[308] + src33[309] + src33[310] + src33[311] + src33[312] + src33[313] + src33[314] + src33[315] + src33[316] + src33[317] + src33[318] + src33[319] + src33[320] + src33[321] + src33[322] + src33[323] + src33[324] + src33[325] + src33[326] + src33[327] + src33[328] + src33[329] + src33[330] + src33[331] + src33[332] + src33[333] + src33[334] + src33[335] + src33[336] + src33[337] + src33[338] + src33[339] + src33[340] + src33[341] + src33[342] + src33[343] + src33[344] + src33[345] + src33[346] + src33[347] + src33[348] + src33[349] + src33[350] + src33[351] + src33[352] + src33[353] + src33[354] + src33[355] + src33[356] + src33[357] + src33[358] + src33[359] + src33[360] + src33[361] + src33[362] + src33[363] + src33[364] + src33[365] + src33[366] + src33[367] + src33[368] + src33[369] + src33[370] + src33[371] + src33[372] + src33[373] + src33[374] + src33[375] + src33[376] + src33[377] + src33[378] + src33[379] + src33[380] + src33[381] + src33[382] + src33[383] + src33[384] + src33[385] + src33[386] + src33[387] + src33[388] + src33[389] + src33[390] + src33[391] + src33[392] + src33[393] + src33[394] + src33[395] + src33[396] + src33[397] + src33[398] + src33[399] + src33[400] + src33[401] + src33[402] + src33[403] + src33[404] + src33[405] + src33[406] + src33[407] + src33[408] + src33[409] + src33[410] + src33[411] + src33[412] + src33[413] + src33[414] + src33[415] + src33[416] + src33[417] + src33[418] + src33[419] + src33[420] + src33[421] + src33[422] + src33[423] + src33[424] + src33[425] + src33[426] + src33[427] + src33[428] + src33[429] + src33[430] + src33[431] + src33[432] + src33[433] + src33[434] + src33[435] + src33[436] + src33[437] + src33[438] + src33[439] + src33[440] + src33[441] + src33[442] + src33[443] + src33[444] + src33[445] + src33[446] + src33[447] + src33[448] + src33[449] + src33[450] + src33[451] + src33[452] + src33[453] + src33[454] + src33[455] + src33[456] + src33[457] + src33[458] + src33[459] + src33[460] + src33[461] + src33[462] + src33[463] + src33[464] + src33[465] + src33[466] + src33[467] + src33[468] + src33[469] + src33[470] + src33[471] + src33[472] + src33[473] + src33[474] + src33[475] + src33[476] + src33[477] + src33[478] + src33[479] + src33[480] + src33[481] + src33[482] + src33[483] + src33[484] + src33[485])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26] + src34[27] + src34[28] + src34[29] + src34[30] + src34[31] + src34[32] + src34[33] + src34[34] + src34[35] + src34[36] + src34[37] + src34[38] + src34[39] + src34[40] + src34[41] + src34[42] + src34[43] + src34[44] + src34[45] + src34[46] + src34[47] + src34[48] + src34[49] + src34[50] + src34[51] + src34[52] + src34[53] + src34[54] + src34[55] + src34[56] + src34[57] + src34[58] + src34[59] + src34[60] + src34[61] + src34[62] + src34[63] + src34[64] + src34[65] + src34[66] + src34[67] + src34[68] + src34[69] + src34[70] + src34[71] + src34[72] + src34[73] + src34[74] + src34[75] + src34[76] + src34[77] + src34[78] + src34[79] + src34[80] + src34[81] + src34[82] + src34[83] + src34[84] + src34[85] + src34[86] + src34[87] + src34[88] + src34[89] + src34[90] + src34[91] + src34[92] + src34[93] + src34[94] + src34[95] + src34[96] + src34[97] + src34[98] + src34[99] + src34[100] + src34[101] + src34[102] + src34[103] + src34[104] + src34[105] + src34[106] + src34[107] + src34[108] + src34[109] + src34[110] + src34[111] + src34[112] + src34[113] + src34[114] + src34[115] + src34[116] + src34[117] + src34[118] + src34[119] + src34[120] + src34[121] + src34[122] + src34[123] + src34[124] + src34[125] + src34[126] + src34[127] + src34[128] + src34[129] + src34[130] + src34[131] + src34[132] + src34[133] + src34[134] + src34[135] + src34[136] + src34[137] + src34[138] + src34[139] + src34[140] + src34[141] + src34[142] + src34[143] + src34[144] + src34[145] + src34[146] + src34[147] + src34[148] + src34[149] + src34[150] + src34[151] + src34[152] + src34[153] + src34[154] + src34[155] + src34[156] + src34[157] + src34[158] + src34[159] + src34[160] + src34[161] + src34[162] + src34[163] + src34[164] + src34[165] + src34[166] + src34[167] + src34[168] + src34[169] + src34[170] + src34[171] + src34[172] + src34[173] + src34[174] + src34[175] + src34[176] + src34[177] + src34[178] + src34[179] + src34[180] + src34[181] + src34[182] + src34[183] + src34[184] + src34[185] + src34[186] + src34[187] + src34[188] + src34[189] + src34[190] + src34[191] + src34[192] + src34[193] + src34[194] + src34[195] + src34[196] + src34[197] + src34[198] + src34[199] + src34[200] + src34[201] + src34[202] + src34[203] + src34[204] + src34[205] + src34[206] + src34[207] + src34[208] + src34[209] + src34[210] + src34[211] + src34[212] + src34[213] + src34[214] + src34[215] + src34[216] + src34[217] + src34[218] + src34[219] + src34[220] + src34[221] + src34[222] + src34[223] + src34[224] + src34[225] + src34[226] + src34[227] + src34[228] + src34[229] + src34[230] + src34[231] + src34[232] + src34[233] + src34[234] + src34[235] + src34[236] + src34[237] + src34[238] + src34[239] + src34[240] + src34[241] + src34[242] + src34[243] + src34[244] + src34[245] + src34[246] + src34[247] + src34[248] + src34[249] + src34[250] + src34[251] + src34[252] + src34[253] + src34[254] + src34[255] + src34[256] + src34[257] + src34[258] + src34[259] + src34[260] + src34[261] + src34[262] + src34[263] + src34[264] + src34[265] + src34[266] + src34[267] + src34[268] + src34[269] + src34[270] + src34[271] + src34[272] + src34[273] + src34[274] + src34[275] + src34[276] + src34[277] + src34[278] + src34[279] + src34[280] + src34[281] + src34[282] + src34[283] + src34[284] + src34[285] + src34[286] + src34[287] + src34[288] + src34[289] + src34[290] + src34[291] + src34[292] + src34[293] + src34[294] + src34[295] + src34[296] + src34[297] + src34[298] + src34[299] + src34[300] + src34[301] + src34[302] + src34[303] + src34[304] + src34[305] + src34[306] + src34[307] + src34[308] + src34[309] + src34[310] + src34[311] + src34[312] + src34[313] + src34[314] + src34[315] + src34[316] + src34[317] + src34[318] + src34[319] + src34[320] + src34[321] + src34[322] + src34[323] + src34[324] + src34[325] + src34[326] + src34[327] + src34[328] + src34[329] + src34[330] + src34[331] + src34[332] + src34[333] + src34[334] + src34[335] + src34[336] + src34[337] + src34[338] + src34[339] + src34[340] + src34[341] + src34[342] + src34[343] + src34[344] + src34[345] + src34[346] + src34[347] + src34[348] + src34[349] + src34[350] + src34[351] + src34[352] + src34[353] + src34[354] + src34[355] + src34[356] + src34[357] + src34[358] + src34[359] + src34[360] + src34[361] + src34[362] + src34[363] + src34[364] + src34[365] + src34[366] + src34[367] + src34[368] + src34[369] + src34[370] + src34[371] + src34[372] + src34[373] + src34[374] + src34[375] + src34[376] + src34[377] + src34[378] + src34[379] + src34[380] + src34[381] + src34[382] + src34[383] + src34[384] + src34[385] + src34[386] + src34[387] + src34[388] + src34[389] + src34[390] + src34[391] + src34[392] + src34[393] + src34[394] + src34[395] + src34[396] + src34[397] + src34[398] + src34[399] + src34[400] + src34[401] + src34[402] + src34[403] + src34[404] + src34[405] + src34[406] + src34[407] + src34[408] + src34[409] + src34[410] + src34[411] + src34[412] + src34[413] + src34[414] + src34[415] + src34[416] + src34[417] + src34[418] + src34[419] + src34[420] + src34[421] + src34[422] + src34[423] + src34[424] + src34[425] + src34[426] + src34[427] + src34[428] + src34[429] + src34[430] + src34[431] + src34[432] + src34[433] + src34[434] + src34[435] + src34[436] + src34[437] + src34[438] + src34[439] + src34[440] + src34[441] + src34[442] + src34[443] + src34[444] + src34[445] + src34[446] + src34[447] + src34[448] + src34[449] + src34[450] + src34[451] + src34[452] + src34[453] + src34[454] + src34[455] + src34[456] + src34[457] + src34[458] + src34[459] + src34[460] + src34[461] + src34[462] + src34[463] + src34[464] + src34[465] + src34[466] + src34[467] + src34[468] + src34[469] + src34[470] + src34[471] + src34[472] + src34[473] + src34[474] + src34[475] + src34[476] + src34[477] + src34[478] + src34[479] + src34[480] + src34[481] + src34[482] + src34[483] + src34[484] + src34[485])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25] + src35[26] + src35[27] + src35[28] + src35[29] + src35[30] + src35[31] + src35[32] + src35[33] + src35[34] + src35[35] + src35[36] + src35[37] + src35[38] + src35[39] + src35[40] + src35[41] + src35[42] + src35[43] + src35[44] + src35[45] + src35[46] + src35[47] + src35[48] + src35[49] + src35[50] + src35[51] + src35[52] + src35[53] + src35[54] + src35[55] + src35[56] + src35[57] + src35[58] + src35[59] + src35[60] + src35[61] + src35[62] + src35[63] + src35[64] + src35[65] + src35[66] + src35[67] + src35[68] + src35[69] + src35[70] + src35[71] + src35[72] + src35[73] + src35[74] + src35[75] + src35[76] + src35[77] + src35[78] + src35[79] + src35[80] + src35[81] + src35[82] + src35[83] + src35[84] + src35[85] + src35[86] + src35[87] + src35[88] + src35[89] + src35[90] + src35[91] + src35[92] + src35[93] + src35[94] + src35[95] + src35[96] + src35[97] + src35[98] + src35[99] + src35[100] + src35[101] + src35[102] + src35[103] + src35[104] + src35[105] + src35[106] + src35[107] + src35[108] + src35[109] + src35[110] + src35[111] + src35[112] + src35[113] + src35[114] + src35[115] + src35[116] + src35[117] + src35[118] + src35[119] + src35[120] + src35[121] + src35[122] + src35[123] + src35[124] + src35[125] + src35[126] + src35[127] + src35[128] + src35[129] + src35[130] + src35[131] + src35[132] + src35[133] + src35[134] + src35[135] + src35[136] + src35[137] + src35[138] + src35[139] + src35[140] + src35[141] + src35[142] + src35[143] + src35[144] + src35[145] + src35[146] + src35[147] + src35[148] + src35[149] + src35[150] + src35[151] + src35[152] + src35[153] + src35[154] + src35[155] + src35[156] + src35[157] + src35[158] + src35[159] + src35[160] + src35[161] + src35[162] + src35[163] + src35[164] + src35[165] + src35[166] + src35[167] + src35[168] + src35[169] + src35[170] + src35[171] + src35[172] + src35[173] + src35[174] + src35[175] + src35[176] + src35[177] + src35[178] + src35[179] + src35[180] + src35[181] + src35[182] + src35[183] + src35[184] + src35[185] + src35[186] + src35[187] + src35[188] + src35[189] + src35[190] + src35[191] + src35[192] + src35[193] + src35[194] + src35[195] + src35[196] + src35[197] + src35[198] + src35[199] + src35[200] + src35[201] + src35[202] + src35[203] + src35[204] + src35[205] + src35[206] + src35[207] + src35[208] + src35[209] + src35[210] + src35[211] + src35[212] + src35[213] + src35[214] + src35[215] + src35[216] + src35[217] + src35[218] + src35[219] + src35[220] + src35[221] + src35[222] + src35[223] + src35[224] + src35[225] + src35[226] + src35[227] + src35[228] + src35[229] + src35[230] + src35[231] + src35[232] + src35[233] + src35[234] + src35[235] + src35[236] + src35[237] + src35[238] + src35[239] + src35[240] + src35[241] + src35[242] + src35[243] + src35[244] + src35[245] + src35[246] + src35[247] + src35[248] + src35[249] + src35[250] + src35[251] + src35[252] + src35[253] + src35[254] + src35[255] + src35[256] + src35[257] + src35[258] + src35[259] + src35[260] + src35[261] + src35[262] + src35[263] + src35[264] + src35[265] + src35[266] + src35[267] + src35[268] + src35[269] + src35[270] + src35[271] + src35[272] + src35[273] + src35[274] + src35[275] + src35[276] + src35[277] + src35[278] + src35[279] + src35[280] + src35[281] + src35[282] + src35[283] + src35[284] + src35[285] + src35[286] + src35[287] + src35[288] + src35[289] + src35[290] + src35[291] + src35[292] + src35[293] + src35[294] + src35[295] + src35[296] + src35[297] + src35[298] + src35[299] + src35[300] + src35[301] + src35[302] + src35[303] + src35[304] + src35[305] + src35[306] + src35[307] + src35[308] + src35[309] + src35[310] + src35[311] + src35[312] + src35[313] + src35[314] + src35[315] + src35[316] + src35[317] + src35[318] + src35[319] + src35[320] + src35[321] + src35[322] + src35[323] + src35[324] + src35[325] + src35[326] + src35[327] + src35[328] + src35[329] + src35[330] + src35[331] + src35[332] + src35[333] + src35[334] + src35[335] + src35[336] + src35[337] + src35[338] + src35[339] + src35[340] + src35[341] + src35[342] + src35[343] + src35[344] + src35[345] + src35[346] + src35[347] + src35[348] + src35[349] + src35[350] + src35[351] + src35[352] + src35[353] + src35[354] + src35[355] + src35[356] + src35[357] + src35[358] + src35[359] + src35[360] + src35[361] + src35[362] + src35[363] + src35[364] + src35[365] + src35[366] + src35[367] + src35[368] + src35[369] + src35[370] + src35[371] + src35[372] + src35[373] + src35[374] + src35[375] + src35[376] + src35[377] + src35[378] + src35[379] + src35[380] + src35[381] + src35[382] + src35[383] + src35[384] + src35[385] + src35[386] + src35[387] + src35[388] + src35[389] + src35[390] + src35[391] + src35[392] + src35[393] + src35[394] + src35[395] + src35[396] + src35[397] + src35[398] + src35[399] + src35[400] + src35[401] + src35[402] + src35[403] + src35[404] + src35[405] + src35[406] + src35[407] + src35[408] + src35[409] + src35[410] + src35[411] + src35[412] + src35[413] + src35[414] + src35[415] + src35[416] + src35[417] + src35[418] + src35[419] + src35[420] + src35[421] + src35[422] + src35[423] + src35[424] + src35[425] + src35[426] + src35[427] + src35[428] + src35[429] + src35[430] + src35[431] + src35[432] + src35[433] + src35[434] + src35[435] + src35[436] + src35[437] + src35[438] + src35[439] + src35[440] + src35[441] + src35[442] + src35[443] + src35[444] + src35[445] + src35[446] + src35[447] + src35[448] + src35[449] + src35[450] + src35[451] + src35[452] + src35[453] + src35[454] + src35[455] + src35[456] + src35[457] + src35[458] + src35[459] + src35[460] + src35[461] + src35[462] + src35[463] + src35[464] + src35[465] + src35[466] + src35[467] + src35[468] + src35[469] + src35[470] + src35[471] + src35[472] + src35[473] + src35[474] + src35[475] + src35[476] + src35[477] + src35[478] + src35[479] + src35[480] + src35[481] + src35[482] + src35[483] + src35[484] + src35[485])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24] + src36[25] + src36[26] + src36[27] + src36[28] + src36[29] + src36[30] + src36[31] + src36[32] + src36[33] + src36[34] + src36[35] + src36[36] + src36[37] + src36[38] + src36[39] + src36[40] + src36[41] + src36[42] + src36[43] + src36[44] + src36[45] + src36[46] + src36[47] + src36[48] + src36[49] + src36[50] + src36[51] + src36[52] + src36[53] + src36[54] + src36[55] + src36[56] + src36[57] + src36[58] + src36[59] + src36[60] + src36[61] + src36[62] + src36[63] + src36[64] + src36[65] + src36[66] + src36[67] + src36[68] + src36[69] + src36[70] + src36[71] + src36[72] + src36[73] + src36[74] + src36[75] + src36[76] + src36[77] + src36[78] + src36[79] + src36[80] + src36[81] + src36[82] + src36[83] + src36[84] + src36[85] + src36[86] + src36[87] + src36[88] + src36[89] + src36[90] + src36[91] + src36[92] + src36[93] + src36[94] + src36[95] + src36[96] + src36[97] + src36[98] + src36[99] + src36[100] + src36[101] + src36[102] + src36[103] + src36[104] + src36[105] + src36[106] + src36[107] + src36[108] + src36[109] + src36[110] + src36[111] + src36[112] + src36[113] + src36[114] + src36[115] + src36[116] + src36[117] + src36[118] + src36[119] + src36[120] + src36[121] + src36[122] + src36[123] + src36[124] + src36[125] + src36[126] + src36[127] + src36[128] + src36[129] + src36[130] + src36[131] + src36[132] + src36[133] + src36[134] + src36[135] + src36[136] + src36[137] + src36[138] + src36[139] + src36[140] + src36[141] + src36[142] + src36[143] + src36[144] + src36[145] + src36[146] + src36[147] + src36[148] + src36[149] + src36[150] + src36[151] + src36[152] + src36[153] + src36[154] + src36[155] + src36[156] + src36[157] + src36[158] + src36[159] + src36[160] + src36[161] + src36[162] + src36[163] + src36[164] + src36[165] + src36[166] + src36[167] + src36[168] + src36[169] + src36[170] + src36[171] + src36[172] + src36[173] + src36[174] + src36[175] + src36[176] + src36[177] + src36[178] + src36[179] + src36[180] + src36[181] + src36[182] + src36[183] + src36[184] + src36[185] + src36[186] + src36[187] + src36[188] + src36[189] + src36[190] + src36[191] + src36[192] + src36[193] + src36[194] + src36[195] + src36[196] + src36[197] + src36[198] + src36[199] + src36[200] + src36[201] + src36[202] + src36[203] + src36[204] + src36[205] + src36[206] + src36[207] + src36[208] + src36[209] + src36[210] + src36[211] + src36[212] + src36[213] + src36[214] + src36[215] + src36[216] + src36[217] + src36[218] + src36[219] + src36[220] + src36[221] + src36[222] + src36[223] + src36[224] + src36[225] + src36[226] + src36[227] + src36[228] + src36[229] + src36[230] + src36[231] + src36[232] + src36[233] + src36[234] + src36[235] + src36[236] + src36[237] + src36[238] + src36[239] + src36[240] + src36[241] + src36[242] + src36[243] + src36[244] + src36[245] + src36[246] + src36[247] + src36[248] + src36[249] + src36[250] + src36[251] + src36[252] + src36[253] + src36[254] + src36[255] + src36[256] + src36[257] + src36[258] + src36[259] + src36[260] + src36[261] + src36[262] + src36[263] + src36[264] + src36[265] + src36[266] + src36[267] + src36[268] + src36[269] + src36[270] + src36[271] + src36[272] + src36[273] + src36[274] + src36[275] + src36[276] + src36[277] + src36[278] + src36[279] + src36[280] + src36[281] + src36[282] + src36[283] + src36[284] + src36[285] + src36[286] + src36[287] + src36[288] + src36[289] + src36[290] + src36[291] + src36[292] + src36[293] + src36[294] + src36[295] + src36[296] + src36[297] + src36[298] + src36[299] + src36[300] + src36[301] + src36[302] + src36[303] + src36[304] + src36[305] + src36[306] + src36[307] + src36[308] + src36[309] + src36[310] + src36[311] + src36[312] + src36[313] + src36[314] + src36[315] + src36[316] + src36[317] + src36[318] + src36[319] + src36[320] + src36[321] + src36[322] + src36[323] + src36[324] + src36[325] + src36[326] + src36[327] + src36[328] + src36[329] + src36[330] + src36[331] + src36[332] + src36[333] + src36[334] + src36[335] + src36[336] + src36[337] + src36[338] + src36[339] + src36[340] + src36[341] + src36[342] + src36[343] + src36[344] + src36[345] + src36[346] + src36[347] + src36[348] + src36[349] + src36[350] + src36[351] + src36[352] + src36[353] + src36[354] + src36[355] + src36[356] + src36[357] + src36[358] + src36[359] + src36[360] + src36[361] + src36[362] + src36[363] + src36[364] + src36[365] + src36[366] + src36[367] + src36[368] + src36[369] + src36[370] + src36[371] + src36[372] + src36[373] + src36[374] + src36[375] + src36[376] + src36[377] + src36[378] + src36[379] + src36[380] + src36[381] + src36[382] + src36[383] + src36[384] + src36[385] + src36[386] + src36[387] + src36[388] + src36[389] + src36[390] + src36[391] + src36[392] + src36[393] + src36[394] + src36[395] + src36[396] + src36[397] + src36[398] + src36[399] + src36[400] + src36[401] + src36[402] + src36[403] + src36[404] + src36[405] + src36[406] + src36[407] + src36[408] + src36[409] + src36[410] + src36[411] + src36[412] + src36[413] + src36[414] + src36[415] + src36[416] + src36[417] + src36[418] + src36[419] + src36[420] + src36[421] + src36[422] + src36[423] + src36[424] + src36[425] + src36[426] + src36[427] + src36[428] + src36[429] + src36[430] + src36[431] + src36[432] + src36[433] + src36[434] + src36[435] + src36[436] + src36[437] + src36[438] + src36[439] + src36[440] + src36[441] + src36[442] + src36[443] + src36[444] + src36[445] + src36[446] + src36[447] + src36[448] + src36[449] + src36[450] + src36[451] + src36[452] + src36[453] + src36[454] + src36[455] + src36[456] + src36[457] + src36[458] + src36[459] + src36[460] + src36[461] + src36[462] + src36[463] + src36[464] + src36[465] + src36[466] + src36[467] + src36[468] + src36[469] + src36[470] + src36[471] + src36[472] + src36[473] + src36[474] + src36[475] + src36[476] + src36[477] + src36[478] + src36[479] + src36[480] + src36[481] + src36[482] + src36[483] + src36[484] + src36[485])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23] + src37[24] + src37[25] + src37[26] + src37[27] + src37[28] + src37[29] + src37[30] + src37[31] + src37[32] + src37[33] + src37[34] + src37[35] + src37[36] + src37[37] + src37[38] + src37[39] + src37[40] + src37[41] + src37[42] + src37[43] + src37[44] + src37[45] + src37[46] + src37[47] + src37[48] + src37[49] + src37[50] + src37[51] + src37[52] + src37[53] + src37[54] + src37[55] + src37[56] + src37[57] + src37[58] + src37[59] + src37[60] + src37[61] + src37[62] + src37[63] + src37[64] + src37[65] + src37[66] + src37[67] + src37[68] + src37[69] + src37[70] + src37[71] + src37[72] + src37[73] + src37[74] + src37[75] + src37[76] + src37[77] + src37[78] + src37[79] + src37[80] + src37[81] + src37[82] + src37[83] + src37[84] + src37[85] + src37[86] + src37[87] + src37[88] + src37[89] + src37[90] + src37[91] + src37[92] + src37[93] + src37[94] + src37[95] + src37[96] + src37[97] + src37[98] + src37[99] + src37[100] + src37[101] + src37[102] + src37[103] + src37[104] + src37[105] + src37[106] + src37[107] + src37[108] + src37[109] + src37[110] + src37[111] + src37[112] + src37[113] + src37[114] + src37[115] + src37[116] + src37[117] + src37[118] + src37[119] + src37[120] + src37[121] + src37[122] + src37[123] + src37[124] + src37[125] + src37[126] + src37[127] + src37[128] + src37[129] + src37[130] + src37[131] + src37[132] + src37[133] + src37[134] + src37[135] + src37[136] + src37[137] + src37[138] + src37[139] + src37[140] + src37[141] + src37[142] + src37[143] + src37[144] + src37[145] + src37[146] + src37[147] + src37[148] + src37[149] + src37[150] + src37[151] + src37[152] + src37[153] + src37[154] + src37[155] + src37[156] + src37[157] + src37[158] + src37[159] + src37[160] + src37[161] + src37[162] + src37[163] + src37[164] + src37[165] + src37[166] + src37[167] + src37[168] + src37[169] + src37[170] + src37[171] + src37[172] + src37[173] + src37[174] + src37[175] + src37[176] + src37[177] + src37[178] + src37[179] + src37[180] + src37[181] + src37[182] + src37[183] + src37[184] + src37[185] + src37[186] + src37[187] + src37[188] + src37[189] + src37[190] + src37[191] + src37[192] + src37[193] + src37[194] + src37[195] + src37[196] + src37[197] + src37[198] + src37[199] + src37[200] + src37[201] + src37[202] + src37[203] + src37[204] + src37[205] + src37[206] + src37[207] + src37[208] + src37[209] + src37[210] + src37[211] + src37[212] + src37[213] + src37[214] + src37[215] + src37[216] + src37[217] + src37[218] + src37[219] + src37[220] + src37[221] + src37[222] + src37[223] + src37[224] + src37[225] + src37[226] + src37[227] + src37[228] + src37[229] + src37[230] + src37[231] + src37[232] + src37[233] + src37[234] + src37[235] + src37[236] + src37[237] + src37[238] + src37[239] + src37[240] + src37[241] + src37[242] + src37[243] + src37[244] + src37[245] + src37[246] + src37[247] + src37[248] + src37[249] + src37[250] + src37[251] + src37[252] + src37[253] + src37[254] + src37[255] + src37[256] + src37[257] + src37[258] + src37[259] + src37[260] + src37[261] + src37[262] + src37[263] + src37[264] + src37[265] + src37[266] + src37[267] + src37[268] + src37[269] + src37[270] + src37[271] + src37[272] + src37[273] + src37[274] + src37[275] + src37[276] + src37[277] + src37[278] + src37[279] + src37[280] + src37[281] + src37[282] + src37[283] + src37[284] + src37[285] + src37[286] + src37[287] + src37[288] + src37[289] + src37[290] + src37[291] + src37[292] + src37[293] + src37[294] + src37[295] + src37[296] + src37[297] + src37[298] + src37[299] + src37[300] + src37[301] + src37[302] + src37[303] + src37[304] + src37[305] + src37[306] + src37[307] + src37[308] + src37[309] + src37[310] + src37[311] + src37[312] + src37[313] + src37[314] + src37[315] + src37[316] + src37[317] + src37[318] + src37[319] + src37[320] + src37[321] + src37[322] + src37[323] + src37[324] + src37[325] + src37[326] + src37[327] + src37[328] + src37[329] + src37[330] + src37[331] + src37[332] + src37[333] + src37[334] + src37[335] + src37[336] + src37[337] + src37[338] + src37[339] + src37[340] + src37[341] + src37[342] + src37[343] + src37[344] + src37[345] + src37[346] + src37[347] + src37[348] + src37[349] + src37[350] + src37[351] + src37[352] + src37[353] + src37[354] + src37[355] + src37[356] + src37[357] + src37[358] + src37[359] + src37[360] + src37[361] + src37[362] + src37[363] + src37[364] + src37[365] + src37[366] + src37[367] + src37[368] + src37[369] + src37[370] + src37[371] + src37[372] + src37[373] + src37[374] + src37[375] + src37[376] + src37[377] + src37[378] + src37[379] + src37[380] + src37[381] + src37[382] + src37[383] + src37[384] + src37[385] + src37[386] + src37[387] + src37[388] + src37[389] + src37[390] + src37[391] + src37[392] + src37[393] + src37[394] + src37[395] + src37[396] + src37[397] + src37[398] + src37[399] + src37[400] + src37[401] + src37[402] + src37[403] + src37[404] + src37[405] + src37[406] + src37[407] + src37[408] + src37[409] + src37[410] + src37[411] + src37[412] + src37[413] + src37[414] + src37[415] + src37[416] + src37[417] + src37[418] + src37[419] + src37[420] + src37[421] + src37[422] + src37[423] + src37[424] + src37[425] + src37[426] + src37[427] + src37[428] + src37[429] + src37[430] + src37[431] + src37[432] + src37[433] + src37[434] + src37[435] + src37[436] + src37[437] + src37[438] + src37[439] + src37[440] + src37[441] + src37[442] + src37[443] + src37[444] + src37[445] + src37[446] + src37[447] + src37[448] + src37[449] + src37[450] + src37[451] + src37[452] + src37[453] + src37[454] + src37[455] + src37[456] + src37[457] + src37[458] + src37[459] + src37[460] + src37[461] + src37[462] + src37[463] + src37[464] + src37[465] + src37[466] + src37[467] + src37[468] + src37[469] + src37[470] + src37[471] + src37[472] + src37[473] + src37[474] + src37[475] + src37[476] + src37[477] + src37[478] + src37[479] + src37[480] + src37[481] + src37[482] + src37[483] + src37[484] + src37[485])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22] + src38[23] + src38[24] + src38[25] + src38[26] + src38[27] + src38[28] + src38[29] + src38[30] + src38[31] + src38[32] + src38[33] + src38[34] + src38[35] + src38[36] + src38[37] + src38[38] + src38[39] + src38[40] + src38[41] + src38[42] + src38[43] + src38[44] + src38[45] + src38[46] + src38[47] + src38[48] + src38[49] + src38[50] + src38[51] + src38[52] + src38[53] + src38[54] + src38[55] + src38[56] + src38[57] + src38[58] + src38[59] + src38[60] + src38[61] + src38[62] + src38[63] + src38[64] + src38[65] + src38[66] + src38[67] + src38[68] + src38[69] + src38[70] + src38[71] + src38[72] + src38[73] + src38[74] + src38[75] + src38[76] + src38[77] + src38[78] + src38[79] + src38[80] + src38[81] + src38[82] + src38[83] + src38[84] + src38[85] + src38[86] + src38[87] + src38[88] + src38[89] + src38[90] + src38[91] + src38[92] + src38[93] + src38[94] + src38[95] + src38[96] + src38[97] + src38[98] + src38[99] + src38[100] + src38[101] + src38[102] + src38[103] + src38[104] + src38[105] + src38[106] + src38[107] + src38[108] + src38[109] + src38[110] + src38[111] + src38[112] + src38[113] + src38[114] + src38[115] + src38[116] + src38[117] + src38[118] + src38[119] + src38[120] + src38[121] + src38[122] + src38[123] + src38[124] + src38[125] + src38[126] + src38[127] + src38[128] + src38[129] + src38[130] + src38[131] + src38[132] + src38[133] + src38[134] + src38[135] + src38[136] + src38[137] + src38[138] + src38[139] + src38[140] + src38[141] + src38[142] + src38[143] + src38[144] + src38[145] + src38[146] + src38[147] + src38[148] + src38[149] + src38[150] + src38[151] + src38[152] + src38[153] + src38[154] + src38[155] + src38[156] + src38[157] + src38[158] + src38[159] + src38[160] + src38[161] + src38[162] + src38[163] + src38[164] + src38[165] + src38[166] + src38[167] + src38[168] + src38[169] + src38[170] + src38[171] + src38[172] + src38[173] + src38[174] + src38[175] + src38[176] + src38[177] + src38[178] + src38[179] + src38[180] + src38[181] + src38[182] + src38[183] + src38[184] + src38[185] + src38[186] + src38[187] + src38[188] + src38[189] + src38[190] + src38[191] + src38[192] + src38[193] + src38[194] + src38[195] + src38[196] + src38[197] + src38[198] + src38[199] + src38[200] + src38[201] + src38[202] + src38[203] + src38[204] + src38[205] + src38[206] + src38[207] + src38[208] + src38[209] + src38[210] + src38[211] + src38[212] + src38[213] + src38[214] + src38[215] + src38[216] + src38[217] + src38[218] + src38[219] + src38[220] + src38[221] + src38[222] + src38[223] + src38[224] + src38[225] + src38[226] + src38[227] + src38[228] + src38[229] + src38[230] + src38[231] + src38[232] + src38[233] + src38[234] + src38[235] + src38[236] + src38[237] + src38[238] + src38[239] + src38[240] + src38[241] + src38[242] + src38[243] + src38[244] + src38[245] + src38[246] + src38[247] + src38[248] + src38[249] + src38[250] + src38[251] + src38[252] + src38[253] + src38[254] + src38[255] + src38[256] + src38[257] + src38[258] + src38[259] + src38[260] + src38[261] + src38[262] + src38[263] + src38[264] + src38[265] + src38[266] + src38[267] + src38[268] + src38[269] + src38[270] + src38[271] + src38[272] + src38[273] + src38[274] + src38[275] + src38[276] + src38[277] + src38[278] + src38[279] + src38[280] + src38[281] + src38[282] + src38[283] + src38[284] + src38[285] + src38[286] + src38[287] + src38[288] + src38[289] + src38[290] + src38[291] + src38[292] + src38[293] + src38[294] + src38[295] + src38[296] + src38[297] + src38[298] + src38[299] + src38[300] + src38[301] + src38[302] + src38[303] + src38[304] + src38[305] + src38[306] + src38[307] + src38[308] + src38[309] + src38[310] + src38[311] + src38[312] + src38[313] + src38[314] + src38[315] + src38[316] + src38[317] + src38[318] + src38[319] + src38[320] + src38[321] + src38[322] + src38[323] + src38[324] + src38[325] + src38[326] + src38[327] + src38[328] + src38[329] + src38[330] + src38[331] + src38[332] + src38[333] + src38[334] + src38[335] + src38[336] + src38[337] + src38[338] + src38[339] + src38[340] + src38[341] + src38[342] + src38[343] + src38[344] + src38[345] + src38[346] + src38[347] + src38[348] + src38[349] + src38[350] + src38[351] + src38[352] + src38[353] + src38[354] + src38[355] + src38[356] + src38[357] + src38[358] + src38[359] + src38[360] + src38[361] + src38[362] + src38[363] + src38[364] + src38[365] + src38[366] + src38[367] + src38[368] + src38[369] + src38[370] + src38[371] + src38[372] + src38[373] + src38[374] + src38[375] + src38[376] + src38[377] + src38[378] + src38[379] + src38[380] + src38[381] + src38[382] + src38[383] + src38[384] + src38[385] + src38[386] + src38[387] + src38[388] + src38[389] + src38[390] + src38[391] + src38[392] + src38[393] + src38[394] + src38[395] + src38[396] + src38[397] + src38[398] + src38[399] + src38[400] + src38[401] + src38[402] + src38[403] + src38[404] + src38[405] + src38[406] + src38[407] + src38[408] + src38[409] + src38[410] + src38[411] + src38[412] + src38[413] + src38[414] + src38[415] + src38[416] + src38[417] + src38[418] + src38[419] + src38[420] + src38[421] + src38[422] + src38[423] + src38[424] + src38[425] + src38[426] + src38[427] + src38[428] + src38[429] + src38[430] + src38[431] + src38[432] + src38[433] + src38[434] + src38[435] + src38[436] + src38[437] + src38[438] + src38[439] + src38[440] + src38[441] + src38[442] + src38[443] + src38[444] + src38[445] + src38[446] + src38[447] + src38[448] + src38[449] + src38[450] + src38[451] + src38[452] + src38[453] + src38[454] + src38[455] + src38[456] + src38[457] + src38[458] + src38[459] + src38[460] + src38[461] + src38[462] + src38[463] + src38[464] + src38[465] + src38[466] + src38[467] + src38[468] + src38[469] + src38[470] + src38[471] + src38[472] + src38[473] + src38[474] + src38[475] + src38[476] + src38[477] + src38[478] + src38[479] + src38[480] + src38[481] + src38[482] + src38[483] + src38[484] + src38[485])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21] + src39[22] + src39[23] + src39[24] + src39[25] + src39[26] + src39[27] + src39[28] + src39[29] + src39[30] + src39[31] + src39[32] + src39[33] + src39[34] + src39[35] + src39[36] + src39[37] + src39[38] + src39[39] + src39[40] + src39[41] + src39[42] + src39[43] + src39[44] + src39[45] + src39[46] + src39[47] + src39[48] + src39[49] + src39[50] + src39[51] + src39[52] + src39[53] + src39[54] + src39[55] + src39[56] + src39[57] + src39[58] + src39[59] + src39[60] + src39[61] + src39[62] + src39[63] + src39[64] + src39[65] + src39[66] + src39[67] + src39[68] + src39[69] + src39[70] + src39[71] + src39[72] + src39[73] + src39[74] + src39[75] + src39[76] + src39[77] + src39[78] + src39[79] + src39[80] + src39[81] + src39[82] + src39[83] + src39[84] + src39[85] + src39[86] + src39[87] + src39[88] + src39[89] + src39[90] + src39[91] + src39[92] + src39[93] + src39[94] + src39[95] + src39[96] + src39[97] + src39[98] + src39[99] + src39[100] + src39[101] + src39[102] + src39[103] + src39[104] + src39[105] + src39[106] + src39[107] + src39[108] + src39[109] + src39[110] + src39[111] + src39[112] + src39[113] + src39[114] + src39[115] + src39[116] + src39[117] + src39[118] + src39[119] + src39[120] + src39[121] + src39[122] + src39[123] + src39[124] + src39[125] + src39[126] + src39[127] + src39[128] + src39[129] + src39[130] + src39[131] + src39[132] + src39[133] + src39[134] + src39[135] + src39[136] + src39[137] + src39[138] + src39[139] + src39[140] + src39[141] + src39[142] + src39[143] + src39[144] + src39[145] + src39[146] + src39[147] + src39[148] + src39[149] + src39[150] + src39[151] + src39[152] + src39[153] + src39[154] + src39[155] + src39[156] + src39[157] + src39[158] + src39[159] + src39[160] + src39[161] + src39[162] + src39[163] + src39[164] + src39[165] + src39[166] + src39[167] + src39[168] + src39[169] + src39[170] + src39[171] + src39[172] + src39[173] + src39[174] + src39[175] + src39[176] + src39[177] + src39[178] + src39[179] + src39[180] + src39[181] + src39[182] + src39[183] + src39[184] + src39[185] + src39[186] + src39[187] + src39[188] + src39[189] + src39[190] + src39[191] + src39[192] + src39[193] + src39[194] + src39[195] + src39[196] + src39[197] + src39[198] + src39[199] + src39[200] + src39[201] + src39[202] + src39[203] + src39[204] + src39[205] + src39[206] + src39[207] + src39[208] + src39[209] + src39[210] + src39[211] + src39[212] + src39[213] + src39[214] + src39[215] + src39[216] + src39[217] + src39[218] + src39[219] + src39[220] + src39[221] + src39[222] + src39[223] + src39[224] + src39[225] + src39[226] + src39[227] + src39[228] + src39[229] + src39[230] + src39[231] + src39[232] + src39[233] + src39[234] + src39[235] + src39[236] + src39[237] + src39[238] + src39[239] + src39[240] + src39[241] + src39[242] + src39[243] + src39[244] + src39[245] + src39[246] + src39[247] + src39[248] + src39[249] + src39[250] + src39[251] + src39[252] + src39[253] + src39[254] + src39[255] + src39[256] + src39[257] + src39[258] + src39[259] + src39[260] + src39[261] + src39[262] + src39[263] + src39[264] + src39[265] + src39[266] + src39[267] + src39[268] + src39[269] + src39[270] + src39[271] + src39[272] + src39[273] + src39[274] + src39[275] + src39[276] + src39[277] + src39[278] + src39[279] + src39[280] + src39[281] + src39[282] + src39[283] + src39[284] + src39[285] + src39[286] + src39[287] + src39[288] + src39[289] + src39[290] + src39[291] + src39[292] + src39[293] + src39[294] + src39[295] + src39[296] + src39[297] + src39[298] + src39[299] + src39[300] + src39[301] + src39[302] + src39[303] + src39[304] + src39[305] + src39[306] + src39[307] + src39[308] + src39[309] + src39[310] + src39[311] + src39[312] + src39[313] + src39[314] + src39[315] + src39[316] + src39[317] + src39[318] + src39[319] + src39[320] + src39[321] + src39[322] + src39[323] + src39[324] + src39[325] + src39[326] + src39[327] + src39[328] + src39[329] + src39[330] + src39[331] + src39[332] + src39[333] + src39[334] + src39[335] + src39[336] + src39[337] + src39[338] + src39[339] + src39[340] + src39[341] + src39[342] + src39[343] + src39[344] + src39[345] + src39[346] + src39[347] + src39[348] + src39[349] + src39[350] + src39[351] + src39[352] + src39[353] + src39[354] + src39[355] + src39[356] + src39[357] + src39[358] + src39[359] + src39[360] + src39[361] + src39[362] + src39[363] + src39[364] + src39[365] + src39[366] + src39[367] + src39[368] + src39[369] + src39[370] + src39[371] + src39[372] + src39[373] + src39[374] + src39[375] + src39[376] + src39[377] + src39[378] + src39[379] + src39[380] + src39[381] + src39[382] + src39[383] + src39[384] + src39[385] + src39[386] + src39[387] + src39[388] + src39[389] + src39[390] + src39[391] + src39[392] + src39[393] + src39[394] + src39[395] + src39[396] + src39[397] + src39[398] + src39[399] + src39[400] + src39[401] + src39[402] + src39[403] + src39[404] + src39[405] + src39[406] + src39[407] + src39[408] + src39[409] + src39[410] + src39[411] + src39[412] + src39[413] + src39[414] + src39[415] + src39[416] + src39[417] + src39[418] + src39[419] + src39[420] + src39[421] + src39[422] + src39[423] + src39[424] + src39[425] + src39[426] + src39[427] + src39[428] + src39[429] + src39[430] + src39[431] + src39[432] + src39[433] + src39[434] + src39[435] + src39[436] + src39[437] + src39[438] + src39[439] + src39[440] + src39[441] + src39[442] + src39[443] + src39[444] + src39[445] + src39[446] + src39[447] + src39[448] + src39[449] + src39[450] + src39[451] + src39[452] + src39[453] + src39[454] + src39[455] + src39[456] + src39[457] + src39[458] + src39[459] + src39[460] + src39[461] + src39[462] + src39[463] + src39[464] + src39[465] + src39[466] + src39[467] + src39[468] + src39[469] + src39[470] + src39[471] + src39[472] + src39[473] + src39[474] + src39[475] + src39[476] + src39[477] + src39[478] + src39[479] + src39[480] + src39[481] + src39[482] + src39[483] + src39[484] + src39[485])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20] + src40[21] + src40[22] + src40[23] + src40[24] + src40[25] + src40[26] + src40[27] + src40[28] + src40[29] + src40[30] + src40[31] + src40[32] + src40[33] + src40[34] + src40[35] + src40[36] + src40[37] + src40[38] + src40[39] + src40[40] + src40[41] + src40[42] + src40[43] + src40[44] + src40[45] + src40[46] + src40[47] + src40[48] + src40[49] + src40[50] + src40[51] + src40[52] + src40[53] + src40[54] + src40[55] + src40[56] + src40[57] + src40[58] + src40[59] + src40[60] + src40[61] + src40[62] + src40[63] + src40[64] + src40[65] + src40[66] + src40[67] + src40[68] + src40[69] + src40[70] + src40[71] + src40[72] + src40[73] + src40[74] + src40[75] + src40[76] + src40[77] + src40[78] + src40[79] + src40[80] + src40[81] + src40[82] + src40[83] + src40[84] + src40[85] + src40[86] + src40[87] + src40[88] + src40[89] + src40[90] + src40[91] + src40[92] + src40[93] + src40[94] + src40[95] + src40[96] + src40[97] + src40[98] + src40[99] + src40[100] + src40[101] + src40[102] + src40[103] + src40[104] + src40[105] + src40[106] + src40[107] + src40[108] + src40[109] + src40[110] + src40[111] + src40[112] + src40[113] + src40[114] + src40[115] + src40[116] + src40[117] + src40[118] + src40[119] + src40[120] + src40[121] + src40[122] + src40[123] + src40[124] + src40[125] + src40[126] + src40[127] + src40[128] + src40[129] + src40[130] + src40[131] + src40[132] + src40[133] + src40[134] + src40[135] + src40[136] + src40[137] + src40[138] + src40[139] + src40[140] + src40[141] + src40[142] + src40[143] + src40[144] + src40[145] + src40[146] + src40[147] + src40[148] + src40[149] + src40[150] + src40[151] + src40[152] + src40[153] + src40[154] + src40[155] + src40[156] + src40[157] + src40[158] + src40[159] + src40[160] + src40[161] + src40[162] + src40[163] + src40[164] + src40[165] + src40[166] + src40[167] + src40[168] + src40[169] + src40[170] + src40[171] + src40[172] + src40[173] + src40[174] + src40[175] + src40[176] + src40[177] + src40[178] + src40[179] + src40[180] + src40[181] + src40[182] + src40[183] + src40[184] + src40[185] + src40[186] + src40[187] + src40[188] + src40[189] + src40[190] + src40[191] + src40[192] + src40[193] + src40[194] + src40[195] + src40[196] + src40[197] + src40[198] + src40[199] + src40[200] + src40[201] + src40[202] + src40[203] + src40[204] + src40[205] + src40[206] + src40[207] + src40[208] + src40[209] + src40[210] + src40[211] + src40[212] + src40[213] + src40[214] + src40[215] + src40[216] + src40[217] + src40[218] + src40[219] + src40[220] + src40[221] + src40[222] + src40[223] + src40[224] + src40[225] + src40[226] + src40[227] + src40[228] + src40[229] + src40[230] + src40[231] + src40[232] + src40[233] + src40[234] + src40[235] + src40[236] + src40[237] + src40[238] + src40[239] + src40[240] + src40[241] + src40[242] + src40[243] + src40[244] + src40[245] + src40[246] + src40[247] + src40[248] + src40[249] + src40[250] + src40[251] + src40[252] + src40[253] + src40[254] + src40[255] + src40[256] + src40[257] + src40[258] + src40[259] + src40[260] + src40[261] + src40[262] + src40[263] + src40[264] + src40[265] + src40[266] + src40[267] + src40[268] + src40[269] + src40[270] + src40[271] + src40[272] + src40[273] + src40[274] + src40[275] + src40[276] + src40[277] + src40[278] + src40[279] + src40[280] + src40[281] + src40[282] + src40[283] + src40[284] + src40[285] + src40[286] + src40[287] + src40[288] + src40[289] + src40[290] + src40[291] + src40[292] + src40[293] + src40[294] + src40[295] + src40[296] + src40[297] + src40[298] + src40[299] + src40[300] + src40[301] + src40[302] + src40[303] + src40[304] + src40[305] + src40[306] + src40[307] + src40[308] + src40[309] + src40[310] + src40[311] + src40[312] + src40[313] + src40[314] + src40[315] + src40[316] + src40[317] + src40[318] + src40[319] + src40[320] + src40[321] + src40[322] + src40[323] + src40[324] + src40[325] + src40[326] + src40[327] + src40[328] + src40[329] + src40[330] + src40[331] + src40[332] + src40[333] + src40[334] + src40[335] + src40[336] + src40[337] + src40[338] + src40[339] + src40[340] + src40[341] + src40[342] + src40[343] + src40[344] + src40[345] + src40[346] + src40[347] + src40[348] + src40[349] + src40[350] + src40[351] + src40[352] + src40[353] + src40[354] + src40[355] + src40[356] + src40[357] + src40[358] + src40[359] + src40[360] + src40[361] + src40[362] + src40[363] + src40[364] + src40[365] + src40[366] + src40[367] + src40[368] + src40[369] + src40[370] + src40[371] + src40[372] + src40[373] + src40[374] + src40[375] + src40[376] + src40[377] + src40[378] + src40[379] + src40[380] + src40[381] + src40[382] + src40[383] + src40[384] + src40[385] + src40[386] + src40[387] + src40[388] + src40[389] + src40[390] + src40[391] + src40[392] + src40[393] + src40[394] + src40[395] + src40[396] + src40[397] + src40[398] + src40[399] + src40[400] + src40[401] + src40[402] + src40[403] + src40[404] + src40[405] + src40[406] + src40[407] + src40[408] + src40[409] + src40[410] + src40[411] + src40[412] + src40[413] + src40[414] + src40[415] + src40[416] + src40[417] + src40[418] + src40[419] + src40[420] + src40[421] + src40[422] + src40[423] + src40[424] + src40[425] + src40[426] + src40[427] + src40[428] + src40[429] + src40[430] + src40[431] + src40[432] + src40[433] + src40[434] + src40[435] + src40[436] + src40[437] + src40[438] + src40[439] + src40[440] + src40[441] + src40[442] + src40[443] + src40[444] + src40[445] + src40[446] + src40[447] + src40[448] + src40[449] + src40[450] + src40[451] + src40[452] + src40[453] + src40[454] + src40[455] + src40[456] + src40[457] + src40[458] + src40[459] + src40[460] + src40[461] + src40[462] + src40[463] + src40[464] + src40[465] + src40[466] + src40[467] + src40[468] + src40[469] + src40[470] + src40[471] + src40[472] + src40[473] + src40[474] + src40[475] + src40[476] + src40[477] + src40[478] + src40[479] + src40[480] + src40[481] + src40[482] + src40[483] + src40[484] + src40[485])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19] + src41[20] + src41[21] + src41[22] + src41[23] + src41[24] + src41[25] + src41[26] + src41[27] + src41[28] + src41[29] + src41[30] + src41[31] + src41[32] + src41[33] + src41[34] + src41[35] + src41[36] + src41[37] + src41[38] + src41[39] + src41[40] + src41[41] + src41[42] + src41[43] + src41[44] + src41[45] + src41[46] + src41[47] + src41[48] + src41[49] + src41[50] + src41[51] + src41[52] + src41[53] + src41[54] + src41[55] + src41[56] + src41[57] + src41[58] + src41[59] + src41[60] + src41[61] + src41[62] + src41[63] + src41[64] + src41[65] + src41[66] + src41[67] + src41[68] + src41[69] + src41[70] + src41[71] + src41[72] + src41[73] + src41[74] + src41[75] + src41[76] + src41[77] + src41[78] + src41[79] + src41[80] + src41[81] + src41[82] + src41[83] + src41[84] + src41[85] + src41[86] + src41[87] + src41[88] + src41[89] + src41[90] + src41[91] + src41[92] + src41[93] + src41[94] + src41[95] + src41[96] + src41[97] + src41[98] + src41[99] + src41[100] + src41[101] + src41[102] + src41[103] + src41[104] + src41[105] + src41[106] + src41[107] + src41[108] + src41[109] + src41[110] + src41[111] + src41[112] + src41[113] + src41[114] + src41[115] + src41[116] + src41[117] + src41[118] + src41[119] + src41[120] + src41[121] + src41[122] + src41[123] + src41[124] + src41[125] + src41[126] + src41[127] + src41[128] + src41[129] + src41[130] + src41[131] + src41[132] + src41[133] + src41[134] + src41[135] + src41[136] + src41[137] + src41[138] + src41[139] + src41[140] + src41[141] + src41[142] + src41[143] + src41[144] + src41[145] + src41[146] + src41[147] + src41[148] + src41[149] + src41[150] + src41[151] + src41[152] + src41[153] + src41[154] + src41[155] + src41[156] + src41[157] + src41[158] + src41[159] + src41[160] + src41[161] + src41[162] + src41[163] + src41[164] + src41[165] + src41[166] + src41[167] + src41[168] + src41[169] + src41[170] + src41[171] + src41[172] + src41[173] + src41[174] + src41[175] + src41[176] + src41[177] + src41[178] + src41[179] + src41[180] + src41[181] + src41[182] + src41[183] + src41[184] + src41[185] + src41[186] + src41[187] + src41[188] + src41[189] + src41[190] + src41[191] + src41[192] + src41[193] + src41[194] + src41[195] + src41[196] + src41[197] + src41[198] + src41[199] + src41[200] + src41[201] + src41[202] + src41[203] + src41[204] + src41[205] + src41[206] + src41[207] + src41[208] + src41[209] + src41[210] + src41[211] + src41[212] + src41[213] + src41[214] + src41[215] + src41[216] + src41[217] + src41[218] + src41[219] + src41[220] + src41[221] + src41[222] + src41[223] + src41[224] + src41[225] + src41[226] + src41[227] + src41[228] + src41[229] + src41[230] + src41[231] + src41[232] + src41[233] + src41[234] + src41[235] + src41[236] + src41[237] + src41[238] + src41[239] + src41[240] + src41[241] + src41[242] + src41[243] + src41[244] + src41[245] + src41[246] + src41[247] + src41[248] + src41[249] + src41[250] + src41[251] + src41[252] + src41[253] + src41[254] + src41[255] + src41[256] + src41[257] + src41[258] + src41[259] + src41[260] + src41[261] + src41[262] + src41[263] + src41[264] + src41[265] + src41[266] + src41[267] + src41[268] + src41[269] + src41[270] + src41[271] + src41[272] + src41[273] + src41[274] + src41[275] + src41[276] + src41[277] + src41[278] + src41[279] + src41[280] + src41[281] + src41[282] + src41[283] + src41[284] + src41[285] + src41[286] + src41[287] + src41[288] + src41[289] + src41[290] + src41[291] + src41[292] + src41[293] + src41[294] + src41[295] + src41[296] + src41[297] + src41[298] + src41[299] + src41[300] + src41[301] + src41[302] + src41[303] + src41[304] + src41[305] + src41[306] + src41[307] + src41[308] + src41[309] + src41[310] + src41[311] + src41[312] + src41[313] + src41[314] + src41[315] + src41[316] + src41[317] + src41[318] + src41[319] + src41[320] + src41[321] + src41[322] + src41[323] + src41[324] + src41[325] + src41[326] + src41[327] + src41[328] + src41[329] + src41[330] + src41[331] + src41[332] + src41[333] + src41[334] + src41[335] + src41[336] + src41[337] + src41[338] + src41[339] + src41[340] + src41[341] + src41[342] + src41[343] + src41[344] + src41[345] + src41[346] + src41[347] + src41[348] + src41[349] + src41[350] + src41[351] + src41[352] + src41[353] + src41[354] + src41[355] + src41[356] + src41[357] + src41[358] + src41[359] + src41[360] + src41[361] + src41[362] + src41[363] + src41[364] + src41[365] + src41[366] + src41[367] + src41[368] + src41[369] + src41[370] + src41[371] + src41[372] + src41[373] + src41[374] + src41[375] + src41[376] + src41[377] + src41[378] + src41[379] + src41[380] + src41[381] + src41[382] + src41[383] + src41[384] + src41[385] + src41[386] + src41[387] + src41[388] + src41[389] + src41[390] + src41[391] + src41[392] + src41[393] + src41[394] + src41[395] + src41[396] + src41[397] + src41[398] + src41[399] + src41[400] + src41[401] + src41[402] + src41[403] + src41[404] + src41[405] + src41[406] + src41[407] + src41[408] + src41[409] + src41[410] + src41[411] + src41[412] + src41[413] + src41[414] + src41[415] + src41[416] + src41[417] + src41[418] + src41[419] + src41[420] + src41[421] + src41[422] + src41[423] + src41[424] + src41[425] + src41[426] + src41[427] + src41[428] + src41[429] + src41[430] + src41[431] + src41[432] + src41[433] + src41[434] + src41[435] + src41[436] + src41[437] + src41[438] + src41[439] + src41[440] + src41[441] + src41[442] + src41[443] + src41[444] + src41[445] + src41[446] + src41[447] + src41[448] + src41[449] + src41[450] + src41[451] + src41[452] + src41[453] + src41[454] + src41[455] + src41[456] + src41[457] + src41[458] + src41[459] + src41[460] + src41[461] + src41[462] + src41[463] + src41[464] + src41[465] + src41[466] + src41[467] + src41[468] + src41[469] + src41[470] + src41[471] + src41[472] + src41[473] + src41[474] + src41[475] + src41[476] + src41[477] + src41[478] + src41[479] + src41[480] + src41[481] + src41[482] + src41[483] + src41[484] + src41[485])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18] + src42[19] + src42[20] + src42[21] + src42[22] + src42[23] + src42[24] + src42[25] + src42[26] + src42[27] + src42[28] + src42[29] + src42[30] + src42[31] + src42[32] + src42[33] + src42[34] + src42[35] + src42[36] + src42[37] + src42[38] + src42[39] + src42[40] + src42[41] + src42[42] + src42[43] + src42[44] + src42[45] + src42[46] + src42[47] + src42[48] + src42[49] + src42[50] + src42[51] + src42[52] + src42[53] + src42[54] + src42[55] + src42[56] + src42[57] + src42[58] + src42[59] + src42[60] + src42[61] + src42[62] + src42[63] + src42[64] + src42[65] + src42[66] + src42[67] + src42[68] + src42[69] + src42[70] + src42[71] + src42[72] + src42[73] + src42[74] + src42[75] + src42[76] + src42[77] + src42[78] + src42[79] + src42[80] + src42[81] + src42[82] + src42[83] + src42[84] + src42[85] + src42[86] + src42[87] + src42[88] + src42[89] + src42[90] + src42[91] + src42[92] + src42[93] + src42[94] + src42[95] + src42[96] + src42[97] + src42[98] + src42[99] + src42[100] + src42[101] + src42[102] + src42[103] + src42[104] + src42[105] + src42[106] + src42[107] + src42[108] + src42[109] + src42[110] + src42[111] + src42[112] + src42[113] + src42[114] + src42[115] + src42[116] + src42[117] + src42[118] + src42[119] + src42[120] + src42[121] + src42[122] + src42[123] + src42[124] + src42[125] + src42[126] + src42[127] + src42[128] + src42[129] + src42[130] + src42[131] + src42[132] + src42[133] + src42[134] + src42[135] + src42[136] + src42[137] + src42[138] + src42[139] + src42[140] + src42[141] + src42[142] + src42[143] + src42[144] + src42[145] + src42[146] + src42[147] + src42[148] + src42[149] + src42[150] + src42[151] + src42[152] + src42[153] + src42[154] + src42[155] + src42[156] + src42[157] + src42[158] + src42[159] + src42[160] + src42[161] + src42[162] + src42[163] + src42[164] + src42[165] + src42[166] + src42[167] + src42[168] + src42[169] + src42[170] + src42[171] + src42[172] + src42[173] + src42[174] + src42[175] + src42[176] + src42[177] + src42[178] + src42[179] + src42[180] + src42[181] + src42[182] + src42[183] + src42[184] + src42[185] + src42[186] + src42[187] + src42[188] + src42[189] + src42[190] + src42[191] + src42[192] + src42[193] + src42[194] + src42[195] + src42[196] + src42[197] + src42[198] + src42[199] + src42[200] + src42[201] + src42[202] + src42[203] + src42[204] + src42[205] + src42[206] + src42[207] + src42[208] + src42[209] + src42[210] + src42[211] + src42[212] + src42[213] + src42[214] + src42[215] + src42[216] + src42[217] + src42[218] + src42[219] + src42[220] + src42[221] + src42[222] + src42[223] + src42[224] + src42[225] + src42[226] + src42[227] + src42[228] + src42[229] + src42[230] + src42[231] + src42[232] + src42[233] + src42[234] + src42[235] + src42[236] + src42[237] + src42[238] + src42[239] + src42[240] + src42[241] + src42[242] + src42[243] + src42[244] + src42[245] + src42[246] + src42[247] + src42[248] + src42[249] + src42[250] + src42[251] + src42[252] + src42[253] + src42[254] + src42[255] + src42[256] + src42[257] + src42[258] + src42[259] + src42[260] + src42[261] + src42[262] + src42[263] + src42[264] + src42[265] + src42[266] + src42[267] + src42[268] + src42[269] + src42[270] + src42[271] + src42[272] + src42[273] + src42[274] + src42[275] + src42[276] + src42[277] + src42[278] + src42[279] + src42[280] + src42[281] + src42[282] + src42[283] + src42[284] + src42[285] + src42[286] + src42[287] + src42[288] + src42[289] + src42[290] + src42[291] + src42[292] + src42[293] + src42[294] + src42[295] + src42[296] + src42[297] + src42[298] + src42[299] + src42[300] + src42[301] + src42[302] + src42[303] + src42[304] + src42[305] + src42[306] + src42[307] + src42[308] + src42[309] + src42[310] + src42[311] + src42[312] + src42[313] + src42[314] + src42[315] + src42[316] + src42[317] + src42[318] + src42[319] + src42[320] + src42[321] + src42[322] + src42[323] + src42[324] + src42[325] + src42[326] + src42[327] + src42[328] + src42[329] + src42[330] + src42[331] + src42[332] + src42[333] + src42[334] + src42[335] + src42[336] + src42[337] + src42[338] + src42[339] + src42[340] + src42[341] + src42[342] + src42[343] + src42[344] + src42[345] + src42[346] + src42[347] + src42[348] + src42[349] + src42[350] + src42[351] + src42[352] + src42[353] + src42[354] + src42[355] + src42[356] + src42[357] + src42[358] + src42[359] + src42[360] + src42[361] + src42[362] + src42[363] + src42[364] + src42[365] + src42[366] + src42[367] + src42[368] + src42[369] + src42[370] + src42[371] + src42[372] + src42[373] + src42[374] + src42[375] + src42[376] + src42[377] + src42[378] + src42[379] + src42[380] + src42[381] + src42[382] + src42[383] + src42[384] + src42[385] + src42[386] + src42[387] + src42[388] + src42[389] + src42[390] + src42[391] + src42[392] + src42[393] + src42[394] + src42[395] + src42[396] + src42[397] + src42[398] + src42[399] + src42[400] + src42[401] + src42[402] + src42[403] + src42[404] + src42[405] + src42[406] + src42[407] + src42[408] + src42[409] + src42[410] + src42[411] + src42[412] + src42[413] + src42[414] + src42[415] + src42[416] + src42[417] + src42[418] + src42[419] + src42[420] + src42[421] + src42[422] + src42[423] + src42[424] + src42[425] + src42[426] + src42[427] + src42[428] + src42[429] + src42[430] + src42[431] + src42[432] + src42[433] + src42[434] + src42[435] + src42[436] + src42[437] + src42[438] + src42[439] + src42[440] + src42[441] + src42[442] + src42[443] + src42[444] + src42[445] + src42[446] + src42[447] + src42[448] + src42[449] + src42[450] + src42[451] + src42[452] + src42[453] + src42[454] + src42[455] + src42[456] + src42[457] + src42[458] + src42[459] + src42[460] + src42[461] + src42[462] + src42[463] + src42[464] + src42[465] + src42[466] + src42[467] + src42[468] + src42[469] + src42[470] + src42[471] + src42[472] + src42[473] + src42[474] + src42[475] + src42[476] + src42[477] + src42[478] + src42[479] + src42[480] + src42[481] + src42[482] + src42[483] + src42[484] + src42[485])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17] + src43[18] + src43[19] + src43[20] + src43[21] + src43[22] + src43[23] + src43[24] + src43[25] + src43[26] + src43[27] + src43[28] + src43[29] + src43[30] + src43[31] + src43[32] + src43[33] + src43[34] + src43[35] + src43[36] + src43[37] + src43[38] + src43[39] + src43[40] + src43[41] + src43[42] + src43[43] + src43[44] + src43[45] + src43[46] + src43[47] + src43[48] + src43[49] + src43[50] + src43[51] + src43[52] + src43[53] + src43[54] + src43[55] + src43[56] + src43[57] + src43[58] + src43[59] + src43[60] + src43[61] + src43[62] + src43[63] + src43[64] + src43[65] + src43[66] + src43[67] + src43[68] + src43[69] + src43[70] + src43[71] + src43[72] + src43[73] + src43[74] + src43[75] + src43[76] + src43[77] + src43[78] + src43[79] + src43[80] + src43[81] + src43[82] + src43[83] + src43[84] + src43[85] + src43[86] + src43[87] + src43[88] + src43[89] + src43[90] + src43[91] + src43[92] + src43[93] + src43[94] + src43[95] + src43[96] + src43[97] + src43[98] + src43[99] + src43[100] + src43[101] + src43[102] + src43[103] + src43[104] + src43[105] + src43[106] + src43[107] + src43[108] + src43[109] + src43[110] + src43[111] + src43[112] + src43[113] + src43[114] + src43[115] + src43[116] + src43[117] + src43[118] + src43[119] + src43[120] + src43[121] + src43[122] + src43[123] + src43[124] + src43[125] + src43[126] + src43[127] + src43[128] + src43[129] + src43[130] + src43[131] + src43[132] + src43[133] + src43[134] + src43[135] + src43[136] + src43[137] + src43[138] + src43[139] + src43[140] + src43[141] + src43[142] + src43[143] + src43[144] + src43[145] + src43[146] + src43[147] + src43[148] + src43[149] + src43[150] + src43[151] + src43[152] + src43[153] + src43[154] + src43[155] + src43[156] + src43[157] + src43[158] + src43[159] + src43[160] + src43[161] + src43[162] + src43[163] + src43[164] + src43[165] + src43[166] + src43[167] + src43[168] + src43[169] + src43[170] + src43[171] + src43[172] + src43[173] + src43[174] + src43[175] + src43[176] + src43[177] + src43[178] + src43[179] + src43[180] + src43[181] + src43[182] + src43[183] + src43[184] + src43[185] + src43[186] + src43[187] + src43[188] + src43[189] + src43[190] + src43[191] + src43[192] + src43[193] + src43[194] + src43[195] + src43[196] + src43[197] + src43[198] + src43[199] + src43[200] + src43[201] + src43[202] + src43[203] + src43[204] + src43[205] + src43[206] + src43[207] + src43[208] + src43[209] + src43[210] + src43[211] + src43[212] + src43[213] + src43[214] + src43[215] + src43[216] + src43[217] + src43[218] + src43[219] + src43[220] + src43[221] + src43[222] + src43[223] + src43[224] + src43[225] + src43[226] + src43[227] + src43[228] + src43[229] + src43[230] + src43[231] + src43[232] + src43[233] + src43[234] + src43[235] + src43[236] + src43[237] + src43[238] + src43[239] + src43[240] + src43[241] + src43[242] + src43[243] + src43[244] + src43[245] + src43[246] + src43[247] + src43[248] + src43[249] + src43[250] + src43[251] + src43[252] + src43[253] + src43[254] + src43[255] + src43[256] + src43[257] + src43[258] + src43[259] + src43[260] + src43[261] + src43[262] + src43[263] + src43[264] + src43[265] + src43[266] + src43[267] + src43[268] + src43[269] + src43[270] + src43[271] + src43[272] + src43[273] + src43[274] + src43[275] + src43[276] + src43[277] + src43[278] + src43[279] + src43[280] + src43[281] + src43[282] + src43[283] + src43[284] + src43[285] + src43[286] + src43[287] + src43[288] + src43[289] + src43[290] + src43[291] + src43[292] + src43[293] + src43[294] + src43[295] + src43[296] + src43[297] + src43[298] + src43[299] + src43[300] + src43[301] + src43[302] + src43[303] + src43[304] + src43[305] + src43[306] + src43[307] + src43[308] + src43[309] + src43[310] + src43[311] + src43[312] + src43[313] + src43[314] + src43[315] + src43[316] + src43[317] + src43[318] + src43[319] + src43[320] + src43[321] + src43[322] + src43[323] + src43[324] + src43[325] + src43[326] + src43[327] + src43[328] + src43[329] + src43[330] + src43[331] + src43[332] + src43[333] + src43[334] + src43[335] + src43[336] + src43[337] + src43[338] + src43[339] + src43[340] + src43[341] + src43[342] + src43[343] + src43[344] + src43[345] + src43[346] + src43[347] + src43[348] + src43[349] + src43[350] + src43[351] + src43[352] + src43[353] + src43[354] + src43[355] + src43[356] + src43[357] + src43[358] + src43[359] + src43[360] + src43[361] + src43[362] + src43[363] + src43[364] + src43[365] + src43[366] + src43[367] + src43[368] + src43[369] + src43[370] + src43[371] + src43[372] + src43[373] + src43[374] + src43[375] + src43[376] + src43[377] + src43[378] + src43[379] + src43[380] + src43[381] + src43[382] + src43[383] + src43[384] + src43[385] + src43[386] + src43[387] + src43[388] + src43[389] + src43[390] + src43[391] + src43[392] + src43[393] + src43[394] + src43[395] + src43[396] + src43[397] + src43[398] + src43[399] + src43[400] + src43[401] + src43[402] + src43[403] + src43[404] + src43[405] + src43[406] + src43[407] + src43[408] + src43[409] + src43[410] + src43[411] + src43[412] + src43[413] + src43[414] + src43[415] + src43[416] + src43[417] + src43[418] + src43[419] + src43[420] + src43[421] + src43[422] + src43[423] + src43[424] + src43[425] + src43[426] + src43[427] + src43[428] + src43[429] + src43[430] + src43[431] + src43[432] + src43[433] + src43[434] + src43[435] + src43[436] + src43[437] + src43[438] + src43[439] + src43[440] + src43[441] + src43[442] + src43[443] + src43[444] + src43[445] + src43[446] + src43[447] + src43[448] + src43[449] + src43[450] + src43[451] + src43[452] + src43[453] + src43[454] + src43[455] + src43[456] + src43[457] + src43[458] + src43[459] + src43[460] + src43[461] + src43[462] + src43[463] + src43[464] + src43[465] + src43[466] + src43[467] + src43[468] + src43[469] + src43[470] + src43[471] + src43[472] + src43[473] + src43[474] + src43[475] + src43[476] + src43[477] + src43[478] + src43[479] + src43[480] + src43[481] + src43[482] + src43[483] + src43[484] + src43[485])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16] + src44[17] + src44[18] + src44[19] + src44[20] + src44[21] + src44[22] + src44[23] + src44[24] + src44[25] + src44[26] + src44[27] + src44[28] + src44[29] + src44[30] + src44[31] + src44[32] + src44[33] + src44[34] + src44[35] + src44[36] + src44[37] + src44[38] + src44[39] + src44[40] + src44[41] + src44[42] + src44[43] + src44[44] + src44[45] + src44[46] + src44[47] + src44[48] + src44[49] + src44[50] + src44[51] + src44[52] + src44[53] + src44[54] + src44[55] + src44[56] + src44[57] + src44[58] + src44[59] + src44[60] + src44[61] + src44[62] + src44[63] + src44[64] + src44[65] + src44[66] + src44[67] + src44[68] + src44[69] + src44[70] + src44[71] + src44[72] + src44[73] + src44[74] + src44[75] + src44[76] + src44[77] + src44[78] + src44[79] + src44[80] + src44[81] + src44[82] + src44[83] + src44[84] + src44[85] + src44[86] + src44[87] + src44[88] + src44[89] + src44[90] + src44[91] + src44[92] + src44[93] + src44[94] + src44[95] + src44[96] + src44[97] + src44[98] + src44[99] + src44[100] + src44[101] + src44[102] + src44[103] + src44[104] + src44[105] + src44[106] + src44[107] + src44[108] + src44[109] + src44[110] + src44[111] + src44[112] + src44[113] + src44[114] + src44[115] + src44[116] + src44[117] + src44[118] + src44[119] + src44[120] + src44[121] + src44[122] + src44[123] + src44[124] + src44[125] + src44[126] + src44[127] + src44[128] + src44[129] + src44[130] + src44[131] + src44[132] + src44[133] + src44[134] + src44[135] + src44[136] + src44[137] + src44[138] + src44[139] + src44[140] + src44[141] + src44[142] + src44[143] + src44[144] + src44[145] + src44[146] + src44[147] + src44[148] + src44[149] + src44[150] + src44[151] + src44[152] + src44[153] + src44[154] + src44[155] + src44[156] + src44[157] + src44[158] + src44[159] + src44[160] + src44[161] + src44[162] + src44[163] + src44[164] + src44[165] + src44[166] + src44[167] + src44[168] + src44[169] + src44[170] + src44[171] + src44[172] + src44[173] + src44[174] + src44[175] + src44[176] + src44[177] + src44[178] + src44[179] + src44[180] + src44[181] + src44[182] + src44[183] + src44[184] + src44[185] + src44[186] + src44[187] + src44[188] + src44[189] + src44[190] + src44[191] + src44[192] + src44[193] + src44[194] + src44[195] + src44[196] + src44[197] + src44[198] + src44[199] + src44[200] + src44[201] + src44[202] + src44[203] + src44[204] + src44[205] + src44[206] + src44[207] + src44[208] + src44[209] + src44[210] + src44[211] + src44[212] + src44[213] + src44[214] + src44[215] + src44[216] + src44[217] + src44[218] + src44[219] + src44[220] + src44[221] + src44[222] + src44[223] + src44[224] + src44[225] + src44[226] + src44[227] + src44[228] + src44[229] + src44[230] + src44[231] + src44[232] + src44[233] + src44[234] + src44[235] + src44[236] + src44[237] + src44[238] + src44[239] + src44[240] + src44[241] + src44[242] + src44[243] + src44[244] + src44[245] + src44[246] + src44[247] + src44[248] + src44[249] + src44[250] + src44[251] + src44[252] + src44[253] + src44[254] + src44[255] + src44[256] + src44[257] + src44[258] + src44[259] + src44[260] + src44[261] + src44[262] + src44[263] + src44[264] + src44[265] + src44[266] + src44[267] + src44[268] + src44[269] + src44[270] + src44[271] + src44[272] + src44[273] + src44[274] + src44[275] + src44[276] + src44[277] + src44[278] + src44[279] + src44[280] + src44[281] + src44[282] + src44[283] + src44[284] + src44[285] + src44[286] + src44[287] + src44[288] + src44[289] + src44[290] + src44[291] + src44[292] + src44[293] + src44[294] + src44[295] + src44[296] + src44[297] + src44[298] + src44[299] + src44[300] + src44[301] + src44[302] + src44[303] + src44[304] + src44[305] + src44[306] + src44[307] + src44[308] + src44[309] + src44[310] + src44[311] + src44[312] + src44[313] + src44[314] + src44[315] + src44[316] + src44[317] + src44[318] + src44[319] + src44[320] + src44[321] + src44[322] + src44[323] + src44[324] + src44[325] + src44[326] + src44[327] + src44[328] + src44[329] + src44[330] + src44[331] + src44[332] + src44[333] + src44[334] + src44[335] + src44[336] + src44[337] + src44[338] + src44[339] + src44[340] + src44[341] + src44[342] + src44[343] + src44[344] + src44[345] + src44[346] + src44[347] + src44[348] + src44[349] + src44[350] + src44[351] + src44[352] + src44[353] + src44[354] + src44[355] + src44[356] + src44[357] + src44[358] + src44[359] + src44[360] + src44[361] + src44[362] + src44[363] + src44[364] + src44[365] + src44[366] + src44[367] + src44[368] + src44[369] + src44[370] + src44[371] + src44[372] + src44[373] + src44[374] + src44[375] + src44[376] + src44[377] + src44[378] + src44[379] + src44[380] + src44[381] + src44[382] + src44[383] + src44[384] + src44[385] + src44[386] + src44[387] + src44[388] + src44[389] + src44[390] + src44[391] + src44[392] + src44[393] + src44[394] + src44[395] + src44[396] + src44[397] + src44[398] + src44[399] + src44[400] + src44[401] + src44[402] + src44[403] + src44[404] + src44[405] + src44[406] + src44[407] + src44[408] + src44[409] + src44[410] + src44[411] + src44[412] + src44[413] + src44[414] + src44[415] + src44[416] + src44[417] + src44[418] + src44[419] + src44[420] + src44[421] + src44[422] + src44[423] + src44[424] + src44[425] + src44[426] + src44[427] + src44[428] + src44[429] + src44[430] + src44[431] + src44[432] + src44[433] + src44[434] + src44[435] + src44[436] + src44[437] + src44[438] + src44[439] + src44[440] + src44[441] + src44[442] + src44[443] + src44[444] + src44[445] + src44[446] + src44[447] + src44[448] + src44[449] + src44[450] + src44[451] + src44[452] + src44[453] + src44[454] + src44[455] + src44[456] + src44[457] + src44[458] + src44[459] + src44[460] + src44[461] + src44[462] + src44[463] + src44[464] + src44[465] + src44[466] + src44[467] + src44[468] + src44[469] + src44[470] + src44[471] + src44[472] + src44[473] + src44[474] + src44[475] + src44[476] + src44[477] + src44[478] + src44[479] + src44[480] + src44[481] + src44[482] + src44[483] + src44[484] + src44[485])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15] + src45[16] + src45[17] + src45[18] + src45[19] + src45[20] + src45[21] + src45[22] + src45[23] + src45[24] + src45[25] + src45[26] + src45[27] + src45[28] + src45[29] + src45[30] + src45[31] + src45[32] + src45[33] + src45[34] + src45[35] + src45[36] + src45[37] + src45[38] + src45[39] + src45[40] + src45[41] + src45[42] + src45[43] + src45[44] + src45[45] + src45[46] + src45[47] + src45[48] + src45[49] + src45[50] + src45[51] + src45[52] + src45[53] + src45[54] + src45[55] + src45[56] + src45[57] + src45[58] + src45[59] + src45[60] + src45[61] + src45[62] + src45[63] + src45[64] + src45[65] + src45[66] + src45[67] + src45[68] + src45[69] + src45[70] + src45[71] + src45[72] + src45[73] + src45[74] + src45[75] + src45[76] + src45[77] + src45[78] + src45[79] + src45[80] + src45[81] + src45[82] + src45[83] + src45[84] + src45[85] + src45[86] + src45[87] + src45[88] + src45[89] + src45[90] + src45[91] + src45[92] + src45[93] + src45[94] + src45[95] + src45[96] + src45[97] + src45[98] + src45[99] + src45[100] + src45[101] + src45[102] + src45[103] + src45[104] + src45[105] + src45[106] + src45[107] + src45[108] + src45[109] + src45[110] + src45[111] + src45[112] + src45[113] + src45[114] + src45[115] + src45[116] + src45[117] + src45[118] + src45[119] + src45[120] + src45[121] + src45[122] + src45[123] + src45[124] + src45[125] + src45[126] + src45[127] + src45[128] + src45[129] + src45[130] + src45[131] + src45[132] + src45[133] + src45[134] + src45[135] + src45[136] + src45[137] + src45[138] + src45[139] + src45[140] + src45[141] + src45[142] + src45[143] + src45[144] + src45[145] + src45[146] + src45[147] + src45[148] + src45[149] + src45[150] + src45[151] + src45[152] + src45[153] + src45[154] + src45[155] + src45[156] + src45[157] + src45[158] + src45[159] + src45[160] + src45[161] + src45[162] + src45[163] + src45[164] + src45[165] + src45[166] + src45[167] + src45[168] + src45[169] + src45[170] + src45[171] + src45[172] + src45[173] + src45[174] + src45[175] + src45[176] + src45[177] + src45[178] + src45[179] + src45[180] + src45[181] + src45[182] + src45[183] + src45[184] + src45[185] + src45[186] + src45[187] + src45[188] + src45[189] + src45[190] + src45[191] + src45[192] + src45[193] + src45[194] + src45[195] + src45[196] + src45[197] + src45[198] + src45[199] + src45[200] + src45[201] + src45[202] + src45[203] + src45[204] + src45[205] + src45[206] + src45[207] + src45[208] + src45[209] + src45[210] + src45[211] + src45[212] + src45[213] + src45[214] + src45[215] + src45[216] + src45[217] + src45[218] + src45[219] + src45[220] + src45[221] + src45[222] + src45[223] + src45[224] + src45[225] + src45[226] + src45[227] + src45[228] + src45[229] + src45[230] + src45[231] + src45[232] + src45[233] + src45[234] + src45[235] + src45[236] + src45[237] + src45[238] + src45[239] + src45[240] + src45[241] + src45[242] + src45[243] + src45[244] + src45[245] + src45[246] + src45[247] + src45[248] + src45[249] + src45[250] + src45[251] + src45[252] + src45[253] + src45[254] + src45[255] + src45[256] + src45[257] + src45[258] + src45[259] + src45[260] + src45[261] + src45[262] + src45[263] + src45[264] + src45[265] + src45[266] + src45[267] + src45[268] + src45[269] + src45[270] + src45[271] + src45[272] + src45[273] + src45[274] + src45[275] + src45[276] + src45[277] + src45[278] + src45[279] + src45[280] + src45[281] + src45[282] + src45[283] + src45[284] + src45[285] + src45[286] + src45[287] + src45[288] + src45[289] + src45[290] + src45[291] + src45[292] + src45[293] + src45[294] + src45[295] + src45[296] + src45[297] + src45[298] + src45[299] + src45[300] + src45[301] + src45[302] + src45[303] + src45[304] + src45[305] + src45[306] + src45[307] + src45[308] + src45[309] + src45[310] + src45[311] + src45[312] + src45[313] + src45[314] + src45[315] + src45[316] + src45[317] + src45[318] + src45[319] + src45[320] + src45[321] + src45[322] + src45[323] + src45[324] + src45[325] + src45[326] + src45[327] + src45[328] + src45[329] + src45[330] + src45[331] + src45[332] + src45[333] + src45[334] + src45[335] + src45[336] + src45[337] + src45[338] + src45[339] + src45[340] + src45[341] + src45[342] + src45[343] + src45[344] + src45[345] + src45[346] + src45[347] + src45[348] + src45[349] + src45[350] + src45[351] + src45[352] + src45[353] + src45[354] + src45[355] + src45[356] + src45[357] + src45[358] + src45[359] + src45[360] + src45[361] + src45[362] + src45[363] + src45[364] + src45[365] + src45[366] + src45[367] + src45[368] + src45[369] + src45[370] + src45[371] + src45[372] + src45[373] + src45[374] + src45[375] + src45[376] + src45[377] + src45[378] + src45[379] + src45[380] + src45[381] + src45[382] + src45[383] + src45[384] + src45[385] + src45[386] + src45[387] + src45[388] + src45[389] + src45[390] + src45[391] + src45[392] + src45[393] + src45[394] + src45[395] + src45[396] + src45[397] + src45[398] + src45[399] + src45[400] + src45[401] + src45[402] + src45[403] + src45[404] + src45[405] + src45[406] + src45[407] + src45[408] + src45[409] + src45[410] + src45[411] + src45[412] + src45[413] + src45[414] + src45[415] + src45[416] + src45[417] + src45[418] + src45[419] + src45[420] + src45[421] + src45[422] + src45[423] + src45[424] + src45[425] + src45[426] + src45[427] + src45[428] + src45[429] + src45[430] + src45[431] + src45[432] + src45[433] + src45[434] + src45[435] + src45[436] + src45[437] + src45[438] + src45[439] + src45[440] + src45[441] + src45[442] + src45[443] + src45[444] + src45[445] + src45[446] + src45[447] + src45[448] + src45[449] + src45[450] + src45[451] + src45[452] + src45[453] + src45[454] + src45[455] + src45[456] + src45[457] + src45[458] + src45[459] + src45[460] + src45[461] + src45[462] + src45[463] + src45[464] + src45[465] + src45[466] + src45[467] + src45[468] + src45[469] + src45[470] + src45[471] + src45[472] + src45[473] + src45[474] + src45[475] + src45[476] + src45[477] + src45[478] + src45[479] + src45[480] + src45[481] + src45[482] + src45[483] + src45[484] + src45[485])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14] + src46[15] + src46[16] + src46[17] + src46[18] + src46[19] + src46[20] + src46[21] + src46[22] + src46[23] + src46[24] + src46[25] + src46[26] + src46[27] + src46[28] + src46[29] + src46[30] + src46[31] + src46[32] + src46[33] + src46[34] + src46[35] + src46[36] + src46[37] + src46[38] + src46[39] + src46[40] + src46[41] + src46[42] + src46[43] + src46[44] + src46[45] + src46[46] + src46[47] + src46[48] + src46[49] + src46[50] + src46[51] + src46[52] + src46[53] + src46[54] + src46[55] + src46[56] + src46[57] + src46[58] + src46[59] + src46[60] + src46[61] + src46[62] + src46[63] + src46[64] + src46[65] + src46[66] + src46[67] + src46[68] + src46[69] + src46[70] + src46[71] + src46[72] + src46[73] + src46[74] + src46[75] + src46[76] + src46[77] + src46[78] + src46[79] + src46[80] + src46[81] + src46[82] + src46[83] + src46[84] + src46[85] + src46[86] + src46[87] + src46[88] + src46[89] + src46[90] + src46[91] + src46[92] + src46[93] + src46[94] + src46[95] + src46[96] + src46[97] + src46[98] + src46[99] + src46[100] + src46[101] + src46[102] + src46[103] + src46[104] + src46[105] + src46[106] + src46[107] + src46[108] + src46[109] + src46[110] + src46[111] + src46[112] + src46[113] + src46[114] + src46[115] + src46[116] + src46[117] + src46[118] + src46[119] + src46[120] + src46[121] + src46[122] + src46[123] + src46[124] + src46[125] + src46[126] + src46[127] + src46[128] + src46[129] + src46[130] + src46[131] + src46[132] + src46[133] + src46[134] + src46[135] + src46[136] + src46[137] + src46[138] + src46[139] + src46[140] + src46[141] + src46[142] + src46[143] + src46[144] + src46[145] + src46[146] + src46[147] + src46[148] + src46[149] + src46[150] + src46[151] + src46[152] + src46[153] + src46[154] + src46[155] + src46[156] + src46[157] + src46[158] + src46[159] + src46[160] + src46[161] + src46[162] + src46[163] + src46[164] + src46[165] + src46[166] + src46[167] + src46[168] + src46[169] + src46[170] + src46[171] + src46[172] + src46[173] + src46[174] + src46[175] + src46[176] + src46[177] + src46[178] + src46[179] + src46[180] + src46[181] + src46[182] + src46[183] + src46[184] + src46[185] + src46[186] + src46[187] + src46[188] + src46[189] + src46[190] + src46[191] + src46[192] + src46[193] + src46[194] + src46[195] + src46[196] + src46[197] + src46[198] + src46[199] + src46[200] + src46[201] + src46[202] + src46[203] + src46[204] + src46[205] + src46[206] + src46[207] + src46[208] + src46[209] + src46[210] + src46[211] + src46[212] + src46[213] + src46[214] + src46[215] + src46[216] + src46[217] + src46[218] + src46[219] + src46[220] + src46[221] + src46[222] + src46[223] + src46[224] + src46[225] + src46[226] + src46[227] + src46[228] + src46[229] + src46[230] + src46[231] + src46[232] + src46[233] + src46[234] + src46[235] + src46[236] + src46[237] + src46[238] + src46[239] + src46[240] + src46[241] + src46[242] + src46[243] + src46[244] + src46[245] + src46[246] + src46[247] + src46[248] + src46[249] + src46[250] + src46[251] + src46[252] + src46[253] + src46[254] + src46[255] + src46[256] + src46[257] + src46[258] + src46[259] + src46[260] + src46[261] + src46[262] + src46[263] + src46[264] + src46[265] + src46[266] + src46[267] + src46[268] + src46[269] + src46[270] + src46[271] + src46[272] + src46[273] + src46[274] + src46[275] + src46[276] + src46[277] + src46[278] + src46[279] + src46[280] + src46[281] + src46[282] + src46[283] + src46[284] + src46[285] + src46[286] + src46[287] + src46[288] + src46[289] + src46[290] + src46[291] + src46[292] + src46[293] + src46[294] + src46[295] + src46[296] + src46[297] + src46[298] + src46[299] + src46[300] + src46[301] + src46[302] + src46[303] + src46[304] + src46[305] + src46[306] + src46[307] + src46[308] + src46[309] + src46[310] + src46[311] + src46[312] + src46[313] + src46[314] + src46[315] + src46[316] + src46[317] + src46[318] + src46[319] + src46[320] + src46[321] + src46[322] + src46[323] + src46[324] + src46[325] + src46[326] + src46[327] + src46[328] + src46[329] + src46[330] + src46[331] + src46[332] + src46[333] + src46[334] + src46[335] + src46[336] + src46[337] + src46[338] + src46[339] + src46[340] + src46[341] + src46[342] + src46[343] + src46[344] + src46[345] + src46[346] + src46[347] + src46[348] + src46[349] + src46[350] + src46[351] + src46[352] + src46[353] + src46[354] + src46[355] + src46[356] + src46[357] + src46[358] + src46[359] + src46[360] + src46[361] + src46[362] + src46[363] + src46[364] + src46[365] + src46[366] + src46[367] + src46[368] + src46[369] + src46[370] + src46[371] + src46[372] + src46[373] + src46[374] + src46[375] + src46[376] + src46[377] + src46[378] + src46[379] + src46[380] + src46[381] + src46[382] + src46[383] + src46[384] + src46[385] + src46[386] + src46[387] + src46[388] + src46[389] + src46[390] + src46[391] + src46[392] + src46[393] + src46[394] + src46[395] + src46[396] + src46[397] + src46[398] + src46[399] + src46[400] + src46[401] + src46[402] + src46[403] + src46[404] + src46[405] + src46[406] + src46[407] + src46[408] + src46[409] + src46[410] + src46[411] + src46[412] + src46[413] + src46[414] + src46[415] + src46[416] + src46[417] + src46[418] + src46[419] + src46[420] + src46[421] + src46[422] + src46[423] + src46[424] + src46[425] + src46[426] + src46[427] + src46[428] + src46[429] + src46[430] + src46[431] + src46[432] + src46[433] + src46[434] + src46[435] + src46[436] + src46[437] + src46[438] + src46[439] + src46[440] + src46[441] + src46[442] + src46[443] + src46[444] + src46[445] + src46[446] + src46[447] + src46[448] + src46[449] + src46[450] + src46[451] + src46[452] + src46[453] + src46[454] + src46[455] + src46[456] + src46[457] + src46[458] + src46[459] + src46[460] + src46[461] + src46[462] + src46[463] + src46[464] + src46[465] + src46[466] + src46[467] + src46[468] + src46[469] + src46[470] + src46[471] + src46[472] + src46[473] + src46[474] + src46[475] + src46[476] + src46[477] + src46[478] + src46[479] + src46[480] + src46[481] + src46[482] + src46[483] + src46[484] + src46[485])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13] + src47[14] + src47[15] + src47[16] + src47[17] + src47[18] + src47[19] + src47[20] + src47[21] + src47[22] + src47[23] + src47[24] + src47[25] + src47[26] + src47[27] + src47[28] + src47[29] + src47[30] + src47[31] + src47[32] + src47[33] + src47[34] + src47[35] + src47[36] + src47[37] + src47[38] + src47[39] + src47[40] + src47[41] + src47[42] + src47[43] + src47[44] + src47[45] + src47[46] + src47[47] + src47[48] + src47[49] + src47[50] + src47[51] + src47[52] + src47[53] + src47[54] + src47[55] + src47[56] + src47[57] + src47[58] + src47[59] + src47[60] + src47[61] + src47[62] + src47[63] + src47[64] + src47[65] + src47[66] + src47[67] + src47[68] + src47[69] + src47[70] + src47[71] + src47[72] + src47[73] + src47[74] + src47[75] + src47[76] + src47[77] + src47[78] + src47[79] + src47[80] + src47[81] + src47[82] + src47[83] + src47[84] + src47[85] + src47[86] + src47[87] + src47[88] + src47[89] + src47[90] + src47[91] + src47[92] + src47[93] + src47[94] + src47[95] + src47[96] + src47[97] + src47[98] + src47[99] + src47[100] + src47[101] + src47[102] + src47[103] + src47[104] + src47[105] + src47[106] + src47[107] + src47[108] + src47[109] + src47[110] + src47[111] + src47[112] + src47[113] + src47[114] + src47[115] + src47[116] + src47[117] + src47[118] + src47[119] + src47[120] + src47[121] + src47[122] + src47[123] + src47[124] + src47[125] + src47[126] + src47[127] + src47[128] + src47[129] + src47[130] + src47[131] + src47[132] + src47[133] + src47[134] + src47[135] + src47[136] + src47[137] + src47[138] + src47[139] + src47[140] + src47[141] + src47[142] + src47[143] + src47[144] + src47[145] + src47[146] + src47[147] + src47[148] + src47[149] + src47[150] + src47[151] + src47[152] + src47[153] + src47[154] + src47[155] + src47[156] + src47[157] + src47[158] + src47[159] + src47[160] + src47[161] + src47[162] + src47[163] + src47[164] + src47[165] + src47[166] + src47[167] + src47[168] + src47[169] + src47[170] + src47[171] + src47[172] + src47[173] + src47[174] + src47[175] + src47[176] + src47[177] + src47[178] + src47[179] + src47[180] + src47[181] + src47[182] + src47[183] + src47[184] + src47[185] + src47[186] + src47[187] + src47[188] + src47[189] + src47[190] + src47[191] + src47[192] + src47[193] + src47[194] + src47[195] + src47[196] + src47[197] + src47[198] + src47[199] + src47[200] + src47[201] + src47[202] + src47[203] + src47[204] + src47[205] + src47[206] + src47[207] + src47[208] + src47[209] + src47[210] + src47[211] + src47[212] + src47[213] + src47[214] + src47[215] + src47[216] + src47[217] + src47[218] + src47[219] + src47[220] + src47[221] + src47[222] + src47[223] + src47[224] + src47[225] + src47[226] + src47[227] + src47[228] + src47[229] + src47[230] + src47[231] + src47[232] + src47[233] + src47[234] + src47[235] + src47[236] + src47[237] + src47[238] + src47[239] + src47[240] + src47[241] + src47[242] + src47[243] + src47[244] + src47[245] + src47[246] + src47[247] + src47[248] + src47[249] + src47[250] + src47[251] + src47[252] + src47[253] + src47[254] + src47[255] + src47[256] + src47[257] + src47[258] + src47[259] + src47[260] + src47[261] + src47[262] + src47[263] + src47[264] + src47[265] + src47[266] + src47[267] + src47[268] + src47[269] + src47[270] + src47[271] + src47[272] + src47[273] + src47[274] + src47[275] + src47[276] + src47[277] + src47[278] + src47[279] + src47[280] + src47[281] + src47[282] + src47[283] + src47[284] + src47[285] + src47[286] + src47[287] + src47[288] + src47[289] + src47[290] + src47[291] + src47[292] + src47[293] + src47[294] + src47[295] + src47[296] + src47[297] + src47[298] + src47[299] + src47[300] + src47[301] + src47[302] + src47[303] + src47[304] + src47[305] + src47[306] + src47[307] + src47[308] + src47[309] + src47[310] + src47[311] + src47[312] + src47[313] + src47[314] + src47[315] + src47[316] + src47[317] + src47[318] + src47[319] + src47[320] + src47[321] + src47[322] + src47[323] + src47[324] + src47[325] + src47[326] + src47[327] + src47[328] + src47[329] + src47[330] + src47[331] + src47[332] + src47[333] + src47[334] + src47[335] + src47[336] + src47[337] + src47[338] + src47[339] + src47[340] + src47[341] + src47[342] + src47[343] + src47[344] + src47[345] + src47[346] + src47[347] + src47[348] + src47[349] + src47[350] + src47[351] + src47[352] + src47[353] + src47[354] + src47[355] + src47[356] + src47[357] + src47[358] + src47[359] + src47[360] + src47[361] + src47[362] + src47[363] + src47[364] + src47[365] + src47[366] + src47[367] + src47[368] + src47[369] + src47[370] + src47[371] + src47[372] + src47[373] + src47[374] + src47[375] + src47[376] + src47[377] + src47[378] + src47[379] + src47[380] + src47[381] + src47[382] + src47[383] + src47[384] + src47[385] + src47[386] + src47[387] + src47[388] + src47[389] + src47[390] + src47[391] + src47[392] + src47[393] + src47[394] + src47[395] + src47[396] + src47[397] + src47[398] + src47[399] + src47[400] + src47[401] + src47[402] + src47[403] + src47[404] + src47[405] + src47[406] + src47[407] + src47[408] + src47[409] + src47[410] + src47[411] + src47[412] + src47[413] + src47[414] + src47[415] + src47[416] + src47[417] + src47[418] + src47[419] + src47[420] + src47[421] + src47[422] + src47[423] + src47[424] + src47[425] + src47[426] + src47[427] + src47[428] + src47[429] + src47[430] + src47[431] + src47[432] + src47[433] + src47[434] + src47[435] + src47[436] + src47[437] + src47[438] + src47[439] + src47[440] + src47[441] + src47[442] + src47[443] + src47[444] + src47[445] + src47[446] + src47[447] + src47[448] + src47[449] + src47[450] + src47[451] + src47[452] + src47[453] + src47[454] + src47[455] + src47[456] + src47[457] + src47[458] + src47[459] + src47[460] + src47[461] + src47[462] + src47[463] + src47[464] + src47[465] + src47[466] + src47[467] + src47[468] + src47[469] + src47[470] + src47[471] + src47[472] + src47[473] + src47[474] + src47[475] + src47[476] + src47[477] + src47[478] + src47[479] + src47[480] + src47[481] + src47[482] + src47[483] + src47[484] + src47[485])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12] + src48[13] + src48[14] + src48[15] + src48[16] + src48[17] + src48[18] + src48[19] + src48[20] + src48[21] + src48[22] + src48[23] + src48[24] + src48[25] + src48[26] + src48[27] + src48[28] + src48[29] + src48[30] + src48[31] + src48[32] + src48[33] + src48[34] + src48[35] + src48[36] + src48[37] + src48[38] + src48[39] + src48[40] + src48[41] + src48[42] + src48[43] + src48[44] + src48[45] + src48[46] + src48[47] + src48[48] + src48[49] + src48[50] + src48[51] + src48[52] + src48[53] + src48[54] + src48[55] + src48[56] + src48[57] + src48[58] + src48[59] + src48[60] + src48[61] + src48[62] + src48[63] + src48[64] + src48[65] + src48[66] + src48[67] + src48[68] + src48[69] + src48[70] + src48[71] + src48[72] + src48[73] + src48[74] + src48[75] + src48[76] + src48[77] + src48[78] + src48[79] + src48[80] + src48[81] + src48[82] + src48[83] + src48[84] + src48[85] + src48[86] + src48[87] + src48[88] + src48[89] + src48[90] + src48[91] + src48[92] + src48[93] + src48[94] + src48[95] + src48[96] + src48[97] + src48[98] + src48[99] + src48[100] + src48[101] + src48[102] + src48[103] + src48[104] + src48[105] + src48[106] + src48[107] + src48[108] + src48[109] + src48[110] + src48[111] + src48[112] + src48[113] + src48[114] + src48[115] + src48[116] + src48[117] + src48[118] + src48[119] + src48[120] + src48[121] + src48[122] + src48[123] + src48[124] + src48[125] + src48[126] + src48[127] + src48[128] + src48[129] + src48[130] + src48[131] + src48[132] + src48[133] + src48[134] + src48[135] + src48[136] + src48[137] + src48[138] + src48[139] + src48[140] + src48[141] + src48[142] + src48[143] + src48[144] + src48[145] + src48[146] + src48[147] + src48[148] + src48[149] + src48[150] + src48[151] + src48[152] + src48[153] + src48[154] + src48[155] + src48[156] + src48[157] + src48[158] + src48[159] + src48[160] + src48[161] + src48[162] + src48[163] + src48[164] + src48[165] + src48[166] + src48[167] + src48[168] + src48[169] + src48[170] + src48[171] + src48[172] + src48[173] + src48[174] + src48[175] + src48[176] + src48[177] + src48[178] + src48[179] + src48[180] + src48[181] + src48[182] + src48[183] + src48[184] + src48[185] + src48[186] + src48[187] + src48[188] + src48[189] + src48[190] + src48[191] + src48[192] + src48[193] + src48[194] + src48[195] + src48[196] + src48[197] + src48[198] + src48[199] + src48[200] + src48[201] + src48[202] + src48[203] + src48[204] + src48[205] + src48[206] + src48[207] + src48[208] + src48[209] + src48[210] + src48[211] + src48[212] + src48[213] + src48[214] + src48[215] + src48[216] + src48[217] + src48[218] + src48[219] + src48[220] + src48[221] + src48[222] + src48[223] + src48[224] + src48[225] + src48[226] + src48[227] + src48[228] + src48[229] + src48[230] + src48[231] + src48[232] + src48[233] + src48[234] + src48[235] + src48[236] + src48[237] + src48[238] + src48[239] + src48[240] + src48[241] + src48[242] + src48[243] + src48[244] + src48[245] + src48[246] + src48[247] + src48[248] + src48[249] + src48[250] + src48[251] + src48[252] + src48[253] + src48[254] + src48[255] + src48[256] + src48[257] + src48[258] + src48[259] + src48[260] + src48[261] + src48[262] + src48[263] + src48[264] + src48[265] + src48[266] + src48[267] + src48[268] + src48[269] + src48[270] + src48[271] + src48[272] + src48[273] + src48[274] + src48[275] + src48[276] + src48[277] + src48[278] + src48[279] + src48[280] + src48[281] + src48[282] + src48[283] + src48[284] + src48[285] + src48[286] + src48[287] + src48[288] + src48[289] + src48[290] + src48[291] + src48[292] + src48[293] + src48[294] + src48[295] + src48[296] + src48[297] + src48[298] + src48[299] + src48[300] + src48[301] + src48[302] + src48[303] + src48[304] + src48[305] + src48[306] + src48[307] + src48[308] + src48[309] + src48[310] + src48[311] + src48[312] + src48[313] + src48[314] + src48[315] + src48[316] + src48[317] + src48[318] + src48[319] + src48[320] + src48[321] + src48[322] + src48[323] + src48[324] + src48[325] + src48[326] + src48[327] + src48[328] + src48[329] + src48[330] + src48[331] + src48[332] + src48[333] + src48[334] + src48[335] + src48[336] + src48[337] + src48[338] + src48[339] + src48[340] + src48[341] + src48[342] + src48[343] + src48[344] + src48[345] + src48[346] + src48[347] + src48[348] + src48[349] + src48[350] + src48[351] + src48[352] + src48[353] + src48[354] + src48[355] + src48[356] + src48[357] + src48[358] + src48[359] + src48[360] + src48[361] + src48[362] + src48[363] + src48[364] + src48[365] + src48[366] + src48[367] + src48[368] + src48[369] + src48[370] + src48[371] + src48[372] + src48[373] + src48[374] + src48[375] + src48[376] + src48[377] + src48[378] + src48[379] + src48[380] + src48[381] + src48[382] + src48[383] + src48[384] + src48[385] + src48[386] + src48[387] + src48[388] + src48[389] + src48[390] + src48[391] + src48[392] + src48[393] + src48[394] + src48[395] + src48[396] + src48[397] + src48[398] + src48[399] + src48[400] + src48[401] + src48[402] + src48[403] + src48[404] + src48[405] + src48[406] + src48[407] + src48[408] + src48[409] + src48[410] + src48[411] + src48[412] + src48[413] + src48[414] + src48[415] + src48[416] + src48[417] + src48[418] + src48[419] + src48[420] + src48[421] + src48[422] + src48[423] + src48[424] + src48[425] + src48[426] + src48[427] + src48[428] + src48[429] + src48[430] + src48[431] + src48[432] + src48[433] + src48[434] + src48[435] + src48[436] + src48[437] + src48[438] + src48[439] + src48[440] + src48[441] + src48[442] + src48[443] + src48[444] + src48[445] + src48[446] + src48[447] + src48[448] + src48[449] + src48[450] + src48[451] + src48[452] + src48[453] + src48[454] + src48[455] + src48[456] + src48[457] + src48[458] + src48[459] + src48[460] + src48[461] + src48[462] + src48[463] + src48[464] + src48[465] + src48[466] + src48[467] + src48[468] + src48[469] + src48[470] + src48[471] + src48[472] + src48[473] + src48[474] + src48[475] + src48[476] + src48[477] + src48[478] + src48[479] + src48[480] + src48[481] + src48[482] + src48[483] + src48[484] + src48[485])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11] + src49[12] + src49[13] + src49[14] + src49[15] + src49[16] + src49[17] + src49[18] + src49[19] + src49[20] + src49[21] + src49[22] + src49[23] + src49[24] + src49[25] + src49[26] + src49[27] + src49[28] + src49[29] + src49[30] + src49[31] + src49[32] + src49[33] + src49[34] + src49[35] + src49[36] + src49[37] + src49[38] + src49[39] + src49[40] + src49[41] + src49[42] + src49[43] + src49[44] + src49[45] + src49[46] + src49[47] + src49[48] + src49[49] + src49[50] + src49[51] + src49[52] + src49[53] + src49[54] + src49[55] + src49[56] + src49[57] + src49[58] + src49[59] + src49[60] + src49[61] + src49[62] + src49[63] + src49[64] + src49[65] + src49[66] + src49[67] + src49[68] + src49[69] + src49[70] + src49[71] + src49[72] + src49[73] + src49[74] + src49[75] + src49[76] + src49[77] + src49[78] + src49[79] + src49[80] + src49[81] + src49[82] + src49[83] + src49[84] + src49[85] + src49[86] + src49[87] + src49[88] + src49[89] + src49[90] + src49[91] + src49[92] + src49[93] + src49[94] + src49[95] + src49[96] + src49[97] + src49[98] + src49[99] + src49[100] + src49[101] + src49[102] + src49[103] + src49[104] + src49[105] + src49[106] + src49[107] + src49[108] + src49[109] + src49[110] + src49[111] + src49[112] + src49[113] + src49[114] + src49[115] + src49[116] + src49[117] + src49[118] + src49[119] + src49[120] + src49[121] + src49[122] + src49[123] + src49[124] + src49[125] + src49[126] + src49[127] + src49[128] + src49[129] + src49[130] + src49[131] + src49[132] + src49[133] + src49[134] + src49[135] + src49[136] + src49[137] + src49[138] + src49[139] + src49[140] + src49[141] + src49[142] + src49[143] + src49[144] + src49[145] + src49[146] + src49[147] + src49[148] + src49[149] + src49[150] + src49[151] + src49[152] + src49[153] + src49[154] + src49[155] + src49[156] + src49[157] + src49[158] + src49[159] + src49[160] + src49[161] + src49[162] + src49[163] + src49[164] + src49[165] + src49[166] + src49[167] + src49[168] + src49[169] + src49[170] + src49[171] + src49[172] + src49[173] + src49[174] + src49[175] + src49[176] + src49[177] + src49[178] + src49[179] + src49[180] + src49[181] + src49[182] + src49[183] + src49[184] + src49[185] + src49[186] + src49[187] + src49[188] + src49[189] + src49[190] + src49[191] + src49[192] + src49[193] + src49[194] + src49[195] + src49[196] + src49[197] + src49[198] + src49[199] + src49[200] + src49[201] + src49[202] + src49[203] + src49[204] + src49[205] + src49[206] + src49[207] + src49[208] + src49[209] + src49[210] + src49[211] + src49[212] + src49[213] + src49[214] + src49[215] + src49[216] + src49[217] + src49[218] + src49[219] + src49[220] + src49[221] + src49[222] + src49[223] + src49[224] + src49[225] + src49[226] + src49[227] + src49[228] + src49[229] + src49[230] + src49[231] + src49[232] + src49[233] + src49[234] + src49[235] + src49[236] + src49[237] + src49[238] + src49[239] + src49[240] + src49[241] + src49[242] + src49[243] + src49[244] + src49[245] + src49[246] + src49[247] + src49[248] + src49[249] + src49[250] + src49[251] + src49[252] + src49[253] + src49[254] + src49[255] + src49[256] + src49[257] + src49[258] + src49[259] + src49[260] + src49[261] + src49[262] + src49[263] + src49[264] + src49[265] + src49[266] + src49[267] + src49[268] + src49[269] + src49[270] + src49[271] + src49[272] + src49[273] + src49[274] + src49[275] + src49[276] + src49[277] + src49[278] + src49[279] + src49[280] + src49[281] + src49[282] + src49[283] + src49[284] + src49[285] + src49[286] + src49[287] + src49[288] + src49[289] + src49[290] + src49[291] + src49[292] + src49[293] + src49[294] + src49[295] + src49[296] + src49[297] + src49[298] + src49[299] + src49[300] + src49[301] + src49[302] + src49[303] + src49[304] + src49[305] + src49[306] + src49[307] + src49[308] + src49[309] + src49[310] + src49[311] + src49[312] + src49[313] + src49[314] + src49[315] + src49[316] + src49[317] + src49[318] + src49[319] + src49[320] + src49[321] + src49[322] + src49[323] + src49[324] + src49[325] + src49[326] + src49[327] + src49[328] + src49[329] + src49[330] + src49[331] + src49[332] + src49[333] + src49[334] + src49[335] + src49[336] + src49[337] + src49[338] + src49[339] + src49[340] + src49[341] + src49[342] + src49[343] + src49[344] + src49[345] + src49[346] + src49[347] + src49[348] + src49[349] + src49[350] + src49[351] + src49[352] + src49[353] + src49[354] + src49[355] + src49[356] + src49[357] + src49[358] + src49[359] + src49[360] + src49[361] + src49[362] + src49[363] + src49[364] + src49[365] + src49[366] + src49[367] + src49[368] + src49[369] + src49[370] + src49[371] + src49[372] + src49[373] + src49[374] + src49[375] + src49[376] + src49[377] + src49[378] + src49[379] + src49[380] + src49[381] + src49[382] + src49[383] + src49[384] + src49[385] + src49[386] + src49[387] + src49[388] + src49[389] + src49[390] + src49[391] + src49[392] + src49[393] + src49[394] + src49[395] + src49[396] + src49[397] + src49[398] + src49[399] + src49[400] + src49[401] + src49[402] + src49[403] + src49[404] + src49[405] + src49[406] + src49[407] + src49[408] + src49[409] + src49[410] + src49[411] + src49[412] + src49[413] + src49[414] + src49[415] + src49[416] + src49[417] + src49[418] + src49[419] + src49[420] + src49[421] + src49[422] + src49[423] + src49[424] + src49[425] + src49[426] + src49[427] + src49[428] + src49[429] + src49[430] + src49[431] + src49[432] + src49[433] + src49[434] + src49[435] + src49[436] + src49[437] + src49[438] + src49[439] + src49[440] + src49[441] + src49[442] + src49[443] + src49[444] + src49[445] + src49[446] + src49[447] + src49[448] + src49[449] + src49[450] + src49[451] + src49[452] + src49[453] + src49[454] + src49[455] + src49[456] + src49[457] + src49[458] + src49[459] + src49[460] + src49[461] + src49[462] + src49[463] + src49[464] + src49[465] + src49[466] + src49[467] + src49[468] + src49[469] + src49[470] + src49[471] + src49[472] + src49[473] + src49[474] + src49[475] + src49[476] + src49[477] + src49[478] + src49[479] + src49[480] + src49[481] + src49[482] + src49[483] + src49[484] + src49[485])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10] + src50[11] + src50[12] + src50[13] + src50[14] + src50[15] + src50[16] + src50[17] + src50[18] + src50[19] + src50[20] + src50[21] + src50[22] + src50[23] + src50[24] + src50[25] + src50[26] + src50[27] + src50[28] + src50[29] + src50[30] + src50[31] + src50[32] + src50[33] + src50[34] + src50[35] + src50[36] + src50[37] + src50[38] + src50[39] + src50[40] + src50[41] + src50[42] + src50[43] + src50[44] + src50[45] + src50[46] + src50[47] + src50[48] + src50[49] + src50[50] + src50[51] + src50[52] + src50[53] + src50[54] + src50[55] + src50[56] + src50[57] + src50[58] + src50[59] + src50[60] + src50[61] + src50[62] + src50[63] + src50[64] + src50[65] + src50[66] + src50[67] + src50[68] + src50[69] + src50[70] + src50[71] + src50[72] + src50[73] + src50[74] + src50[75] + src50[76] + src50[77] + src50[78] + src50[79] + src50[80] + src50[81] + src50[82] + src50[83] + src50[84] + src50[85] + src50[86] + src50[87] + src50[88] + src50[89] + src50[90] + src50[91] + src50[92] + src50[93] + src50[94] + src50[95] + src50[96] + src50[97] + src50[98] + src50[99] + src50[100] + src50[101] + src50[102] + src50[103] + src50[104] + src50[105] + src50[106] + src50[107] + src50[108] + src50[109] + src50[110] + src50[111] + src50[112] + src50[113] + src50[114] + src50[115] + src50[116] + src50[117] + src50[118] + src50[119] + src50[120] + src50[121] + src50[122] + src50[123] + src50[124] + src50[125] + src50[126] + src50[127] + src50[128] + src50[129] + src50[130] + src50[131] + src50[132] + src50[133] + src50[134] + src50[135] + src50[136] + src50[137] + src50[138] + src50[139] + src50[140] + src50[141] + src50[142] + src50[143] + src50[144] + src50[145] + src50[146] + src50[147] + src50[148] + src50[149] + src50[150] + src50[151] + src50[152] + src50[153] + src50[154] + src50[155] + src50[156] + src50[157] + src50[158] + src50[159] + src50[160] + src50[161] + src50[162] + src50[163] + src50[164] + src50[165] + src50[166] + src50[167] + src50[168] + src50[169] + src50[170] + src50[171] + src50[172] + src50[173] + src50[174] + src50[175] + src50[176] + src50[177] + src50[178] + src50[179] + src50[180] + src50[181] + src50[182] + src50[183] + src50[184] + src50[185] + src50[186] + src50[187] + src50[188] + src50[189] + src50[190] + src50[191] + src50[192] + src50[193] + src50[194] + src50[195] + src50[196] + src50[197] + src50[198] + src50[199] + src50[200] + src50[201] + src50[202] + src50[203] + src50[204] + src50[205] + src50[206] + src50[207] + src50[208] + src50[209] + src50[210] + src50[211] + src50[212] + src50[213] + src50[214] + src50[215] + src50[216] + src50[217] + src50[218] + src50[219] + src50[220] + src50[221] + src50[222] + src50[223] + src50[224] + src50[225] + src50[226] + src50[227] + src50[228] + src50[229] + src50[230] + src50[231] + src50[232] + src50[233] + src50[234] + src50[235] + src50[236] + src50[237] + src50[238] + src50[239] + src50[240] + src50[241] + src50[242] + src50[243] + src50[244] + src50[245] + src50[246] + src50[247] + src50[248] + src50[249] + src50[250] + src50[251] + src50[252] + src50[253] + src50[254] + src50[255] + src50[256] + src50[257] + src50[258] + src50[259] + src50[260] + src50[261] + src50[262] + src50[263] + src50[264] + src50[265] + src50[266] + src50[267] + src50[268] + src50[269] + src50[270] + src50[271] + src50[272] + src50[273] + src50[274] + src50[275] + src50[276] + src50[277] + src50[278] + src50[279] + src50[280] + src50[281] + src50[282] + src50[283] + src50[284] + src50[285] + src50[286] + src50[287] + src50[288] + src50[289] + src50[290] + src50[291] + src50[292] + src50[293] + src50[294] + src50[295] + src50[296] + src50[297] + src50[298] + src50[299] + src50[300] + src50[301] + src50[302] + src50[303] + src50[304] + src50[305] + src50[306] + src50[307] + src50[308] + src50[309] + src50[310] + src50[311] + src50[312] + src50[313] + src50[314] + src50[315] + src50[316] + src50[317] + src50[318] + src50[319] + src50[320] + src50[321] + src50[322] + src50[323] + src50[324] + src50[325] + src50[326] + src50[327] + src50[328] + src50[329] + src50[330] + src50[331] + src50[332] + src50[333] + src50[334] + src50[335] + src50[336] + src50[337] + src50[338] + src50[339] + src50[340] + src50[341] + src50[342] + src50[343] + src50[344] + src50[345] + src50[346] + src50[347] + src50[348] + src50[349] + src50[350] + src50[351] + src50[352] + src50[353] + src50[354] + src50[355] + src50[356] + src50[357] + src50[358] + src50[359] + src50[360] + src50[361] + src50[362] + src50[363] + src50[364] + src50[365] + src50[366] + src50[367] + src50[368] + src50[369] + src50[370] + src50[371] + src50[372] + src50[373] + src50[374] + src50[375] + src50[376] + src50[377] + src50[378] + src50[379] + src50[380] + src50[381] + src50[382] + src50[383] + src50[384] + src50[385] + src50[386] + src50[387] + src50[388] + src50[389] + src50[390] + src50[391] + src50[392] + src50[393] + src50[394] + src50[395] + src50[396] + src50[397] + src50[398] + src50[399] + src50[400] + src50[401] + src50[402] + src50[403] + src50[404] + src50[405] + src50[406] + src50[407] + src50[408] + src50[409] + src50[410] + src50[411] + src50[412] + src50[413] + src50[414] + src50[415] + src50[416] + src50[417] + src50[418] + src50[419] + src50[420] + src50[421] + src50[422] + src50[423] + src50[424] + src50[425] + src50[426] + src50[427] + src50[428] + src50[429] + src50[430] + src50[431] + src50[432] + src50[433] + src50[434] + src50[435] + src50[436] + src50[437] + src50[438] + src50[439] + src50[440] + src50[441] + src50[442] + src50[443] + src50[444] + src50[445] + src50[446] + src50[447] + src50[448] + src50[449] + src50[450] + src50[451] + src50[452] + src50[453] + src50[454] + src50[455] + src50[456] + src50[457] + src50[458] + src50[459] + src50[460] + src50[461] + src50[462] + src50[463] + src50[464] + src50[465] + src50[466] + src50[467] + src50[468] + src50[469] + src50[470] + src50[471] + src50[472] + src50[473] + src50[474] + src50[475] + src50[476] + src50[477] + src50[478] + src50[479] + src50[480] + src50[481] + src50[482] + src50[483] + src50[484] + src50[485])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9] + src51[10] + src51[11] + src51[12] + src51[13] + src51[14] + src51[15] + src51[16] + src51[17] + src51[18] + src51[19] + src51[20] + src51[21] + src51[22] + src51[23] + src51[24] + src51[25] + src51[26] + src51[27] + src51[28] + src51[29] + src51[30] + src51[31] + src51[32] + src51[33] + src51[34] + src51[35] + src51[36] + src51[37] + src51[38] + src51[39] + src51[40] + src51[41] + src51[42] + src51[43] + src51[44] + src51[45] + src51[46] + src51[47] + src51[48] + src51[49] + src51[50] + src51[51] + src51[52] + src51[53] + src51[54] + src51[55] + src51[56] + src51[57] + src51[58] + src51[59] + src51[60] + src51[61] + src51[62] + src51[63] + src51[64] + src51[65] + src51[66] + src51[67] + src51[68] + src51[69] + src51[70] + src51[71] + src51[72] + src51[73] + src51[74] + src51[75] + src51[76] + src51[77] + src51[78] + src51[79] + src51[80] + src51[81] + src51[82] + src51[83] + src51[84] + src51[85] + src51[86] + src51[87] + src51[88] + src51[89] + src51[90] + src51[91] + src51[92] + src51[93] + src51[94] + src51[95] + src51[96] + src51[97] + src51[98] + src51[99] + src51[100] + src51[101] + src51[102] + src51[103] + src51[104] + src51[105] + src51[106] + src51[107] + src51[108] + src51[109] + src51[110] + src51[111] + src51[112] + src51[113] + src51[114] + src51[115] + src51[116] + src51[117] + src51[118] + src51[119] + src51[120] + src51[121] + src51[122] + src51[123] + src51[124] + src51[125] + src51[126] + src51[127] + src51[128] + src51[129] + src51[130] + src51[131] + src51[132] + src51[133] + src51[134] + src51[135] + src51[136] + src51[137] + src51[138] + src51[139] + src51[140] + src51[141] + src51[142] + src51[143] + src51[144] + src51[145] + src51[146] + src51[147] + src51[148] + src51[149] + src51[150] + src51[151] + src51[152] + src51[153] + src51[154] + src51[155] + src51[156] + src51[157] + src51[158] + src51[159] + src51[160] + src51[161] + src51[162] + src51[163] + src51[164] + src51[165] + src51[166] + src51[167] + src51[168] + src51[169] + src51[170] + src51[171] + src51[172] + src51[173] + src51[174] + src51[175] + src51[176] + src51[177] + src51[178] + src51[179] + src51[180] + src51[181] + src51[182] + src51[183] + src51[184] + src51[185] + src51[186] + src51[187] + src51[188] + src51[189] + src51[190] + src51[191] + src51[192] + src51[193] + src51[194] + src51[195] + src51[196] + src51[197] + src51[198] + src51[199] + src51[200] + src51[201] + src51[202] + src51[203] + src51[204] + src51[205] + src51[206] + src51[207] + src51[208] + src51[209] + src51[210] + src51[211] + src51[212] + src51[213] + src51[214] + src51[215] + src51[216] + src51[217] + src51[218] + src51[219] + src51[220] + src51[221] + src51[222] + src51[223] + src51[224] + src51[225] + src51[226] + src51[227] + src51[228] + src51[229] + src51[230] + src51[231] + src51[232] + src51[233] + src51[234] + src51[235] + src51[236] + src51[237] + src51[238] + src51[239] + src51[240] + src51[241] + src51[242] + src51[243] + src51[244] + src51[245] + src51[246] + src51[247] + src51[248] + src51[249] + src51[250] + src51[251] + src51[252] + src51[253] + src51[254] + src51[255] + src51[256] + src51[257] + src51[258] + src51[259] + src51[260] + src51[261] + src51[262] + src51[263] + src51[264] + src51[265] + src51[266] + src51[267] + src51[268] + src51[269] + src51[270] + src51[271] + src51[272] + src51[273] + src51[274] + src51[275] + src51[276] + src51[277] + src51[278] + src51[279] + src51[280] + src51[281] + src51[282] + src51[283] + src51[284] + src51[285] + src51[286] + src51[287] + src51[288] + src51[289] + src51[290] + src51[291] + src51[292] + src51[293] + src51[294] + src51[295] + src51[296] + src51[297] + src51[298] + src51[299] + src51[300] + src51[301] + src51[302] + src51[303] + src51[304] + src51[305] + src51[306] + src51[307] + src51[308] + src51[309] + src51[310] + src51[311] + src51[312] + src51[313] + src51[314] + src51[315] + src51[316] + src51[317] + src51[318] + src51[319] + src51[320] + src51[321] + src51[322] + src51[323] + src51[324] + src51[325] + src51[326] + src51[327] + src51[328] + src51[329] + src51[330] + src51[331] + src51[332] + src51[333] + src51[334] + src51[335] + src51[336] + src51[337] + src51[338] + src51[339] + src51[340] + src51[341] + src51[342] + src51[343] + src51[344] + src51[345] + src51[346] + src51[347] + src51[348] + src51[349] + src51[350] + src51[351] + src51[352] + src51[353] + src51[354] + src51[355] + src51[356] + src51[357] + src51[358] + src51[359] + src51[360] + src51[361] + src51[362] + src51[363] + src51[364] + src51[365] + src51[366] + src51[367] + src51[368] + src51[369] + src51[370] + src51[371] + src51[372] + src51[373] + src51[374] + src51[375] + src51[376] + src51[377] + src51[378] + src51[379] + src51[380] + src51[381] + src51[382] + src51[383] + src51[384] + src51[385] + src51[386] + src51[387] + src51[388] + src51[389] + src51[390] + src51[391] + src51[392] + src51[393] + src51[394] + src51[395] + src51[396] + src51[397] + src51[398] + src51[399] + src51[400] + src51[401] + src51[402] + src51[403] + src51[404] + src51[405] + src51[406] + src51[407] + src51[408] + src51[409] + src51[410] + src51[411] + src51[412] + src51[413] + src51[414] + src51[415] + src51[416] + src51[417] + src51[418] + src51[419] + src51[420] + src51[421] + src51[422] + src51[423] + src51[424] + src51[425] + src51[426] + src51[427] + src51[428] + src51[429] + src51[430] + src51[431] + src51[432] + src51[433] + src51[434] + src51[435] + src51[436] + src51[437] + src51[438] + src51[439] + src51[440] + src51[441] + src51[442] + src51[443] + src51[444] + src51[445] + src51[446] + src51[447] + src51[448] + src51[449] + src51[450] + src51[451] + src51[452] + src51[453] + src51[454] + src51[455] + src51[456] + src51[457] + src51[458] + src51[459] + src51[460] + src51[461] + src51[462] + src51[463] + src51[464] + src51[465] + src51[466] + src51[467] + src51[468] + src51[469] + src51[470] + src51[471] + src51[472] + src51[473] + src51[474] + src51[475] + src51[476] + src51[477] + src51[478] + src51[479] + src51[480] + src51[481] + src51[482] + src51[483] + src51[484] + src51[485])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8] + src52[9] + src52[10] + src52[11] + src52[12] + src52[13] + src52[14] + src52[15] + src52[16] + src52[17] + src52[18] + src52[19] + src52[20] + src52[21] + src52[22] + src52[23] + src52[24] + src52[25] + src52[26] + src52[27] + src52[28] + src52[29] + src52[30] + src52[31] + src52[32] + src52[33] + src52[34] + src52[35] + src52[36] + src52[37] + src52[38] + src52[39] + src52[40] + src52[41] + src52[42] + src52[43] + src52[44] + src52[45] + src52[46] + src52[47] + src52[48] + src52[49] + src52[50] + src52[51] + src52[52] + src52[53] + src52[54] + src52[55] + src52[56] + src52[57] + src52[58] + src52[59] + src52[60] + src52[61] + src52[62] + src52[63] + src52[64] + src52[65] + src52[66] + src52[67] + src52[68] + src52[69] + src52[70] + src52[71] + src52[72] + src52[73] + src52[74] + src52[75] + src52[76] + src52[77] + src52[78] + src52[79] + src52[80] + src52[81] + src52[82] + src52[83] + src52[84] + src52[85] + src52[86] + src52[87] + src52[88] + src52[89] + src52[90] + src52[91] + src52[92] + src52[93] + src52[94] + src52[95] + src52[96] + src52[97] + src52[98] + src52[99] + src52[100] + src52[101] + src52[102] + src52[103] + src52[104] + src52[105] + src52[106] + src52[107] + src52[108] + src52[109] + src52[110] + src52[111] + src52[112] + src52[113] + src52[114] + src52[115] + src52[116] + src52[117] + src52[118] + src52[119] + src52[120] + src52[121] + src52[122] + src52[123] + src52[124] + src52[125] + src52[126] + src52[127] + src52[128] + src52[129] + src52[130] + src52[131] + src52[132] + src52[133] + src52[134] + src52[135] + src52[136] + src52[137] + src52[138] + src52[139] + src52[140] + src52[141] + src52[142] + src52[143] + src52[144] + src52[145] + src52[146] + src52[147] + src52[148] + src52[149] + src52[150] + src52[151] + src52[152] + src52[153] + src52[154] + src52[155] + src52[156] + src52[157] + src52[158] + src52[159] + src52[160] + src52[161] + src52[162] + src52[163] + src52[164] + src52[165] + src52[166] + src52[167] + src52[168] + src52[169] + src52[170] + src52[171] + src52[172] + src52[173] + src52[174] + src52[175] + src52[176] + src52[177] + src52[178] + src52[179] + src52[180] + src52[181] + src52[182] + src52[183] + src52[184] + src52[185] + src52[186] + src52[187] + src52[188] + src52[189] + src52[190] + src52[191] + src52[192] + src52[193] + src52[194] + src52[195] + src52[196] + src52[197] + src52[198] + src52[199] + src52[200] + src52[201] + src52[202] + src52[203] + src52[204] + src52[205] + src52[206] + src52[207] + src52[208] + src52[209] + src52[210] + src52[211] + src52[212] + src52[213] + src52[214] + src52[215] + src52[216] + src52[217] + src52[218] + src52[219] + src52[220] + src52[221] + src52[222] + src52[223] + src52[224] + src52[225] + src52[226] + src52[227] + src52[228] + src52[229] + src52[230] + src52[231] + src52[232] + src52[233] + src52[234] + src52[235] + src52[236] + src52[237] + src52[238] + src52[239] + src52[240] + src52[241] + src52[242] + src52[243] + src52[244] + src52[245] + src52[246] + src52[247] + src52[248] + src52[249] + src52[250] + src52[251] + src52[252] + src52[253] + src52[254] + src52[255] + src52[256] + src52[257] + src52[258] + src52[259] + src52[260] + src52[261] + src52[262] + src52[263] + src52[264] + src52[265] + src52[266] + src52[267] + src52[268] + src52[269] + src52[270] + src52[271] + src52[272] + src52[273] + src52[274] + src52[275] + src52[276] + src52[277] + src52[278] + src52[279] + src52[280] + src52[281] + src52[282] + src52[283] + src52[284] + src52[285] + src52[286] + src52[287] + src52[288] + src52[289] + src52[290] + src52[291] + src52[292] + src52[293] + src52[294] + src52[295] + src52[296] + src52[297] + src52[298] + src52[299] + src52[300] + src52[301] + src52[302] + src52[303] + src52[304] + src52[305] + src52[306] + src52[307] + src52[308] + src52[309] + src52[310] + src52[311] + src52[312] + src52[313] + src52[314] + src52[315] + src52[316] + src52[317] + src52[318] + src52[319] + src52[320] + src52[321] + src52[322] + src52[323] + src52[324] + src52[325] + src52[326] + src52[327] + src52[328] + src52[329] + src52[330] + src52[331] + src52[332] + src52[333] + src52[334] + src52[335] + src52[336] + src52[337] + src52[338] + src52[339] + src52[340] + src52[341] + src52[342] + src52[343] + src52[344] + src52[345] + src52[346] + src52[347] + src52[348] + src52[349] + src52[350] + src52[351] + src52[352] + src52[353] + src52[354] + src52[355] + src52[356] + src52[357] + src52[358] + src52[359] + src52[360] + src52[361] + src52[362] + src52[363] + src52[364] + src52[365] + src52[366] + src52[367] + src52[368] + src52[369] + src52[370] + src52[371] + src52[372] + src52[373] + src52[374] + src52[375] + src52[376] + src52[377] + src52[378] + src52[379] + src52[380] + src52[381] + src52[382] + src52[383] + src52[384] + src52[385] + src52[386] + src52[387] + src52[388] + src52[389] + src52[390] + src52[391] + src52[392] + src52[393] + src52[394] + src52[395] + src52[396] + src52[397] + src52[398] + src52[399] + src52[400] + src52[401] + src52[402] + src52[403] + src52[404] + src52[405] + src52[406] + src52[407] + src52[408] + src52[409] + src52[410] + src52[411] + src52[412] + src52[413] + src52[414] + src52[415] + src52[416] + src52[417] + src52[418] + src52[419] + src52[420] + src52[421] + src52[422] + src52[423] + src52[424] + src52[425] + src52[426] + src52[427] + src52[428] + src52[429] + src52[430] + src52[431] + src52[432] + src52[433] + src52[434] + src52[435] + src52[436] + src52[437] + src52[438] + src52[439] + src52[440] + src52[441] + src52[442] + src52[443] + src52[444] + src52[445] + src52[446] + src52[447] + src52[448] + src52[449] + src52[450] + src52[451] + src52[452] + src52[453] + src52[454] + src52[455] + src52[456] + src52[457] + src52[458] + src52[459] + src52[460] + src52[461] + src52[462] + src52[463] + src52[464] + src52[465] + src52[466] + src52[467] + src52[468] + src52[469] + src52[470] + src52[471] + src52[472] + src52[473] + src52[474] + src52[475] + src52[476] + src52[477] + src52[478] + src52[479] + src52[480] + src52[481] + src52[482] + src52[483] + src52[484] + src52[485])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7] + src53[8] + src53[9] + src53[10] + src53[11] + src53[12] + src53[13] + src53[14] + src53[15] + src53[16] + src53[17] + src53[18] + src53[19] + src53[20] + src53[21] + src53[22] + src53[23] + src53[24] + src53[25] + src53[26] + src53[27] + src53[28] + src53[29] + src53[30] + src53[31] + src53[32] + src53[33] + src53[34] + src53[35] + src53[36] + src53[37] + src53[38] + src53[39] + src53[40] + src53[41] + src53[42] + src53[43] + src53[44] + src53[45] + src53[46] + src53[47] + src53[48] + src53[49] + src53[50] + src53[51] + src53[52] + src53[53] + src53[54] + src53[55] + src53[56] + src53[57] + src53[58] + src53[59] + src53[60] + src53[61] + src53[62] + src53[63] + src53[64] + src53[65] + src53[66] + src53[67] + src53[68] + src53[69] + src53[70] + src53[71] + src53[72] + src53[73] + src53[74] + src53[75] + src53[76] + src53[77] + src53[78] + src53[79] + src53[80] + src53[81] + src53[82] + src53[83] + src53[84] + src53[85] + src53[86] + src53[87] + src53[88] + src53[89] + src53[90] + src53[91] + src53[92] + src53[93] + src53[94] + src53[95] + src53[96] + src53[97] + src53[98] + src53[99] + src53[100] + src53[101] + src53[102] + src53[103] + src53[104] + src53[105] + src53[106] + src53[107] + src53[108] + src53[109] + src53[110] + src53[111] + src53[112] + src53[113] + src53[114] + src53[115] + src53[116] + src53[117] + src53[118] + src53[119] + src53[120] + src53[121] + src53[122] + src53[123] + src53[124] + src53[125] + src53[126] + src53[127] + src53[128] + src53[129] + src53[130] + src53[131] + src53[132] + src53[133] + src53[134] + src53[135] + src53[136] + src53[137] + src53[138] + src53[139] + src53[140] + src53[141] + src53[142] + src53[143] + src53[144] + src53[145] + src53[146] + src53[147] + src53[148] + src53[149] + src53[150] + src53[151] + src53[152] + src53[153] + src53[154] + src53[155] + src53[156] + src53[157] + src53[158] + src53[159] + src53[160] + src53[161] + src53[162] + src53[163] + src53[164] + src53[165] + src53[166] + src53[167] + src53[168] + src53[169] + src53[170] + src53[171] + src53[172] + src53[173] + src53[174] + src53[175] + src53[176] + src53[177] + src53[178] + src53[179] + src53[180] + src53[181] + src53[182] + src53[183] + src53[184] + src53[185] + src53[186] + src53[187] + src53[188] + src53[189] + src53[190] + src53[191] + src53[192] + src53[193] + src53[194] + src53[195] + src53[196] + src53[197] + src53[198] + src53[199] + src53[200] + src53[201] + src53[202] + src53[203] + src53[204] + src53[205] + src53[206] + src53[207] + src53[208] + src53[209] + src53[210] + src53[211] + src53[212] + src53[213] + src53[214] + src53[215] + src53[216] + src53[217] + src53[218] + src53[219] + src53[220] + src53[221] + src53[222] + src53[223] + src53[224] + src53[225] + src53[226] + src53[227] + src53[228] + src53[229] + src53[230] + src53[231] + src53[232] + src53[233] + src53[234] + src53[235] + src53[236] + src53[237] + src53[238] + src53[239] + src53[240] + src53[241] + src53[242] + src53[243] + src53[244] + src53[245] + src53[246] + src53[247] + src53[248] + src53[249] + src53[250] + src53[251] + src53[252] + src53[253] + src53[254] + src53[255] + src53[256] + src53[257] + src53[258] + src53[259] + src53[260] + src53[261] + src53[262] + src53[263] + src53[264] + src53[265] + src53[266] + src53[267] + src53[268] + src53[269] + src53[270] + src53[271] + src53[272] + src53[273] + src53[274] + src53[275] + src53[276] + src53[277] + src53[278] + src53[279] + src53[280] + src53[281] + src53[282] + src53[283] + src53[284] + src53[285] + src53[286] + src53[287] + src53[288] + src53[289] + src53[290] + src53[291] + src53[292] + src53[293] + src53[294] + src53[295] + src53[296] + src53[297] + src53[298] + src53[299] + src53[300] + src53[301] + src53[302] + src53[303] + src53[304] + src53[305] + src53[306] + src53[307] + src53[308] + src53[309] + src53[310] + src53[311] + src53[312] + src53[313] + src53[314] + src53[315] + src53[316] + src53[317] + src53[318] + src53[319] + src53[320] + src53[321] + src53[322] + src53[323] + src53[324] + src53[325] + src53[326] + src53[327] + src53[328] + src53[329] + src53[330] + src53[331] + src53[332] + src53[333] + src53[334] + src53[335] + src53[336] + src53[337] + src53[338] + src53[339] + src53[340] + src53[341] + src53[342] + src53[343] + src53[344] + src53[345] + src53[346] + src53[347] + src53[348] + src53[349] + src53[350] + src53[351] + src53[352] + src53[353] + src53[354] + src53[355] + src53[356] + src53[357] + src53[358] + src53[359] + src53[360] + src53[361] + src53[362] + src53[363] + src53[364] + src53[365] + src53[366] + src53[367] + src53[368] + src53[369] + src53[370] + src53[371] + src53[372] + src53[373] + src53[374] + src53[375] + src53[376] + src53[377] + src53[378] + src53[379] + src53[380] + src53[381] + src53[382] + src53[383] + src53[384] + src53[385] + src53[386] + src53[387] + src53[388] + src53[389] + src53[390] + src53[391] + src53[392] + src53[393] + src53[394] + src53[395] + src53[396] + src53[397] + src53[398] + src53[399] + src53[400] + src53[401] + src53[402] + src53[403] + src53[404] + src53[405] + src53[406] + src53[407] + src53[408] + src53[409] + src53[410] + src53[411] + src53[412] + src53[413] + src53[414] + src53[415] + src53[416] + src53[417] + src53[418] + src53[419] + src53[420] + src53[421] + src53[422] + src53[423] + src53[424] + src53[425] + src53[426] + src53[427] + src53[428] + src53[429] + src53[430] + src53[431] + src53[432] + src53[433] + src53[434] + src53[435] + src53[436] + src53[437] + src53[438] + src53[439] + src53[440] + src53[441] + src53[442] + src53[443] + src53[444] + src53[445] + src53[446] + src53[447] + src53[448] + src53[449] + src53[450] + src53[451] + src53[452] + src53[453] + src53[454] + src53[455] + src53[456] + src53[457] + src53[458] + src53[459] + src53[460] + src53[461] + src53[462] + src53[463] + src53[464] + src53[465] + src53[466] + src53[467] + src53[468] + src53[469] + src53[470] + src53[471] + src53[472] + src53[473] + src53[474] + src53[475] + src53[476] + src53[477] + src53[478] + src53[479] + src53[480] + src53[481] + src53[482] + src53[483] + src53[484] + src53[485])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6] + src54[7] + src54[8] + src54[9] + src54[10] + src54[11] + src54[12] + src54[13] + src54[14] + src54[15] + src54[16] + src54[17] + src54[18] + src54[19] + src54[20] + src54[21] + src54[22] + src54[23] + src54[24] + src54[25] + src54[26] + src54[27] + src54[28] + src54[29] + src54[30] + src54[31] + src54[32] + src54[33] + src54[34] + src54[35] + src54[36] + src54[37] + src54[38] + src54[39] + src54[40] + src54[41] + src54[42] + src54[43] + src54[44] + src54[45] + src54[46] + src54[47] + src54[48] + src54[49] + src54[50] + src54[51] + src54[52] + src54[53] + src54[54] + src54[55] + src54[56] + src54[57] + src54[58] + src54[59] + src54[60] + src54[61] + src54[62] + src54[63] + src54[64] + src54[65] + src54[66] + src54[67] + src54[68] + src54[69] + src54[70] + src54[71] + src54[72] + src54[73] + src54[74] + src54[75] + src54[76] + src54[77] + src54[78] + src54[79] + src54[80] + src54[81] + src54[82] + src54[83] + src54[84] + src54[85] + src54[86] + src54[87] + src54[88] + src54[89] + src54[90] + src54[91] + src54[92] + src54[93] + src54[94] + src54[95] + src54[96] + src54[97] + src54[98] + src54[99] + src54[100] + src54[101] + src54[102] + src54[103] + src54[104] + src54[105] + src54[106] + src54[107] + src54[108] + src54[109] + src54[110] + src54[111] + src54[112] + src54[113] + src54[114] + src54[115] + src54[116] + src54[117] + src54[118] + src54[119] + src54[120] + src54[121] + src54[122] + src54[123] + src54[124] + src54[125] + src54[126] + src54[127] + src54[128] + src54[129] + src54[130] + src54[131] + src54[132] + src54[133] + src54[134] + src54[135] + src54[136] + src54[137] + src54[138] + src54[139] + src54[140] + src54[141] + src54[142] + src54[143] + src54[144] + src54[145] + src54[146] + src54[147] + src54[148] + src54[149] + src54[150] + src54[151] + src54[152] + src54[153] + src54[154] + src54[155] + src54[156] + src54[157] + src54[158] + src54[159] + src54[160] + src54[161] + src54[162] + src54[163] + src54[164] + src54[165] + src54[166] + src54[167] + src54[168] + src54[169] + src54[170] + src54[171] + src54[172] + src54[173] + src54[174] + src54[175] + src54[176] + src54[177] + src54[178] + src54[179] + src54[180] + src54[181] + src54[182] + src54[183] + src54[184] + src54[185] + src54[186] + src54[187] + src54[188] + src54[189] + src54[190] + src54[191] + src54[192] + src54[193] + src54[194] + src54[195] + src54[196] + src54[197] + src54[198] + src54[199] + src54[200] + src54[201] + src54[202] + src54[203] + src54[204] + src54[205] + src54[206] + src54[207] + src54[208] + src54[209] + src54[210] + src54[211] + src54[212] + src54[213] + src54[214] + src54[215] + src54[216] + src54[217] + src54[218] + src54[219] + src54[220] + src54[221] + src54[222] + src54[223] + src54[224] + src54[225] + src54[226] + src54[227] + src54[228] + src54[229] + src54[230] + src54[231] + src54[232] + src54[233] + src54[234] + src54[235] + src54[236] + src54[237] + src54[238] + src54[239] + src54[240] + src54[241] + src54[242] + src54[243] + src54[244] + src54[245] + src54[246] + src54[247] + src54[248] + src54[249] + src54[250] + src54[251] + src54[252] + src54[253] + src54[254] + src54[255] + src54[256] + src54[257] + src54[258] + src54[259] + src54[260] + src54[261] + src54[262] + src54[263] + src54[264] + src54[265] + src54[266] + src54[267] + src54[268] + src54[269] + src54[270] + src54[271] + src54[272] + src54[273] + src54[274] + src54[275] + src54[276] + src54[277] + src54[278] + src54[279] + src54[280] + src54[281] + src54[282] + src54[283] + src54[284] + src54[285] + src54[286] + src54[287] + src54[288] + src54[289] + src54[290] + src54[291] + src54[292] + src54[293] + src54[294] + src54[295] + src54[296] + src54[297] + src54[298] + src54[299] + src54[300] + src54[301] + src54[302] + src54[303] + src54[304] + src54[305] + src54[306] + src54[307] + src54[308] + src54[309] + src54[310] + src54[311] + src54[312] + src54[313] + src54[314] + src54[315] + src54[316] + src54[317] + src54[318] + src54[319] + src54[320] + src54[321] + src54[322] + src54[323] + src54[324] + src54[325] + src54[326] + src54[327] + src54[328] + src54[329] + src54[330] + src54[331] + src54[332] + src54[333] + src54[334] + src54[335] + src54[336] + src54[337] + src54[338] + src54[339] + src54[340] + src54[341] + src54[342] + src54[343] + src54[344] + src54[345] + src54[346] + src54[347] + src54[348] + src54[349] + src54[350] + src54[351] + src54[352] + src54[353] + src54[354] + src54[355] + src54[356] + src54[357] + src54[358] + src54[359] + src54[360] + src54[361] + src54[362] + src54[363] + src54[364] + src54[365] + src54[366] + src54[367] + src54[368] + src54[369] + src54[370] + src54[371] + src54[372] + src54[373] + src54[374] + src54[375] + src54[376] + src54[377] + src54[378] + src54[379] + src54[380] + src54[381] + src54[382] + src54[383] + src54[384] + src54[385] + src54[386] + src54[387] + src54[388] + src54[389] + src54[390] + src54[391] + src54[392] + src54[393] + src54[394] + src54[395] + src54[396] + src54[397] + src54[398] + src54[399] + src54[400] + src54[401] + src54[402] + src54[403] + src54[404] + src54[405] + src54[406] + src54[407] + src54[408] + src54[409] + src54[410] + src54[411] + src54[412] + src54[413] + src54[414] + src54[415] + src54[416] + src54[417] + src54[418] + src54[419] + src54[420] + src54[421] + src54[422] + src54[423] + src54[424] + src54[425] + src54[426] + src54[427] + src54[428] + src54[429] + src54[430] + src54[431] + src54[432] + src54[433] + src54[434] + src54[435] + src54[436] + src54[437] + src54[438] + src54[439] + src54[440] + src54[441] + src54[442] + src54[443] + src54[444] + src54[445] + src54[446] + src54[447] + src54[448] + src54[449] + src54[450] + src54[451] + src54[452] + src54[453] + src54[454] + src54[455] + src54[456] + src54[457] + src54[458] + src54[459] + src54[460] + src54[461] + src54[462] + src54[463] + src54[464] + src54[465] + src54[466] + src54[467] + src54[468] + src54[469] + src54[470] + src54[471] + src54[472] + src54[473] + src54[474] + src54[475] + src54[476] + src54[477] + src54[478] + src54[479] + src54[480] + src54[481] + src54[482] + src54[483] + src54[484] + src54[485])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5] + src55[6] + src55[7] + src55[8] + src55[9] + src55[10] + src55[11] + src55[12] + src55[13] + src55[14] + src55[15] + src55[16] + src55[17] + src55[18] + src55[19] + src55[20] + src55[21] + src55[22] + src55[23] + src55[24] + src55[25] + src55[26] + src55[27] + src55[28] + src55[29] + src55[30] + src55[31] + src55[32] + src55[33] + src55[34] + src55[35] + src55[36] + src55[37] + src55[38] + src55[39] + src55[40] + src55[41] + src55[42] + src55[43] + src55[44] + src55[45] + src55[46] + src55[47] + src55[48] + src55[49] + src55[50] + src55[51] + src55[52] + src55[53] + src55[54] + src55[55] + src55[56] + src55[57] + src55[58] + src55[59] + src55[60] + src55[61] + src55[62] + src55[63] + src55[64] + src55[65] + src55[66] + src55[67] + src55[68] + src55[69] + src55[70] + src55[71] + src55[72] + src55[73] + src55[74] + src55[75] + src55[76] + src55[77] + src55[78] + src55[79] + src55[80] + src55[81] + src55[82] + src55[83] + src55[84] + src55[85] + src55[86] + src55[87] + src55[88] + src55[89] + src55[90] + src55[91] + src55[92] + src55[93] + src55[94] + src55[95] + src55[96] + src55[97] + src55[98] + src55[99] + src55[100] + src55[101] + src55[102] + src55[103] + src55[104] + src55[105] + src55[106] + src55[107] + src55[108] + src55[109] + src55[110] + src55[111] + src55[112] + src55[113] + src55[114] + src55[115] + src55[116] + src55[117] + src55[118] + src55[119] + src55[120] + src55[121] + src55[122] + src55[123] + src55[124] + src55[125] + src55[126] + src55[127] + src55[128] + src55[129] + src55[130] + src55[131] + src55[132] + src55[133] + src55[134] + src55[135] + src55[136] + src55[137] + src55[138] + src55[139] + src55[140] + src55[141] + src55[142] + src55[143] + src55[144] + src55[145] + src55[146] + src55[147] + src55[148] + src55[149] + src55[150] + src55[151] + src55[152] + src55[153] + src55[154] + src55[155] + src55[156] + src55[157] + src55[158] + src55[159] + src55[160] + src55[161] + src55[162] + src55[163] + src55[164] + src55[165] + src55[166] + src55[167] + src55[168] + src55[169] + src55[170] + src55[171] + src55[172] + src55[173] + src55[174] + src55[175] + src55[176] + src55[177] + src55[178] + src55[179] + src55[180] + src55[181] + src55[182] + src55[183] + src55[184] + src55[185] + src55[186] + src55[187] + src55[188] + src55[189] + src55[190] + src55[191] + src55[192] + src55[193] + src55[194] + src55[195] + src55[196] + src55[197] + src55[198] + src55[199] + src55[200] + src55[201] + src55[202] + src55[203] + src55[204] + src55[205] + src55[206] + src55[207] + src55[208] + src55[209] + src55[210] + src55[211] + src55[212] + src55[213] + src55[214] + src55[215] + src55[216] + src55[217] + src55[218] + src55[219] + src55[220] + src55[221] + src55[222] + src55[223] + src55[224] + src55[225] + src55[226] + src55[227] + src55[228] + src55[229] + src55[230] + src55[231] + src55[232] + src55[233] + src55[234] + src55[235] + src55[236] + src55[237] + src55[238] + src55[239] + src55[240] + src55[241] + src55[242] + src55[243] + src55[244] + src55[245] + src55[246] + src55[247] + src55[248] + src55[249] + src55[250] + src55[251] + src55[252] + src55[253] + src55[254] + src55[255] + src55[256] + src55[257] + src55[258] + src55[259] + src55[260] + src55[261] + src55[262] + src55[263] + src55[264] + src55[265] + src55[266] + src55[267] + src55[268] + src55[269] + src55[270] + src55[271] + src55[272] + src55[273] + src55[274] + src55[275] + src55[276] + src55[277] + src55[278] + src55[279] + src55[280] + src55[281] + src55[282] + src55[283] + src55[284] + src55[285] + src55[286] + src55[287] + src55[288] + src55[289] + src55[290] + src55[291] + src55[292] + src55[293] + src55[294] + src55[295] + src55[296] + src55[297] + src55[298] + src55[299] + src55[300] + src55[301] + src55[302] + src55[303] + src55[304] + src55[305] + src55[306] + src55[307] + src55[308] + src55[309] + src55[310] + src55[311] + src55[312] + src55[313] + src55[314] + src55[315] + src55[316] + src55[317] + src55[318] + src55[319] + src55[320] + src55[321] + src55[322] + src55[323] + src55[324] + src55[325] + src55[326] + src55[327] + src55[328] + src55[329] + src55[330] + src55[331] + src55[332] + src55[333] + src55[334] + src55[335] + src55[336] + src55[337] + src55[338] + src55[339] + src55[340] + src55[341] + src55[342] + src55[343] + src55[344] + src55[345] + src55[346] + src55[347] + src55[348] + src55[349] + src55[350] + src55[351] + src55[352] + src55[353] + src55[354] + src55[355] + src55[356] + src55[357] + src55[358] + src55[359] + src55[360] + src55[361] + src55[362] + src55[363] + src55[364] + src55[365] + src55[366] + src55[367] + src55[368] + src55[369] + src55[370] + src55[371] + src55[372] + src55[373] + src55[374] + src55[375] + src55[376] + src55[377] + src55[378] + src55[379] + src55[380] + src55[381] + src55[382] + src55[383] + src55[384] + src55[385] + src55[386] + src55[387] + src55[388] + src55[389] + src55[390] + src55[391] + src55[392] + src55[393] + src55[394] + src55[395] + src55[396] + src55[397] + src55[398] + src55[399] + src55[400] + src55[401] + src55[402] + src55[403] + src55[404] + src55[405] + src55[406] + src55[407] + src55[408] + src55[409] + src55[410] + src55[411] + src55[412] + src55[413] + src55[414] + src55[415] + src55[416] + src55[417] + src55[418] + src55[419] + src55[420] + src55[421] + src55[422] + src55[423] + src55[424] + src55[425] + src55[426] + src55[427] + src55[428] + src55[429] + src55[430] + src55[431] + src55[432] + src55[433] + src55[434] + src55[435] + src55[436] + src55[437] + src55[438] + src55[439] + src55[440] + src55[441] + src55[442] + src55[443] + src55[444] + src55[445] + src55[446] + src55[447] + src55[448] + src55[449] + src55[450] + src55[451] + src55[452] + src55[453] + src55[454] + src55[455] + src55[456] + src55[457] + src55[458] + src55[459] + src55[460] + src55[461] + src55[462] + src55[463] + src55[464] + src55[465] + src55[466] + src55[467] + src55[468] + src55[469] + src55[470] + src55[471] + src55[472] + src55[473] + src55[474] + src55[475] + src55[476] + src55[477] + src55[478] + src55[479] + src55[480] + src55[481] + src55[482] + src55[483] + src55[484] + src55[485])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4] + src56[5] + src56[6] + src56[7] + src56[8] + src56[9] + src56[10] + src56[11] + src56[12] + src56[13] + src56[14] + src56[15] + src56[16] + src56[17] + src56[18] + src56[19] + src56[20] + src56[21] + src56[22] + src56[23] + src56[24] + src56[25] + src56[26] + src56[27] + src56[28] + src56[29] + src56[30] + src56[31] + src56[32] + src56[33] + src56[34] + src56[35] + src56[36] + src56[37] + src56[38] + src56[39] + src56[40] + src56[41] + src56[42] + src56[43] + src56[44] + src56[45] + src56[46] + src56[47] + src56[48] + src56[49] + src56[50] + src56[51] + src56[52] + src56[53] + src56[54] + src56[55] + src56[56] + src56[57] + src56[58] + src56[59] + src56[60] + src56[61] + src56[62] + src56[63] + src56[64] + src56[65] + src56[66] + src56[67] + src56[68] + src56[69] + src56[70] + src56[71] + src56[72] + src56[73] + src56[74] + src56[75] + src56[76] + src56[77] + src56[78] + src56[79] + src56[80] + src56[81] + src56[82] + src56[83] + src56[84] + src56[85] + src56[86] + src56[87] + src56[88] + src56[89] + src56[90] + src56[91] + src56[92] + src56[93] + src56[94] + src56[95] + src56[96] + src56[97] + src56[98] + src56[99] + src56[100] + src56[101] + src56[102] + src56[103] + src56[104] + src56[105] + src56[106] + src56[107] + src56[108] + src56[109] + src56[110] + src56[111] + src56[112] + src56[113] + src56[114] + src56[115] + src56[116] + src56[117] + src56[118] + src56[119] + src56[120] + src56[121] + src56[122] + src56[123] + src56[124] + src56[125] + src56[126] + src56[127] + src56[128] + src56[129] + src56[130] + src56[131] + src56[132] + src56[133] + src56[134] + src56[135] + src56[136] + src56[137] + src56[138] + src56[139] + src56[140] + src56[141] + src56[142] + src56[143] + src56[144] + src56[145] + src56[146] + src56[147] + src56[148] + src56[149] + src56[150] + src56[151] + src56[152] + src56[153] + src56[154] + src56[155] + src56[156] + src56[157] + src56[158] + src56[159] + src56[160] + src56[161] + src56[162] + src56[163] + src56[164] + src56[165] + src56[166] + src56[167] + src56[168] + src56[169] + src56[170] + src56[171] + src56[172] + src56[173] + src56[174] + src56[175] + src56[176] + src56[177] + src56[178] + src56[179] + src56[180] + src56[181] + src56[182] + src56[183] + src56[184] + src56[185] + src56[186] + src56[187] + src56[188] + src56[189] + src56[190] + src56[191] + src56[192] + src56[193] + src56[194] + src56[195] + src56[196] + src56[197] + src56[198] + src56[199] + src56[200] + src56[201] + src56[202] + src56[203] + src56[204] + src56[205] + src56[206] + src56[207] + src56[208] + src56[209] + src56[210] + src56[211] + src56[212] + src56[213] + src56[214] + src56[215] + src56[216] + src56[217] + src56[218] + src56[219] + src56[220] + src56[221] + src56[222] + src56[223] + src56[224] + src56[225] + src56[226] + src56[227] + src56[228] + src56[229] + src56[230] + src56[231] + src56[232] + src56[233] + src56[234] + src56[235] + src56[236] + src56[237] + src56[238] + src56[239] + src56[240] + src56[241] + src56[242] + src56[243] + src56[244] + src56[245] + src56[246] + src56[247] + src56[248] + src56[249] + src56[250] + src56[251] + src56[252] + src56[253] + src56[254] + src56[255] + src56[256] + src56[257] + src56[258] + src56[259] + src56[260] + src56[261] + src56[262] + src56[263] + src56[264] + src56[265] + src56[266] + src56[267] + src56[268] + src56[269] + src56[270] + src56[271] + src56[272] + src56[273] + src56[274] + src56[275] + src56[276] + src56[277] + src56[278] + src56[279] + src56[280] + src56[281] + src56[282] + src56[283] + src56[284] + src56[285] + src56[286] + src56[287] + src56[288] + src56[289] + src56[290] + src56[291] + src56[292] + src56[293] + src56[294] + src56[295] + src56[296] + src56[297] + src56[298] + src56[299] + src56[300] + src56[301] + src56[302] + src56[303] + src56[304] + src56[305] + src56[306] + src56[307] + src56[308] + src56[309] + src56[310] + src56[311] + src56[312] + src56[313] + src56[314] + src56[315] + src56[316] + src56[317] + src56[318] + src56[319] + src56[320] + src56[321] + src56[322] + src56[323] + src56[324] + src56[325] + src56[326] + src56[327] + src56[328] + src56[329] + src56[330] + src56[331] + src56[332] + src56[333] + src56[334] + src56[335] + src56[336] + src56[337] + src56[338] + src56[339] + src56[340] + src56[341] + src56[342] + src56[343] + src56[344] + src56[345] + src56[346] + src56[347] + src56[348] + src56[349] + src56[350] + src56[351] + src56[352] + src56[353] + src56[354] + src56[355] + src56[356] + src56[357] + src56[358] + src56[359] + src56[360] + src56[361] + src56[362] + src56[363] + src56[364] + src56[365] + src56[366] + src56[367] + src56[368] + src56[369] + src56[370] + src56[371] + src56[372] + src56[373] + src56[374] + src56[375] + src56[376] + src56[377] + src56[378] + src56[379] + src56[380] + src56[381] + src56[382] + src56[383] + src56[384] + src56[385] + src56[386] + src56[387] + src56[388] + src56[389] + src56[390] + src56[391] + src56[392] + src56[393] + src56[394] + src56[395] + src56[396] + src56[397] + src56[398] + src56[399] + src56[400] + src56[401] + src56[402] + src56[403] + src56[404] + src56[405] + src56[406] + src56[407] + src56[408] + src56[409] + src56[410] + src56[411] + src56[412] + src56[413] + src56[414] + src56[415] + src56[416] + src56[417] + src56[418] + src56[419] + src56[420] + src56[421] + src56[422] + src56[423] + src56[424] + src56[425] + src56[426] + src56[427] + src56[428] + src56[429] + src56[430] + src56[431] + src56[432] + src56[433] + src56[434] + src56[435] + src56[436] + src56[437] + src56[438] + src56[439] + src56[440] + src56[441] + src56[442] + src56[443] + src56[444] + src56[445] + src56[446] + src56[447] + src56[448] + src56[449] + src56[450] + src56[451] + src56[452] + src56[453] + src56[454] + src56[455] + src56[456] + src56[457] + src56[458] + src56[459] + src56[460] + src56[461] + src56[462] + src56[463] + src56[464] + src56[465] + src56[466] + src56[467] + src56[468] + src56[469] + src56[470] + src56[471] + src56[472] + src56[473] + src56[474] + src56[475] + src56[476] + src56[477] + src56[478] + src56[479] + src56[480] + src56[481] + src56[482] + src56[483] + src56[484] + src56[485])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3] + src57[4] + src57[5] + src57[6] + src57[7] + src57[8] + src57[9] + src57[10] + src57[11] + src57[12] + src57[13] + src57[14] + src57[15] + src57[16] + src57[17] + src57[18] + src57[19] + src57[20] + src57[21] + src57[22] + src57[23] + src57[24] + src57[25] + src57[26] + src57[27] + src57[28] + src57[29] + src57[30] + src57[31] + src57[32] + src57[33] + src57[34] + src57[35] + src57[36] + src57[37] + src57[38] + src57[39] + src57[40] + src57[41] + src57[42] + src57[43] + src57[44] + src57[45] + src57[46] + src57[47] + src57[48] + src57[49] + src57[50] + src57[51] + src57[52] + src57[53] + src57[54] + src57[55] + src57[56] + src57[57] + src57[58] + src57[59] + src57[60] + src57[61] + src57[62] + src57[63] + src57[64] + src57[65] + src57[66] + src57[67] + src57[68] + src57[69] + src57[70] + src57[71] + src57[72] + src57[73] + src57[74] + src57[75] + src57[76] + src57[77] + src57[78] + src57[79] + src57[80] + src57[81] + src57[82] + src57[83] + src57[84] + src57[85] + src57[86] + src57[87] + src57[88] + src57[89] + src57[90] + src57[91] + src57[92] + src57[93] + src57[94] + src57[95] + src57[96] + src57[97] + src57[98] + src57[99] + src57[100] + src57[101] + src57[102] + src57[103] + src57[104] + src57[105] + src57[106] + src57[107] + src57[108] + src57[109] + src57[110] + src57[111] + src57[112] + src57[113] + src57[114] + src57[115] + src57[116] + src57[117] + src57[118] + src57[119] + src57[120] + src57[121] + src57[122] + src57[123] + src57[124] + src57[125] + src57[126] + src57[127] + src57[128] + src57[129] + src57[130] + src57[131] + src57[132] + src57[133] + src57[134] + src57[135] + src57[136] + src57[137] + src57[138] + src57[139] + src57[140] + src57[141] + src57[142] + src57[143] + src57[144] + src57[145] + src57[146] + src57[147] + src57[148] + src57[149] + src57[150] + src57[151] + src57[152] + src57[153] + src57[154] + src57[155] + src57[156] + src57[157] + src57[158] + src57[159] + src57[160] + src57[161] + src57[162] + src57[163] + src57[164] + src57[165] + src57[166] + src57[167] + src57[168] + src57[169] + src57[170] + src57[171] + src57[172] + src57[173] + src57[174] + src57[175] + src57[176] + src57[177] + src57[178] + src57[179] + src57[180] + src57[181] + src57[182] + src57[183] + src57[184] + src57[185] + src57[186] + src57[187] + src57[188] + src57[189] + src57[190] + src57[191] + src57[192] + src57[193] + src57[194] + src57[195] + src57[196] + src57[197] + src57[198] + src57[199] + src57[200] + src57[201] + src57[202] + src57[203] + src57[204] + src57[205] + src57[206] + src57[207] + src57[208] + src57[209] + src57[210] + src57[211] + src57[212] + src57[213] + src57[214] + src57[215] + src57[216] + src57[217] + src57[218] + src57[219] + src57[220] + src57[221] + src57[222] + src57[223] + src57[224] + src57[225] + src57[226] + src57[227] + src57[228] + src57[229] + src57[230] + src57[231] + src57[232] + src57[233] + src57[234] + src57[235] + src57[236] + src57[237] + src57[238] + src57[239] + src57[240] + src57[241] + src57[242] + src57[243] + src57[244] + src57[245] + src57[246] + src57[247] + src57[248] + src57[249] + src57[250] + src57[251] + src57[252] + src57[253] + src57[254] + src57[255] + src57[256] + src57[257] + src57[258] + src57[259] + src57[260] + src57[261] + src57[262] + src57[263] + src57[264] + src57[265] + src57[266] + src57[267] + src57[268] + src57[269] + src57[270] + src57[271] + src57[272] + src57[273] + src57[274] + src57[275] + src57[276] + src57[277] + src57[278] + src57[279] + src57[280] + src57[281] + src57[282] + src57[283] + src57[284] + src57[285] + src57[286] + src57[287] + src57[288] + src57[289] + src57[290] + src57[291] + src57[292] + src57[293] + src57[294] + src57[295] + src57[296] + src57[297] + src57[298] + src57[299] + src57[300] + src57[301] + src57[302] + src57[303] + src57[304] + src57[305] + src57[306] + src57[307] + src57[308] + src57[309] + src57[310] + src57[311] + src57[312] + src57[313] + src57[314] + src57[315] + src57[316] + src57[317] + src57[318] + src57[319] + src57[320] + src57[321] + src57[322] + src57[323] + src57[324] + src57[325] + src57[326] + src57[327] + src57[328] + src57[329] + src57[330] + src57[331] + src57[332] + src57[333] + src57[334] + src57[335] + src57[336] + src57[337] + src57[338] + src57[339] + src57[340] + src57[341] + src57[342] + src57[343] + src57[344] + src57[345] + src57[346] + src57[347] + src57[348] + src57[349] + src57[350] + src57[351] + src57[352] + src57[353] + src57[354] + src57[355] + src57[356] + src57[357] + src57[358] + src57[359] + src57[360] + src57[361] + src57[362] + src57[363] + src57[364] + src57[365] + src57[366] + src57[367] + src57[368] + src57[369] + src57[370] + src57[371] + src57[372] + src57[373] + src57[374] + src57[375] + src57[376] + src57[377] + src57[378] + src57[379] + src57[380] + src57[381] + src57[382] + src57[383] + src57[384] + src57[385] + src57[386] + src57[387] + src57[388] + src57[389] + src57[390] + src57[391] + src57[392] + src57[393] + src57[394] + src57[395] + src57[396] + src57[397] + src57[398] + src57[399] + src57[400] + src57[401] + src57[402] + src57[403] + src57[404] + src57[405] + src57[406] + src57[407] + src57[408] + src57[409] + src57[410] + src57[411] + src57[412] + src57[413] + src57[414] + src57[415] + src57[416] + src57[417] + src57[418] + src57[419] + src57[420] + src57[421] + src57[422] + src57[423] + src57[424] + src57[425] + src57[426] + src57[427] + src57[428] + src57[429] + src57[430] + src57[431] + src57[432] + src57[433] + src57[434] + src57[435] + src57[436] + src57[437] + src57[438] + src57[439] + src57[440] + src57[441] + src57[442] + src57[443] + src57[444] + src57[445] + src57[446] + src57[447] + src57[448] + src57[449] + src57[450] + src57[451] + src57[452] + src57[453] + src57[454] + src57[455] + src57[456] + src57[457] + src57[458] + src57[459] + src57[460] + src57[461] + src57[462] + src57[463] + src57[464] + src57[465] + src57[466] + src57[467] + src57[468] + src57[469] + src57[470] + src57[471] + src57[472] + src57[473] + src57[474] + src57[475] + src57[476] + src57[477] + src57[478] + src57[479] + src57[480] + src57[481] + src57[482] + src57[483] + src57[484] + src57[485])<<57) + ((src58[0] + src58[1] + src58[2] + src58[3] + src58[4] + src58[5] + src58[6] + src58[7] + src58[8] + src58[9] + src58[10] + src58[11] + src58[12] + src58[13] + src58[14] + src58[15] + src58[16] + src58[17] + src58[18] + src58[19] + src58[20] + src58[21] + src58[22] + src58[23] + src58[24] + src58[25] + src58[26] + src58[27] + src58[28] + src58[29] + src58[30] + src58[31] + src58[32] + src58[33] + src58[34] + src58[35] + src58[36] + src58[37] + src58[38] + src58[39] + src58[40] + src58[41] + src58[42] + src58[43] + src58[44] + src58[45] + src58[46] + src58[47] + src58[48] + src58[49] + src58[50] + src58[51] + src58[52] + src58[53] + src58[54] + src58[55] + src58[56] + src58[57] + src58[58] + src58[59] + src58[60] + src58[61] + src58[62] + src58[63] + src58[64] + src58[65] + src58[66] + src58[67] + src58[68] + src58[69] + src58[70] + src58[71] + src58[72] + src58[73] + src58[74] + src58[75] + src58[76] + src58[77] + src58[78] + src58[79] + src58[80] + src58[81] + src58[82] + src58[83] + src58[84] + src58[85] + src58[86] + src58[87] + src58[88] + src58[89] + src58[90] + src58[91] + src58[92] + src58[93] + src58[94] + src58[95] + src58[96] + src58[97] + src58[98] + src58[99] + src58[100] + src58[101] + src58[102] + src58[103] + src58[104] + src58[105] + src58[106] + src58[107] + src58[108] + src58[109] + src58[110] + src58[111] + src58[112] + src58[113] + src58[114] + src58[115] + src58[116] + src58[117] + src58[118] + src58[119] + src58[120] + src58[121] + src58[122] + src58[123] + src58[124] + src58[125] + src58[126] + src58[127] + src58[128] + src58[129] + src58[130] + src58[131] + src58[132] + src58[133] + src58[134] + src58[135] + src58[136] + src58[137] + src58[138] + src58[139] + src58[140] + src58[141] + src58[142] + src58[143] + src58[144] + src58[145] + src58[146] + src58[147] + src58[148] + src58[149] + src58[150] + src58[151] + src58[152] + src58[153] + src58[154] + src58[155] + src58[156] + src58[157] + src58[158] + src58[159] + src58[160] + src58[161] + src58[162] + src58[163] + src58[164] + src58[165] + src58[166] + src58[167] + src58[168] + src58[169] + src58[170] + src58[171] + src58[172] + src58[173] + src58[174] + src58[175] + src58[176] + src58[177] + src58[178] + src58[179] + src58[180] + src58[181] + src58[182] + src58[183] + src58[184] + src58[185] + src58[186] + src58[187] + src58[188] + src58[189] + src58[190] + src58[191] + src58[192] + src58[193] + src58[194] + src58[195] + src58[196] + src58[197] + src58[198] + src58[199] + src58[200] + src58[201] + src58[202] + src58[203] + src58[204] + src58[205] + src58[206] + src58[207] + src58[208] + src58[209] + src58[210] + src58[211] + src58[212] + src58[213] + src58[214] + src58[215] + src58[216] + src58[217] + src58[218] + src58[219] + src58[220] + src58[221] + src58[222] + src58[223] + src58[224] + src58[225] + src58[226] + src58[227] + src58[228] + src58[229] + src58[230] + src58[231] + src58[232] + src58[233] + src58[234] + src58[235] + src58[236] + src58[237] + src58[238] + src58[239] + src58[240] + src58[241] + src58[242] + src58[243] + src58[244] + src58[245] + src58[246] + src58[247] + src58[248] + src58[249] + src58[250] + src58[251] + src58[252] + src58[253] + src58[254] + src58[255] + src58[256] + src58[257] + src58[258] + src58[259] + src58[260] + src58[261] + src58[262] + src58[263] + src58[264] + src58[265] + src58[266] + src58[267] + src58[268] + src58[269] + src58[270] + src58[271] + src58[272] + src58[273] + src58[274] + src58[275] + src58[276] + src58[277] + src58[278] + src58[279] + src58[280] + src58[281] + src58[282] + src58[283] + src58[284] + src58[285] + src58[286] + src58[287] + src58[288] + src58[289] + src58[290] + src58[291] + src58[292] + src58[293] + src58[294] + src58[295] + src58[296] + src58[297] + src58[298] + src58[299] + src58[300] + src58[301] + src58[302] + src58[303] + src58[304] + src58[305] + src58[306] + src58[307] + src58[308] + src58[309] + src58[310] + src58[311] + src58[312] + src58[313] + src58[314] + src58[315] + src58[316] + src58[317] + src58[318] + src58[319] + src58[320] + src58[321] + src58[322] + src58[323] + src58[324] + src58[325] + src58[326] + src58[327] + src58[328] + src58[329] + src58[330] + src58[331] + src58[332] + src58[333] + src58[334] + src58[335] + src58[336] + src58[337] + src58[338] + src58[339] + src58[340] + src58[341] + src58[342] + src58[343] + src58[344] + src58[345] + src58[346] + src58[347] + src58[348] + src58[349] + src58[350] + src58[351] + src58[352] + src58[353] + src58[354] + src58[355] + src58[356] + src58[357] + src58[358] + src58[359] + src58[360] + src58[361] + src58[362] + src58[363] + src58[364] + src58[365] + src58[366] + src58[367] + src58[368] + src58[369] + src58[370] + src58[371] + src58[372] + src58[373] + src58[374] + src58[375] + src58[376] + src58[377] + src58[378] + src58[379] + src58[380] + src58[381] + src58[382] + src58[383] + src58[384] + src58[385] + src58[386] + src58[387] + src58[388] + src58[389] + src58[390] + src58[391] + src58[392] + src58[393] + src58[394] + src58[395] + src58[396] + src58[397] + src58[398] + src58[399] + src58[400] + src58[401] + src58[402] + src58[403] + src58[404] + src58[405] + src58[406] + src58[407] + src58[408] + src58[409] + src58[410] + src58[411] + src58[412] + src58[413] + src58[414] + src58[415] + src58[416] + src58[417] + src58[418] + src58[419] + src58[420] + src58[421] + src58[422] + src58[423] + src58[424] + src58[425] + src58[426] + src58[427] + src58[428] + src58[429] + src58[430] + src58[431] + src58[432] + src58[433] + src58[434] + src58[435] + src58[436] + src58[437] + src58[438] + src58[439] + src58[440] + src58[441] + src58[442] + src58[443] + src58[444] + src58[445] + src58[446] + src58[447] + src58[448] + src58[449] + src58[450] + src58[451] + src58[452] + src58[453] + src58[454] + src58[455] + src58[456] + src58[457] + src58[458] + src58[459] + src58[460] + src58[461] + src58[462] + src58[463] + src58[464] + src58[465] + src58[466] + src58[467] + src58[468] + src58[469] + src58[470] + src58[471] + src58[472] + src58[473] + src58[474] + src58[475] + src58[476] + src58[477] + src58[478] + src58[479] + src58[480] + src58[481] + src58[482] + src58[483] + src58[484] + src58[485])<<58) + ((src59[0] + src59[1] + src59[2] + src59[3] + src59[4] + src59[5] + src59[6] + src59[7] + src59[8] + src59[9] + src59[10] + src59[11] + src59[12] + src59[13] + src59[14] + src59[15] + src59[16] + src59[17] + src59[18] + src59[19] + src59[20] + src59[21] + src59[22] + src59[23] + src59[24] + src59[25] + src59[26] + src59[27] + src59[28] + src59[29] + src59[30] + src59[31] + src59[32] + src59[33] + src59[34] + src59[35] + src59[36] + src59[37] + src59[38] + src59[39] + src59[40] + src59[41] + src59[42] + src59[43] + src59[44] + src59[45] + src59[46] + src59[47] + src59[48] + src59[49] + src59[50] + src59[51] + src59[52] + src59[53] + src59[54] + src59[55] + src59[56] + src59[57] + src59[58] + src59[59] + src59[60] + src59[61] + src59[62] + src59[63] + src59[64] + src59[65] + src59[66] + src59[67] + src59[68] + src59[69] + src59[70] + src59[71] + src59[72] + src59[73] + src59[74] + src59[75] + src59[76] + src59[77] + src59[78] + src59[79] + src59[80] + src59[81] + src59[82] + src59[83] + src59[84] + src59[85] + src59[86] + src59[87] + src59[88] + src59[89] + src59[90] + src59[91] + src59[92] + src59[93] + src59[94] + src59[95] + src59[96] + src59[97] + src59[98] + src59[99] + src59[100] + src59[101] + src59[102] + src59[103] + src59[104] + src59[105] + src59[106] + src59[107] + src59[108] + src59[109] + src59[110] + src59[111] + src59[112] + src59[113] + src59[114] + src59[115] + src59[116] + src59[117] + src59[118] + src59[119] + src59[120] + src59[121] + src59[122] + src59[123] + src59[124] + src59[125] + src59[126] + src59[127] + src59[128] + src59[129] + src59[130] + src59[131] + src59[132] + src59[133] + src59[134] + src59[135] + src59[136] + src59[137] + src59[138] + src59[139] + src59[140] + src59[141] + src59[142] + src59[143] + src59[144] + src59[145] + src59[146] + src59[147] + src59[148] + src59[149] + src59[150] + src59[151] + src59[152] + src59[153] + src59[154] + src59[155] + src59[156] + src59[157] + src59[158] + src59[159] + src59[160] + src59[161] + src59[162] + src59[163] + src59[164] + src59[165] + src59[166] + src59[167] + src59[168] + src59[169] + src59[170] + src59[171] + src59[172] + src59[173] + src59[174] + src59[175] + src59[176] + src59[177] + src59[178] + src59[179] + src59[180] + src59[181] + src59[182] + src59[183] + src59[184] + src59[185] + src59[186] + src59[187] + src59[188] + src59[189] + src59[190] + src59[191] + src59[192] + src59[193] + src59[194] + src59[195] + src59[196] + src59[197] + src59[198] + src59[199] + src59[200] + src59[201] + src59[202] + src59[203] + src59[204] + src59[205] + src59[206] + src59[207] + src59[208] + src59[209] + src59[210] + src59[211] + src59[212] + src59[213] + src59[214] + src59[215] + src59[216] + src59[217] + src59[218] + src59[219] + src59[220] + src59[221] + src59[222] + src59[223] + src59[224] + src59[225] + src59[226] + src59[227] + src59[228] + src59[229] + src59[230] + src59[231] + src59[232] + src59[233] + src59[234] + src59[235] + src59[236] + src59[237] + src59[238] + src59[239] + src59[240] + src59[241] + src59[242] + src59[243] + src59[244] + src59[245] + src59[246] + src59[247] + src59[248] + src59[249] + src59[250] + src59[251] + src59[252] + src59[253] + src59[254] + src59[255] + src59[256] + src59[257] + src59[258] + src59[259] + src59[260] + src59[261] + src59[262] + src59[263] + src59[264] + src59[265] + src59[266] + src59[267] + src59[268] + src59[269] + src59[270] + src59[271] + src59[272] + src59[273] + src59[274] + src59[275] + src59[276] + src59[277] + src59[278] + src59[279] + src59[280] + src59[281] + src59[282] + src59[283] + src59[284] + src59[285] + src59[286] + src59[287] + src59[288] + src59[289] + src59[290] + src59[291] + src59[292] + src59[293] + src59[294] + src59[295] + src59[296] + src59[297] + src59[298] + src59[299] + src59[300] + src59[301] + src59[302] + src59[303] + src59[304] + src59[305] + src59[306] + src59[307] + src59[308] + src59[309] + src59[310] + src59[311] + src59[312] + src59[313] + src59[314] + src59[315] + src59[316] + src59[317] + src59[318] + src59[319] + src59[320] + src59[321] + src59[322] + src59[323] + src59[324] + src59[325] + src59[326] + src59[327] + src59[328] + src59[329] + src59[330] + src59[331] + src59[332] + src59[333] + src59[334] + src59[335] + src59[336] + src59[337] + src59[338] + src59[339] + src59[340] + src59[341] + src59[342] + src59[343] + src59[344] + src59[345] + src59[346] + src59[347] + src59[348] + src59[349] + src59[350] + src59[351] + src59[352] + src59[353] + src59[354] + src59[355] + src59[356] + src59[357] + src59[358] + src59[359] + src59[360] + src59[361] + src59[362] + src59[363] + src59[364] + src59[365] + src59[366] + src59[367] + src59[368] + src59[369] + src59[370] + src59[371] + src59[372] + src59[373] + src59[374] + src59[375] + src59[376] + src59[377] + src59[378] + src59[379] + src59[380] + src59[381] + src59[382] + src59[383] + src59[384] + src59[385] + src59[386] + src59[387] + src59[388] + src59[389] + src59[390] + src59[391] + src59[392] + src59[393] + src59[394] + src59[395] + src59[396] + src59[397] + src59[398] + src59[399] + src59[400] + src59[401] + src59[402] + src59[403] + src59[404] + src59[405] + src59[406] + src59[407] + src59[408] + src59[409] + src59[410] + src59[411] + src59[412] + src59[413] + src59[414] + src59[415] + src59[416] + src59[417] + src59[418] + src59[419] + src59[420] + src59[421] + src59[422] + src59[423] + src59[424] + src59[425] + src59[426] + src59[427] + src59[428] + src59[429] + src59[430] + src59[431] + src59[432] + src59[433] + src59[434] + src59[435] + src59[436] + src59[437] + src59[438] + src59[439] + src59[440] + src59[441] + src59[442] + src59[443] + src59[444] + src59[445] + src59[446] + src59[447] + src59[448] + src59[449] + src59[450] + src59[451] + src59[452] + src59[453] + src59[454] + src59[455] + src59[456] + src59[457] + src59[458] + src59[459] + src59[460] + src59[461] + src59[462] + src59[463] + src59[464] + src59[465] + src59[466] + src59[467] + src59[468] + src59[469] + src59[470] + src59[471] + src59[472] + src59[473] + src59[474] + src59[475] + src59[476] + src59[477] + src59[478] + src59[479] + src59[480] + src59[481] + src59[482] + src59[483] + src59[484] + src59[485])<<59) + ((src60[0] + src60[1] + src60[2] + src60[3] + src60[4] + src60[5] + src60[6] + src60[7] + src60[8] + src60[9] + src60[10] + src60[11] + src60[12] + src60[13] + src60[14] + src60[15] + src60[16] + src60[17] + src60[18] + src60[19] + src60[20] + src60[21] + src60[22] + src60[23] + src60[24] + src60[25] + src60[26] + src60[27] + src60[28] + src60[29] + src60[30] + src60[31] + src60[32] + src60[33] + src60[34] + src60[35] + src60[36] + src60[37] + src60[38] + src60[39] + src60[40] + src60[41] + src60[42] + src60[43] + src60[44] + src60[45] + src60[46] + src60[47] + src60[48] + src60[49] + src60[50] + src60[51] + src60[52] + src60[53] + src60[54] + src60[55] + src60[56] + src60[57] + src60[58] + src60[59] + src60[60] + src60[61] + src60[62] + src60[63] + src60[64] + src60[65] + src60[66] + src60[67] + src60[68] + src60[69] + src60[70] + src60[71] + src60[72] + src60[73] + src60[74] + src60[75] + src60[76] + src60[77] + src60[78] + src60[79] + src60[80] + src60[81] + src60[82] + src60[83] + src60[84] + src60[85] + src60[86] + src60[87] + src60[88] + src60[89] + src60[90] + src60[91] + src60[92] + src60[93] + src60[94] + src60[95] + src60[96] + src60[97] + src60[98] + src60[99] + src60[100] + src60[101] + src60[102] + src60[103] + src60[104] + src60[105] + src60[106] + src60[107] + src60[108] + src60[109] + src60[110] + src60[111] + src60[112] + src60[113] + src60[114] + src60[115] + src60[116] + src60[117] + src60[118] + src60[119] + src60[120] + src60[121] + src60[122] + src60[123] + src60[124] + src60[125] + src60[126] + src60[127] + src60[128] + src60[129] + src60[130] + src60[131] + src60[132] + src60[133] + src60[134] + src60[135] + src60[136] + src60[137] + src60[138] + src60[139] + src60[140] + src60[141] + src60[142] + src60[143] + src60[144] + src60[145] + src60[146] + src60[147] + src60[148] + src60[149] + src60[150] + src60[151] + src60[152] + src60[153] + src60[154] + src60[155] + src60[156] + src60[157] + src60[158] + src60[159] + src60[160] + src60[161] + src60[162] + src60[163] + src60[164] + src60[165] + src60[166] + src60[167] + src60[168] + src60[169] + src60[170] + src60[171] + src60[172] + src60[173] + src60[174] + src60[175] + src60[176] + src60[177] + src60[178] + src60[179] + src60[180] + src60[181] + src60[182] + src60[183] + src60[184] + src60[185] + src60[186] + src60[187] + src60[188] + src60[189] + src60[190] + src60[191] + src60[192] + src60[193] + src60[194] + src60[195] + src60[196] + src60[197] + src60[198] + src60[199] + src60[200] + src60[201] + src60[202] + src60[203] + src60[204] + src60[205] + src60[206] + src60[207] + src60[208] + src60[209] + src60[210] + src60[211] + src60[212] + src60[213] + src60[214] + src60[215] + src60[216] + src60[217] + src60[218] + src60[219] + src60[220] + src60[221] + src60[222] + src60[223] + src60[224] + src60[225] + src60[226] + src60[227] + src60[228] + src60[229] + src60[230] + src60[231] + src60[232] + src60[233] + src60[234] + src60[235] + src60[236] + src60[237] + src60[238] + src60[239] + src60[240] + src60[241] + src60[242] + src60[243] + src60[244] + src60[245] + src60[246] + src60[247] + src60[248] + src60[249] + src60[250] + src60[251] + src60[252] + src60[253] + src60[254] + src60[255] + src60[256] + src60[257] + src60[258] + src60[259] + src60[260] + src60[261] + src60[262] + src60[263] + src60[264] + src60[265] + src60[266] + src60[267] + src60[268] + src60[269] + src60[270] + src60[271] + src60[272] + src60[273] + src60[274] + src60[275] + src60[276] + src60[277] + src60[278] + src60[279] + src60[280] + src60[281] + src60[282] + src60[283] + src60[284] + src60[285] + src60[286] + src60[287] + src60[288] + src60[289] + src60[290] + src60[291] + src60[292] + src60[293] + src60[294] + src60[295] + src60[296] + src60[297] + src60[298] + src60[299] + src60[300] + src60[301] + src60[302] + src60[303] + src60[304] + src60[305] + src60[306] + src60[307] + src60[308] + src60[309] + src60[310] + src60[311] + src60[312] + src60[313] + src60[314] + src60[315] + src60[316] + src60[317] + src60[318] + src60[319] + src60[320] + src60[321] + src60[322] + src60[323] + src60[324] + src60[325] + src60[326] + src60[327] + src60[328] + src60[329] + src60[330] + src60[331] + src60[332] + src60[333] + src60[334] + src60[335] + src60[336] + src60[337] + src60[338] + src60[339] + src60[340] + src60[341] + src60[342] + src60[343] + src60[344] + src60[345] + src60[346] + src60[347] + src60[348] + src60[349] + src60[350] + src60[351] + src60[352] + src60[353] + src60[354] + src60[355] + src60[356] + src60[357] + src60[358] + src60[359] + src60[360] + src60[361] + src60[362] + src60[363] + src60[364] + src60[365] + src60[366] + src60[367] + src60[368] + src60[369] + src60[370] + src60[371] + src60[372] + src60[373] + src60[374] + src60[375] + src60[376] + src60[377] + src60[378] + src60[379] + src60[380] + src60[381] + src60[382] + src60[383] + src60[384] + src60[385] + src60[386] + src60[387] + src60[388] + src60[389] + src60[390] + src60[391] + src60[392] + src60[393] + src60[394] + src60[395] + src60[396] + src60[397] + src60[398] + src60[399] + src60[400] + src60[401] + src60[402] + src60[403] + src60[404] + src60[405] + src60[406] + src60[407] + src60[408] + src60[409] + src60[410] + src60[411] + src60[412] + src60[413] + src60[414] + src60[415] + src60[416] + src60[417] + src60[418] + src60[419] + src60[420] + src60[421] + src60[422] + src60[423] + src60[424] + src60[425] + src60[426] + src60[427] + src60[428] + src60[429] + src60[430] + src60[431] + src60[432] + src60[433] + src60[434] + src60[435] + src60[436] + src60[437] + src60[438] + src60[439] + src60[440] + src60[441] + src60[442] + src60[443] + src60[444] + src60[445] + src60[446] + src60[447] + src60[448] + src60[449] + src60[450] + src60[451] + src60[452] + src60[453] + src60[454] + src60[455] + src60[456] + src60[457] + src60[458] + src60[459] + src60[460] + src60[461] + src60[462] + src60[463] + src60[464] + src60[465] + src60[466] + src60[467] + src60[468] + src60[469] + src60[470] + src60[471] + src60[472] + src60[473] + src60[474] + src60[475] + src60[476] + src60[477] + src60[478] + src60[479] + src60[480] + src60[481] + src60[482] + src60[483] + src60[484] + src60[485])<<60) + ((src61[0] + src61[1] + src61[2] + src61[3] + src61[4] + src61[5] + src61[6] + src61[7] + src61[8] + src61[9] + src61[10] + src61[11] + src61[12] + src61[13] + src61[14] + src61[15] + src61[16] + src61[17] + src61[18] + src61[19] + src61[20] + src61[21] + src61[22] + src61[23] + src61[24] + src61[25] + src61[26] + src61[27] + src61[28] + src61[29] + src61[30] + src61[31] + src61[32] + src61[33] + src61[34] + src61[35] + src61[36] + src61[37] + src61[38] + src61[39] + src61[40] + src61[41] + src61[42] + src61[43] + src61[44] + src61[45] + src61[46] + src61[47] + src61[48] + src61[49] + src61[50] + src61[51] + src61[52] + src61[53] + src61[54] + src61[55] + src61[56] + src61[57] + src61[58] + src61[59] + src61[60] + src61[61] + src61[62] + src61[63] + src61[64] + src61[65] + src61[66] + src61[67] + src61[68] + src61[69] + src61[70] + src61[71] + src61[72] + src61[73] + src61[74] + src61[75] + src61[76] + src61[77] + src61[78] + src61[79] + src61[80] + src61[81] + src61[82] + src61[83] + src61[84] + src61[85] + src61[86] + src61[87] + src61[88] + src61[89] + src61[90] + src61[91] + src61[92] + src61[93] + src61[94] + src61[95] + src61[96] + src61[97] + src61[98] + src61[99] + src61[100] + src61[101] + src61[102] + src61[103] + src61[104] + src61[105] + src61[106] + src61[107] + src61[108] + src61[109] + src61[110] + src61[111] + src61[112] + src61[113] + src61[114] + src61[115] + src61[116] + src61[117] + src61[118] + src61[119] + src61[120] + src61[121] + src61[122] + src61[123] + src61[124] + src61[125] + src61[126] + src61[127] + src61[128] + src61[129] + src61[130] + src61[131] + src61[132] + src61[133] + src61[134] + src61[135] + src61[136] + src61[137] + src61[138] + src61[139] + src61[140] + src61[141] + src61[142] + src61[143] + src61[144] + src61[145] + src61[146] + src61[147] + src61[148] + src61[149] + src61[150] + src61[151] + src61[152] + src61[153] + src61[154] + src61[155] + src61[156] + src61[157] + src61[158] + src61[159] + src61[160] + src61[161] + src61[162] + src61[163] + src61[164] + src61[165] + src61[166] + src61[167] + src61[168] + src61[169] + src61[170] + src61[171] + src61[172] + src61[173] + src61[174] + src61[175] + src61[176] + src61[177] + src61[178] + src61[179] + src61[180] + src61[181] + src61[182] + src61[183] + src61[184] + src61[185] + src61[186] + src61[187] + src61[188] + src61[189] + src61[190] + src61[191] + src61[192] + src61[193] + src61[194] + src61[195] + src61[196] + src61[197] + src61[198] + src61[199] + src61[200] + src61[201] + src61[202] + src61[203] + src61[204] + src61[205] + src61[206] + src61[207] + src61[208] + src61[209] + src61[210] + src61[211] + src61[212] + src61[213] + src61[214] + src61[215] + src61[216] + src61[217] + src61[218] + src61[219] + src61[220] + src61[221] + src61[222] + src61[223] + src61[224] + src61[225] + src61[226] + src61[227] + src61[228] + src61[229] + src61[230] + src61[231] + src61[232] + src61[233] + src61[234] + src61[235] + src61[236] + src61[237] + src61[238] + src61[239] + src61[240] + src61[241] + src61[242] + src61[243] + src61[244] + src61[245] + src61[246] + src61[247] + src61[248] + src61[249] + src61[250] + src61[251] + src61[252] + src61[253] + src61[254] + src61[255] + src61[256] + src61[257] + src61[258] + src61[259] + src61[260] + src61[261] + src61[262] + src61[263] + src61[264] + src61[265] + src61[266] + src61[267] + src61[268] + src61[269] + src61[270] + src61[271] + src61[272] + src61[273] + src61[274] + src61[275] + src61[276] + src61[277] + src61[278] + src61[279] + src61[280] + src61[281] + src61[282] + src61[283] + src61[284] + src61[285] + src61[286] + src61[287] + src61[288] + src61[289] + src61[290] + src61[291] + src61[292] + src61[293] + src61[294] + src61[295] + src61[296] + src61[297] + src61[298] + src61[299] + src61[300] + src61[301] + src61[302] + src61[303] + src61[304] + src61[305] + src61[306] + src61[307] + src61[308] + src61[309] + src61[310] + src61[311] + src61[312] + src61[313] + src61[314] + src61[315] + src61[316] + src61[317] + src61[318] + src61[319] + src61[320] + src61[321] + src61[322] + src61[323] + src61[324] + src61[325] + src61[326] + src61[327] + src61[328] + src61[329] + src61[330] + src61[331] + src61[332] + src61[333] + src61[334] + src61[335] + src61[336] + src61[337] + src61[338] + src61[339] + src61[340] + src61[341] + src61[342] + src61[343] + src61[344] + src61[345] + src61[346] + src61[347] + src61[348] + src61[349] + src61[350] + src61[351] + src61[352] + src61[353] + src61[354] + src61[355] + src61[356] + src61[357] + src61[358] + src61[359] + src61[360] + src61[361] + src61[362] + src61[363] + src61[364] + src61[365] + src61[366] + src61[367] + src61[368] + src61[369] + src61[370] + src61[371] + src61[372] + src61[373] + src61[374] + src61[375] + src61[376] + src61[377] + src61[378] + src61[379] + src61[380] + src61[381] + src61[382] + src61[383] + src61[384] + src61[385] + src61[386] + src61[387] + src61[388] + src61[389] + src61[390] + src61[391] + src61[392] + src61[393] + src61[394] + src61[395] + src61[396] + src61[397] + src61[398] + src61[399] + src61[400] + src61[401] + src61[402] + src61[403] + src61[404] + src61[405] + src61[406] + src61[407] + src61[408] + src61[409] + src61[410] + src61[411] + src61[412] + src61[413] + src61[414] + src61[415] + src61[416] + src61[417] + src61[418] + src61[419] + src61[420] + src61[421] + src61[422] + src61[423] + src61[424] + src61[425] + src61[426] + src61[427] + src61[428] + src61[429] + src61[430] + src61[431] + src61[432] + src61[433] + src61[434] + src61[435] + src61[436] + src61[437] + src61[438] + src61[439] + src61[440] + src61[441] + src61[442] + src61[443] + src61[444] + src61[445] + src61[446] + src61[447] + src61[448] + src61[449] + src61[450] + src61[451] + src61[452] + src61[453] + src61[454] + src61[455] + src61[456] + src61[457] + src61[458] + src61[459] + src61[460] + src61[461] + src61[462] + src61[463] + src61[464] + src61[465] + src61[466] + src61[467] + src61[468] + src61[469] + src61[470] + src61[471] + src61[472] + src61[473] + src61[474] + src61[475] + src61[476] + src61[477] + src61[478] + src61[479] + src61[480] + src61[481] + src61[482] + src61[483] + src61[484] + src61[485])<<61) + ((src62[0] + src62[1] + src62[2] + src62[3] + src62[4] + src62[5] + src62[6] + src62[7] + src62[8] + src62[9] + src62[10] + src62[11] + src62[12] + src62[13] + src62[14] + src62[15] + src62[16] + src62[17] + src62[18] + src62[19] + src62[20] + src62[21] + src62[22] + src62[23] + src62[24] + src62[25] + src62[26] + src62[27] + src62[28] + src62[29] + src62[30] + src62[31] + src62[32] + src62[33] + src62[34] + src62[35] + src62[36] + src62[37] + src62[38] + src62[39] + src62[40] + src62[41] + src62[42] + src62[43] + src62[44] + src62[45] + src62[46] + src62[47] + src62[48] + src62[49] + src62[50] + src62[51] + src62[52] + src62[53] + src62[54] + src62[55] + src62[56] + src62[57] + src62[58] + src62[59] + src62[60] + src62[61] + src62[62] + src62[63] + src62[64] + src62[65] + src62[66] + src62[67] + src62[68] + src62[69] + src62[70] + src62[71] + src62[72] + src62[73] + src62[74] + src62[75] + src62[76] + src62[77] + src62[78] + src62[79] + src62[80] + src62[81] + src62[82] + src62[83] + src62[84] + src62[85] + src62[86] + src62[87] + src62[88] + src62[89] + src62[90] + src62[91] + src62[92] + src62[93] + src62[94] + src62[95] + src62[96] + src62[97] + src62[98] + src62[99] + src62[100] + src62[101] + src62[102] + src62[103] + src62[104] + src62[105] + src62[106] + src62[107] + src62[108] + src62[109] + src62[110] + src62[111] + src62[112] + src62[113] + src62[114] + src62[115] + src62[116] + src62[117] + src62[118] + src62[119] + src62[120] + src62[121] + src62[122] + src62[123] + src62[124] + src62[125] + src62[126] + src62[127] + src62[128] + src62[129] + src62[130] + src62[131] + src62[132] + src62[133] + src62[134] + src62[135] + src62[136] + src62[137] + src62[138] + src62[139] + src62[140] + src62[141] + src62[142] + src62[143] + src62[144] + src62[145] + src62[146] + src62[147] + src62[148] + src62[149] + src62[150] + src62[151] + src62[152] + src62[153] + src62[154] + src62[155] + src62[156] + src62[157] + src62[158] + src62[159] + src62[160] + src62[161] + src62[162] + src62[163] + src62[164] + src62[165] + src62[166] + src62[167] + src62[168] + src62[169] + src62[170] + src62[171] + src62[172] + src62[173] + src62[174] + src62[175] + src62[176] + src62[177] + src62[178] + src62[179] + src62[180] + src62[181] + src62[182] + src62[183] + src62[184] + src62[185] + src62[186] + src62[187] + src62[188] + src62[189] + src62[190] + src62[191] + src62[192] + src62[193] + src62[194] + src62[195] + src62[196] + src62[197] + src62[198] + src62[199] + src62[200] + src62[201] + src62[202] + src62[203] + src62[204] + src62[205] + src62[206] + src62[207] + src62[208] + src62[209] + src62[210] + src62[211] + src62[212] + src62[213] + src62[214] + src62[215] + src62[216] + src62[217] + src62[218] + src62[219] + src62[220] + src62[221] + src62[222] + src62[223] + src62[224] + src62[225] + src62[226] + src62[227] + src62[228] + src62[229] + src62[230] + src62[231] + src62[232] + src62[233] + src62[234] + src62[235] + src62[236] + src62[237] + src62[238] + src62[239] + src62[240] + src62[241] + src62[242] + src62[243] + src62[244] + src62[245] + src62[246] + src62[247] + src62[248] + src62[249] + src62[250] + src62[251] + src62[252] + src62[253] + src62[254] + src62[255] + src62[256] + src62[257] + src62[258] + src62[259] + src62[260] + src62[261] + src62[262] + src62[263] + src62[264] + src62[265] + src62[266] + src62[267] + src62[268] + src62[269] + src62[270] + src62[271] + src62[272] + src62[273] + src62[274] + src62[275] + src62[276] + src62[277] + src62[278] + src62[279] + src62[280] + src62[281] + src62[282] + src62[283] + src62[284] + src62[285] + src62[286] + src62[287] + src62[288] + src62[289] + src62[290] + src62[291] + src62[292] + src62[293] + src62[294] + src62[295] + src62[296] + src62[297] + src62[298] + src62[299] + src62[300] + src62[301] + src62[302] + src62[303] + src62[304] + src62[305] + src62[306] + src62[307] + src62[308] + src62[309] + src62[310] + src62[311] + src62[312] + src62[313] + src62[314] + src62[315] + src62[316] + src62[317] + src62[318] + src62[319] + src62[320] + src62[321] + src62[322] + src62[323] + src62[324] + src62[325] + src62[326] + src62[327] + src62[328] + src62[329] + src62[330] + src62[331] + src62[332] + src62[333] + src62[334] + src62[335] + src62[336] + src62[337] + src62[338] + src62[339] + src62[340] + src62[341] + src62[342] + src62[343] + src62[344] + src62[345] + src62[346] + src62[347] + src62[348] + src62[349] + src62[350] + src62[351] + src62[352] + src62[353] + src62[354] + src62[355] + src62[356] + src62[357] + src62[358] + src62[359] + src62[360] + src62[361] + src62[362] + src62[363] + src62[364] + src62[365] + src62[366] + src62[367] + src62[368] + src62[369] + src62[370] + src62[371] + src62[372] + src62[373] + src62[374] + src62[375] + src62[376] + src62[377] + src62[378] + src62[379] + src62[380] + src62[381] + src62[382] + src62[383] + src62[384] + src62[385] + src62[386] + src62[387] + src62[388] + src62[389] + src62[390] + src62[391] + src62[392] + src62[393] + src62[394] + src62[395] + src62[396] + src62[397] + src62[398] + src62[399] + src62[400] + src62[401] + src62[402] + src62[403] + src62[404] + src62[405] + src62[406] + src62[407] + src62[408] + src62[409] + src62[410] + src62[411] + src62[412] + src62[413] + src62[414] + src62[415] + src62[416] + src62[417] + src62[418] + src62[419] + src62[420] + src62[421] + src62[422] + src62[423] + src62[424] + src62[425] + src62[426] + src62[427] + src62[428] + src62[429] + src62[430] + src62[431] + src62[432] + src62[433] + src62[434] + src62[435] + src62[436] + src62[437] + src62[438] + src62[439] + src62[440] + src62[441] + src62[442] + src62[443] + src62[444] + src62[445] + src62[446] + src62[447] + src62[448] + src62[449] + src62[450] + src62[451] + src62[452] + src62[453] + src62[454] + src62[455] + src62[456] + src62[457] + src62[458] + src62[459] + src62[460] + src62[461] + src62[462] + src62[463] + src62[464] + src62[465] + src62[466] + src62[467] + src62[468] + src62[469] + src62[470] + src62[471] + src62[472] + src62[473] + src62[474] + src62[475] + src62[476] + src62[477] + src62[478] + src62[479] + src62[480] + src62[481] + src62[482] + src62[483] + src62[484] + src62[485])<<62) + ((src63[0] + src63[1] + src63[2] + src63[3] + src63[4] + src63[5] + src63[6] + src63[7] + src63[8] + src63[9] + src63[10] + src63[11] + src63[12] + src63[13] + src63[14] + src63[15] + src63[16] + src63[17] + src63[18] + src63[19] + src63[20] + src63[21] + src63[22] + src63[23] + src63[24] + src63[25] + src63[26] + src63[27] + src63[28] + src63[29] + src63[30] + src63[31] + src63[32] + src63[33] + src63[34] + src63[35] + src63[36] + src63[37] + src63[38] + src63[39] + src63[40] + src63[41] + src63[42] + src63[43] + src63[44] + src63[45] + src63[46] + src63[47] + src63[48] + src63[49] + src63[50] + src63[51] + src63[52] + src63[53] + src63[54] + src63[55] + src63[56] + src63[57] + src63[58] + src63[59] + src63[60] + src63[61] + src63[62] + src63[63] + src63[64] + src63[65] + src63[66] + src63[67] + src63[68] + src63[69] + src63[70] + src63[71] + src63[72] + src63[73] + src63[74] + src63[75] + src63[76] + src63[77] + src63[78] + src63[79] + src63[80] + src63[81] + src63[82] + src63[83] + src63[84] + src63[85] + src63[86] + src63[87] + src63[88] + src63[89] + src63[90] + src63[91] + src63[92] + src63[93] + src63[94] + src63[95] + src63[96] + src63[97] + src63[98] + src63[99] + src63[100] + src63[101] + src63[102] + src63[103] + src63[104] + src63[105] + src63[106] + src63[107] + src63[108] + src63[109] + src63[110] + src63[111] + src63[112] + src63[113] + src63[114] + src63[115] + src63[116] + src63[117] + src63[118] + src63[119] + src63[120] + src63[121] + src63[122] + src63[123] + src63[124] + src63[125] + src63[126] + src63[127] + src63[128] + src63[129] + src63[130] + src63[131] + src63[132] + src63[133] + src63[134] + src63[135] + src63[136] + src63[137] + src63[138] + src63[139] + src63[140] + src63[141] + src63[142] + src63[143] + src63[144] + src63[145] + src63[146] + src63[147] + src63[148] + src63[149] + src63[150] + src63[151] + src63[152] + src63[153] + src63[154] + src63[155] + src63[156] + src63[157] + src63[158] + src63[159] + src63[160] + src63[161] + src63[162] + src63[163] + src63[164] + src63[165] + src63[166] + src63[167] + src63[168] + src63[169] + src63[170] + src63[171] + src63[172] + src63[173] + src63[174] + src63[175] + src63[176] + src63[177] + src63[178] + src63[179] + src63[180] + src63[181] + src63[182] + src63[183] + src63[184] + src63[185] + src63[186] + src63[187] + src63[188] + src63[189] + src63[190] + src63[191] + src63[192] + src63[193] + src63[194] + src63[195] + src63[196] + src63[197] + src63[198] + src63[199] + src63[200] + src63[201] + src63[202] + src63[203] + src63[204] + src63[205] + src63[206] + src63[207] + src63[208] + src63[209] + src63[210] + src63[211] + src63[212] + src63[213] + src63[214] + src63[215] + src63[216] + src63[217] + src63[218] + src63[219] + src63[220] + src63[221] + src63[222] + src63[223] + src63[224] + src63[225] + src63[226] + src63[227] + src63[228] + src63[229] + src63[230] + src63[231] + src63[232] + src63[233] + src63[234] + src63[235] + src63[236] + src63[237] + src63[238] + src63[239] + src63[240] + src63[241] + src63[242] + src63[243] + src63[244] + src63[245] + src63[246] + src63[247] + src63[248] + src63[249] + src63[250] + src63[251] + src63[252] + src63[253] + src63[254] + src63[255] + src63[256] + src63[257] + src63[258] + src63[259] + src63[260] + src63[261] + src63[262] + src63[263] + src63[264] + src63[265] + src63[266] + src63[267] + src63[268] + src63[269] + src63[270] + src63[271] + src63[272] + src63[273] + src63[274] + src63[275] + src63[276] + src63[277] + src63[278] + src63[279] + src63[280] + src63[281] + src63[282] + src63[283] + src63[284] + src63[285] + src63[286] + src63[287] + src63[288] + src63[289] + src63[290] + src63[291] + src63[292] + src63[293] + src63[294] + src63[295] + src63[296] + src63[297] + src63[298] + src63[299] + src63[300] + src63[301] + src63[302] + src63[303] + src63[304] + src63[305] + src63[306] + src63[307] + src63[308] + src63[309] + src63[310] + src63[311] + src63[312] + src63[313] + src63[314] + src63[315] + src63[316] + src63[317] + src63[318] + src63[319] + src63[320] + src63[321] + src63[322] + src63[323] + src63[324] + src63[325] + src63[326] + src63[327] + src63[328] + src63[329] + src63[330] + src63[331] + src63[332] + src63[333] + src63[334] + src63[335] + src63[336] + src63[337] + src63[338] + src63[339] + src63[340] + src63[341] + src63[342] + src63[343] + src63[344] + src63[345] + src63[346] + src63[347] + src63[348] + src63[349] + src63[350] + src63[351] + src63[352] + src63[353] + src63[354] + src63[355] + src63[356] + src63[357] + src63[358] + src63[359] + src63[360] + src63[361] + src63[362] + src63[363] + src63[364] + src63[365] + src63[366] + src63[367] + src63[368] + src63[369] + src63[370] + src63[371] + src63[372] + src63[373] + src63[374] + src63[375] + src63[376] + src63[377] + src63[378] + src63[379] + src63[380] + src63[381] + src63[382] + src63[383] + src63[384] + src63[385] + src63[386] + src63[387] + src63[388] + src63[389] + src63[390] + src63[391] + src63[392] + src63[393] + src63[394] + src63[395] + src63[396] + src63[397] + src63[398] + src63[399] + src63[400] + src63[401] + src63[402] + src63[403] + src63[404] + src63[405] + src63[406] + src63[407] + src63[408] + src63[409] + src63[410] + src63[411] + src63[412] + src63[413] + src63[414] + src63[415] + src63[416] + src63[417] + src63[418] + src63[419] + src63[420] + src63[421] + src63[422] + src63[423] + src63[424] + src63[425] + src63[426] + src63[427] + src63[428] + src63[429] + src63[430] + src63[431] + src63[432] + src63[433] + src63[434] + src63[435] + src63[436] + src63[437] + src63[438] + src63[439] + src63[440] + src63[441] + src63[442] + src63[443] + src63[444] + src63[445] + src63[446] + src63[447] + src63[448] + src63[449] + src63[450] + src63[451] + src63[452] + src63[453] + src63[454] + src63[455] + src63[456] + src63[457] + src63[458] + src63[459] + src63[460] + src63[461] + src63[462] + src63[463] + src63[464] + src63[465] + src63[466] + src63[467] + src63[468] + src63[469] + src63[470] + src63[471] + src63[472] + src63[473] + src63[474] + src63[475] + src63[476] + src63[477] + src63[478] + src63[479] + src63[480] + src63[481] + src63[482] + src63[483] + src63[484] + src63[485])<<63);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62) + ((dst63[0])<<63) + ((dst64[0])<<64) + ((dst65[0])<<65) + ((dst66[0])<<66) + ((dst67[0])<<67) + ((dst68[0])<<68) + ((dst69[0])<<69) + ((dst70[0])<<70) + ((dst71[0])<<71) + ((dst72[0])<<72);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hb555680f6bd582028342d7df7d29fd98ce0dd5da752bd088b592f4eefd02e94b31589aeeb4fc180e87d13585c3d373987b3e6c01414bd0e9675203a6428cddebada46a176b3e6116b5422fc8833fec7301bc5ab2656b3934d88031e8db318feaa3ede383f3029d73eba0bfd2c24f5c6b46e0dfe290edcdd36d9142378fe074dad9217d08facf0575a8e24c48669f47385488c10c749cf230a7ea01153fc742a6c000eb17911ea660d3223c1d6c5920f74d4e92a776b694e0a71dbb2e3b5e0fd456d4e7b6bf6d937ce413fa6c316a6b8a6c916c15f1a1437c8e0a93aa99a2f23447041ceb942f51fb732cc5520e2e1e1d709fe77c8880ee57b78cce8d5163c1eb01d37e9b0fc8814d56b75e5ef6ec8d13cd299076a7e18219f1825c8e8d0ce038cba4d6a5b356856f7bfbdf63069aee2a2a7d843c2ef90a5ac2c0006e406c651c14a071f0f4b18aa3b20fb8f7eae1d4a4684d6a56551ce23922a3bb5fee51899394439804797eeba2a0b1d310e2893bdf8ea1fd0784945516d14fa7fe1ad096078742f493f49790543298bb677eba95328ac3ba3aae85cd76af69482791103a390fc0855353261c773262c90955693abf86d0b7add28e2da0dba43a2178ebefc167fea122c529650f2da92e4e79dc91703f242cbaa257dab4aa60061a9e1b43344a473ac9e9ab4de2f3b84e84f6275007b4e8c790fd47416ca237ee76e00bac53288e3cd3ced5f2bceafd08392bd098e90b001077f1b7981cb2c8180e75ba1ededd5597e5f9e568119e3d9067a1dae5720070a7b7e6c49863c4906bedc46efa1611a432eef67d4b71558e60d0604c7bfdd3f1837762be5977e188d9461f7a49df967148db1d2b6a9b18c3d884dd765a798f52aa7786b5328ea37438dc0396c9df4846b10f6456f2098c38d68c48a525f65b30576bae46060a929b8d6bc4e531f9a3f68da87b9e6b319ce24f85284e6af6bc7c0e4cd7293d5e4c2b92e030b6634aea3d7d8bb8975347b16a8ccb349e126890a6d30d82bb53a9e97fff1d4c84e266529c614e92758613c9461f1521da0192c47ac557332352c6cf84d3a59a6668ce754c39e60d9d5abc10d2deb08b5fa80abb78b517482c3315831f106834c8d2eef2a8914335fddd7916ced3b139c2ead192bdc881d2d035fc2d5001e9d5ff23fc07f4eff2d4548f6cbbbf8df04924b68eaec7eff0f90a7231500a8b62e6b2fe37dcf3528380f53666697f3c303cf1d73ef7b1787f748c99f2e718c9b26bf6302e91f13dec0b39a8df88fcbb930333c3f8fd0cafba2e0dca1ddc1a8ded1fe5011d7c92a7cb4408248f75b225616fe7872f705d3c8ae8165c578be65229dbac5da9eeb5a51c38266a124a41ab8b3a1570f7020ccdd9ab635acbcd26e7de524dc06433424fe8bb65393b95af86083637ab55ae59cf9e800a14dc5da219e767de9d77acb20f22fe22c85e1edcc05c9f6cf45b6321e6480269d1e1c9c9926def35d5447297680da722462e97011fb7986b6f96492a9496b62492ff94ea59ef0bfcd7488f939e9c293c61c36dc03c0669f910ffcaad715180d90983e1fce967b0655cd0067c6685cec4483e5b5d7390bb8aa9f8fec32bdf37f52647694bcf72ba7d37f778941f97bb25017b06df907861e4b935750a527faf95074ff9353f1317d53978f54f5cb5a2ca81d4b7bc49b1e0143758b1f2c033969ed0b2ee9a20ae246b14efe5c87622ab591bf978456372e96702490141b3f79c5065956b4691f5208cfeca14b0dfc0b1af5d8d3690dc38a42af9c6ce80d0cb3bf89c84ba36914ce3f77beae298ddc4f61a152ea32d70de64530d14d3d576f49105c636df15e644a61a58d0d7855e6ae269dc0be01cf18d2d756dd9a4456d41ab82f3a6271936d3e1f6a5cefc532b67fb1002aef2bde084a705121da066fc45d648958e25f80ad7fb6e08641d1e897bdc7b47d9457e7793641608624f36f65c7b3b6694e0865f9b90ca7b94a0947b6efc0d9ecdddd7fd98707dd5bffd97cf7de02d842b98891f1fc0486edc527439902f1528c31f8c58da497a8cca32477662a0930b883e2c9f87dfa4cd489cd781c48c02d6ead574cceeb6224c1553da5f2dff80479862c7fdd07c0221bd7984de0f953bf6b2f22941898c19aa64b679af92d781f29b9279b0a7fe7d0323a29b12e1364d93a5156d8c10aecbafd8caf92ee2669f7772e645a4255012f5fa448f842a7abbf10e57102bfbbb6461c225ca9f576451d8950c52f4a2742ff27afdc3aaea79a06132ca41300681dccae575bfd9600478298f195ed7a09f30735015cd5ab2039520a65ab0384811b18377281284f5350b6c8967a95a409f530fcfce082752f6614759ac484eecb42b32a41ae7b95c6230af3ecd819b675432e469886fe94f8df254a44d8d901ef649cdfee5957b36904433f851c44f55c5add486635baa15e16a077be61c65d39354ea1fc91d37a6bb1c3c35a7bf53bd9fd6a1024751360d136e13fb39fa0217ea87c126000ec024aaa43285e54c10c8222166a20fc94007ce43239411acc43402c4b09d19f98d644d3ade955f7de7cf82b392233c5fe5da83f25f03f59f9d435f14e8d646b71ccc324eac124c8e9396fe51fd88ab4c2a0d2e148ebde334740474954738cff625cae723bf9f17fe407ea22e86242d13616a651f337e6dcd0cc7f5acff2bec3b6657e1182954876512533c9dfddf5a5647a241ac07e30ce1fa6d661edd96b1a2926a3db691e6ad57b2d400f566d2a26ab84769cb3310ba55e461b6e216b0e821326d0110e2051d3bfda942dabff25532d23dd1c18a8b961552228087b086b69ca84ee5a2f342aca483687af53c1e3c6b7f1e8609ce9c4d787c5aaa071ff4ad6da1c560b6cf4b318d1a55a76d8940474b2c9443809a8294e3a561e1280fa0124e296fa52e1eb5f88b80801f8b09620bd7db4293aca1a608ff6386953e47795995beb0f95dd458ba095bbaba5dea8a70cf3f90edca87c2d5a11d586cadc32b64610ad61c952eb77a1ee4424bbf5c9d3ce7d856b127775ede328ebe0684e571d315bd98dd929903c191d57ef1b4f2d103d1daf7fcf56a7dba58c29277c4a4aa756191d53e14a12182b89231256bb1ac7da8033d33e156172fb6984c622e42f019ac5ea6ffe2e13196bba9b2d0948667e3d81753752e92ddc01ccd1c7624947ad69b24970a561af3abc61e6f9dc3eda5bc842884c8f294c46ff6e41655a61e03c91145ecf0aa7fd11459997d0bebc12258580b77fead782e653734ec74b4122ff5b8b07a37d3d2cdbfdd17f3dcb404f981a718125c83fcf13c51b5962e7c55c3806f3f5d0d1b3e6099563be0f1d77fde615d18cbab5c9408cc4e200c237d9281e817ef4fdeafd6d2d54c3bde0f34fe4094e1af40769abf13fcc121a1b16d89bcf5cc5fbfba1823596db45ac2d6dedd648eb40d971e83ef0eef41a8a7278ddd727a93f10a606d50e33eba1d268bd05f5941b535f276c11e217f4b8a13e1d8517cdf678e573d1ec1680bf91620e1c75e2ca95b53d8efdd24473dea060883dabb1eca2d124306d35a3bb4e090a63d20719450bdf464292c4d0de5f1859637dfd5fccca6853d465004c7cf8b6bd6b2ad39214b641fcc0cfceda8ea5bc2d3011e558124d7fe8a73c416a5c75ba7ce4f670b0b128bd74685d2c1af5bdf428b83850c469a0e3cdda2c374ba36a5653bdf6ca5c99e8befaf07ade47c2cd976b7e73f0c1318c90acd43bf74eecd5f9e0400fe5d1abf553eb17f4c3007fad5e34fd4053d948deefa906154680dcb3fec362e29780fb7de695eef8ed44adde2f17a5de0e0887de425e4a2a8ff7671f686d9f9ba791d78d1a798f1017b062e2e4b75d48021d462adc2215e4b56ab0160f0a0504eebc73874748b90fc330cef66c9a7056d0f39ce284716e86a42989fc5c83a1b814143293b9336ad15a9462a656310a3d83f4973c1528bfae24c5aff524f9d90d675a54bb8323f413bcca4a426db79f82cf8c1e8d99080e02e4e3a33dbb3d38f5d43f5385dd2a990f0b431c2a092c320a58bd810c9f711150bf2c991a917a724462b84e216f576916c3db63ac2218a9e8f2c9ad45977aeb2ee2970f72882370b89612d206b1854aeb1221114f0d4dc87e5ff3f760914f0b40aee46fe88b402c237b78f2fe4f1d8542c44e971a4cc265a6b9690893a43749b053cd9322311670a5ccbe9b240f2b1160621e108a545d3502d7692b7900589fe7723e4a3174eae2424c43bbc34dcae7ae7a1f5c38346a0fa485f60e02c3161cfa0a61dc413e2053bdd31ac1a092726e90952ca2f13dac706a2b13d9c47e9445ec3eaf67b5ac1aa7016a8b0b85d86eff7d66d630d8d057df9027dbe7590cf1bb8adf009e2233f9ffcd2356d70faf9162b1a72d9eff350471ea5f697e86c08526642d56c6e766afe4a3e2ce64a2bbc8baf7aad63102fbb5c5ca98e1981b1c3c9907f22579fe7429596acd82413fcd38bfc5b556e9708bb773ee1b1fce89f0aba947368fd74add45bbb42846ec60ac9ca6e8268b397990096dbe6aa9ae79aa2eb97716edebf48d006f8de4a413c74ace3d8b7c7a1a8a8f4370215eaa03e08403ec01b048d66f067ee7ad79011078ff79fc8f2dad162928710305f12dd2eb9953ad9bb28934b5e8a9596469f1a50f68284869bc970625e050f094531c4db5e3953eabbaa85c9e397c58be022f3e50cbde1ba1c474e6244d7a828303d609ac85b670c7e300dd97430aa560672633248bb79fbb7e2788c60bab8857b2cbed9cf983b7b60cdaa927e1a154547faa8ec7ef209fe1a64e9860b04d9d9fb6300435695f2b5d5b7dc1c26e91b2b547d2d5ea5ede35de5aee03214d7c290a9e0a9e69c7cbfb37a4c9c523d338ade09165b7dccd32bec5b6e1c65741d3ac8f484d7d8dbd8de8e09745f1ec342360b91781487c5ec943468fbebdb142df3719cc18712e7c5f9419ea1e8c79a9bcdd2e76f8779505dfc78c4ccf1890154d01427ded7801401498e3eab66e07889e4e34964811ce0cb3e9896c7db71b8f2ab796bb6f83f8e7ced88eeeff53aa35a091dd207ca51a529a3165ae43d67cb9cf322ab708a67a49b8bd5cc4b7fc355255c0a9f2e6a9ea3540b0c27c64b81432a896d9ee11d1fd3b11f41278fde251ae9b68de7745b52985a3a2647f4724ac4c76d76cea7c93a8a1e8b3f52f7e128e7e3c3a1f2ffdc782c2e6df817f326e57d4f86bfdb4ec096e53a544689e653f32016c38f9f5d4734774a4d5124ccab87c496480519ab6dbd75ee81441102e3d45192b1b610697df06c95ffe1febc0893009ded5d9e1fc9b739272f809097b4d9f9fbd972301dfe65e493a103d7dc16479a244a74df9bd9e2c8876050000bcf14fbb3d0b866bdf96cf33b84c29dbeb315e148c9f9c5c055a313a602b29d4e2081e8492ac55ce9c5375beff2305f4d0cb537125b4025478973960984ba06d630af61e9f198901d9bcb4ed70daee9b1c7eb204bc3e442bc03;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h9b84f72b1d83246344bfac0513203e09c2b01722080ff2f9b96de8cc6b5357f70922022b7e917054045ddeaf098f6748d4dee9076787cd95eb3b52cca25fc3c5088f5918baba24355460671176e75522583c9c8c762cc9160d6df82fa75cd406dcc36c6c7ca57e52619ce3763bfa46648c148e2ac62794ac4266aa28fefd1730c3e38c6b46a2ae34a507c242ec84b29dafe41190ba754a55523a0b1b4ef5f9b9c5bbcfcaaf432585a129e80a1844ffc6fb72585e6a292c083d0a8fbd9c40c41595b3214d15e31b8d93ac3e8a12f9a5141d8f86cd8bad52d75824dcbceac7246369a4f6e51561707b68f04f2d6fb93a73a0831683640bb772bba996af758906c1a3310acd795bf0dc8e90b714f80c2d6f80e1061b52435b8c1fc4dfe5a428682e1033100ff4f57bbdfd9fb47303b0cc8551417534138dee761b2136d3db0b7be43210c797c48c0d642802c1974cc3cdc46df65f27b35af1ba068f20cd86d16f027f1492573c62ac9f777ef7729c5790d23d8f3c31e267190f202a3194f58dac3c4ed67d10e740e07ff8fcca43c0d2f7731afc5b56090ac3ff8af1ef47098514866f058436de8d51dddccb6c518e12399f4adfe49ead4a672a4ce6b2aca5884cb698b10cf4959b95ce9140109f04fbb0572e0664f469d88514809f1b7e9e051ed6694144ab21e9f7522739d2cd72db090ff62c15205c2a7350092861f5f6aa3db76fa68c9e60cbaf352c048f6b18d68dd403ee4ae2a09872a5127a642131b3c8c3d5d33013de526c7a7a89e082234ebc61b014ffb2c711b0c6a836594a5572dceb7fa736dab563a94001c3543a355571071e4865e4d52e9e79eb0b5cba073c344e634e77b80255bdc6ba638e239ffd6453a57a058d9b116fcd73cbc69467a4bcb3dd5c033ffdb0b920190c1a298a079729ed947aa0c2548af8838d367707ec5304d19098fc16cd753ecaf339c9b885f3ede3819bab37d23eb8c376f8a3993f9e5afccde08630505a9dd49c46cc9672e0b6de9d2d95e2bea131b1ca2523ceb79386fb9fa9724a352a970ce8c6530d5450d84851acb8171d7107668a94aa2679058c011170bd892974d6bd94e0b3b0b7d379f39ce86e9b1ea2015349677ed536cabc06ece5f1c275164821f6341e67711543bd05239da5ada79ba0da23da3996005eb2e5d4444bfea006821cdb4d1f500fa201a83eac3d8aaf9f2df15bf6a5c8e7ecd26e0e26f445ad6a80a29e57bc5722ee4e43ac17f2a0f571e3c00b72fcde1241e4b8b0edfc01da95badbfd535c688f47bc66c785618a1efe39744c667b7d3ee943e952a6650e07fc0775ebfa642bfa17065a1ed3f0a3406b234b99e021f574d73638b9672d40fc76e4e4e69ae58933c7791e67de04ec7a890f0cc0da4c483bbdfdaa3032deefc01bb4a501c23f2a243859cf84eb6ef345ee368d6308930c107f37ad06a92a915d235b457d7305b4fb3462f5e7410c5d06e9148e82d9c8f4a30bb4a5834b5ab52b25f7b174998157fcee85e1228b8a85eb215fa86f65a5db7bbfba6537b855891c434f23e8d7a55177cb31a6384c50492cac684a165f949524473b24343f57c1bedd608519ed8ab78ccf2fb88de893fa52ccd25b5ad2c2ba8e61b761094e269ba0afc7e5391f8f3242533032b981f58950275e71152d6ceb4e4ac537d34c3ebd6320880921327b0b9e04ba15c0ec100cfaf639af2746cca6a2bd6de174ab9ee83cd443a2e7b6aefc070dd63b57216818dbd8f395539ce34ef1a35a33e98c6ad4549f4613f22e7ebd7a7bc98bc6fdd7b8c37cf85bf8d95e66c791747969354df9fa107e8402e07d58fcdfa4364f7c6d32ff603fa2c3de3be8c1347d5f255b41617b704188a6ff17bdbfcd949961eb96a26ca391ce1c496a34fcec057179b9206c52db982fd43ca7016ddd27b0985f47372b17d8e21fd352bd6930913fd1d860323ad8667dcf508d3fdfd7bd4c7d1fc1a870ee3a239ac366906bbe7057533a725f94fb5a40fdc8c4feae1d715abfdf2f010c777df4bb612770875264453131351bc3b3a45adaf61e133ce1a849dcf1f1917c39b56ac993f08cae55d46f5f38470f104c461522aa9400d8e143e7744049875b88ab544c70abb9a7f8df8dafd7a5dff955f7286be7332a16f1dfac3bee3d4603f0410447219c6f9d73926f321d363fa341fac4b8e49cb659cf0fd23aa227a634e1ded822a29410a3df901e5060c1c2c24f2735fdd417dbc86d3127131861649bdbfe25e0adc3954fa6d15ec7cdd8a62567b40bf38cd8bb0aa766e35655406b67d21eb329275324c69230231e3e1102511322afcc9a9abe3156760150f05bb00f2b0379ceaa0ceb7b8e833ddbb24b539eed43c9b890b55119f508fda1b60da930c83d857779304f84bdbb5c9c6adcf21a4579504d4eb83631ea3fd72a404f4824ecce9012fce04c2f4c7686cd1502a874c3390774974c3d59e8be91ac766c8ac7077dde75999c663985b8f8d917b553d753c60bc2268a1c2a139fb1b2040d4f6573e66c542e37234cf48087cb443325e19a8f4deff5589b1473d43e3f209c80acc7381581f127a2176e3b1a6855691494fc2165046fdabd4f44de4b2bdc4bc60d5bc54c0c106d96bd09a1a046d35a460d55f53f1e837d5f38d4ff8e7216cc22a642a2fd657cf86de7dafe29715bfda85cacab7ade3afb8ade4f4f448d80670560e3409693ab79364ff9aa7e82d76567571ce06e540e85f3cd371128b032b1f5efe06f190add5ada09d4eb2f9e5991b17b377d15ad23cf8b9c192e652fcefbc8be9d6c2d24139b9e157ad32ef20a557025f8413268ed714afb039fdafe19785052ce75a07461f029ecb4386d4bc1721e76ba35401c30887eaedfe361ecc7f68ab655a5c8f299a4e8c6edd9822b402509181691d01d0ede507c2fbe991e45a470b2290a1ce8569bf8ba5f1878cac43c6c1bb41b6dcbc923791d6b53cbfdec8244dbe90b49a0236d6d1ce3027d3e99d9adc3c4fc053dde15caafa52a158193a76b178f25cf4c59f371bb3ad60dc80b731db3912e2e805f71cd5c039a7f3869eef9808d8b15a26d7050d17a6de10a0a82e3d94093780a00c7efbacba9da4d72238c6e6feb8f89ebe194fc0e1817b64463d767d5b176ba5c41db6248ff71e5890fefc176aa148d059ac723c8297c855c256b4baf49e1a8d454992e6f2f9ca7434d838326aa09970cc269a7167d40abba3c04e567cc205653e88dd15d5b5a1862a52a78ed02c373e3cac09c182b70021c163ecb54cf95e112fa55b6266d00a4cf3b9395d4992fe4a8ba72b8e0217b8a64c87b7f3a2d7c77a37b228ebd655b32e5cf5aa191c95fbda9dab2dbb94470f7c3e75622ceee07357faaa003b84ffd4d370385304d063b8c647253c6b093479e6181d936fbe88dce551bbbcfecf171689c55465ae9de31d8c98f0bef709667cbec0b636ab594ad9ac75248a539d84ff425543eb19b6bda88dacac67d1d0908a95777a294b0a8811a949e6641a04c6ecd0714ceafd207ed37c60eade096c3f2df50b009e96e85962a101e82b05162afdfe7257cf29dd6de18ac702da0f76a91a95cc4a46ecc2121797a0869d9af86c2f90b3b54738ebe82374207523869388d8934a8c602c63d859a65a6c545e98d6ab6426b00d3683ffd970a15fc4e2353c0f325528efeb7fd4ac2b1a1046b740404dddc736e972529ec252162f45f29c7eed1ba7cead852d5126b492328e667da586a5054e2c8029cdef3476676c62298429fddbdef9fe809223beb6f4fdb56016e7c9c9fae8d4410c82e069e6d4bf421ea8d5b2b83774dd3366f10da29ff1287bb1de852e64f89899e065b2e2864d78ca4077035a6e8aedd5cf1e5c72f591349708683aa38401618ff82a6904839afec100e8b4b74f3a559910fcd014156e54eb6b3845a09643551a5e352c4a559a3393d369d609292e65bacff70c4ef205a793835d1eed5ffcd8e984c451d6de998f4c10b724ea8ce38ca51580fb29c7f617b19510d7d9281ecaf0a0ae987d6d06af28a8a92baa1ce44d474df0dcd1acc601a03f768aa5018679009263eedb26a27d7c7904d1f7b146d10d780c4bf1ccb1bf91bf8a59430583816925cc2d9334ff5332d19be859e6db77318f905d28a5c32498e62d80f52476de59975a0fb23c1d0044fbbb7e7cdd74b4431a289099fae21f2c9fb4b78714715b4896a9305f8c5ab18985ffd53a120e6f8e3cfdcb9b8aa0c19fdc2867c4d9bb5b5653a521ad7a48d5b8fd66d2197565e66fc3fc4e4fba31097af803fe05e4d117bcfd87e205115822b38ba46e0c9bd497321242d09e0c07b6eba0f7eaf0e06537df3724c81095be6e30ebb13895e3a908ad0645ae68787e08d2447c48a64773e04f30df63cbcb50e09d1325904862087c45db39ce4164c600b36b6d35d27358b517ed9c0667d6598791819e0d4d17662ee74a1f656b4e203839fb6728225c25ea122e497e4831b35abec2dc2fd5a3eabe7abb7a87031ac9daa4b793e83b1a60dff92e9d2e676a47732d13deeeddff3a31694907554180fc7c6c0edf37e71c68bd3bd8549c3b83b25ed42bb84f9bb2d32877400bd8b2db6fb843e64e7ba329d6fe9a2619bea7f89bd7ffa0746f1a8d71010da213cd9d74ea9b37ebba8a2a2c483f3670e8e6959c40cf95458143f07a3e9fd3427c32ca75c3c9302d8c97840e09bb2caace944cf6f869460eccfd8d612eb2b70576db61554a358070aba3df95364731b3fa1c248fd4170d96703c1055bff3eafe6a5473bd7b80162fda11ab8899e46f0e08eb6a2cb9710b202caf2b48e28f5223b9b20049da7dc791f924dd7087118445e90011a44285b5a623422288983f2c5da0d85d29935711ac1b63059eb7b3482d1ec88916ef0b4d86883d310c8162b198598298b12d2812ca98dc2b72a13134814d60aa5acc2a4f68bdf1fc8e560dd151fbd4048ddd817869047640dd14df048a4c108a226297d8da31cb2cfc74cd579a1da3ed6379ae689137a91afb429caf2249dd0c02e025c891c0e1e4aec34f117d803822749465c82c823587e2dc86e0944418f9ccc95e4b95233ddb47af4dbd4cb5885a5f3de408be9781a3bd97d5d0f56545d742aa3dc76fbf8ced19cc2eba1bbe9ba40acb33b35a9fa70d0f21486511ffe9d8a50b9670bc216f95e29e289b41de2fbf84427d14d6c6dd887630ed45f67d330f953d7746907382700d24323819c1caa41a8320ed692401f433c55113e8a4b73f4f5677ca747d9054d18c4d94a7d62006d038964bb50104adf3968f8901bede72e5438380a77ba4758b9656bdecb1c6c5619f7b720619a8ad6ef5ac1ac7c5594874017464d67c60e0bde0b9899e5b68adc1f90bf650d91243e1eb18e15b808d01a96e30e9d985da3fad05f2df3f1aad0ac074351a590f873a4a2f65ec584b9c36b7c910732ee96cd5f65270d1480f1ab9ffe0bd54c7a2045519fcf64dd8b2d674b2e9250034fd3ab402f131cd43031b52d3402;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h32d7babef945181cd2fe7e05089358a12a5a24826b821e0f38d0105992fd73a1370df148593b3a00429fd4ad08359c41d6d8f20ecdde5f6ba51b7c8d6b601360f75a7b8df0943107421786c2f03bf6db888b6f4fbd4723f5463748023209a44a917c868e84ba6ebd362595dc53ad6f6fdd61fa3e291410cb051d8305ff26418a045161381cdf3e20dad4e45d199f9d754abc7fb036caf6d77569d7fabe76c35fe913a363136b1ef30b9b0608efbd1aec7dd9dfd93d39c91b1d7f3f1949bdec0ecd47cbecf708bb80788ba7a0e933d91470e573cdf209968ca6aea79f66ca9a08a8d25498e3b000ea139411d9251c98c660a1153b3c3b449944e94f76748fcfe0d54bfbb783961db99c88c3404b2079ddb2a26a999dd0e6d7da3b456e2e886844f7e41a0026257c0653f53af3c8d583ff38ee5a7d22cd64f21098d460a4761f7c8086b83f5be25db3c34083d58f7634878b2e13cf59feb67e9844e405bc16f1b668979392d0ef710fa72573d6e9061e4b058f871651fca9b3e56d64a93af523c877c3087727c2d13d331b921369940ecb80879e894cb5b051c7196a2281d61f92d97b6b874c856a047a633b3a89e5f59bfc36f100d2a4b97a9397719c2e2b8a3750a2d80b3263ad782915e7961f1d5ab113c65b3a2b179a7561239ad9d362c585f3a41be8939b9a6b3e24362e6532488a251d9e7c77f703c9e224a7e4fb768a44edb268592d1ac027f7af2fdfc4a7b761a088d63e1d6f54a31c014d42ce7d4c5877588e6231161649ba2db3ee472f2bec22b96e8007996cd9f076346d2c07b16ecb48fcaff5925f5ad1614d0125a27bf97192e7f5818c955c142da4f8c002dfe74b959fad06389cb9e325bf9082e5e14d9e213b37f076c211191cd35a051860c427f0d543a51c5b2e58e02522db663f5b58ecaa5bbd2cb596cc6efaac51bf058c272500eb55a6d015d2196172a0b4451b46e98226e5f0e7d031b41e148ba29223035ce47c20b69ea940189150f050747c4624435c07ef02c9c56c000530386d5741f6e0a0d0f8a8de628262dd9a6cc3e8f01ec6376a658cdad86a73bf22612d945281fe13987aa8be41b0f0f807c447086d29d60f0ab961b8ba04782698dbf1352acf3b6e91fed3834116e6c6e92aee4aa42f29736a2438fc3888b740c65c73e2ed5a0227cacef727ad1ea226c553de3f35a91315ffbe57ec805ceb3784df37fcf9c9bc0e1de854ba9a58e1fb48ad962cc2fbadbaa451c8964ecdbe052a821a754b99c42ce29818a38dd1ab225588c2045861cc8f3a805e0c69903dce26c81b6879c2cc8c934648217c6fbe437a38ae0680cae7b5bc587a6263bd58770a60f7f289fa0dc43cef97472b0d232e38449d26d2155b1d691152c1d4feb593488b3055ab58b313a5d28e25e27e295059f33aa5388d847a3870edc5194ff7991d75f7632652cb7012fdfb7003bce4dfd7cc2c90a32d4da4e74acd29a127025dff5afa632121dc7643a7e2bf62fb9bed49f3c34778b09f1e9af66313bb6ad1d758a8472e188dc86903dc5ba6ff65187eba8c637d0ae886dd093e98a37d22e5c4f1002a834843b106f517fbb2d3be73520f57eaf35bb8e5495869c3311e29c5714aee0d9ad7e646406908353521119ecd217b6a9d99f49317405139a8c89afa1c7424b06807615df8b7487e3e3cd2120e2494e7871676e8ec85679408ec908ef7e524ad1f5f2b6ca4496a04d6e7700fc0908e487bfcd0bcb423ac36d5613a8512f1933fbf0a3a02f984e1add86a8bff8ba4ba04fe478e562535032c5206e6100c9e84b117b4a6b78ea7fb7b195f1fe7d2097cc0473d32b3afd34cdedcdcbc82dc6559a604edf4272e582bde8d902ecfb9dc691fc6949b8095d97fdd9acd0fb4db90a0ba6d2b46642f33348056d5710bf806e79addc0d4b1192088b006dc12770106ad4924e1c610b2b4ff50802879b7ce8001141e1128278734cb6c42003ed49b66819456bdcf39b058919307192b2b8938ee9ed53e6275753462a1df5bf5914890a0b76d4110d9e9ade9320ae9bf5a0b896303984b53748a12980ec62513b65df2e022a1c25eee734f3dee97169b29376900be954d8aa2316d49d8ab41e683898623a1645a532f60309dd394e71313467a4d461f2bf72d1f0a8acb863752e5988aa48d92db24c969b02a052d103dc6357e19ebf46bd2e7a7e8029861431d46ba9577223130fd9faf8074272e5b897af6348922e3967a75831d2ac17e745f61f3d1877c45ee458fc7a32f480174b711dcc98c52f98760ba01726373b1a9699b9474f77b70fa856e69e35e9e4fa2d5629ae7f0990f42e8b4053876fb4678c8577379e4ab185e7316d440db0e7dd854adef88a9d89f26c23ce4b02ec6062275c8a85fc14b65611ceb0ab9ff628db8a11436a4ea5cb3354580d389cbbf98c02736ee503eaf437ad07230adc2ec62de2e4caf405bb775f30534f94a688beaa8dcf54bde198b01a3f5eaf79c381b146bd3927240f1264655268878fdc6bfb2e578cfaf680a0583e7177ccd44e20788863b9549920209232e29662abef3c8dac3bbd5a04d931b39e0b0b310246771920a96f86a8035776df159fff1680896c72904d6fb980d48086ccf957d22678f960bb078b5ee02e3a723afcff8464e1d9c3ea63a457fb0c005cc3ae2e3b601928b5e368a17c686a0c8891efadc776244cd0a100a5d7e95a55ab866912562c09fda332e15f1d7e61602b6cadf1065db28a3e4d5f24b20e476c9a6884d112c256398899f5826d5b3b9c4057bfd59ca4255b23029c82b32b849d633eb70f754a8fae15aef75675732e5d88289c1741b89bdb9dd3642bf9aacbd03f1ae77fe1dbed790a9818be75a4c1f9d4eea95173e56dc9e4e2fe0b0801d31be1bf489e4c0d8bb02f83e267ee51bdfaca3cb9bb5bb930025d7140d7cc8c2a9011c67dd80b9429680f71c1d6f7ca0295b9eb89b28204e46753d104753fccfcf81571b9f6779eb7fc4a5a9cd0764e48c241a63ea63cee13cec0e5a2f619e2b41250f2fbda98da66ff224106985369d58265c449a679ad266e37822a04502f2a0eeeb819c67f000425b45c26282cc91e0cd224503586969097ffd3cf1e1367f67725c71f232758785bded8ad05510d4177e37a42ee3223d062bf677fe6a06332de64f89217e5f3f1e20569a4b7ca07c6e3be18b5a115ff50656e8f42f33226e85cf5797bab2ba4bc232f777ced33d0a2e6f84c6522bc04956e5c68cd44da43bcded369ea487692816a38fd2bcbaba7e4407363983e59a64548c3476cbf6849b9f3e0a7a9225ea343393891c1c2328328548484c151887ddc7b033aa064e7b04bb1095ba04779bc7a3a0147869cf319e6b88959a3f9e091e027a68b5a00c3c00395b40379acb3429ed10b39b831f2ea7d69cbeae057ad58159a0bd31e86d0b5b5d5643aa0985a8193d3ae906e67d4664b115e8af5e32d88b9eccdb98edd28292f97c7252c924d80cda04f1b7a608ebedf5692a86079a74d92bb1c6248c4283120b9f3b732de9e9ae1cc636ac5cf5644eaa0e7ff04348c977ad746c13b58872fc07b93e1f9194c181681da3b226d6e8528db06f1a3e0bb2c8e74ecf7aa2748265e2c0ad7c54aa27bc15f928066772853ae5fbfbbbf52c3f564bfb501de50912171095bcc20d36ed7127d69a3c1b001af7471e0d83d9b49128d650ac408f647d94267ac34b93313e6db3aeea135a0902449857e96cbfed94fea652b25981a747dc994ea969876c0d6da2c819b5b0f0727d14c908f6898275a448c692f355309f96cd30b100890ac5141d99f5d5bd4f592857a5fad834078be0f07e87d849eb3b11ab51d48183e37b9e6e5b4093af42c02b457dedc461ac8b7c7ba9a466eb0c6747639d9187068cd55e17f8646c97d7a5cacc4089e51a7fdbca7eea7a6b58316b2f537d3e0ea76c78abf394afb5d94d9b22d57a26168cdb72483894c837a8e49990effbe31c81c38aa4e0cc552c605449234fe5a0eb1ad678a910d1f7e3b3dfdc0aff5e46d0e650f4f04226c68d024f8cd441b3a15e8d00675ff5ee7581c721e1a58c571c2d86449c7377bb2a0af2aa0e1599621e9eb16bcde7f6bff92547e3f877368563dc5049adbf5420b82d976dc587bae2b1de203e15e2372ea01dcfb458bb1832200281190f1bb83bd488fcc4b92523d269419937b893faf9d119c7ceb9d493ca98843fb2afebaa47eda8005c370312c89be244976f2465557ca5771cad8094c55cddfcae972d2bac96385ff58cf8200dc16fd5f1f025cb7ed2f54b694fe06482ce1bfa3106ffae346984498fdcb7175097967ac165afdbbaaa73fde1a8fc57ee801a0c4e0c31d64c846902d8922948639d6575cf57a3cafaaf10239c11a56f6048d8558f1ac663ca8842c9e17c9c9bbdb45fe55c6ba0bb8f4dc08f929e895c2b9420626f921bfdf18edb845bae4b550b5c2ecc9156c66b2b8d8aab0d82ae0e6dd33dff0de7c0bd63d163a6efd4d13a44fdb3738bbf94f9024cb6324af7c2e7810764c2e2805d076866b62b73be9ede16a98a7796378483ff87f80593f3f5d5b25b9ebd5996ff19f3c6c838c55d3058ee17a7a07eef3c6613ae0da4ee0f122149a9e6ce8269f016cfa86bef821dc1f4d0a385d3d670d19a8d040d42b831a9b7505faffa85d2a168e844d9d779df1371ac038b8f9214b089cc64e3d989ce451d34368f3efb1a8bd49307acf2441dbad90c75cca372870496a604d1f42f63e011e79319c824023625d1876f55247e331b0749b7d1f80c3d7782d1556e71e63c45cf9c51fecccad7bf473f4a4382fa1c3200c02117a9607a075c301d4d2dbc00df2b2c9986882b912b4c8de9aa8cfa54869e137188a8aa73b6b2e66794fff7aea8c243fd26323a17c452a66f3fac0c5cf1e6dd1b6d96d558691894645051b157f61e0a45541643365bf82645228255a5b5b7120fbf5a886a6fdb5320a552ae6011b5a9f6d9a7f3bc95b7b5ff10c41beb495631996477b033cb941c18ebfd36914d9bcf8b9d53b88717c3e8ae0a1f1d4bc547682f295e86c6c2bc7915c0e625e34c56baae3bb6bbc1ef0859ff2d3491f533f0031a38a62a6dceefa090653e0dd42cd7d9138f628a60da66decbf91a1bc2bb5e3d9fea91119bbf6ac5b46f4c1b8a9cd6086469eb2b2932dbd690fbd16371fc796e2a3f523039644882f972adb1d748c056dba162af34d5759f5a382ec1a448ef7c9c9046f1c81e3af7430534bd29002d70e11bd6461e2b969a768cc30fba0122f2ac078146fbf1b1838fdf4427af3314fdafcd54686e49f4295a57fece6a0fa1b5c133db04e634649ab9ac265287afaf9262bc454a8de4c387d68a992081aebd57feaa3c3c3b9d43e022714354af7089dc548a1c6451c138b7c35027a32a016b7731767ec100bc3c875cd87bd3addccd464724c0dc158189fa7d484bc37c50ae30b8d1c86357601ed50543437296e57945414e09ad145d997aec2e48422db456;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h9bd1d9367ae33ee1d3b29564377afd8635063fea2d4f2c769d0176d57aac32877dbced1504ab1d2d48dd6c1a3571911102746e8a27d269538b6d7c1ceba7aa309b0ec9c1d4e2ba9db8b7700efeb446c95fec9be6bc7a5233769177c75f2204ad0bc117a0d7b83e2e180b4f032d468fc704f867cc789e8ba62c3328d78c23886983782349653f0172f68b39362d9a4db349c3923660052438eba050f5cf59f003277167d5991d87498571b89027cafa4df698d87c05a95c2eb33c65df890f46139bc0b3c30764944e28e0a944983684af3ad5b0ebf32be6fbd2d33168d2804649cef759da462bad0fc1b7fde8b265ba3be347adacdc99f539befac783a70f558ecb84f6008c8cf783e3a5eda91353df0cf5df630f26c633033a2898f9f927023afd0d0cc413e200608a7636cca487a0de41cc42c3bbd3d3016eac67ce3f39f2cefbde350182b91dd1833d0f2bd33139256c3e8270f814da712195dee05fe9f631793426d813d6840eddddefc4524dfde1e6e10bb80174af5196b928713e7ce74a6bb403749ad28a20a185dcd7716183d5b341ff2c70207dd3c8f98e972b89507c75766c155627278376ed453fb0920f5a1416f4b8ca32e96fd832c72ef91939c9c24e05acc1fd01c07111388d27b2c00b30dc6057abee6a2675913383c93ddcbe6043380c4cf77f969a2f8717723b89bfe6c003978d95621636c606b18320d739a7fe5028313b058031d01e06e92ea55a5714db838b0ce99d62eda9c717cd51d2c9154f06bd96375519c299a196f342e4afcf9760d6a7a422484f0fd34357f7613e1013f32a9a15b036c9ea050327293b0d0c03c91f0b94333140312098f4a4f633c1093a0378f174a94c65d41a4a41d0cbc0f1a0de2b8a6b3cb6fdd26591184e27bbdefc21017d15d92f4bcd366c7497648a4b4222d1722add4e2019be5575cbb7c8772cfbd6953e0a3d2212e89e270666aa38f066101ea267e7913fdf736717af6b6f277e11687f254413c2f5ecc3da1e076aca0fc89d31476b2ee1c3fa4217a52ae9e38a8a7135ad914b023719c4b7a006e89b4d9a22aa49b38c9489f2fd596229684abe90e687959d59c5b4ac66d89daed91e6e2e0d6e3f39d3ace62b0c6a1783a3eea9ba937046b3918371cba4883a970e5dac180dbe7ddbe806276aef61cad5b14b27eaa86b14aff95bf16eb7ade1ca5f585f0f8d8b6cb3e600a9b5b50875b043afd087715cdb436fd70a9fa267e3da9902627cb900609dbb298b9c5c05e85d7e7b5919d40131a39e81cc784c6c080fe04fb31ecbfd53ea0ed44493ace1b000caecdfe6d9d3540127d55942b1d5de4f63aa782af8f0933aef0d58f6c7227a8866df1d0e766234a8842d82c0217b0fcc4ba0a5bd3a86a581c9e9aa36921b49b109937e0774fc11bdf4c281c94ac334d9aa26f1566f6678bc4760f6005edfc794b0bcc13a01c9c78c162172770bfaa3afabbc1d4f754e065e34a65f922d46af408ee9c01e47b5e4b6bf4b508e17f2ef4a747c0d8508ffc9a8cf3c68264aab50e95fcf2b770fc741e2187d138e49c8be7d1d973f505e4137257ce07da7d12fa52da21d4af14162bdc10680489b00c8a8adf0ee80ac0453c16f217512226f01d70708ba651cf7ed1e9f6adecb2a062627e3d54ac52e78479a7748de8fa8abe4136f73bfe3a9b9c13475dddad18efcd50c1063ae70b54c66e4c92277b0de5b3483d2bbeee125d4b58963bfed7ca6694fc47b9c37e30d4ec6f626fa1430257d02cb0731d7ea178f8855a7afbac15a44deaffc502c40131fc73b64e9213ef8396ffc665acb6f0d1e0f0139d6b1b1fb4236411ff4324e87a773cb268822a34a6e4db3b5b9c5e11f852a41d16873a30d8222f4477151619bd7cf0d1a8e63d4aec198e944b887516bb5731e98720c77a6dacfc76be967a1c972e7ec89382aadec1d04514e9fe182be7046b04abf706d00f15b8cbdf8e24b96ad115b918514594b1925628ea0d98c88cc6c12e4832a51fdadb91e23052928a80700a35625dbc0224b3ada4dd231fabe7ea5da2e77789297de918ade77b66d0c2ba91be700b34e96ec753a740b8b9fd2eed9e26bf75cd4a1a6536c87383706540c839c64c5dd6b6771a3f107ef6679a40de70a5e9a38e93e541a902bd1a4c47aff0d70f919d9f8da27aebf96128eaa4228c04ef93401b3bb47dadbee258992ba9729fb9c0875270c4c473a4862a8eb2f724e285249820643f08c7e79410cc5e548079525c1334f53e7a7a5afd4e00d5d8c0b3ff779b17166e941d05b31c09e11b8fc0891177ef77298f3285a5b65878bc1ca038b2b2e13b015f4f5d8fd485fc33c7a05cda6871380b618cd31c6aaa00bc6465357425d5b90985651b6590191df980090cc74cc0e8d8427ca65c157a1353f36266e9e89250dfe02891d6914b0476b34503eae46947dfa0c481d31be7f6807b1a6d6a9748b8514175c1392d49acd857fc34832ef9ae49d28f2637478acd848cadd3764d0fb776227a8d96c4c356d0e3896a24c6a3e1d915b7e5744841d9f328415ddefb385587ab0fe5224df25fd88630162f02cded6eb0da829f1d4bfebbeae31beb4cf59d36baa275b7b0962e000ad2797f9e3347ae56c93c5a876e11ac823b5a58895c32bc1866fbabbf1d04b6ec78ced6e3b08731b25809e7db8846545ab43cb78863e54dbbb37353c7158936b499eb4bc26fbb6864088154c0a961d1b546927726e7d9f9a6e204c4589ec3ea498f54692f0902a92cb73cd4facb69a0f5a848b25a6ca1b99ddd5a711de7409f028617598e76afef2938a23b152b32c331d43f940acf4e79d22debcb68164c429aa88a22ca067e3e452ade42ca514b30b4fd0413b0c9973481f91f012ade8349783cde866edf8ecd90e91dbd4ec437064af7a1114569c14033cc00e51ad741f6740742442f1af121439b3731c01e22c5a5841b487b760b8d78d708ab7ae4018d41db52109f4dfc7617ce8f936112c4d5806a0f16cd32ea6d673c136f20a27a869cc943b8eeb924935e10c3e689536dbde039653aff4cc64e0bce26c18842c99aa32c8abda3293dacf6185e68b0375763d2c486777f407a4caad5a5a114ab141461202cc487dd929e96e13286eb6b450ad2ede749f3b72c75890ccb4143d60707cd9113f108cb7ea5c6178ed463598c5ee36639dec3a96dbb09fb73c6bd2e91726d5a7200bbeb1aaaff110fb3b60cda531af0f9c2175c43634b52dda892d8bd0e2bf60f66be505edd9aa2b8d67d0420ab8bf4a3e6a5f60cfa37c5fe7b27ca5752d59e6feb2d2a425734300a90116baa8e3b8ea35cbc0c61a52532229cc00b30be7dd9bb9ac11456fb0ddfd1d359c44d9a1abc73f1617b2cebbfb23aaf62298020c27d7234b4a5d40c0b1a341f46e45e108b26425e88ee794cfa7ea38d1a0f1a7df89dd8f104673c321a8a45cff3bae09fe47dee20a9c96efd24ffbf1989a7ab1a1bc68c01f076e58f131c4efc4ce46a70d7e59b7e7d68642b317770c6c2599a7bedb79e02c926603a8e00b19176d2ee957cdee439dfdc17144803503c7d2153541b2c4d275477476cde3b6c6874c73ca1dce9e2b6185833d56df6dbaf0daea17e4db64a793861bc2f1f079ac0094dd5e66c3af10120d5aa917afab0756f794723da150a4782ba0b4b6ef0110ea7642a816ce1d7de5ed4f38311526eb9b98e3a927c0376e548e350ad4a2303f505a419797e5034f64085964e0030d3c525cec0148ccd3ffef0b867141be8d7c3d8d04eb771f50eb037a035512a4b2443072143bf4887899749f2ac1a280522e23a6bf8da3b0664ed696b4d8d58759ce57bd21f5c5eb01f94cde3ec39430798ff1f0a79b831c061d861e13186a3daf09b50a90fd59026b876b9a5df17e66f48c3f86fae82d318fb3535b40b9ce43afa30157024a76227ec1765924002d711cc2fdd55d2be6ec77c382844b750929505fd15b84687aba66a38a50d2c45f9134d77f99fcf0edfec9c8b50897e0e6824c01bfc4f56872cb26d0a78492a34600ccde8ef52599d7861caff32c99b67e4e958c094db2baaf884c072646833a9e6cbcfdbc6fde54d7dc78a836677a81d766392af7bfbd7b8fc5fefb001eb36bb20951faa2ea72359bd71c4ce337a23a2813bc8b4fdac8db7ab23e0529d839da105784b892b8957fe2753ab9f0f145fe3e41382810c75634e391c2efbb0fd4b2413199a32a25be6a7bcbd3371b5c6422232929cb71e15350f5da1efa85fb2d30797d13199a0baee84d8bcf6f8c641a191c6e4dfab40788c5b25ce190c1417683e04e28f342cca227cd7e970af567aa606f1ec82f023138f3ce676b4a38b7f22b2a13bfe93468e08bcce192958048a9516e26b35a7f7a5af2b14039445a189ff78851254562cb9c9ad71ddca693639a9e38a58f65a84c1257ce4a5ed3288d97777f10bbdf22aa54486b827cba1a93d308fb0ac0d1de6f50ef83b675a585ea07d2f7e274e72e0a8a72f2db872e6b6eaa2b2959bec3f36b162e90bfec59168a295c6b8e2c7846c5d0d637f0fa1592f2f1fbccb603d64c077447303775856db957b5870e6ece767388a85d736f5cc7ddd06eb25e81aae12d83eb1a9194707c55edb2d61a33d7cf6b8855f23e76cc23abb9e6ac9ba88a2867f4d53286ee5eefe110826d3f3ca322b260b39c38658f4c9768f8adfb2dce8071c13a16ea8ce5f6deb82e2f08be06a682689c1ddee52402cc65879b172c72655f7793f0c58dea2199f25281e61799e37aec5cefdfb839be0a021135c76c69640642dd546d2c6262c6a0a7feaf717cc55496db104f95c45aefda86bb49ef1aa28ffeaa30cc0f298b92cf0254b7e00813fba8e2bfb8416cbc5d0cc1b0a6b63200761322d184e800b0c63c97ac47f8c0c5de93d551d0b6679c1cb38787a7eca7b6578cb4f348055e21014cb8be1ea653be05f809e5030ac5da4427160f3e4fae5193962a7233b7b5200ed5a50e5b1204653a0162c2e15851a5983bdb94c9dcc154a755f710f482f31d62eca0456dd0b213a7aaa5d7a38939cf19e4f897a89f5d57de138e22f0125996e401333d11606443e3b9c5a6df393dc91af06b01dff1f0596ffee1e8be7624a6af94597ebd54a85434275618bb4bc906925f01ff33fe1e175041c603cbb2983510aac3392744d66cafce0a27fef49b989cfb1d3359dffdf6cf9ff2aedccc9bbf9dff4d0d5d22b47e621fd2f64ce325eaddfb58f198aa8cf26b1befa5c97d229011941b0b95e42b3c6f41c69b4469fda27919e8475c601b5baa34b20dfd35b473a89eb2d6d9aae1129c63ee6cf4cef79a1c6c5d7b1e84b430cd3ead8938586288603844a22e65ae0d4bf6097d798a58ed1b606bdcabc1a244a6c6fb768eb2222a68face76b2a43c87673f04f4c471e4212ebfe00fcf876b2d9485f8893ae48f30ecc15307b9437c8da46d70f32807399b6ed927c197e369db5fa516e058566855c10d1c76c1a93c5eb9275f6517806f501c10fc1a86;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hbf9de0bf160e22ab86ac6ef0ce22ad172e50291f538cbf74a31c15e7b9c9c592595db0ca6b273135a584e22c89ddd039acb741ba87de9c38c5362ab516df14debf9b13b99faffb2f4cede5c27df051403d9b3f3a1ac990e540d08c161db330759de591665b0a3094b20cdf4f3f89f326f34836e9ecd4e318bcf4e5e326eb5b799c18d016e627acac90fe6d2324a6c645352375abfea1396c1e62da42e1e422812a5a2579b58c0e59a1325f10fc91c47f2bb994514848255425659c761004a3267b1b27b53a943a625cd2781955763d7c50709616c0a0694521a065ec4700bd7566d256005baa54af8a5886ad7c2bb4612328904cb164db03731f8dbaa63d80095ba9e9fd5dc9359b0bbe674ebbe532139da58160be723daa21cd13edc0eb0924664af45f7a1e57de1987f9f53923b46f622a5408e6bd353196e7400732d4a05ae25bace06bd8d80970a3fbeecc830ec0035f15e51c3023c7e107161a30f647a9a0719c8b9f50d33f53fa5934ea767f336bcb3c4b1e51340cf4fd81cfc3c2723acb8ffc23dce215dc01e25313fd36fc85dac38615730713bfa634ca6eda1f486347acd7bd260577aa4b503df80cdc2851caa61d82d7325fb6e8b456cad2697cc5a65e6da29f2157dafe738959506d9a17b1c375875817a1dc2473ca9e501b1f0e5afed6bf00cfd537285b478a1d9d43a1a08981a5ee8773b06e45bf8f9d235021d60efd491b60d774469944c4b220c4f580d2ab33d891733d4f41e013779a6a11014d6df2fa5c63fc008d4bdd8bd93ca00b4f6a1ffea13c5e53cd7281c3766e9dbd8a55f686db83c2bbd6918f8d48a55de10d95a4008cd2705a755f22b1c6debbeed60505bf8ba450b18db7aff8561bb138769c84493a5a9442599f75e77b7c1543a2fa52c5fc0f999f623ab33d353b1ec21aa0f0a72e24bad3ea68a58ba66ae4ea1922d94f752f01c58f747caa7393735351ed4aaa9d5a0eb85c7e66450ada4d1d370f19caf161d801aee2761eb1a18f5ffb0542278d86c2317b70ee719a031b6efc4097d157bce3d0624d76b2b738c80dab9db47a88256598caa85c2f7fd934ad3a22883e4c0f05b17da7ac05f7144956acb9b5fe1b95b213f27549b23bb3a77c7e037252ba3f24059ecdb144bce03d573bf309544d9fa96bd829cf3e73cd8ad96fa206cc386e10c6af0818ef6dbca68340ef21e04398871f5d8f7b8ba82cf33d1e6e1cdc88f96c620f13c14177e6140ea8cdaec93c54e6d10bfb80d73da17ec9ad6b39b3e8c7665e71370e16031b957700ee4a530086115bbe37a7a39824ec14a7dfb964883da1ac8aace9d9d23078e6582ac7b6bdf6380fa8ce467c717bcae6e0e483e0b1ecf50bac7147642adc37a7f2182b1cf3136338ac1f3cc3b9bd7c79cd0f9d67cb45a59e6acc63ab6af0ca5f11978b088c84b0c775ab78b07452d5287fbda45e455aa7634099f35258eac47a16a3b54add78eeabe034caa9b116a5ac4f7b3c5469533e8883caea16b064183c062f4c64a52faeec6c996122db932ff8a3b95dd4efb5638a36674e36c00b8fbface7763919d42d197444e07eec0bfb80b733640b3626116837cbcf97ac75a0af70e143f10632550c0dd61534e0ceea72bd38963484132b5eaf951469501c8586bf9080b7ce6608c652482e1d817d16a0fdfec4d14384d26f74f8e47485397e71192865da4d66de8193f470dadbc8c0c504b7495ae6c77767da83897beaa443e449a06a4b980450eb979203c58bae359dc056f76661a50019b128d7d268a6e06b52d49cddca717be7c0b866b29044cb5e3819b19334836aa3ccaf5e712a173019bfde3883266d8629a98ca663902efad977635830b0b8a16ea85c079efeb6f748af3d9f24e4dbdc586bba978a183397cd4c2ae13b79502d29b3d00fa4bc79b696216d6f97da8a7dcf9e6e73c37e18e3b294118b5d21254f9e5f584c0b1762c29a8500c6b08e8ddb3e734b7b884467ec14b1d2ae9af611b39181f373cb36354bfbff11e7e29356723f828155e6b5a3532cc24b6098b942e0970403c877cf65822fe7a3c2f00879df316f99ae147a72467884a4b28a830173414c0ac074f4d10a42687ef4e12b966e5913531505c7bbe6159f8b464b8092d82907dfc8c3af4d889b62156762135ce51658a1847b6d7cf5240f092113d8123f487e58f0aa07efb940210454faa7c231a1ad27a5d69bdd249692169c6e5a1f12323ddf7ad9154a4770bec2f54850bff9e1972fa9e4ffcf52a611cfe3fbe0f3ef12afde4226a0d8b5eec4ff6ee185221c010ba2cd9232d0911f70cb863899bf8d43c598cc7c57e90a06b37e6cdcfe92eda9725433ecf3b9736532716381215a9fdc86f5f7df02e90264ec8b867f7d0b86650df0fe17590e588d86e47dded455fcd716b45ef221d8739e301369891cebb75ace5f1826901267a78b65c53763c0f3dbe1ca7bc59a8838e5859454f24adf8257920111ed2dc26f03ddab3116ca1dfeed7daef82dc438be49d54198586ad58469daafbe0aa68a00c3cc37e6bf8515ae3f2a3297bde442ba93a7d591f9087d3995ff67ccff90c009a6a5f498caf53b442988b1014f2b7fd3c72830d64eb557354c386264c4a9c84ef66bfcc174f5564fdd1557cc7478ea37fca965f4f6dce0a0184e40e6c557e0a629ceff1cee07cf3c999bdf9d77de8af4f8860ead8083d0044ef08b64bb11f32eb5e57bd1e966901ad829f3e7fc42bb285ea100965dffa07a8732bbaa3bff6bdeffdf6b7200066aaa08613dbef000dd4a670b039e062f59b6cd247f688c773657a924147eb4538a9b5e9c4565872c6c73a2bfbdb93e6733caf9ee1d9f9fbe30feb4d30dc257fa9c062b4efd090b562ec6c902d7a75968dea5628aac2410564295ff4f2b944d576b2e007fb0b710019033ab6604a8b3adf291e73c2fb2153da128a6757df51b892f07c4a643a525d51a81137991fff42a7e1c26aba434a118ca6a8dde700c013dd75f8bf04383b03349c31c5bb9b1b4c9636e9076905c7bb82531adff2d6539e66658b6a7757c4a49741abb1c93fd925716296c1f3e92ca348173319ba7c5b8382b89f9f68f1a7f3de36882b6b4e04d45dd73d33213833f15117dc4aadf5b1d825b24803551ed204ebfdcdbb299983d224ae8ae4627894895de4c1214321c5f3f4f6f25144d2ef2269807d495464081f333109ef0eeb09036d17d507760f1ee13e9b0cf5746e37c0b7d9b14238d0fb7053ec7577088707de1d899df360abbbe46315ea2a1c939fe6f0d943868807157ead37c2400f4545142d6c2a8518e9d5128ff4265332c71f9303d0322ad464aa6eec830444885b9f62a2b129d5fbea67885699c99885fa8301d31457f558cfd4512bdd03edd411fae6ac8059cbc2cb09e68692a9121eb3fae1061659ef6c04efd17e5358e60547b7a9fe83583b8c97fc91607150c65c069b1685e7b8da0038b8ee16dbd511363202bf60eef1b899b9900804de3307c759a80ae7bbc7afdfb6d96aa257b584d40fa27a162f31d4b0c97da030715b89f0208bdd310e4d6b454229eaa37ec4e9b03e3ac18183709f539345e2cecbe563bebd861afa6fa24fb5b4408db3df539e1e9e129f6f9aa9afa0c0ac7a835b5d322219e2bd8d8794a9124d6aff75a17780024528f1313c94138a6eea6ea18049d1c0a851129fd3e4fc73dcea6dcad74d85771543b653d4e5525b7707741f9498393d858122ea65e9a46e047c009fdfeecaded4fb65e6aa0d071a2600db0dbda529d64773965450699929611ba92f74a5455305c04795495174ba76653b13ce1f6cf131962d41d32a13e9c865d87bec2a688204c79d13918aeabe01eb743d28e9a4340f8336789e3f771781a49169cb8bd7fa33e13c135fd415896c955ca1347f6adc4995bc3558f3260af9041615ee107ad16a56f9d1ac3aec3c8d6897d24edbcd6405322d39d5c8931a56009371a2cf6cfa380976f50d7a307ff5deff0ca0fd97f1ed24dde852fbb4faf58914f42543e246ed7e56d7e925511201111f2507b1d25b739deb0788116745dd39140c17fad9b4229910115b51a09c0651d7b7884046a8b12f28a69c7813e6fb9b0f58b73b025f4090919d5e8c4ca898dcd76e2dc25420e14920662744a903d341a0d11b86d5e64bdd58cb43b0ce003d2c7ab2a65ce4c6fb07b33d5c87b721b21e8a2bbb0a399f1534396b0f8e5d05fa11828ddd1091ca305fb46ffb74d5c5c62d237022cb09c75c016ceb0383afc20459434e2e4f96c3b4adb126c36a1d988767539ba54be9515cb3da797da3813b425037bdc8bdc0860d66d6eb4f2dd4cc78a9effeeeea7a2f3cf855b6f108d9ac24123b47051221eb728f137013f3687a456238efbfe5383fa7578c7a984367ff4049512d08cbbb8fc109e95f54a1b266f393f5d170257e948203b7cd35a4bd4fd81e77989b98d7b2ef6f6623c70b3c09962c6bedb982e9ca744a0e03982fd129adad1cd1797fe6fc05c648a75c44653f6891c2f5fc7dbef94248e043b81f4a129dfd5d0c6a7759bdf2d1a67eadb3d2472bff41f3cb0591c1b55c356ba2938bf9242c196520eb543905756743d3e6f9f37248a9891c73c7e96e4fe759114ee78d75a690b8f97fdbaac6f6478a5ac6e12e955ecb7874718ebeacc648d7a0fccdee6681af54d6320ee235a5e73ed15c1b2c7c48df6aecb757712e55bebac6e0fc548a7f909a80426e3a629699945df8dfce45c4ed8b1e4b542c33f73134affb8da55e23f874659dc8ab120a633ee44d56b2d31c9a5d0f23113b79cd3c12f4099cef33acf0e9d907e4967cdd6b6ce63220e77438536412f6cd99c658bb146fec61d022b0afd5798b005c35f88b424d5db07a84a30e1db05a7f5995088126420d7e7aaf7f5bc388b9632898e623bf8c64f1be1a6ed8a39a4c44b53523dff6ba514d7e411a8b92787a128655b7ec485fb88ea5a5f2ee3ebe689ac96b33e2f081f9373fb5ee958741a0af0fa55f6131c279ccbe11863838bc1003eedd1c7c8d1aa58ccd6c32aeb18d5177b2c6690f3aea074b5dfdfb71d343e9a116fb3f42482805d5d14d81d82644033517ff01e8a53a90dde8c5eff7a0b476adc24902bf82ecbe34062b59b72ada6eee5bb23bf97acdbc850d533ecfaeb76dda7c88e50477e056e9de3c34680e92ac2c4b9689feb26791de02b5e418f084fd810dd71632c7a4707c269b67343f78e247a380ef2991bb8a5937e1bad0c2dca758faa71e47ade8364d22e677cf114fb1dc7811337a6083599c2afa984c680ac035f0dd3df2ff147f41fff504e4aa81dcae255f413fa4d923c997e72fdc2c5c004d1bba53dd011d6528dfa64f97bc55382d4c9dfee68be57a2c0375e1dec597803e716971a0d0917e098765547d89cec7d2575e9022efda36d6ec8b078015f5a4b42c2a5e01a19ec3e49a52c974f3c4c64be58163e6e0427df7e018320e8d4698eaff0aca75fc6aaa6923eb7f4ebde120a25d2df831c0259;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h291dd61f88e930f01156712117035c8e7ff2e55e910825996a8144054ed6681a1a58a9138508efe0c2cba6c6281e5d9ee5323d4d07752bbf991c6b4d44879d0d24ea827d30f956710ab553fda6a1a8b7770fb36fc0bfcacfe65b1d0347d9c4901b087696ab4b7c1fc3cdbbadf45520eaf99e059b7850ecb9676bc35c7421aa64bd68a19897a1697f68c63ce92f38283f4796814654318126f69a47132671adbbf9e04f0cde083ab464ef155632c534889a4be8f64cc25e6a03ef1118ae8d3d0783959c6edaf2a713d9c2809f2a07470686a0e4c90a4768538615a5e2c5c42be86282765bfc0427ccc8eb4bb1b081d552313418143c7a4b4139be6897c3467c118deb506004a8057eff97c60dd9b09225ddfd3448ef887e2ccfec66d3d7d7c166af3171fa9bcf6235d181ec369d588cf19f78d4667d76ac31e7249b9bc2d8c0af571bc8b7f1a75e6a9a109beba8dfaaa403dad0e564cd51c77690849174d9a7de735bf64786198527722690bd9efab07dabd9b683e8275d68235d649ea6a13287db1fceca84c9a79b6e7730f1fb39801bd0fa0335aa6890516ab783628757da6d7e0522d8beff4c4d4702cb6c6d4ec54198883cde44adaa5b5a1a542e321305925c6062e977f19cb6e2388708946cc8f16c273325a14344a8fbc6647284f931c0932dea96a00aab6f7e8b6d2b0fd2468e38413edccf17528668474398b4c88f13c869a7c9298dd25304495507c05c3b7d6d598596cd195ec42c94a0e831ad4a43d63b2eed1340605f3f640e177d46bfe69513c4d806ddb49d616de5d9ac12925b0353426b196f7775ec2b2a43edd0945eaaae074c4f489b13aa92b015d3ad25bddb698d2d477dee6949b5eef3af34cbd1406441f234099b4602670970c8f62a16dc59b075f69adab9630ff7bb576fcdb38e430e1a33cdf719c4e1803a68aea554e5aed0dd5edb1ca0bee193246dd4464392b68ad96852bfd1f573c6492e5316ad09380fd66740f29a2e761449567b137935b5240a61668899fc5cf853563b27d707546a84e6b6e360357cc7749ee91472058f70482e63656a186832a3f8547413058ae821f952083728a61b7aebaa801f55440b655e806affa7ea4d23bf6bc345d49f341d2ea76d1f165042c1460d502feeae60c07b7c4f4514e79c0e3af6295e474e19991cab2096a7b304725dac7f9655bda9e271efeaf721279f0a8c7d0c100325523c12762141781ed54ace46d9c517b5f903253bd662143e58ce1ba78fb4baacaef10403f2ced1a5ec69ac829d018c7fbdc681dc2a2044d01f135887d23299958cb3f0ee8001a3e7f5de61243eca0f23af8daf10da9725383e75b471799bb1f635637d32ff7e67549613bc0e1ee6d543e5db3d6f05cf821c4f2e6c2c2277dcffcd4a8a434b3b42d9e51149cb06a5ce624352a5b4175919a35b5b71beadffbd06269713f9725e33b06603cecd52e38f217fc30338a003a794995cc05110045feadac72225b834f611d5c97fe0ba1ef0ad7e940b8f27c613f3c67725648683f2c912aa89100ae51c0eb9031ea6cdf0e436e6f40126e1385a8b1c3486fa1c29dc0b1f92483c6775dd7bd167345ec409cc89e5d38719e238e9346a294fb526c8b5bc9482cbd2c74ca516016d4385144176aab720af0bbbb4afb26ab0f208e468ee9ba39932872b80039e9b96736ca28524d800ce684a8e506399c3440bc04f9b1a9dd0a0239c7111431e47a17be7ec99b0b580bb48be1df48f1a0ce155338648790d1cacbbdd5c78f2f6b1e655c270ce35bf5bf614fd7e0e27d7ecd767e0f1ed5c069f2dcd44bb3c33c04eb86cab8a8d340152d55007285a1b65d38ec2aa4146d8f70c081f58600dd1e28aaaff7e7d53099e27d28748a953c89a8af899baa2fb0c822f3837f5014e4808cd353c350c5768b0e435a3adf219bd744285dc22595e2c3c044447bc3a9f31ab112e8466177be50ed3f242bb7db73734dc2ce2b075dde1e840d672ceb5459925daa41688b953d2dd2f8c1dd97f17f15786848cf9f393ac6fa649159098a616db3c463591399d22516c10fd52e642925e9ccc5e9149a1f8294ee6d4e5b294ea72653f5380d75a11584bf8dba78fd9043d125341609bee231820e8c971b7bf57498f83f6b57e5303998a93823c8c499750fd50ac29fbfca30259c0e7fd4bf38e315aabf0e97a2e1b4eabe5e13f316fd18bc66842382b0659c9d327b669fdcb5182bccb9b2a0f9b4813ebca7c12f2218dad49a301dc5d0b0eabf8f1c230836df696bbdaa187cb40c2b9cd9fa3847903ed8b60674ad3a7b79836c0d7ac2114b34b185a1dac2820dd0058af59d94217069ab58b2257a66a4ad7e3b996ac6679dba411f111ac1dae529e880af8a097597940a8dc21af0b26dcf59d2bc58efdbc0f649a0124ce252aa0809119cf8b5aba5356dcfcfbce7ddfbd6f5fd4da725fe1adfaaf6cba1117e8a227f6a11c78e424a440b0aded2cb04c1c998e8b21c01b9ecb153e2199638212c625d639f2a08d85b53a76addd67488a1a340e09d0d01e672f35408f9c3dfd9a253f2c1964efc49d8a79bdab7a37793871b5a6d5dd2bfe86bd5a5c7c640961545ae15178de0c9a0e1997e61eb71ccc16a4ce5d957b19a19da0d9bde3266ff76d55b05085a92296f4dc6d623649f680ddf40f51bf387815226e4b894999ff11881198cac5da39684ad3b60254a9aedadfed70f768ed72d7dcf2df316e37fea3b6716ce09c308f6f523d3e52c2f8387fd91b7bfd4d06241e1971493812d844091e669dc0b6359b9c70cb916e1304ff1a1fe3a4273c3e889840c0e232a814287cfb1e45e57c8d304e2a8404054f2490757ce65bfe378d7a9eaea5645cbe09e01889118629e78df5716bdbd4ba448e5440b734ae728021ff3d1d7c148cb15074a592dba16b21d14e68120329883bd578a67eaa8591ade792879b178b81837cff76584b1b3992d493cd493d013651a9305e5f9144f2516003dd89c8da2334283a46eca57efb808272b43fdbf02f07bf1f9a96c20ba6673f986ab6bd08774bdb01a6b057eb04c8dc04482d0a25e382cd1aa168a1bd93136373fe22c9ac69d8aa3c88a74dd51dbc3b1a93ec3081129bca64071ece48055961a36b1e54dccb5b454d36decf8c14c04afd834865b6ca750f32465b52d1d1fa3363de168191c7e4cd553a50fe093dd38e2d0d8f6a09522189ab57df040ce050377a3869db1e2cce7dca31aefa0cf817915aa9564d5d2f41f1d0f21935d7c52229aafc943eacb8716381a160752b9cc22ae25aee991239bb30b82936bc6c88b53bcc5e4ae52061a66d67fdbe05134a6b887f76c5baf89a8a289f3d5d32660333142833904d0bd31a07a62a6e8d2113e9cc391589c236a0f7ce86a905dbe97175188bbd65128ee5d003d0e7cbf708c4f267737a78fdc561f7fdcffbcfb05f33603d6da56a9ac98462dbfe077759f1f918091afa61dd98eecac7a6863d901a2865612f3d4ba400081df7f932e85e05d492024a3c3908d9c47bf0c2257ee9e04cd02654552bc15c7e50cd55e93a0b5070a81592c6991d331bc9d655bb05e39e53e249b9e720a5d52e568e7a843dad768d60c94225727805b8ecba48bbc56a2dd2bdef1be4717181ea2c05cd13cc6530a77f10758dde8d08476180af70e1daa8f4e5b27e7e7cd997b06c749caa38e1d9133b334c5369d9bbf596fb25da274141ebca511b799b758d154dd5b12d7e2dc33411e32a73960d877db018dfe06f4ed492a336780b678193b8001890e77e56de74b398ad7b78482827fbc042b74c1af68ef30fcc3565a3276b756a5dd71499a1dafe534548097b6a4b43d2231d268cc8a4f5c3cb55b73f33be2f517e2e25f2e25c1261f8d9583704c820e2c90104a68bc8c6dcc8f118928cf17897ec27d5321714ac3423dd06f6e61367d215d3a5255c83d4ce5465fe220c95013c94870b8727db4bb2fd964bbf6cd0cd5833fba04eaee1a792593dc3278cefcc534da765d57e5e102072e5714c92f878d8290edc8fd961eaa93453629f67fa9d3c010688008feb34e1dde0bc23fc406e5f2e5672c1f78df71b2f769632a98a7f66af26c507a396b00ad85cb9ad8bd7a1321712abefa6b3053158481bc905d004ec764aab5305f0243eb90429f6a55447855c10d1d3e0937610aeb9f255d19465126ef78edb3ebb98dbe356a8330f09c124da697d6540241b30a6d3e506ccb0628800bda1464f97282867ad029400d2752d31a07cad35c863f6bd14072cda5e0d7305d8742d24dd1816af05af4d3e634bba202ecd3f8afca9a9de315e3c8a9b986d21ad6e59baaf67279cfe78e0e6f90cc74a90f23ce9eda4e98502eba1e1ad3287393993ec51a85d26518078c4c0bcc63221f212fc9c3e8f0884b9ba8d80e4c988bde0d75107238f407563e8000255a99e9844346d91c37ab00c4997a224ea3f7f22f026b8efa27d96acf23a9a8eabbf90f06cbd47f70a63e014ddfcd71ad8934a94e9cbabb91f6ae98bc6431983d9547a7297f8d73b68d92c1c45caef22a6516d643e22d4e93dafe9320586fe6c346c889b2d065512fa6dbab89101ded33fcb41e11aad56917d79e6ad517fb1c41986a151ffbd40b3dfc096506b3c1785d95599eac03665ff21f22109931d37840bd1386011d83184f446064c117c254e64c1cbb8e8ea3a14d12b1a852f03c358940f40271be91d3563ca63c2cffea68431b3f5e1e7f6038e8c5e3fbbf1b4729fad0acbf3ccde55147d97ba93dcb2c066209ba0497b8d8098a5ea568cd8576574a9789a15414cc2930c6c12887825698f3e152675c85a8d7b57981332dde97de024e6dadb9d1f4f72ec36c8c950e9f653eb0573f71ef7f17c108bfb7f3256b81487ccbdda645b741f4a9f4d926af8e4522bbef057282ff5d24520e08ef7252a01b847e125c8323269c1cd77e7ea12b539f82f82e1e5205b47c66439c4bd7bc79d067f054362f8540f5f48060a62bd8a480772798dd4dd78ec0c8ef90eab09b5f8a0fd24741b40b43011d466a008d6d3c9664db9d1406b64c622432d758cd72b3dba736bce147725d4890d9bcda4725436e81ed06866758f74331e0a19bc80d57576425cee126899eb97a51f816bfb26b2f7e7400091db9dbec35fa49c57f229b6c61e8fda2fa2270b722aa95eab165a0aecfb95d6624b1861a0500308e6767f47c7f28f98849360a664977db2ba9942839f45933ab5a342c08ce10cfe5483af0ffbb47b1340dfb6dce5302cd960cef97b763e662c68c2ffe27b0616dad5c93443cb6776c0506724c306c077aadfab31a4a97ebd040ce0a2557dcaa1bdb4ea56823555d4ac49cb06db95c655b79ba45e3ecef26011e5cd5e43be4599dc16caa482bf630b33c2b38dc26acaa1f641fd3e4ba89788ce75c6e34d933f7a881684c777855f21f5eb25396097d0c17054b029e63c7b00e625858bf507573a9c441b8a40ce9c6033d7938f0fd5445861c280367109666007a13619;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h5663a1b82a7d9b184e03190969329741aaf9d4475b2ae135c3057a1619b9ec58941770fc1121535824e171f68fbfb3c59b841229e566dedbec3593ffae4e66882240ff28b7c2d89a8eee907d4b40ad76013bdba68fa6c7d7bb251732df3cc9c5bd0d982adcca409809b672ee4811e6419007db4012a5461b519f2c508d3d6576cd2a03e7ba30815ba619f9e86bca069e920f4414e9698c0c64c42d90a3e143a803db10fc01c3bf3fdb30a9162298f2bf9cce1f7098e870ecc5a5382963282d4266a6fbbe40a1e36cffe129e1c4f354f4aae4059614e27ac5a1027663a657b5bec6ceb9803bb3b8e494bbc67a928625846a2fbd716419807a074b929febd4f13039315d3a22102c5d983106c579bbf1c3c845b32e797639ebda71f805c123b03c58a591eb387e8bd2ea9889e3fd3f486b1c62dfd573371319fb023128f12aa94e9ca69d168fb0035c9c17c24cf4a158d80537e3caabe27c8e16c30a0b1f5d2fdf6c018fd4ff7578cd04cd882765ded8be8bc78a5e3593e9f498be86d700922273faabdb20bf112c2080874b1dca6c2575b43b06fab01964b052397ca297a61d833b727f18aefa833d4f7769f83dd7c43bf98a5df43ceba4b536b8116a594e4a5c14dbec5cda4fbf55b1f8531dfb3b80e68f521da591e8eca682d2cfe97cf4e9a704dea71ac97732f156d706f123f857d5ca556dfca20e46d9f75600ee51bcf558e58f521132751584f27123814df0c85e893077b96647aa5854eba2648f6a27c7585e7bbc05ccb5b0154d2fbb3a11d5bfc3cdc64abb51aaf7caf6c8d510e114b25251aba411df4d8bc8b0f8a9eeef0a5079b012e9fce994304a60063ca81635c02431ed2b57caa61a8ee12db7500e43de6667cc1ce94e3ca6339b51281d2032c513a136e5d466f8e1113711208612e5ecc77c420966968793c4fbe406403be754eee56ef35ccc2c514490a3301976d52a32fff8c952963cacd5dd13bfdc9abb9e9d337693fa4d9b662b3002eb7e035552d84d1e6d690f56464c4510a420d26ef83105d4296e915fbc2a1d8b5f5e39cb6e9f78678fe763c0b40df42c2324bc59268741c6de2bd691a4377dbfda72d56ffb9ea3a0436ba4f826b5ec96e232cfb1cd9b2e4d4965b3015d0591b4369146cd8fe39c35a60d6bbca3620c2c5fa45f8309f05678531845ba94c2591a6b30bce5cc332687d24661f576d799fa88e4faea27ce3b4424ffaa381411ed439ef6fa4d4ce6cf65a96a5312d5f4bd5c0a6e4690b5db474ff5d25ce97cfbc854a67408d0bb18afbed0ce0c5f43f74335398230de2b0e2a9968fa300069991064958321b3dbdb5cd160ca35d682866eba351f5f3b94970843e036a82a8cc9904b8a6b744227b94bbecbd23b2bcd68e57d498e748eea2c1011e14676c25b2d83b2f0d58dbc6054e5b3a9171e98049aa6d5eb035af6f0e36ca14b667ab7ddb2a70ea8b4de8510e95cec4a1923189930af55f95f92ac573667dcdeae956d11a649c539de103c7cd31a9d43cc196e9a3413b1653571264cdb798f409c3e337a36a022962ddafe778759f31abbb4e89163e5d294e0aa233a7fac94abe3042b59bca027b6651fc9200dcfc628d3ec38bf3c4b2b334bc1081a6e6abe7013e35f9e183b21978923887055d8be8719439a7b065f417ef121835b58dbb5a1f079194103a0ca0295b999feb26954971c6a40ca602187715970283bd9decf524c7ca89ade1196a930bf6c964a3b5e44df56111759d9540c9b20b860dd01958a19f69625cb1af5e7bb4d41c02aa241c5e9a3384162be4706ed3b7852a847148c902064286ca946289157146b97c05b8fe512c9e5cf613437befef4475ea8d3108c55ef859d0d34a9b824d425da0192eceb9844b3aee91764e68024948615b79c145503a39465176e1f9996ec28d0a38dee302efab2c6537ff419c5f63753c08bec4a6ffddca434ac7b493c9bd8fb9f3e6dd67f05b4deb743fe76a27816ef17e9770edcc9df7aeb87144483dfc75ee3cef12d754d4c7aa3d20fc09748a4ee1a29aea61e1bdfc5a4b7c4409269bc30a371673be601988ef96cdd6b8db5fa8d768f9c3fe84d313c15c17fcfb103103a6edd921cb1e9b295a2d6fe0c967790ce2d34be15a7f479452b6ff44b162b01a9b6ec884a3c88502034c3be013f8fb4c6f7fbdb9b5d989f93baff4f8c1f3528b4fb8fbd7cb55529ced4f07a457e92581957bb0e873509b740150cd79c37bee7f2d637137059bea3e126a6eb3f66cb6433d4cf07df708745bb04324e181272912c0eb7a772010caca2cecc6b1c4521dd48b2d37d9baa45942e0186824f4c041ffbc14fb88536fd49f162b391a7337dd075465643b8017586e0a018651e8adc31acce714c4ec335c76dde083951732b6358c57b307e84c9ce277abdcd91166a58be8b00bf41291b6f334c59c9a3240e47e7c354f7dc7394ec1b02e554152d4177149a697dbeab546c622c9cfbed7389207000fa75de261d70aeb17263a9e2ad0f6a0fc8dcd718f3c35fac5bd18537e44d8e0c2a98968aae389cb686d3aa023620eda07cd94f24f25fdf333b98dac2d532f322ca1e26e4bed0a43f01d4bf8275458e16f163c83ae031bf47c8a70d11342250011d0f347132107459ce79672dc2e2e4528fc2a5dd44834f69057daafbee994d9b109a3a728ae54c11ef87ed969241a0cbe02330d3e9140da1668f4ab0840ca5df3de77c5600cd2326b40ac9a3a100b565cda81f037b54292c93fcdb85389567d34bec9c8e6e8a351828a21b4070538e4483b159869dfe3468e0a77bac036bf5df48b00e409c4d8a78601427e53ab4f146bde140f43788deb9ff15373d7f6640fe898fd2dc447b05fdd8c1e42db8c6657d6c8aa668cb0dd39e3c2b79cb86a9f5d88ac142af715be89300273828cc30ac292a7cd5c612796ed968f175ad6924bb2a314417820e8d9196e76476bc39a999678ebc80eda6eb806f1a91f83c06022ee4b258ce037f4b0e1268aa59c453fa14f558186fd6d04e588e79ae75fa9b31495ee3ee7fc165dd87113a7a5d313c36eb2deedd05fe1d375abe72a2e4ec78c88d20602b3e5227052d08e871b01a67997151052911fa857ea2800d93f4f0d1f6aa6ad5992339a948e19a2d26df86d606fb539b22dab47a2ed381cca7e63f2a067be7e95e543c661dcb5a9cee87fceb85271154e1e0f837ecb740694b8e054cb5471b53ea5238b87a2aad1e9ffa87e90ceaa385b3c0691f0afb07ee70222d4a5bed5882c1f9856ff37218dc4346b0703cc3e65407d65d3461acca8889ba832c6fb526fcae558ddbc806e96823b1388ddc156d3b535b709915b82ba6b973116d3c4cea830f9f3d82b3c3dfb146c3a534528dabe75328f312991a4dc6d1251cd9a51eda53ad0c881a0887c4ba884fbb3bab587198743d48cfefe5b59f5d48b85e9773b9f03f598db5883144c18219dd207a2b384ced90e6eea4fce77c60d10cc534356cd449bc7c1f4899ec77096a29d8766c4e26b7d6eb1b9b2b56be737af66d6998301f47f6146fdd10bf1e738c46deccb87014c65ceb72a546780de3c03cb680be01f3e78a22f274a28aa105cf78f7a83aea5dfe3ff02751bf6f17bb1f3243bf13f4311a4f5e189ffe27c18a34d43254c7b3871f4b6a290324157ccedd467004e6fadf3935944c6b5ff44b6c78ea51d791a121789f42cf7d1cefb6a840f29655014fc7f918fb2bd2276667aa9cdf7dd8e86999ef124eee02cb74c56f63bdaeff5fbbd10c51c598a4e9be58a75bbf6328fcff3d46e29ad2dea5d357a35977e9efdcf066777b5c14ec7e26c7c936e1b2c89281cc2d31c8a802dc7bce50e2f4111bfd50cb05cbcf52f0491588d1f95e5e6a77922344df2a616c50f8bfd7bcee6063992eb65724ed9fdf0a4a59ea170d4f0edfaa7493733150c3ff5c5189fd65c84dac4b7957f68e45fa81379bebb83ea9ce90ccd43a558f4f2f39a98f86311680256cab2e24eae63f312daa4c4c84407fbe181d6c8c0a1cd7c327479b1d6bb35560d19a5c10e6c8d192957865e6acbede616525c255a66f4b258226ca21ed1313c7afb24fd0f71a867f8abe610ae7eaa1788c6da9d2a1c5d0f8818a334ca1ecf8e7db28bac42d2af8705963364bd52e23867dab21ddd8711397c9e211a8f4ba7c81909b9adb8710d8d74e378dd553b956e54752440aa4a45f330b7dfcd22b5cc3e975c1056576c7356bd74bca094b0f4a54aae53a7ef2354c0e41705f0418016de7a0ccfb5b2221fe462a2cd7c73d7a55858d7bd5b387c139557283f9519c38518a718a72116b0d14e82a4263940aef2f403303129f1f0480421d619c0d6ce05a6574f48286759658ce9dd497cb9d898435f3c0e7798815dbaebf66cba5afad572e7b08d0b6217e3037dd924957871474649b1a580074dd7de905f96d80e0060f66de3b0316b69b70ec9106606b550fed4d22c4ccd08963830af11fb000d35e016212fbc5a210e7fa24007941b6e30f5c0bc660f7f4bb494dc543e298d4d83e6011acf06a9bc1770dab7546b19f9a50d6219f1b6fbecbd09e25684c59f76f2f25c2ee7ffabb311cc4e82bc9d5e03a570507afb4248e2c1f807ac2f7f1d94ace78e18d22e63c8468e65f1e546f192200f222397759f02df286e25cf910c42624907ea66c864d5d6de4aef6ff3884bcb461bd9bc6dd3c5ec1692e0555fad447ac0609e9be3b8f99dceb4a9c2efb724f794143bca36dd9ebde72908c98a3f7ed4f212d2b9781573105186bc6db1e5b1eb278d0157106b6ba7f609fa322f1d0d25345b4ad0de1fe49dcea964f067991a28458170b513c3a02602f38248d857402fef1aeceaa5d56f5f4a9378a6f99e5a7c7e9985a1c09def2570dd791055641b1e10d8a6bcba942fdbb38617a1206d88d248b922a0318fa794b65555c3653bc83fc38ac05120fb496d94f86917afa699fd07997e4f557ed9a784ffe2a412d411f01d3edaaecbe5bacf9909de1be854b5f3a633bccffe7942a842f0dba70d0b2be0d5fa322d560a624c549d06bffa2c74d52f19f55be06fc82074e7bb48cc92e7091c680aa2f434d9a6fc7e057cf15c5b31e9077efdd2265d62b4ee4e3402a6c453792155a520d8aa73cc390a57664884dca87e8d5f4534f2365c815572b7558edf76a9c8f5b7f9a00026e8820731e72fa28b5677234a777743b0a3787ebd25ddc29119422c7667abb0565f2bae7e806655360ba9263e4b80f8b697663cb13381ac1c6760bc6a07b797c80e71ef2f99272b496803f587b178a97f1bffd2d98063dfa4de3f03376edf6de06a8f9a050f0958bfcdd027d945b94d967f9f29002c12bb075e9edce1b2420729dd7017177436cf46ee6eccf14b9da14ebf3059108d0979b01add9271c5fd96b3b38cebe9bedd606186d8509a43ea288f29c987c1320411aa5b91e6890fcd080576d84e66fffcb515f19795324e00e2146bbd1bb2f547a878ed382efd273c2fa24033bb4efe5e14bfc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h15272935a3307e917a4b80e77ce0224c83255281adf87d156fe0e92cdb7b0f5364f4beb939a726987bf3cf9c333147d66f49f48893cc03e03d3eaf081ef86e49ee5668f1d241543a71f8bfc504f28c42c9b79f5002871ece5c901d42c5a7fc476ab32e25395104af0d05db31bf0a88f032fb214ff4ee3d11684665e2aaa469ff9c3e4f466e444c1e12854ddfb2d3f0488eacebc9ee15664db8377f92fb4782910196a5e512951b217eb1da52efe35c938f19c5215ac88450cdc256b5ec91987bb99b3d666e01f27633d558197935ae4b695fc95272f241160cda5b742a725a267bdbbbd6982055718a1d012d42788e49cac1d9e2e43d7ebc5156438e96504dc03a5dcd1d1b80cb20d197ea9b41f16026b8562cfcd807ce8a492d0b1d6fa89b1587175090105ba3a3db05b091b23ef153147a9e4957108053d1631f016077bdff319762cae8137f334a6d4ac0b76f166c56d0ad1c47595e17f45b246df9a37327ec05bac0b2aeb992b9b57ea1d9a9edd88a4fbfe274b293afb453685a213153315bf32afe7be3bb709535a44e1a7cae2d1a681afe0cda21b76b007474b98903b19c2147ac0a1cf3f2d5d267d248d07911d3e79e9f0f65c48ca8fa982da5996250ffefd6feba46815f154e2bf33f2981a93c746758432a03e1ca124f4771865cc69d23a398e1c7e10ef153277d2af39ac0295bb627d6a7de1f007041a328751eaa6a65ba714e4df280e41165e5d2f109d97d5e88c3ec521bbc665c7c79b9525ae834f2c911ff0792883f3879c726f6874f659b743b1b8a5d91fab8b2054b6c12a40e0ff34ecd9f69de0c79ad3bcceb3f8f38e4bb0e54d73b4db96ee0f1400eb9d775958674924442b477087f26087f9d769b55efa3fd67a492a983acad852febd7a0b1d3bffe2b30d6980c0a22027f7aa661866c20a54ebe5b573b0c92a538bd36aaba6dc1a8ece43ae43cbf98f652e1918d7ba4b387e7975a266cad7b2bdfd9cc8b700535752e4372017901b5016c00bafa78bc1bba4aeb49b9568dbcbe7102d4148329c798490aab3ab6274106d248fca5962a0c74864db6783977dc9a87ecd9aa030ef8bdbbbd9ab71ae98258e73d9cdf3294629039f2de008d6d3ced4782b44f95b1094385d7e4cc60ea52fc881c4aef0069f46b178c11b10d6811bcc03a00afc74815e2c2c21d706c50b45d2b2881f537b1cbd00d2ad825a1be01424209cb7aeadb6b440d93fc3b7476602c6dd7489013eceb4cfa3b823b02bd014a679648da9b30e50e0ee6f95a7ff0f58e6f5455b7d854dcf141f6014583ee216a1ef4fd99d6ea4e8b8a1076b6eb31dd5e10502ae533f8cc537bca401a0c814941bfae6c1999c43f9e183a0f22d64bfcb199c009d3928e1a846e9a84e3ffa6a14f151188ac6fb76878d626aa0003d3f9698f1fde610776c0a65a2fdf7c7048af000c7c3fa3bc5b28c8af82e97741b39d2c1798abd4d2a12a41321c5abb605aa754cfbadc607f0126df50a0cea8cf52637423535ac3feb63af8b4e571f930211d6a6c7e6417ea0c40a222303d5c05a974483dd422a8c853840c91d9c9171276910d949eb8ae79fa44847126ab16089f680dda743084fcf63a516140f55b7bd21f290f4b72ae9870814db2311d63850641de8a8d2a05f96348325a2f15c57978fa4cee2650fe51396aeb089d8422a5f7f5795bad3858c9f443493d3c87785fe17b00719956185a5f3a22244ebedde7be611a36170d92107e7d22cc302fa969986be069d11b3fde2f8d9560afd8e562feaf6e7fa7f3514b0bcc22ea54318eaee7099cdf2b697ce95d1df2fbb3170d022a85a7b7c9e6be18d86e70cffaa16c436dd0adb99b7414fda1e50b80cc884bf80524bbd05f554cb6e665a476031602999a340e4025bb28e6fa789930ed3c529f806270ca360c7103cabcc8e0ce4bebabcb0455113e113ba348128efbe23b948e7f14cb2b58ed6fa9468189c3de3c92669c27d942c1338a8159ccc959d9cac53a7a38f7e02ade5753423b5aafea48254e9e7c1425ba8c04279a9223dd3a75eab20a99b74c8d33b4d920858c7d0e5e932041c792c43ba77c406bf77326e1f41fc98fcbea76b28956edaf57cc27056f672a10444795196a2b3425e0df3e349cfa1a3bb0fdd306244bac9af5f23359776b5f278a65139d26d1c209c9c0ade449157a9526beec0696a1d961865867cf65c08ff8906ad7f459dfae966f0ba713a57425fd4d51ab577d956242c6d01d36e5307905d4cfd1cdae4e8db68be98c9ca6767b7600003ba0f691bcc96bcf3840a3d54c6dbe015692f13b77b2d6289436abae23e0207771d5c5133949bf91a997f299e1c20b593e1623b0bee1f813bb101a0a6fb3b74dc003852f26ba2cf54d310fac152b4cba836b5e356f79f8571e698ff65a0cc1b6a2fde6fdd2d44e492eec790b6df3c73e49d7171ba5f44ddaf3d56e4abe0db4205110d5e27195b781e347fe6679cfea11f1fcc915a698d3bc4ec75d4b2b262fd85f4651b7d9971880c0b112fe57e59bcf44285ee73232b8dfe34efd8b87676305864c1a337ec1de05e8836dca561679540c843c71c8ea2ef15621db0a05c256069febda934488252fc91f02faf491720b55eb0311777be0971649e0fd60c65aea2701fba00ec0539f0633051c3cd7fb11073b64e7b7a93c3c2e3fe0b2ecfd4820045d907f42ed1b85601c57296eb4a5cfbc9fe7c3568581be918d51ba0405cdf7fbcc63b5b447c3bd865df3ad5aedde80739155615b8a26343ad68965b6cdf68225f43b426727ac75591240b75660ee1949a79372158f327f72be05beee075b97e72e7cbb9ccdac9da31df9a70aff838e54d28ebdccee743e776c89ca435d9d34160a900bebe0ebb1a6d41930819789dc8e0e0dcfa0e064fe88dc27e36e4e3c3f9c5e87f2e9e1816597cd73dc3837298d6cf56fe4f28280a2e2a4e514b4c0996f74b2082f106eae3286f384dd7388f66f023cb4e972b5be1e49300eef3b74280fb367af765484dcfd4b86c008b9ddc365ea729f613a35efe7e620a125ae6c2fbc43d8ab6ca3f134e684f5870f319785626d26de05043a73bffac13a7cf0667a6233a0fc8d22dcd4140c82d8a1c9e80db7c19a52b4cb4a2030c6e6f3dc0ecf3cfdc9e9067dfe99b6547ce049ba1afb5732f63c2aee7caf7a81233c280f5522b80d6318563ce577a44d95350571fde3084e625830bbf6c1684ad33a5ba9a925ad779d2c058634d127d859e5fee798ab78ac28a5a616d0c7cf9b68993d17a2aec143b53bcc1d73cb068050885ebba01ff1c63903833393ddd501f161efe8a96a273aabcd9f62e2eaaf0bdfcdefbc379cacd69dd0ed80039a45fd0c4d90d642ddfa9ee67b3d01421e77f1d621b8b550dadf0286af39005c9cbd250b767152104f5ea4173ea95788089a80b3aafacf72521c2fbc322adc3e08e1166b29d175d34e74ddbffb61efc3f8a49188019122aa3a65e004b6a8ee8103742e359ef2265a9c548a60b87184cd693350070ded07ba5c1261257e3e6626b4e6265081dc19b050946461137cfa5d5ab662c5d831b8fdec79d0f7dee8f37e7c2e1e4ae2ef932f6d6b019718c438d18e219777944113c5881fed25cede9c50a02e7b2c0e835b1a1086a98667927d6a6071de302bff988e488d100856eb9d71f63a87804781b6a2aeb9da85bfa99618ab5ca6f065cdf1861ec57ee18b76d11ac1f60ac183731f3236589f9982efbe10d7e741fcffe785e2da4b09fe64495547e6d3f6fbc1e9b3c8e686e7e725c98eae2e08c103d93272856fe69785263a3cc36fb0965db895106a322e24792fbd14a40e5ba62584f1dee5f319fce69a67b5667eb2614e755d0cb3c692246fbe5cc64e983ae4b278f9362973f0512b87dc7832d072146306e2763e94731056e9909ebe49d7d7c83ac1804b9f47395731a279305545c2ea9a1877058bb2c9caaf48b10f8eb44453c25a1e4aa4e701a855b5a84cdf0e53e09676dd0fa6cef4eeb7e8f913b9a0d0a968dc5ccfba4392bb1566efae6e37fc8f87bebd4a01f3d458df5bdf546d0fa2d3de7a89fd1c1c22a65aa83a51a947e150e6f7d49e985169c9388ed47281b9298af0c993f9ba7e1e95c7bccd9c821d51e4cca28621f167d0708695fcc5228b34761cdb758bd1847ac523c7841f82f18cdfd59135acfbf0d53dc07c6231813db7b51761b4a7eb9b0bb7ac03327e77a43b8521aa9148b7574e97f413c5b4a94bf6a1caee4bad8f7ac7c6f7ff4e5586ecfa1f7c024fb66e6abfb18ddd2aaeacde105ac24fadbfc86e0bc4826b7883a5d4f796c37541b6dd8432b740a983f0efd4e61e48ab2b4958df5d1ebf745e4506ba5b7fe5d8b5afff8f038bc3921e56d43fc869d06917b8dd39fcdad9267c8c1bc7c2bca5914686065b566ffca0f53d03abc7d2bf2bdbfa6336605264fa5fbc3236f17f0f6474dff2a2897f3e8407b8e4f631380c6ebd12ffbd55cd0690d8441dbd0397f98eb4ddcda930a6cc47214a24445d10b20ea1b978a5fff4c3cc19d9d90c66a07ea4be5c970e2a2be8dbf9ed7e4974a4a3f4629135e52c785b70f68c3633e76f7d33d09dd5513127e8501e821e33c0c58b6e3d47caea7c991c2f6a3dae3fafe3a3c82588b63b40a0ef1aad4f9c34f7f4ccd25e29b46f2ebb2f78bc04ccfe84e417c9da7c8164af030fa269b7c11fb37e804dadc5f7b56d2b2f1371703150a245b4d071ec9716366a567dea60be4943580d98761f9fe8597a0d633f18ee65d6709e30ccfce685a1ffee3ebd0bc3c10ec356b9ca4363b79f7689ad35b9c50afac60f4b183082482fae29d25c1d858f47159f5be58e4d393e13629a0b895ea39796274aabde78a77f597ee8c9bbd3a9bd2cf086b66a22193e6435dcc072e13cc12896d1490713e5a9e17ace498c0e7e12f00b440b4a7cbddc62254e0fdea4cd66b136405d61a2de56eb9929164299b91d02cc5eec14e5e50c363e2b658ca6a80d55e16ab4dca57b6bb483c2dc220ad7f0cd9b4275c29b98633f88585c769fd104adceb46336f79e3afd23a4398cf434581a8084ee395ba3e6d486cbc2033d7cef09d28bc98519aa45524a9c3aa4d37d275ae854da68602962e21cb47e43765d08625d2cd65d87c87f0f68145ef0dbede292362cc6a48c84e9daed79ca6ae59ccb80769f1a7c3bd2a55d43d2facfb54c4e5882f6890b98fc4aa1e7fea8cae5794b9aeb952e14d28ca643221b6c5610d3a4da2bc5042a6741f3cfce3e17ebc106b466c68c4cd766eff7c847ca5193e40dfc04e3c0c0bc8ab69abfc82d905d1ebd0feb26ca808bb2fa41b208daeb93af85eb6d6f047d818e436af05e018ea511d01b3740f1a8dc1a5e93bcee7be6bed93da3ea716c8aae136085466e0d649bca7753d23a7e89a11a0975ecae576bc8eebc6433e6692c3c470281b53d72d6b058e40eb547e75f4017d06b201373336ec996b6211e0b9ae19e0e2604ffb147d7bbb83b9625c96edbd3459776a2c1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h749fedccb043894189575a7ffb8acc482dd761c6c39ae74bd13125a6b4742c639cfcf7a79527233bdd3cadfddfc2c783d5a47984305caa0169d1ea63d4ec901ef6e3bf36f125125cb3f2c39d27702ebcaa6e078ba1908c9c9c635db07e774a9e4c434586e84bcb516f7c3bd0492949cda8b8704015375924d8430e0e1d9043532156a2a7ec5d3f2c4db76ac832d5c54154261fcc3db5e5acc43108fcfdbab6dd1938b46930cef0c4f59e5b7c60c96de1bda11689ab97d66c6135c6f7abd34ba3e21d222be6d6c0b4a1704724ca18e5f527be5a61173ea91a991318aeb6bfca64fdb1b69efced35952648b41c7a7f44cbe3622428a0183248812b1fe2095219f6fb9c2a3e7625d0a210afa483ce042fc14a9af9113f7b4645c48552a4b550578104b8e08713b356527207f61a1c92ad38dd7fb74fbd15ff3ce279014fda8f4de2eeaf7ea05d428ee9858d5b978aae203b638e90a399e4644606281dd31ec15a5e07265b419c37e7ccbc9a38a0417330df4313814a5af5c17be0bd95e2ed35eb9a22b8a646117b2c022566a4260c751e4f70c79105271bacffe4139ba2b06e0ff3bfd24a3f8a800e2e4d66e81437965fae4f826d45a1c0e1f4414170b0c818f59b7489546e07151777e4ad6514274a748104b135c5a732f1c5a06d418c92e54f5e3488b157a6c3c935497af311eebee3f30267555887687911925abf145edcb6305d8a5404f9ecbc8be47951c6722aefa1c4cd47ddfb340627f68318fc9f855cf823fd873fbbdec2e49e1701749de5bf919128dab9661ae8835ba0cd37e8297ebd1f2076cbd9004a23c23b36f23e9a96c5b7137760a2247739228264d9fd87164e851568180a8139229da2e9a4a44db64be9d8b48eb17e97774e6800e4628adb1b59bb04abf44de969f2456063f96ab623e451cf8c1659c83e866ac052d582293c4c49e90d6fc37632cc883fd0deb2542a4df55eab7f9fe23edd771ae2cb0802c97a570bc1012e6cd05b67e9ed7861f68bcf5d958d6fb5450a7055b017a5904bf6da5b9e5507104d6de502d15b2639e0a00186d8e990a6861dd40097d20c4b73cdd6c4103370b03fdbc1e97b2dcb0eaef9e5815812cc2b5052dd0cd533d4e1f49467270718ecd7619f7c8348a1dba72ca964484ba028d7b6ed89f7641cfaf2b0c46362499ad6cd41076d46b5e333fa0422904a28caf2bbd3eeb0e1e3812badd3fc34c19563ea5f579391e728524e2133bbff450491e50e0f36a87958a97404f0535a832810aba038fe429bd83429735e1a19f85d084e376e6f1677d20a7378f28997edf5c5e931e8db954c6dcc7597bbb258087755385a44a6ba8a9427502f7c6c548a01544ce642faf545e61f87feebcb6e2f41057012a3de89afbd358182df6efea4241d4d46e115c9efca090633dbac86071d514b8292a71e2b5fd7b0b12b26f4e93c72b4436ad296496264a67c7ce4e73b0cd7d5b9f07d805392f3c936bd091048c119cf072838c6376558cbf6a792e8a2725e21b195a1f0214997d3477a41b26cd1b79f11bda49613c36802eef8bb36d35c848b3e407528a5a158beb17f9db0a2e03c1e11f96104dc21fdff779d2e5b3338c2f01e5b68ad4688ea8a371aa6d6d1886f4ca3e1b6f1d45f51ed4302c125307ae78e0e7e7f0e8420bfe6b4d6b152da2238ede3760444bd3061c89a95500296a559207d88124725827d22a18517f5305643b7680bad84d4d307bbd8775bbcc758f695b0b8c12be230fd6036358401258bb65cc1b1e283d88646bcd2c98515948098e53ad91a503904481f81111cbf783b63593a56136d64114de7ba9e526e7dd9d182be37d6becee6ecaf84a6d14ce543ac040b591c6ccdffee2f75604ebb5c80fed1b6b4939b5494ed71bb84e49a81b2ccb1c5d510d049af4ba67ecb5273ed3519ca30d6f88a7562983b257efd9eec909f79603b40a46201c872f69133a85b8e8da4f56af0abd2b638b120fdbb5c9b6401ddee069c90ed919b689e366c4f65cb097f77db5924337c0996ef093b61699252559720d46710607f5927f5aa9f79cc8dbb165f848a0b4eed1f78d4fafaf2a9980f61576a97b631356987404cc961306eee451b4a4d09a935f36c7fd5d6df41e9cfa61d5b6f90bf9fe7d3a9833071cf9be41523b8bd404da250ff42e14b927550d6674398284b061ebaee8d27d9e8cbe90df002f78d5bbc28a5d7bd8703573f7babcf690a545b92de26712c28ddfee14f606b3672968d2fb3a2455290df672ef5b33c8a798f93d45dd74b371fe5c322ce1d376cdae4e2b7f626e69df342c5ff38b1be7204894110d120359350c8b4b3bc2f3ebb413d3814fcc51b6d5ba57c260ed5cd199ded0b0e66d2dbb698ed1effdb19c6d3e8e5af4a4bf78ac8960da80e8ae1475b6fcd2df9d161a751e0100dc6b41a55ec214673d23d664a05b5261a4ea1ee2f1d17e79a367b7f2453b6512f54fc66d0c5c295d8f3e8e0e883370354531897ac8679b0eb7bada7178f7b0f132be1432c21d6ab1e0ed16935520ca7a5601ed227191a51e408d4b119e70d3793c03d504289234a74e9d6b62965666c500971b124986ac1e837b6aa06ac746847754826e4aaf80f538a6592aa902b4f1cdb091e00975b5a7581d68f8e3b488da24ebe07b0e7698dbb24f1af66d72d8c8a23e15c8570282bf0a0817de966463d2a2cd18216b739f6e9c2fdb0cdbb4360db1a4f723f7db434475dcd7b33e9370c4e89169bbde0da57ef630966eafcc76a30a8e4c6bfe26816318dc3eec5ffdcf5c5e4058863ba51f70da2e9c941679e94a96d2a24e8a2eadf524d7e2189df275da4c9c4b21c4830b6ee4094dc4c1ea73504d4b68ac813df5efbff9496cfc19f6b4f9e76d03bb9f3e0a38ced09aa4e3231fce214a52a1a05c55c7ce1751cf6e40e38748c2b25ad5b41813bc8c8b0da160b827e8e308f29710edd9a91f8e7d03d9c19593f67a66b662a6294dd879767f644eea109796f3774b7a193eb4df934ccdc41f3396797f2d23ec429b95ac60531f5fe58a6d6972c432620317dfc1e59d3b40a9137b7fb4f32037883bf707e08175bccfc04ab584b195be656e3b5ac6d63c9651a51f796aacfa1482f9c205d0ec8e0f0f5469cdd4f3a997933bae269dec030726214284da310440ff99159b1ace687c8c3a2dbcfca1296445423bbe3a4a60a638360199e4db4008e3c77a2f0d6bda21b2536edca8cb981b1f493db8b840367164544064e4db848757e728ba27a7c1df12e329a59e42dc72a2b1e869675b1d099467b076f1d5fb12213f628989e9cbe6936987b585911e00549f08eb7cc5c00ce01c670cac6a4299d9ecd3c8850db871d39bdee26f21de93071bd13d55b85f5f772f05adab9b02517e59fd2f5ff71c1fa6afbe7f0198fa7aaf35970fc4d107ecf2e1891434a93b7f3605776a4bd17ce1a5d1020d56ea32b3be35ec1107b862b167af349f0b788e6c644c9a50639dde2f9f7150e977b525aa66c996bd56f6d3bf68671d78e5898814d7416b5314d970fc15cbe6ec8d822b402de7a5aac9cf104cf7e069a9d59dce447a8c02a7c2d805fea78b0df38f6d9a7652d26412cd3de5fcd13330f5f907fb55f59132274236827099866965ebf60e5d173894270cd320ef656b7c117c91c8b958907d950feaa755f9571ed3650ceefbd85482f06d10993df5c2706782626be62691a30bdfa3d09be42aa6bdcb2881c19013332f5063e1977f0dafa77901d67baa23129436fd3a6ca22a3dada7088a39c607f2b38152c9a360446b3e51cdf721b28f0027c0ed4e9bbdb8d1d2dbddcfd5cc5d236d0314bebd8baf5c7db3a6987432ed2cf3ce44c037f8a8c34daba66389d967856500722c4d00c8c3ef0c4c3029910b9a6c63b217de881692090c11e14cd429cf7961f320ce66c137ad359d47354b062b1cefacd3c8ac03463213c764ef5ab7ffe260fd728ce6d4dd474a851fa75dffa72f887736bd6df9b45c306437a8f1d9a257e685f54c346b0a97d544986aaee058f01e2b218b9d745ca370f29b8d36dad923358e9a7855496907b6fbf9ec6b2a526444b39f788985470936a2894af04b035316e5781320086bc5d62e65a644ae0aa466ea0e68c7cfeac12efe31a67357fb43e29c30bda51267b2e4fda47b668e4a60f7f00d723787b2732d149e0af7394f1e0ec431304739b188094bfa98c1f0d31b57788b49ddc89978a8174e47b432d68d920d3f29a83ff5f7ec106cc43dbcc8a3736c452a5e37bb6652d21ac8e6e6c93ad99a5ca6ed6cd720337c8179fc13198f53ee94cad3eb819f17a8e98ccafaf1b160eeaf964531b64ec8d7383a06bb7ed7047005d9159ddd7fd38a2cca106135af08f69ad88963f7531b0488d2b6963f464c65ea1b63af52e0c31724a2143dce8bacb718791005dfce40ec730e0c141b1a0f4c97ab6247fa4450971b043e28cae85e6663f2fe9463c0c9972f614f93f431ce782befec9483bf8d14b5abb3410e496058bcb058aaa39fcf27e49d64c834c174624166e4ad115770f9a7a59683f4aa1051ae98f32bf729c72660b8752d481f2ddc11f01a5b006b8a1844d7f6ee604587aae0da6dbb0888306584b5ae2a1cd07d4985ce7326ec2e2a437f939fa7abef66623e6893fc1522e3f853a2d49f49fefb2d98fdee9de9549ee38a379fa9d2a67e5a02592e689650ca1b9b8414c5b481491fe76c59525c35c155f79b4837bdb166b7cf8902dac2e2078dedcd9aa36b5e35ab1865c0a5499f06e91055dcb8f74007a83d1c72a66ce4fcec8502f8c74ee78c8fa8e5ab41b16d1ece58d1097cc27fcb4cbe468e595a7965e8d6a68b1bf415cf6c15bc7a76d083f0fb3f6be01e2ceb42912c3934e99c43a3f33823a95441677263452cb9e8bd55005433ea6dc6d02f9364aa589ced1d7e716d68f227a2e63f6556cd5b0ae4079c80b6f0ab5c8702ba5fd285ced29c6c1fd43a0dcaa4a860c43dd76782aa59794dc06234a7d3f1f90e3e471afe83e0c21b8ea2ed233d20851ff17a05ffef8f6d406572a9c76f2979639c5edfa4ebf9bd7594248aeb71acae63684de2045ab988c269fac9b8ba73d240e780ba88995397fc733c9177beee8cf5138b7da6be1884969fbb52a5977680df7f6432f95196c6c7ea9e4272efbf152c2c0c16688e908d5426d2f29fff41e4d265678463ac02b5d5e53cfea1f8fe02465320db3448b5b5df6f17ebab58cd8220ac74f9b7f9eb2436b7e6d787cc16754bdd6c7dc3da93231b1dcf410ccda798c034b1c70ed9c52d64811d530645ee1b49d5cf067f32c21cbe8a11117977d5659e22700548940f645d998f6dc8878eea9cbd10b695e1bfd0a08616c2470586a94c5bd92970f12c54655013196ebc4124054559870630127e4ed1b941692e1b5f94c341563751492844986326cd3f1c5f77550aa47479a7145f13ae95929b278beade36dbfc05fea31f24a72f2645d1c0f0a494884f7a89dc355e130dee795fa1bbe1663;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h6b57b9bef20c36ba24f080dce227c6095cac39276c3e29f4895e71b510396c6673abebcfc4a39a3daaa38472ad6dc6ebcc425c2174f916b07a6d982bcf65f19a44b3c091fdf2fb074c6398a9ab39177f7e01110e9e460d386f537128ffe3a62a4e8a1226c60247795c41be233d7e300d1e9d0110661b8a50603a4bab3f8856ec334a303ccd7feb11d7e7d4a50155de71da9292e8bce6477185bda2218db65041f5cb8af485074e21235b0d9dd83845b33079b5a696b857ae696023b8e5d82522ba6d56b370bcb4ebc0f49d149aeda2128639c776815fd9b5e5e5352fe3fc0933bb5eb60692ccc58982757ef08d41ae93cd2775c10c9e6819b50eb9863217583f09e192017b3d25064db075ce4633bd384760830d79d45e9497391ce3ab88837c12c6dae176b0d87f833249e14669a8edb50bde47dbf887f3d67764a38f38991d318e03b40abf129ca07470792eeb030c7ddace3dbbd1ab93e67c06bdcfdac1a86049edc2f5e5e730f9035c75eb6c0bc9271e4a1e66fbc2b7063137a6190e1c225fb1ae12b65bf2f8af444b9bbb03eef5f131d309fea9aca458b5daf5d3e245008ab2016df99f065bfae9395bd6de46284596e03e6291a4ff96fd11540aacef11a4f706b5770d4fbc6d781aa3cba21ecfef0a2ed707d1e9e406852cdaeb18f51ccc6bfbd68eb8b48927e2bfe267a67fc9c284d86bbbc15e63ee417940fd6437b77c2f8e45be507fad81a1e312428721317a2ddf81519b1b3917f3a777ab36451c07c16bf8a11bb188c66648f5e9685c909fe5b59f5d70e86c0c165bf96e17af3d656fe381038e758e0bb47315569939ab74a1db8346f71ce3f9fe93678c70b71f5b5c28c25f86cbec62d781f3e08c0caca7324f7dffbe4330fa7c994daf323b0092722872bdfb7bb321c46615676cc7823652d24e9b6ef3a79eb4bc3da107c604c92f999e40ebdebfa3ec01d333f8decd90286bc92372c4d31fb55457cac12024928efdcb508e630d01cc4b21efdf0be15c58242f0c33d77191f6cf7c97aae2032c22b5568a4c6c9296f0fc362ebbcdaf067a6df3a7cf3d7edf18502b062ddea714914f70536bcee5a09e9bd0a6006874e6d80e6251a4959fef61682fe6db3d6d1902810859549b2871cb55a5be8c614f0aea70f31f352858cb1eb7cbd1f13ba364ff8257d695126bebb7076e03bbf83f4486f4b12e03c30964bbc46515559645befe8012fed554b1224d80357092ff457e5c9b1104b97e393a87709a357afae7e2f096fb53b208a561a5f069ef1a6a9bb2382822c9e6c9f09d230b45c561d3fcfca6ed97617821476b84c840c0e8ec29fd8a80278a7dc7ba445db912536f9b9f0283a157eb1f1c96c0df923d4b81cded87caa7a6e35fa0e65af0794a37a3bc0f8aa774362f651d47316626e3f4599d19c770ae8db6ba4730b218fb5a5b65d21bf0b5668881a2a168528e046e03877078594a0050339167ade021c4c4ccdf5d96c57107a36218e5b818c8f5a6308b70357ef7917a14234aa4dbb758d189260862f0bb1f190719b2aac4c49ddb57a0ebb6ed0bdfc199bdedd8fd7f135e19f8f7be0d80054250bd7297ecce5eb936248d523c4cc8e3158b2916a62a03d99107a42e031c3a16bd1f9761d14ebe4bb77062880db00be65aa63e74454b0d34a9ea51b5a31e249d1459cf365d65c8fedc9e7ed2c058081fe857ccb346fc7c867fe93e7f078b86a8710d7c5c6b6ff180f57eb08e41b20baf510a9a36e2d5df0eba7811b9098f57ae6b1e4f945d789d5c7c8c8f479c124dd4950904435bd3dc18c1db93b1bf73ae6e09d3683a746df114ed8f1c5af80186e14fc737a69b9c9fc5aed5065a711e56ed934516367185b274c5eaf4988ce4725c03ff5df919a05f77941375b4e7ee76509c8416857b5fa9df4946d3d4319495af8391ed3c7c05ba3148a063f1856a0d161c55eae89339961d5dd79c1c627e6ef64b0faf05c2e7db44e276296c43db4e90c78e73eb46bf72daf69c6a7f091cc98c535e51e583f4822a3e58464d698319f8fe63e71c706da37706be3edf3e17dde45eecb0f2bedf8bfe63481a7009c963175f4810b9f43d002f3e4a5ea2ba5fc3e7ecb17bfabffdb0b3920346e8b63f8dde8e42c89f892e81876c7e7255bb0a8fafad08f47917197f7493478ef463fbbb9fb1f61ad11d5e5dfd5b6d2f5601f1fb236845791aa26d4155481d5b7bdfce43e5830cb534b9380b8cb0d75cada1653d6959c0df31eabd93aa692c1ccb408a29dd042ec2b158a44643e1a7f18b96cfe62ad689ee27851316d01bc9a694100bdf6799b933370262a4f95350d4a8e4e8001c443a8e48eb6de0e45b9f9c2fa91af39a04730098a5a83d6ee1c3b53f9e95fca34f4e40a9bd80da3ca758235c8f8c115f10a6e009bc25ba836befcbc9d10e97849ab63fd537359feb481cdcd9235917652f2316b493dc29ff66e1cf852da4d4b5173884ad83e4b8605dfebecffaa9d6958cfd148af19fbee3037c41c0cee07c29cad8f78051e62c319d735f223f51e7927ce7fa11295abe91e723db43751a69db40e5fed8a5cee32da8d8c250ac001ce07fa9788b0ec6b9bec989fd2c903bbb2498f9a5b7b52e6a5ab70d8fe4397245b798ea1bed430dfdedfbbe444be093a4f7294da4467fc52b0f6e06ddd722664f6cbcc04f4bbaa7a111c29b4481be6cb20da35568ed22e5cc2b6f7f313c1d4f85bd4389df2b886b858e9b6fc9040e32bfcb7420dfe5b7d89aa5fc38d661dfed01ecf10ef01bde723a367161351c46ab8242a5c8216547c98dc0c6e93576744fac79583f52a41e31c42184dcd726b298491d52ad815d90d4408746ae39ea634005f25e78f8403e0d602832a11ed9faca894c7acdf6d7c084f25a2defcab2fab7780438fb73b3d7308a9f2abc41b29d0581ef6ecd3e5be2ed99179dd776e729c61aedc1af990a7c3fa38e9129f48a389aa9062b2f413114d64bc7c183322a08d0939ebe67e60c259b641dcceaaba9970142a23bf572234326c9a31a907bff289bd8704de0f51e143be564ffa7e842f6515372ef20ea147e762501cce3bb92198709c5b8cd687840cd803784d7e007ce642b9e22e278bd67c4226af7132b311f1ee56f3b4743c48ef41d0a2217a27fe7f32b4a9813d30ffe9100808419a9e00c3322d0c3eafc09a815517c48d5f4d20becb5ee569b7915a39b4f8775bb4d12f6741787ace13a5b2f20857baf01a70f088ac8658621ef1466aed85da7eccb673d26323e7a7815d68ce394218aaac8590b14c451c8a2e8c4b0c0597ea66bc76d4fbedeabdf8ed978390fd821134b6693976eb9a6af137ed7bd6293eac69a3e0c0dab9ff1047f459115cdb59b490da99f846fb889598479c94509fb47965388f9304a86850d3112cb42c6fab89bd8b760f13aee0bbdb66d5f3f6ff0e5cfe40b1b0d1a06ef79f3d87e733d1837d70cb6796e04619e9179bf9fff32362810df1f905fc9a9a9da17fad1c4a51bee4752a746ff839177285d3e2cd4196ed316b9d343aaec26918c802e73ca72fd95f0246e4ae3d1397e5105d92544204e89cab456c16b066261c295bf485a53cf6c51eb25112a19a7f502f243ec758814f0dac7f8431ffe28a1888fe63013e70064c74ac51397e4ef1491addd3d8a804fe255ee3effc4d94a66d6ccf87bd7f36ee043c60689eedf5ad0f9a1baa3d1dee470031c6ba88373f444083d87258433ef4ea5b0b6a5c15fdd2a562e99eaee56e17724a6ec995ea494f4c3d5a5289e7d7e0fee8a6c979e3355f19958d8dc9547fe2d772a00b4711f24da50a843168149d902268a1fd2c29b0fa7a59e163aa585a07fa75d70d0bc6aa80ff140416235e3d2d91387eaae843d8ac29e237edc92f53b78a2bb3ff499e8837dcfe654075d64c7ee5a6bdeae921e8670d47d5a05ba8518410cd26eec124c46b564b64ea91f61e5c565325fdeeab7f6b1beb38ffd1d554fd728046f9f5ded930974f9a19f589541be81caf7b9bbe3252dfc641a7a338fc7c956fe6e56c6e42a9872a3c95293a64a064142a97f0c79ee7ba9279113405af5d9fdbb41e097a98266088e13193b2b0cf75ad739e16c886bf8c01b77f9f7e088317757721207bd694e6959af0afc9cea27a5126200f77849ac7e68de0495b422881e2c31032814cffdb0f07665252aeb77276c08c2246fd9a37c147f1aaf0d3b43adb88d247614f60ab0318026e54b7be894fc0f5afc80134b9e359d2ef3ef93deffc643ce3d6ca92daae76ea87275f9130bdc21c7dd010e5cacce54ac8ddcd81e3741bc339dc69b2f6dc106bba1bdae6984fca3a4dc10b93c977a89f0fa59b5277492c362046fa821786456c404dec5a66ea3112ea63bf81102597cab1756214bb7de58c8fb9bc73572666963ae056de803ef09d3e2813ddcacbc1041cd7da680ec88b2e43dc4a1465f6f85973252132888d9ad7aa83f02db561189d838ad9a25a78a356b712af9b21a124c452a0fad7d13ca5574bd3257bfa6806ab3e284475d3e5ca402b4c214cc905956b8b279c2895dadead51e8f62012940cd72495b3ed4cb658f0f8aee6ff545dc54ef12a606d5946fc9d0768835925fd951b66657a7c5a93f3f79d7c7ed115feabcf3e58e9ba19c7a07a2853f0ddbe33904e141da80c7d1c0e2845d2993ac486498c64dde0371944b4f3ce50d189dd17b743f887f172364a8520140a6911e808cdaf0ad25c0cabc53f4c6428180df11a32b15b323fc7294734af9e7de61dd107e0fbeb26533cb35670c288715dee653b4d2d8931ed8baeeee6a2329c7684b621474c66e8ccd3758fb052b814551024918ec9e05c09ba793bd8c9d22c694c47151f596fa3869992f18538306759680c59eab5123baa6bb2ae96f9d4e3be40b3eae8c144bccd587769a9f235780097b680f6f8be9e29d47fee3a15aa75f3746ea146d008b80f2da04cebb44546cd6e81cb2a68781c9d74c44cf01c7e221e215530d90838ef5662934fa797663e2f844d73ec4e761f4556bf5aa391ca50026eced14acd18c92217d1154f8503bbf3163a8b26c02ccaa01357e6ef445f332a171b1492579fca5e27095aa1dfde27f84344291cc1a35d6b9b08e84d88668edfab7e85dcb4a0d102685608ead515c849b1acfe846469d1661bca92c01d3362cb81a1294c85660e45eda3165c5fbb0d7fea47e7ff610af468cdf9625063cd6f2efbcb44ddc2871f1f2617d54a852c681942ab81fcfde71ee7f060b5a64e58877b675b3466149df8dc607fe8b090047648b9d59b64cd7abf83e77ede43e27833e66a511190a684399bd97a18d9616b9e852b1c7eb0b3595de01f119bf64fd7a35500cb7151fd1e867c24eba51623d29ce9f1f314157bf510e6af38f73b3fd256bfbeb60c5d71e887276028b9ef1f2c44571b6ee6a9bd0faa020bbf9bc47e48cf27c4d624794e7ba9f836feaba7850051a6fd1f688e596fa6baacfde25750e65238fae7dca2cec787c90a033a15483;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h5b48182e2cdf8de6264d21670f7a605b2578646771d2ccbe635a9797c2be51aba62f9d5f0f2d543e3615bf8fde55d95c822c7d7e552fefe23b97ac3b59b6abb9d2af6bb4e5b048dc89e61300ee5a2ac304e74313fd6f496126a58f4b8d6fd2d38ffbb059743e224c75385f1c9e72b870a2edc42f8b003cec72532bdc03ae8418c59907376db07ac8d3092e9d2a1660485ae73268c4711220f7ab6ded135837a95ee02ac8b805919c693bc8cb601d0fc56e7c8ebb49f2eef089d91582f7589fcafde06051c477ab4a018421115b1d436d45fbba3640c3988e35f4257b9c9f3e9a7ae98aab1a582e4132c2f89db80a3d04802bfa49d8b3630eeae4344ef69e34b320648791caf88769b627502854d24bbd3999d4f1a3596b6ec45101f071d7997b0287ad1a3babd589908bbecb4ee302991d0879ecc37d65bd596cea41a176a8b0a2b3d9b5837bb660fccb253d2ac4bee02a1511c75505b956aa5f9a1cdffbe9944cea2160d4a163e2ebd06a33f493c81fc878fbd80f2031219a6aae86c25a12eb65dfb73ecde734afa33888f69aafe04eb3c374c7aadc79bba2b909447857ac69a47a7d96c0a71978ac2d3949ea6a6c6a9b720f9f4e208b47f4da22cde59710fe76a483c67d3abd22a0d1cd7b4b37dd230c6c5c2c42c61d7fd339efde9db092e4ae90bf1a2227d7ef291bfa23fb46451c7fc97c400607665536f8c172d7cb07503d2bc0022b10707e3e32f3e0eea5ac61193fc5a62c1c7f7d5fb30ed0d8db5057a97cc63ae91be5a62a54857246864ab5fd86ceeb9e4e253f80dc740e14500bb2021e8769389f943c4f532eb1e981ec668ce7d0ecc80c206e28afff40c5f97f3cf123a46a42a7749c735ccb26819ff9e6ddde1f29bb4927e4dc00e1f4d47502f7905a3698645c204093de3037924a7c3466f906d2eaba6b47fd745b199a2413742da68cab6f933ccb77902f31985cd10dd9e02fe6bdd16a7e0ba6c2cb49c06b7f65eafdce879e40b99975a79ee2df6e1d4c7e7eb527c9d8172f3612e2a659d4269c75f77422005a4fc3aa64029790b1e5a1d4c8b6cb776a3ea017c4d1f4781e3362be97d9b6366aec40a9f49de566e790416bff6a5cfdaa8cdec4f02dde6307d5ce8a49a849a7a671842de0c3bdacda52f75950f321679ac3096fa25d1cef75d34a6c83ef1af0925079179ed9c74b932ede4647baa20c4a873a53b722fe95c17018ecb88af41d47b1d53ead96c89c32ae19743a19324524da58eee845cdceebfa4e7e3771787d121b0847943e943e488fff5a701751ffda6486ab9859cf7b3feb41b2599c28fabb94bd325c8ce205006da1f0c90d0fd9260edaae2ab202c631fd799cc2313e6f9113e708d0ec28c146eb762ce79407bb82ed9bc0d9f3b5d7bf6e1f37f556a5f250c17544f0417e78ce5e129a8cc786e25f36c3e492c05523011aa4fba2fbc4891d3469502c909971685bd16518123e4bfc914dadef48e1de01f90f724566426168bfc99082972dddb3276b553ce4ac40ce331f3c0631b338165bccea303d282036e910024619c8b45018e8b993d9a90ccbdcbc890727ecfac7150560482d301f04be6fc094762c346572a13a349c07aeeae8aa29c1e9aad7b8008b9a240103b276e51e177944ffc21cf37d4eec01c61af90a0fc3fd84f79aa9a0af3200877fdbdb380b8b59424c0fd5abcabd45e86f88f4ec78b7f59a1415b9322541640869c041f423fc8647f388aadeada74d35b73cb1201e8ee01907d2f5dd4142b01b1c7eaca5b138d5008a4ff2fd5447205f480ef3462ce44f4edd46866d42c4327baaad7b1e2d7cca0170b14af26848a97c301aab1c1d7a43472b8273e749d52428a6f52644ead7191af64826b5a8a48084be21d11f9b332a1eff7f21b9782a804091e98d738138d5af9a66e225a866176928c91add833c12420d3290082238756d1927154aed9a467e7412fb65114938ead18ba110aca12438d0fc030ccd1c174b84463c90b47a0b48b6c58e4ed2fb0a6ff895494c3852222c3cc31036cab3a57382eb44ea537f5f9fcfe03201f57871972e7c3c62ac8acea8b85d3c553f23ebb77479380d3ad1d3a20f0c4c11bc262d24e2fcd06d6874c1fc1d1a4bdc45df45146a777d99a60dfc1186036988d276cebc640a1a157c2d1ce588ad3d2109a64a78cbd767ed235079d490168c1462b0b39e035c4767cc78b045ea78a59785a6a7e39dbc053d7548215c65fb27dc373a611da14fd2cbf8fb2cf46503d95c30b52da82e261ca09c652b7bab0dfde18817f24c5318902879b69ba125f5b61b519ab72b5e3eb7d16c2267a96179e67d0bdabe5c059f6e2c95eeac61f828a84b809eff5cf8448e9bc3679c04fcfc1065225b9a8ef35b22ce1209de933823711909ed6c21e6046cf3000921b4b265a1225334e524179a0a4a281e07dd0bd6d7aa50c9c0be5eda41ba580e1d35bef378c40a137fd5c0dd719a34e04e1d4a4d0e478e416773a949349675ae8cfe07551852dac8c71fcda9c1db43185b6727e30c0307f1b957548da634ced3cf2808bf7ecc327e233c582dbb7c26d43fdb9c97112a37860366f2d77379a33afa979f9873a18d8145184b47e71492c5c566ae7c31417c9c5b72b47eb02a0d1f1802a37dcf8bd409f94a538b7f468a2ec9790821923e81ca5597b3aa3e9dee3baa573a8baac8cc61aa29878dca99ee5d4ff1673ed145ecc1b3dbe101326ab4536960b0f0b09a168df5074816e36d99d211e6a5ddbe8897ba4bacab71c96cfa4fa13b102952551824964aa337daa856a425494bc91aa648cbf1e7ec46f467fad1791406c8c128ee58fe5745438469053c05f52067b2895ac927c8465865890f24a3b4b1e2106a5893b4798e06e9965bafd4873dcd1b48f3ca79a7d357f3aa0ad7cfb7db37b6883be6998f4b9bc9383049005ec19066dce5a5ae6de205417aa2ef825a195c2ea3255bf3addc09f81f424205746459ece11cdba4c1b8bde3b45d4f93c5dccfcec77360fc7a0ba1d59c790eeb91303f5aa8cf36e5d0f94fb67d604d0af9adda62597273bd4177340feca2a6b6369ee14ae05664c72fb60623afc36691ed90e12baa82aae81e72f973f3f03507f7c306e2bb142fa99b1f7138656ce99e95a17248ca78417329f9c62994f0361ccbafbab1a8addaa2665f7b67f8119659c8fe4e6eb90dcbecc47db84b44f6d77a38f95ad174a6d043b80bfb7f4a6ef45d68e5f1e06ce9863f8356a065c183295329ad2db2f0b6d302f7eff29d996eec05d40ee1ce0d7fdfdd366fb0fef51436a34f2dbc64cf1a040895c1b95bcd7125b3854934667fd4c41ef0e647fc40ed700bab8f5a804784a6c735a9466a45cb407e6fbc9442c2a25c0a5595a25eb94f854127a5bf76754a4c9761471f7eadf9a755cfa816137606062dac7a2e4582f5441c7bc0d2aa87f1028719dde4c629a7e1cb553a77366bcb4681db0bb830c84bf79ec8ca0f09963d1638635a4c2f8b20f6adcd2fdb7f195c9d41ebfbf56766b2b72b0f9827fb638cacc2996edfbd698f4686af556adf42ddcf3f0722ea1eeda3ffaee5a4aa6ac802dfedbf2e9fd6437870482e273ce9bdf1dc0a08b486078da2767be888dcc5bf24e735e68a225feece03bd2c92b1354fc6c27a605645302f25b9cb4d03d4673bdac819e593dc85ce292f4373b6ff1e334ed832f6d8ba5a13a2a89cd72445c8ae79d78d3976a99712b5ca89bd88e8c38474c737afcf0320935d6afb51436f3a9bda5aceddf2c0f17dc50a25bb10da09c69d2cb0cf0e95e79cae156a8fd090561c0fbcc42e5a9ffc795635a6412a9447e2233ea3cb83685aa41282f0449522d8870670e81753256307534066889c4d276d9dd2c1fe8b82299deaa684033e003e04615ff7cf1793c6be372856a21b92ca469e74857be69898602fa31cb4f2151ab04a496a5b4c07f8dc179b62cab540d2715fe13e9f0e33d6b04180ddca6165140088db21f2f8abd36bfb1af2109165118f036123733b35eabc74e273f1aa2bdee245ac56e21228861c8d8309f851121fb04cadf37e52438ec291af41ac1188855fb437fc7d0d422f14c210ae6f11a276080d117b7443d9bcc31e741428ab09fd8f910bdbba0c1ae8bf5c07e2d79549890b6e7774059001bb657355de2144f19408b8b10814e2f2106e44166b51e13b532915504c0e57af16cd04a2639a84aa9f948bb33f509ac67f1e3276bc274959d9c67f9d23c5bb16264cb69197de367ae771b95c4d00ce28c793f6cfba537063cec6ea08bfdb0e7ff2d5ffecc4382da62b42e9ecd6bb156f6f6f8d84a7cfc89b3d37c62dafacdd64ff8c04031660bccee4583d866e9fcd6ec8a7892c5a8573e6ca7433bc8a72563fda51bff9c85e75f8f4b836e72110d11c1c192c0c37ce113559f6891c0388681496ceaa504dc13b676066fb59fb1c39e3bb0a8a1e8fefd874b445a3af65ace2c6a69d574a75b5037c710cfca933c1c4236813ae2b302a0d3251da3f85aeec928b01b4dce234636b0b8cfdcf16a179d9b5f6240e66a44620ac06219d6d09991c56e765d580c551f9d54bf29701188b963f125bdd81f545eede54b3dc3cc32cae5baab8a52bc6aa964e2e59f5536e2758fcabf381d6f1c580b6c2fd3aadc0792a9fc57b271a5130c4dc8cc73eb2f54e0e2bffc33670fc4961967103e64aa73f19b6836a7fac36574e90f42e0edc8a5fb3b27c9d64ab831904eca344d49b787a2513352193b5d9ffbd5553393565806f90b5fbeebde3f23bcf7718319dce85a0574e6680c3698ae3d24e0d0834b469631ea8291ab88a73fe97037fce2fef12c3b7137a3b457ca61503756ba01a161832237f8554bc4f26e40e50bcd9ebc1b3b9dd5a7e9c50e9aa3ba3173f53086b04088b49adc62227efdb9de65aaa7e85106ddca19d41d2daf1327facc388324b450b476f141c4cca99ecc421b84c2db306a6af8e8bd65b15f79af83790d877f875080e8524f93e118ebd9711e2ac24909134d46e19bc95554b988766611397fb95b7b11c3bea33b3ad8ca38c952903a79c1608ad17baced11bcd94d9bb8db2269dda9170c90f90aae2b5c47ef450f85bfe5dc1a892df5eaafd063a0564dd3369b993efefc2ca2376a0e8308517e049187ff9f8331da6fd61d025654db696bdb075006ca3ca9773ec89e41ec7a6e4bc36189c54b07221305c525949522e2ae3f4f597bf9d3f9d8920afc39199910663c99b92a02c4c53a41479478f05a218aa337e412bb671f450323951a29e32d0175662312a51262ee189b6e4ff418d999c6fb3474d004d0cfc06d3620eb9c2910f6617be71bf32ce0c5c2b078572236da39f9b64754ab167037cfa97dabce4068864bf8c79812a3353082600efc4dd6759481353be480d06be5c39d419920c339df7a8e15ea41ec077abb2eeac9dd566b98e981d7218778290b3934e9f6bd17ea267ddcd5a1631f7f95984748d927a10722133599a07aef13c61a69d9fc88d66;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h8cbb38afff531b24ec25478ed4b4427f8eaf29ecd53ce8845e4b1c755060a986af564c8c9ae4dd39bec15d0e0fec4327c6b1b2f4f0ee135badc7dc5df8a51ed2bb7af18cdaff345a8dcfe35a5084b1e1e6381a3cf6c0c3eb1c8f8fd4bc3117874e160f64b6e2ea7459b5af6164a58f7faeda3614cb30a88a8cb0f628019bd7298f4e085ddf46a70ec8d255087f50a735488a033ae29e3533ab74e840218e2c70bbb86dd130d1b62c35f856c6af4dcab10f8de60ddf7354f723fc2381313270776a7be186426f850ef2217aef1ce02a5c836745158be9f3e8f289a8c8bd71c57205322a9ebc19a1514268c23162ff69a916664b0c521468b757451f02d891232b49f91a36cdde0d647b1b3f5ea2e80bfa39edfe4071a3cf556b8330f76addd3bcbfd4acbeac6cf16f70a7c356f5d3e9876239c97d11f686b5ed1b7bb25b98d8f38b8fca9b7e854af4c343e54ae6573a7c18145fc6bf4097711aae8cffca81696ddb430af7d9e074baa6bafbc019f5e0516969f1ddd74dca75e57c1cb94f04d06f98c68b77f19141c87ebf048448fc22d72bfc025ff1569d9ea3dcb521303495149ad434e9ef7252b23c5020fe80d2e71845243535859bb0a79f429d0aecf47b4d4a3262290ae17a78167f4f919d3e9983b6cd2fa3441b7c8159afbc27f130d946b30627e7949da726b4908c5ac8bd44cc9e580bfcd0487be4a20b1878568665216874db55e32b6b334e3871d367b7de8e77b10daddb39ef58d02491fe9a8710165d7ef10ea4394d700d3d49ec0616c13f35dfceb92c7bc34cbf18ae4af2bc9063941abff16007c500f3ca792f0783489733cbd1d93a02e314dbd322871ffc5b384912fd4afb175ecf4515f85e9c4eb304e61b2bc52cd8292fa7782649e906dcedab8817ca0c0fda51bec9a09536c84def59f5f5455a2d60aeed75e58d6903238c3119c7e192b0f7b89db52beddca7a50a5513d802709f0c7ae44386a1c8aa7970aa9f344e7d8d9ef483d0a1ec16990ca1a33b0720e83de4a5139bcc61505934789f74b1934c3fe79cea484827becc232f8c4e0057bfb0a32bf98944e219a715e7d35560a8ca38896db12a70df1168a866dead429be9416e30686107300b8e1d3b0e829ace078bcb8baa5fc08b489dfe76923d0d551e7de8111196672171d21dbf4e22a9f2ba909c403fef3113e82d9a9b0ced41ec98ad8a6aca2b98f9e860534ab8b64d66383206e0bd802186dee5210e06a34bfe12e05f7fe4ecb08143f0f06de6715147a28e2aa5cab1b2784e0ee947212d637f3cc472949fa99670113d91dd8d7bf73475a5c5ef0f357c8aab0b91d523af67b4d5412dad147718ac849e49b1d338f187a3f57970ce0847b89e9f6455e8ef2b273c854489475870cafb1e838766d64e6aead42aad80e9304b69d23c9c8be847ad3ca8be2759d18c23cf669298237469e42b7645061e6ba56af66eb803a3f8f70f86d50eeccae63885354501f9eed7883fb88d53729ae8998e6315767dc0920d43a256500a2fbbceeeef6426a5b166e11f82408c993870173467d1155492e4d29be9a5df52f43ca9030fde6476e34e6b7bb6418b4e0f7e4b5fa0bce96ea09c56408b4ed1899723dc178681abef23c896e4c8b545a38e1802ef76f4e1529257c9839d3db2f57d66a0c983a5e8a83a9ae0dd95ce4a550bc8b20fcd2f3f8b42d12e93f9b9dbfd11657a1f9ad25f5a263d886cc2de46a756d9303524979c1d9434ac455d639d54a93c959a5c5f664358471223251b38032b4d855a135ffca2aecdc9e1e2fcd8094e51e8ae85dc8a9d9b667448b456950fac9fa089afceb8e4a1e578ac58ba57094b2fa1922a28891d616cf7f266609f02da92778dc6b6bf45c40e117976d00d58a62d57504c37871aa20176ec1c8526a0ccca9f958d483b6b81a81715a8172bca9827f34546f242abe5724bc79eb1b82572ba6919d20dc5d8365d93d14db25e8532cf9697a76c2092499c7159ad738d6a96da52e2b5daead5789dec6fbe3d0998aca3b9be287b437355ff3ab267bf61acf486cb3bb87f564d599d931ad2e9f0bf23dce3850a840f453816d6a4bd4f2c61a5ded8d0b668f89bd7f9ee50a7f7697b2abc2be000abe3afd3fa0d2eb9ab444293c766a33ea524a457987b88a898288366e61f9c15b64c17fefe253f7007948e4983138e986b49cb5b450920fd3f0d64bf7bf04f1560a208d5e8eefdc89ddd0e2f55fa77ba3e32720ca585cb6cb6c5e2a5f59b25358f064220d049b4866704c71fb5a6192fa988dd1040e38e018d05193da2f6a6c2a562d870f952f49b32700f832e9168c2a059a9ebcab988fb54977627baed61fc5fb4cdc68abe0d52618b0671257bd4360e6bab7d6d433b65c1729aa9a0f4bf5afc795ed0784db69679ab22b45b36ed7c63e81ed41062b65e244cb9e503621c5d46ae279e44b66ca8404157351cb2b70d4506c7da3b005fcffd5226cf3f6d76f93d5a278cafac648a5eb7cbc5570c10a7c27163da00436c95a39eea2c5044130e348ca4200699069520039cbb11afbf653628cdda0ccd18ba8d8c26f1de674341e8a881f234950a8ebfb30d491be34634e08f9bf0c9c652532136866d4a27e19082e6a5d208de836cf3ded4eda8979b64f8d9efe5a7322c7acaea99962d69d6d2ea332be4c0e4b0c350f1246d2e4bdaa6807f2f5dfc2fd0c119c33fd35118061859573217ae96a9cb3436c7e4330489d57898782041a570afd671a5d0a213a3cb598d0a6b600e225b0521feba7e437827b8b1391ad6ad4b57844d89feb80f9b5f96c84a0a21f6cf23347f18d84d3168979540ba78e9c0ef351638cc6d8a763779ab370510130e307567d24be886b52b67705ae85c4add1970e538a09584db245b439ee15ce30cd7df7ca2ef5befea46c13c580058208e0b6d21a7784e773f1a9d33f14e32848a5fcf0d48965c5e2d9ac12cbbbc2ee5057f871eb8394c308e437501c1969e0a9ba1eb47eda11d86e487a4ade58a0895d8742e1e0d911ee56881f976fa79845750fdc190be191fc40d650007e5e71d99caf387b41cf7e77844092de10e23f5147691c233c4b2b0eed387a575f47d1a316857ca1d84bbbadac8942464c1f080476acee29d93002b2075f1b7ed2fa1b1dbf4cf9f2b6bebbba6ff906a0e9e6d064cb2d631727a7516786caac7acfb35a29bdb138541244d16e939bda36303f5a131ca660dc39add052e50b7b8ae205a92efa7b807f84bfb036b4168a101644280e341432fcb7ee102180baee2122789aae82947d0f7ccfc52fb8bf84c1503e420f35fa912beac1ac2d88f61c095c66d1d879806a7307925e7ed61f4281cbedc0eadec447d443e6cacefa74eca798ec370f762e5dfeaba813e9cb872656cec4d59c8ce30351779501a6e8a7ff1323035209e81b0a0216c5905b9f93c67a6696a368b51be78a1622c37d8c817dd2d95241e287e6a59cb44fdfdc159760ec640cac5c66725a705b4e8caf2da2ba5ec1afebb7cefde11dd230ebadbb844687c7a07f4a862a2819000a1f1d41af601160d7d331e3e858bea06aab18093c192f1d6a1c0fa219312e2133ecaee616164310490a7f6373d1ed16bf6da29bd9a12df9d76de0b0ae26c050d03c1f161c4cbbc9e996abaaa3450294e55948e8ed79f74dacf535c2973abbabb6d38cbf4a2f82847df81904e08f4b430018c1af37877d030cbfa81e9ef77690f035d2648e00a6deae8ac1e2e2870cbabaa2db8fd33394b354f2afa9cd2c019b65ba69a03621da164cd3564db11a4bfd440717245fb439a240423139f38b39251cec332498efabef3b495e6f99fdba0e301aad6a6fac0bff6882e9cb855b64b7ce2c32568daed620b7e672e9e11cbef72d3b7242784e24a91cf64933e2edb6b7c9eefbeb15ce30951a422a35337314e37b092ff4640c19a47e2319d17c1e8a7c4e2419d748c1c7bcea50d48ae04a8aea7e37cb15a006214a205a00c6aab49e15c4783bf6016a69308997ce9759d043c853e572a9e511788bc55833bf1ee7ea0a218945e0d3b94012fc97646976dd4ea95d1e826aa889ab48b0fe0409be27df1c0778427176be28cfe5f05859c3711347ad5c71db1a7e4c1b0d9dcb8b5062a667614ffea5c86ea3ed24a6badac30d7a6bb4c499b9849c2d8798ebaafe947d850e09665a52d7a9cbc06a0ff2d7a6192980ead9fd93f0d9d1c492f9216df0bdfe3fd577bb4e7f11d698d8ed3c0a5e16e4e9d18c40b8db93cc66966b32a3d3ae440fb05821b997f016ff91048c04695b8c446cb77cfb5a9bed590b3beab6e2d5cffa873a70fd540d0bd82fa36ff3ccbe0e18744794e4f048b152c3a409155e84657a33073e5971b9b1d9288eb12b1debbed6adf274546e8835e48c272bd03f53bd2001a4c1305e116c60ac3bef0478e03107566678af675541ac97507f4cca81d2216c2ee6fcc0396c5a6f3d54aaf05719b65878db3d9b0aaf2bd1bc08b0a5c92994bb9110abfb4aebf44e03fa596405f97493bce414c4d7b67ff65b4850b2020ad626ecf3cf8cf503197a00f7e200c86075d09319405ec62e44e345a4290429b8ce15df3b81c5a265dc2ab728f1160f60c8eaca04530a5b34699faea4df6957bcbe81f482e9cddbfc52840b75abe468c96f79f11cbcc27e8ea8eea11fd64c979db542e0d2287c0cd5cd99df623517d1a99f6325237d37add50c39f8274fa653c4763e1b23a1acf401a66788bcd0d7d70a7aa64aee81094e6949694fa40c4116b94733e9c2a24ebf7422f3da7cd7cf2e2446f5e19ac2fbf74007437edf9d144ae7fdd2e17d1b695d5b2bae18650c8428c5059e5fdcd0744e249bf924deab4b6e0a00b3ae7c796b9acd6c99255bf0816818549521d0c0f9e0788925372a861bb8305b16236195a4ae9257d402f346c8ee23d91572a32e3bc2eec591b6305193da3cde662fb5810237533e53833a283765643f02a8f08b9592f8308deb0c1d2c738ac3cf90a8cb61712fe6de5cb886625dd60cedf742f7786f302f3fbfe8ada6e9ce1b1802235df8478827022b1508ef784ef1591b0909b2a2a5bc3250e2e3e3390685c5837f1dc8427477e4b38303880bee88386cb5fe8c1ded7ed1f71a294c29a2904abfee322a34b89ac4e04abe140b2e3fdf4c5ba2e8ab1411963aa93fc3f394c8ef26a1bd256861f243dc6d534afcd03fb4bc69b1c3e3b144d5c1d76241c5a0ec70494466e9dc75185b73a916e567b901d1a1c5258960281bb377984e4f0543e43254295e4a5d46ba450c859255f2d64c088d046039178466eaaad9661574bb607592cfec1e9c01614850ae336fd34d0133cd985af5ff15471a56b1bf6c518c58c065cdc4cdc1c5f0fee521198e6263ac2f3fd2b6c1609a5aa8f5b576a80ae3a391f46f4bf9f1665dcb1c7623c1864ecfa5e46794859175d9e32c82da6e2dfcebd94bd385db3fb8054c51eeda171030cf880aa3644dae06548de6901cac63745a3a696864e60b0f9c837;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'haceb6151560045af1ed61d3d8504686119f1815e78d9847fa72757fa80e04cf3a4a45cb543df6d8c7373d77e979388c9efd1f34b143d445089eee232edf955d688abcfa08fba283f2d1cb1908db09bc39070706a214548f4f9453b303bf4f66af21c5cf7109bc99a5471d6375b6f599d044e01e90126fb998477d7d199d4be22ef594ff3f1909e5ad51a6aa001e129ad70fa883ac7bfc5567bdf186c1dcd82ba2d1e364e20c36a19a69223cf842e4a51c86809f60cc3cad626355a701699f57765b8cb9cdf28fbdeacb731eeb2f53025d13d44617d7a7a4ba699dfb580e723b9be11ef44dd7b6a5b61b483746c0cea75420d9c15b004867242548a1656492120ac6174a5ec64ed46d246d6d2a157ed680fa15742b133b54681eca7c146646bf8d9b0486a2d7cd66b5c72bc413dc97a2cf586bbb925ed911d26ae4dda83cca4d6af917eed7e29afb4a1e232d5a1bcf19897b5b1b746ed4f34331ee86223937f9c206eee8aa4a29e39893defc2d9aaa8f40eaeeda4ede5bdf357f2484d8f3f5a4c62294b53821296800ca1e7fe4f7a09b79db7fc891bf3a482ca99a43f0ecbb9d4d75bd2658ddb404b702ca2dfcfd9f7fadff9aa4bc6c0abc59466bb6d265cf9122bda4ea3022f6b65f8b14a13b3a9f84d0c33953203b13becea3c83baa0118723485a04bb8cb0a97cbc520f0dc8d8e048532d5263a54e7032c2c6338d49013aa779ca4594f24fa9d52a91cc48f46acab10d0c9f6a226c9e827e837aa5a983d5b7d630e2d0457aaf5754e9712def1b6e190a782c6b4501d9adb43e1f846fcfcf77fb9456cfb6ce743bbc9db974bcffee52127bd5e83860c111759957a561bff6d3d1201ad8ea238a48de43c3a037378305248701b13912057643e4ea4d3a325c904488ac4840bd76bf0221244a4480d75c02b60fe6b488df4dcf8b072f7ab5d3ca86529d331812b2aeda7dc0d238adc07018a0c9045051b3a990d3c8a8a154a5b74479d9fbe1e7fe0dfc60362b6d9c546b52a48d25adc13bf762a7f992eaa8aee5b992ec8917ee5560bbab1eb62a84503f166432edfa41adf32cca1c2abb9a19cceb32b29e481ea25ca2c339a671708c28252a44f435299cdc0202971891630f47cfba959b01a60236d78c8c7e58b4e76ba9df88a7d368e52f5d4320a8376cf66d14479801d52b21e201e41742193393c062c3fc9b9216bea8bfe1fbed6c57388fef7fc3694bebf61ea17c4458e6452c1c86f99adc3aa3b3e0fafe10f5337c9eaf589173a700662cfe8725551fbf6b1500ab5c921957a217825824bb91c18618bc9eb9e2eb89dd71cdb536969848f245545e06263f578292b3879ca82696d7d5ec306d62f2a41801430d840a12ead1f5afad73f25b34cb2cf134b16e47b53b781fa1b3038c4f9e37c0ef7295b338cb89fa91a0237054254c51d84fe5c331c522b6b0eb3d24902c81e7edd4d6e7d64e5ae6e7603463838be8a219c9b85b7971b104ab6c9bfa1eeac393c0a5b4c7856c2e499d019776936d18425425ce929fe5a4ccd571cd6941b53148ef6015d1e4fdb2c440cffebfd527a694eb32e674a24cef23030a4cbfaab68ce780c2e4fe1c54c1ac52b9b4f2a94e60af9a9ccd2afae35a3decb41951d68f77de4c5fc1e295ca9a5098480077e050119a583da98de8a1ca1ec8f7d6c0a42abfbc0d3d868d8f7a1e1777226f800505551dda09d1d8a20b95031a0666d9d4c48cbfa6dadf7aaada2ea9f342c2313a3b23f29ee4a9e506f59f792d58fab736722aafdaf5a92d4898bd54c6bd653414e71a662cbabe58e7d60f07189c93522876323094a506ebdee0e125e2b01871b84f24ce81cd3fa81f9c5bb66c7b74195e8873d15a38cb6b4a56c2193c39c7b1f3a4a383baed55e3062dcd47a5256aa88064ab6b92aa21b4041e97bce30c9f2c68b79898197543b5ed8dea5aba165c6dafdde00aa1df20c44d18e124be8f78a2c8691a25162da075feab8b5eaded4eabe2f24b1550ca1d66f4c9a861cb424b0fb598a769645d6fdfd6f43c2659719cfa1d17f6c2b555fe87332335ed9936714397a7cf4af773d055dae722621db8e6cadf45e24b38e9b696b7593cd008edfac59814f708d3ada54674a0b078d61634dc6a4b8b2e79e8c4e3d36910fd08f2f8ecea11b8d1e9dbf441361197cfba7922c6aa2ac13bd33786fdfb679f43b31bc54a5a6fb100450a30ad4292ad0dbd38e96efd83131aedee651763967954b63ed2813830a78fa41089ec728b687b7c7e335a3c0d794119b60f8f2635f927943415eaba122720a30d507ee4b143368db1b518a45681efe6f74886cf0fa604d3e7b99d4a48536c6f7e1fa4b3b69efab32f019644cd05bd7cbd49263e92c8d113245d8a29eadb5fcd02180c4f259ff75c56b2033b1ca2f00d04441bdab23529243eff11d6eb4d634ede1e5f774f151d672148c09f09f15349c802ffd4327db1f608f5ba96af822a716c8e132cb4e2f85585bc60def322130fc40da2e18a6b283e18d238c9ef7cced3130acf7323834f56d11ce440721e962cc80f70ad45ffba53af4b307c455ebbd46859ddf6b9a9d4a5ff09f896d533701af852b976901efb1cbe4b5d58686100dfce6da56a29905c338d01fac4e15195a76bb9d8d1936e92c2afe135cb50213460b02b7d872bffa5b9a0ac936abcc428326c1f722447d75c855e9d719b0b12d0cf2622ff73dd91266f6882f8bd8fb5feb9032ed9f6777a6e63700da3738559b07fd21f367e4c76474335a9790177ad67924accb1adb9257f0c209b929d82295f21b140e63a05d7bb0d9256d2e8cf749af8e6fc88f1a7b86595c8f6fe7fefa356c916b299e4fb93c0b9323dd93b9d3d5636a32e45a7f33c0853ce259381723fadb657ab57c203226f774bbd416c7e05b8dd55508e68ee28b4bfd8e1305b55b91436ee6c8aa3b9964462c34d9b4ccc110aaeffa4c081ae6e6c4a27574622e05f8be0e30a456ed5132bd72b9434b7f9097d35e217d021f3c8430df0d733e8b91809443a6c59c6b90f6d38bd4d9db674d19bc83289b456954236bd0643f49ab370353bbcef3b7d91ae8d778099bb4fdc9914234267f19ee7a0d2a9735a38dded17dbb061182ebf11e7d744d051dd6e55bcd75a2b131dea4722d138ae5cb0a18ac78443c617aec976bed6018dc1bcad6e32cd8c2403d9338adea77f5d18b10b6a3ecd51c4fe419973a66e23f1ed40cb33319e0e1b85abe044d4dde7d9ca158fa93dddf5400669d2f64f0c3a83892f167beb5718253f14520fe3f07c362bd1b864b47d59332cc4a7718aaf028bb3271e3e6a1423d9b07c47e97a7f39861af3467152b62fef85872234fb3d72f3ef5d8a4d64b1da003ec14d8183315cfc22f04cf9d329f091dc12c886da0809a60680566c714155468a314452bfff14c49ac76e99d8d579fccac041ff34eccc033abfa38e7d20e1b339ac31b2644c60b67e717e6ede1b9d3bcdc8ce38cc845340140fa84e02b2f5519f22e782befc587fd6d12a889d8feebe15a3bd079cb1da4986d1e14d88847a296f7b92e263d4583fc30459bb27eedea78314b4dc985ebe91943d6e8190d0cfd1f1be81c9d02c0fc6ee9df96685d3c6e7c61cce146726357619e2a0086d390fe417622214a94a614c0f586dd41bf955e3239b72876bd1ef370e04d3dc9083d3e0fc46a409afeaa31254ca9911c3965813df9d416e76fba35576dfddc2d92f4249c76a0c8d4e091abe159fa49e7dd17ba5dcb429fd96dba0fc74933d88900739504dc536a7259a8a7171a8173c38fea6fb4c8f59e14ef85a55a837fc6f37a69e28e4581c99f21ad08c0ef3cf924a56a4e68eb60bf5949d43da5057a3d2892dd8be7858ba3f6d287c48e79e5da95c17fb3c52d3dbf9ec415d67cdace606840845cdbc9f868e9309403e98e15d775ed788e29d6daebd84223e624a73615b67545d91336cd401f9a1c3f9fa037bd8fd1bf637d24cb2849c0c365ccb292e0635a2cf3ab7194dce9c4ff5510909e73c4f7192167e46f0d9afe320f626bb48f7659984abfde9ee9a90ce729b234b91207770c343264158303f16d3cd40c0a8901ea059cfcc85277454a4816e20ba7aaa72ec01f7afe9e6178f698cb7f6294ec989dddaaa7b1147344abebe3c6f35b95206d9de07c7b7223024c22dd31276559011630227e9172c4d650eb80255d0781950854ff9ccd6a1d8c97abfab44484693407a626914896d86c4ca06f249def42fae3293933791bfc3839a7bb3de5f382397ddc45ab3c366e7805cee175ae830d8c421f948e7580f68453b5b3b47c0647ed7640d44426f9be71b377e29e78a95437a720424f1598af6f8e5d475057041ffa75124e468b9d3678d86f40e9231ca3b7ff167edb3a280b765506a05fd333aa760f19a16dcfa9ab3589b866b26dc2f1ca84c5d67ff01849ae84745b274c67e11c0360a54bda0d7ccd124c0da93a8f1255d34decef9b6f278f7a134bf59f5bed05a28936ba92e69f71c16b1a4a00b80a3cf94d3c13cf03d91d7e9f941c0762d3619e22e71366c820975aec3802d15a862f89a3f3cd634d930b299147ea67339b44fa83f30d3878284aa7403a74614b41cb8aa48bc73e8ccd60e7b9049eea37c264ffd6c7e367c9b0f25c3a76da3494bc24e2f592a0fc0c082e8d311324e5ca7cfeb7b79bf4db210e8299441a80b02ce3918dd3e4001f59d94c62c3bf444ce74f9c64a15bacae6fe43bd7fbe4a614b816b19afc269411bdc20fb625f2f5c6c91a3b09e239edd6ae310108fc03a23ac1bcfe4e10a7f1cfb779517b434eed343c65f40fd05295763da49bc68e306149a4a0fbdb8cf6173fedabec38857698159db77e4c20f95400bd9944ba6e8b6072b8f30fa86042179adb616debb5f81bfd79c2a012c00f9b2aaf64f3850934c39b0c763a281cb0164a33fa6aea063b6ca7d1d88a90a9b6692364f802c61f295c651ad0c705810f6028193e0e0a3531b66e0b0513e92d0ded859df557799fffb4f84e6be8c891e4b11f634cf43d298f5cf48b1cf68508e0557a246d3a8bf7d40660ecac32ad40f0600c9b1a30e0917e0aa38d6b8d3741da3d135ef89a294779036e6e2b76f3e4c670222d47e8f8cc90c55857e4871ff3c3f176bb8301bf876a522f6deaff7ff42224c3433765e3b528255c538c7a74a3d78436b6b8a036f18d2de7e37ae2e0f5e442003fc2af3edab2016a8c0dc8747b0668371c97b7660737b559af32de2f8c63bd6dc3beece26328c96a0265dcb41cb1bebc46312d993c6c1453f62a9c50d18e634c1790a4334f5aa28e7c8f64abd87f97da1fb2f86ae753848d4d6685bb01a4d85a7364f50bce931004cbbd24a30d5eddb2dd79a4d695289d358ebdd5244536c65d6f92970d71274814d0496e6230ab7fe0b4d7dc824fbd6b21eed8f576d199ca5cd781f9d4f59671e71677ce2cdb41edf905956006efa931aa561214c2f71cfc148a246574ba9d123da0a5fcc0d9f980dc23f71852e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'he4670ce42a3c77e88d879f3da84529934ad8bec546c3edcd0110d7a5b35a4adfba3ffd14a5cf10c22c165d418dd735756c7ab19de778e3f3f5ab33fd512dddde9a91687e5c9a63beaf02efe669d9b02e17c619cfc16601131026aa6c1fdefde4a9a8ebbba79983c50cca0ebaedcfa014ec649ef2c0aebea86c81d80d1a7b6eaf677c5fd67ec323e45e7f26c90af12303325d61f65f9491215e136d26b3642f5ef1f1e3b6a0bc15e1b4fce825643036319409e71500609b9d92e603eee4323de270c139ef07c70f44eced713cdfe5e23b8ef152262b05a9d2e72b7a3dff8d6aef5c5b75434157e67d2045fa4c864700a49f288e48863cf10b310fd06bc766303bd5d7fdc0443fdd94ddf8a27752513f529ebda6783bf15bd669a6739da5dfaf5172064c7a72a1f9ede7d92210285d097f1dbcd6fb1f5189ad79667faf76ad50d93b2a629cf88a0233805f33b3c4ac1d5a0aeac3555f8cf50c71e350d331df5a34a2625935183598b792a6665becb036d549ef15c2f38798effdb17c3a6556cc24ad533976dbcde1b0883e24b4d676e0bd6e5f250edf736c1b6943a2a433d7e0168bdae618683598af446184f7e10e0ba6563e961907b051d89379dc41935b8ab8c0c84de551856b816e0cdb294f87ce04a208fcb69e0d911f59769ec3d73e3d7f13f63026e1cefbc36471dbc4c2eea73ddb280774de70004ca00ce932deae103f6bbeee989d687a0a37861832c97d88f00669b1b0ab10e2a194b5fc40deff8d2068af9dd6dea4bcde4f0340880848cafadf1f00133ae30d1f1869b02d4c8bff16be79cefaa0b985b18a22bd62544ddabdaae314ee1b97da8aacf6b0c967aaf524490c8ba8758623327b90d2e2a57d2dbccd152a35fe4f1e697e343d531c5aa7f2217f3a46f4f9d5dfecdebf86f26324daf20776047cd9818ece9d9531193650475ce89d5a97d5eec351754e2362613d20d4dc6cb692618692e327ee31741844488baa2185d09a6e87cd2d1843475d8d536175852cbe15cd6569a6915b485c912d66fbb480056806abb79e982283a5681ab4696916b5c3c1e5a8cff9948b36c60160bc57edb2e3c6d57f361235ea4f4bb5a84983e52c0eb0114f5967c11047ad547163c1cf23e8f1ccc6aabe520c567316576b69cbd8ebc65bc838ad28c60eec018a8e2cfebfefcc39472fb17161410aa231594fd6eba97c2242fec28948e48e5f5c6ed3fac5cdc1cac2e7a14ed4ff2d11329c69081430f216ca483b734cbdd23dcb6e39a96247ff83698ffc47024fca5090024224c8761534033a1fe46de24a7b8065e51fbffe95c5445edc7f984b703b5b321685ec559e88c0a1c967a1ce9b3137f657fc1decf85b999b11307fad78d9cd99e5031e93dc1283edf01707bab867385ee85cdb63856f59e4675eb5dae6c68d5fa78d7c6be46750cfeee5aebc211fe177974c16aa4dfba50e76ac1ebd5b0d3637df09c812a9bdde37b9d599271f97e3d1059adb3401300b39616fa6e98abc4157a2e0182430bef9aca965da8d397e69ed89cc23c4f8edb8a2207a2fe63377d85067a5b8b1fb89c9f2d3b68bb278ad208fa04ac7a9c0022d74d158a3de409f9ba4cb1d0e3ad6995c8bcdfcddbcaf08d1a46d22ff0229f13f690f89c13aee1083df91c0ac65e470781cace7b28fe01d174c623aacb1670f2320c9063f2469f9025dd96ca835cb9f6126f5a045b7da0b8965864e72ff46cfb18c7c0dd9b6473ccf167b8a8c1cdfa4e79dc5f9a6b158f781812e10bce53b1fb962096f0a03ed4f76b8100114c68d6b14d5914fc29ed8c834172cc7e3f9eb53fd96620bc5f7b76cc81fd7b4d0357cd14e267fac88a26a562704c20369ee0bdfe6cd709201485ebba6dbe6d1d434ce46091e2b605035043535a031237e5b93aada9881f785a500e368055706897c47fc68c38848d95ca231760aaad6e853b8dcc1749ab2796bcaebe02f27063986b933c2aece06901a200d654b89c20438ecefb11cf647da46907b2e0ae4c806cb969305a904f256655317ef96ac0f1f60730a6c2661b36184402306090026a73f2a31f1d10a50698e42ce5d6530e89f542e6f2431b67f10815d266d26523704bd170ed1c7aa39a396cc0f5c94499b34196f54beabd92c13202798a87a32eb9ab326622853de76ad1a9775023b63a6d39ff14532b9da45305c2189292040b7b4d99105475d4b2756c92f800c59cbe3a7e91d06fcc8e07b9e90404800db370d43026158df794f85780929fafe82885afbb115c96db30c991f3a5ea3ab945bb74b8a15e5347c35fb1d05290a6e514b5fdfd101ceb3910e140a309f3f886e24019bc932bb86882e88b75bdb7ef3d5a26b9648c8af47ff64aeb87e75b71ac8bde630cc397e4c8da8e27af76d12e5d1902d8ad5370fc9c4c09fb214a309df2a439dcd3f89d246b581579702341bafe95afe37fa2d04af6a31410753f64a6b8fc4e65b3cbfd4cb88414d432d3561f694fffef25d2f644f27b60681065ee83b0e5d84a3d76d4899c8a801c2527a6c53a368e78ab797f7cd8fe429b7ab897713ddff8da92e65027a136053d71cacfb6c52f52ab609b455c8acb5b13aaea64a48d39fc3bda94b6a017b5e86af608034ba3d61be3ee6db8f7f0bc273d85a9ebb60f0b1157a87c4ab016af16bbd7f73fe1e8cab279b4fe5405f053f08bdb1910e335d41b8f6cf36daf3b3dabdc8406c20c0309a372b74e89360a656eec5b66fad4d1982fe21f4de208b89a36c27a019c4c41844abea723b620044b4a52b828b0782a8aae5eb90635fc95fb0d04b2f0e4eea71aedbe263f6e74942b6f64a6d6a00c831fdc2f9155eacdf1ef1b68b750adb3379c47a92380b068e675c1f8a39c5287af0ba7ab00c0c34fff1cd05075eb541d0cc8d0bb3a6fc12c163c555df767c36ac00342cfe7fb44f4813946c1f0f452fd76a6510fff776b7fc6b4cb4a072ad7eeafc8e0736b47bf7fa36ec51449da949225e2370a4fe6482588144d995e9492b278a766779a1c387709db036757a31f916046ae1fc4ebeb96cee62c7b435650f03eb2eec7c93d3940ff7118abe5d5eed880fbf3e8679b70b645439042371db1d6b4bc9f9db82b9e765c8a583ab03f4d46d63c08f6188dfb7f313ec34a4f4cc4d122349d6e6a4db5423f0c99fb9c18d06a845b6331414d2200e6b75c85bb9eed02bc3232999fc4caf268f1158e03e3b31fe0f38088c1f6ce739ba7371d3bc99a94933df832a0eadd9ad0a3a82ac9ce55cff9e6ba9263c0b39214dc32777b728e2f68438e40e45b3320cc23ca3f4cc5b608180a9cc9f0ba08bfdb7b51f903778a4113e7642d55d09cd4c1af066b54f27b07417dbcf8c6a975a1b6814989dae1d7bf2445cebe43cdb36357e7d13fa487b4a643f83cbd1faed371752768801ffeeef40d1ab84e4eba6b589a13eec0381f6c780becba58117d5a3a429035eb7b2103de217acd96e1c6a86fb241bd5bf09b71a2d32cf0567bff9c5a593e1cbcd4136315efb2899e54dfd53d4978196719cbb080d5995c3f463faf205b6903d58019c61d6a2bcdffe66bf2f844ef54301efb99ea496a254b32b92787b470bce03e872f927e642334c2dc3e4882cff1f82149bd42bbb369596668ab98caf05d125f8120300424c014c3b99b922824d5a5e74e25fdf74132ff010c37cf2b0ce4f62ecfe9f0b90d341790b70ba2a67dc3665eb64be7b2a707986351f53202b34454f3e81b1aa4294d7c0631234fc3fbed170582d8eafeaad1f49fabf37e29bfb4174534c80d31816a2b1df4960577cb8a7cf2dbbfb8e7a9d965b58e8811b1666d584282d3db2bd23c99a5cbabae29ccca61671cbf5420d9ca9f873591a8437bddb916f458200af58345f6079787d294e3b35404b07db0f0609f8cd8961c69921ea9c5b3756edc81d75042f7a37c2f657ecab596fd290258466075ee62cb553f1d7ecf39f4a0db15ea34100e5cdb90a0cfbb6ee94b55852a429747140939e1a0f4b0197d18cb4168ca922c0b0aa0cfdf2c446222c5fa02cfcb3e0cd0563c8090285fa225037cfce93f98d0f7934de4fbcad84dfbad05773e3ae5c90686be611ca0f5b1c98882d2faa412adc6b854bb4f87a68a7ada637afb4f3cbce4f3a0d62f45dfc59b24a297d4ab2eb459305ef48b2ac5bf514d5e2455d4c2e09c8906eb7fe05f94d8f659db58fee6aef3f85479ced4a73a2d52f9eacc4c267231b4e6d6e628c0c673a605fa47a7a02abea9809e60a42f96c82e0f5eb434ea47ebd69c0e89e47d67d7856ba31f9003d116f3a2c94497c042ae6673b7e2beb272a1a2726ec5f30aa6d6e7a60cd218d173410450a510488626469cfb49b85e43d163441f2467d5de1f735052dd75fd7e9ad6ba6871e5dd6af5006b1d4dedafa0d5f52460e2ac09baea9a22c3dfa585b526fa263052c66d41c6758049b6a1b746a2ce90e8d3e14aa5e89a65e9bc843684fb75d3922c8ba274299433fd6b544b76cccaeffefb6e32b1ae540582a92d1c509d5a04e359cab119c3291897f49582765b4ca73c737190deb7805b9f567f20ffd302ece9112cec36acd113bbf3524899f648fd2a5759cfcfe15facdfbd25163a593adc208f85b968ade6063a97d523e01b32394c857c45a1d86884347879d640753889d0f7ffc9a72c740943701f602ea39d2571e3bbffdece82a2f2c728b44094ac6783e01183329eed96f1f363f4337a63fab94895d0ac335b58a16fd1f9940c7d2bb3acd3773041a5e851f0ed92c79cc9ff46d408df9002a8da4e000dcb81b154432187c722e71c64bbcdd6c678bc418e94e447a0aa49eb2a20e2b9b0b4963ff6c847405a9b2d9308e825b4553d958832cf03ef06fdf4c15654feaed47e315d1c5149f8bea1781656d0126b02cbe6ef6fa9781eeec6e8b7a944514efba4cc23d8ee3a66f4b9af852274620f24e1e4a28ac972b8153317021435de8e4da342acdc0117f1507b9fac4ef81820c99c3ceb792c93296fdeee47314cd9ec6888a006ade45b4dd5d62a5b83a6f60e8b24d5fcb1ad5d98c74e092722bef8b7cf4adc6e9114b4f86dd04cbcaafb98f9c8ec22994ec137cfcfad21e0fa4feeb5481d7ba24931e87bb4af274e6c9a7c8b8b2f30534a43a812867fa0ef6d3797eb10f60173dd39693d494a0efa4be28486ffa3289bf36690c108168880f9eb5ecc927f55b5e2890875a2ce5c1c3fee796c2ac9577fa81c5725d9dce858790d9d3f032840376736681546b7830ecbd258fa97a13b9cf34716d13e145124746d30df367fac2d27b5d1c3c35414e2eedee443c556f27b6bef0512634ab8089eb1a69b3b0b1283107c1c22cb964f3883876d281d4bf3a0220c09b4eb313773d2a928d738e4a9fdae30523dad078606194ee87c062044508fd689a9cf0a0d8c07f93914a0301a7d4b4e29bc680a43fb77686a985002a9ceafeaa1243e4617fae3a1845cafda3930664e2ab31013ef03e1aaaa546345ff27016f6e90741a32bd2b90b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h8ff920a0f1995037f722dbc351c11b8aa394fa7c7869baf66fc9000bae2cfee22e8a5b9b396870a191659e1e5917005514d17571890bdf840e9c8fe2787f044309f1dfdc531411ccfe71f6649081f6e0182e42fe56b635a158265ffcdd2177d7e473b4eddc0481361b65e5934da3ecb1e01cd4e09408642712e2a334b88574b1cd36a917af6c9d1c00f836d26787a2b51939147de5d644dd01f48c8eb16a90451efc855d3a0add0c00b2df848103d0e4d96e89ba04491dd8e235b7978f9de8bb92dec16c959a7d51efa4682e484976508d1020b8a100d2b6e50650a15c4310ac72e8696915eaa43f2e9b400f91d330692dbf3bd15334f9306d02475e2710837181fe0d6fc28262ac0249c7eec3d96d09420e61876109ab5ce734d0120e646644424be116bf259040411ca175bdc71d0d2eda977cbae78e5e6c1f05a59a1665f7c6029a9214509cddcb4f555bdbfda75066b4acd2af45b58f12c049d14d3cce6066c0f80b07907354a08bd42ef18fe6758335d7031f22b370551773cf387f9ee628257fc8a5634b075fb006e61f8cf7728466a2ce615922decb0d72291b910cb0ef4e95cd6a34cfcf413971aa4c60ecc0fa04eece0e5cf2120dc654883f183a6ff1d90ae6f846a4a7b6ed4f5c42e3530f30af0d47b97d4361005b4e38d649ababb321a6d9f26a6fd43078f0622af230eefe9e08b2948f61cf1e0fe3bc0f9d1856979ae6c2e29b0eb98b7213c736a7b013585f087cd16b4356b63b147f2c17bd54f29f3e8773e724af914d31388ce131f57face013743eb99d3d9b493cf4ab6d32987dd8e44ebf6274c8992548834528963328b16f9cb14f4ed5989c177d9a51e1a1aa1d1636ff8f97770c2afbe79f24531ebb716d204efdfae02a760f99ed42eecf1cc6f89a816680251280b9864a18ebac19c7b99019e4f18eed1ab322a1f6328799a4aa20237216092702c31a434a2e3c0d3c2fd6390ef1d86658882f10bc1a6a65043f67912af17300814ee0215127df933b91e522ad941bc70411d9714ff143fe73610bca061ccaaeeb0304c3cc91dd664eac676e1549fcdc122053d64d4935bb8917cbc0bbf94a609f1d356a8b761e960376c2697e229efa4fc1ae173d194e1e6a32392b80523410a9a61051e18490fbd16dcaec305ff15def680b6f2d60b12885d2ef696875173dddff42bcfdb98d51f788502364ce28f7dd19105e6af6f2b73abf0790c333937998bea9236236b381f4fb25b4a9af4589f4ce80e0fc682063e49994c0adb3d79a71181fe0319e53f3731434115c26a292a5b7d01ccd66734d71a5e456b37625d4c5561e949df63ed44a850f049b0fd4ccf9a88c8520fe072c5fdd019003e2f2adbeb6477e979e99347e32ffa12004e3e9395d61ddb05c867a1bc9a16df0435f8e5103acea77a7187c0cfd06cf9d2ac51e2ca6c75e0f9c944fd167e419ff46d0e44693e860d528e3ed0d0dee0a845f2d8086dc208ea4f1b8746618026d970594d1010b3a8cc31fec36886b63cabe221ac34f5058b95b342c208ba3820521a6ac52e6a09ff6ba19b81f44e5a2ee0d924e6d9cf7cff1330cd9560b8579c6b72e308aec84c557c1e25c3992959a1a07bd7d34dc115014cb19221f079d256d1a6e49e6649b7afb27df317db734926e6b6f55a7c036d722153047dcabb966e477e30d1b3beafddb4e4a7df090e4e4ecf3f28180d6709a3987bde1907cd7a8f5b9d82e81e6d49ed61e764ad015da9e9ecde4a6755251fa637623c9b31226baf439b7543c8ca625fd1f8a5b5c4eea3b65da179ae1620b47aba031910c533eca51fa1ccacf17ef4236b86d4b53269d5e376910d9b0455359743bebf64445a149192409d8c2778f7d9a2ecbd398c9bfbeb38a413606fced01968497a2cd5f7f47413e67101ba71ad9bff29bc086e59b9344ee076ad8d0936af784ae5ea442d0fb85ed4c380704b4a1c41ee4d403cd6c97c26a8c5fb422a2062a23b80cf14a548a49deb7651469a8d6a1957dbb85d96685ca9d10b18a1309db35041167ebfa76886aaa6d9d62df7ee9b96c39986091b4504f448e920e773b96b0dc9bfd3d10c4b6b0833e3496fd3a7d6c2c7d304e9445f882073e4c783a6c60c5673f724972be25def764d58264e0021288df7b35115cbde8d6549b38c1ab555182366a7a4fcf09317f8fc68dcecc1e024b5aefddd5be98bbd8acb7bff2dbab358ad465163e0ec35aa26952eb9fa8563adb086862233afb709fc791431d7da449c3998c3db390d750e948985aaa4e907c910cd03780551a70c400db5001f84a4d4e5bbdfb17aee784ab2444b425010c414bec3e7bab83c6f5d99dd8cf37b245b2e56ce3a6f1b07ef28768cac45034b55f560211d35c96018186f3e7d695b8326e280802ab83d8c8e4b459d22ac3d2062e8e79b16eefb0611571e07252fbe8e43122cbfa9498dca2495760f6a16aae15b7e44347ddebbd0aa3a1354a53fe5bb0e319326baf78e15c8befcd6685ef977556a575bab11166d8541d37f8e9ce142ccd26c8584ca710b0c4b3eb3766b4884686d3f96bf6a6f1a9699dc76ef2b3767e5aa2c26ade0fffd5a2ca81f882529b637b5e41aeeca8ebe781abb1ad394b8b5676b6c08fb1c323dff0d80fe0357bbfe4a4e4b8fcb2ad143294a001c3927baff755d58070a0d4a167705c693ca8d66b2327fcfec47496b5be8850dfc9a96604ae989a4e2ef221b2bfe30ad597e0cd0f53ed5b91df3810e01bc35fdbaadbffacf74a48e2da1fb204f7c9cb53367c9c62002aa73568cf440bd45d4e635d6e24f05b482f5f081427ffe46f23e795fe02b0d202cbdd7bee35dacc3e4d108bf64ab7c1ab25ec1944c9e385c8da6841f16e39a2982b2a89deb6a053011e3ac6d2ef9e8951d98746a331ca1df195778925fff27fadbd5953ea970f94a96c0bc03094a279d775c06dc60d1f256569687b0ebef83b1d730f5eaa53a6a35864680a82c57905385e00a6ce03cf3592150018e889407d89e41fbc9d5c28385e2e63b777ab581359a7e57e1ac63711940366dd2f17ce3eca747568612027fd10207cec8f9a00ed96ad26ecc4a3b4b43eccf9ea744e4fb88ac368f12f80908dccec608e1ff8b7e886284183714b527925a76e5c636a1dfdbc69c1ccfc70e005031d96c0f802afa38af13d00e4802a700e3188020197eca3d7ae6ef661989ba54bf1dd9f13eb2973786197ba99abfb33e02c880440cd4270d2fb8213c6f1a87fdc066a5722585eedf1482be8e80729ad58360d4caab0c402e3f0b492d0bc24cd71b0a80a1db997ad3a12ff4bd1e24b8af0a5a3d4c2d104d3ec9a5acadc2629afa8b3eeeaedd617ff3e88c724ffbfa364029cf2673ba8bda767988f3dd1c5c33f6a576e1394240a92ca8b20d4497b0f50cd8d34afc4fd363b3b54118a22cda1556fe6104156bc9ae61ad88d9ebc876333587216b858ab8b02779c20f4f4cf0d031e0d1f6ebf310aa4efd040df39c9198cebe24ff198a982cee903c88204ae36d2d6c6c76fbb02e4110a563260ff555eff389b8f4f8c1ca3033caf3f75f0775b6961a36c8abe5a3beb33c418b6961133b7d902f7afcef6f645c66cc45b7f817fbf9f73e0c375c1de0469b44a2b06c2ac3342d3eb37f42ba11fcd04cef016d3b341bc392763738c31823fea57b605052bae15e4b1bee0b05a1ec90a6bff3b846c8c9a28be564b1cf575d69d20f0938bc7933587afe1c1de32c08b2ce0211b298ed8aee9f1fe904c766ffadf42caa3786bd02bdd68ab467b4a37b6f008afa091b806a9a4d080c6c56045fe5a01c4fa059443ee1727af77d7002c796615575cda881a4fbced59a9c2df688c13f87bcc8dce878705d68e1b4c04bd61521c6852dfc970a34aecac0b00aca92990bb85ea732661e4e2fb6eadaaebf6b30547ee5d1a2489752cd6df9d1f161f6dbeab581ae7a554a9fa4e7f709c9654c97452bb8bb6cb66a4a3b5cbee0f650fde14462ac7147e8f69734c3ee3387ee08b032b577e1ae401a65fbf714617dc1041a08c93647842f659cd01e65925dccde82ed1b8dde8bd1deb59ff7fd555bf03e31b3bc5d1ecca094fad6ec1d0febadc918ae663662528987b8947029f9f623c6f03fc12e6cf0eb72a4fcbbe7fe1654fac8310125ca297af87f26ecd744ca5ce5ad44ddf98a17f2eb3eace9e35a6a9e36bfda5b1509f5be6cc62272232ca065eefee32c8a146ed5d0571c00204873aa6eea074f25fc40d33d22641f899d38d09c6b493f46126a9f9f9dd8c03db54d583724ab29ff2edefae91ca292a9b065be13d00b217e2839ee30241ad72e90cc27de259e6777cf1fe713b05dee43e991245ebd341da4fec08e5b5761ff99acd0c21e2c5bc5c5d3219fd3d9098a541f74d3270b6401d1d25359478c8a0e848fda3b525cf0bf855c7e4aa548f98cb9fff9232dd1e7d8a4197c38b4f54bf0c53060fe55e021b072776b1192a01b6100b04016fbf2568b169f13149a8235b8ff6dbdb0b1b920956dec1e5e2c1d52bb901b8de5b83708a0962a6d14ff6bf5800d35c219770bda6169b55be8907a38a90f9dd2f355c3912c3d1029343dafbe612fadfed932d4ea082ec83bfb3ab046c64d8d6443106b90a240ea2c6319008c965c8acb071c01c71e6cf68274f2037e51f5b04dfe397176b981ccee1e27a42020d0aee9a07562f6f68be29872cd11baeeb60f2a2093c2123fbc90cb9a3c0f6aa1e125d3610e07606a3a3a6634bf565f953c2154d1bf54899a5bb4ad500aa0fbd3de52fd962ad13ea61d719655a4ff3ed0b4f2a43ec723f2feb96587a8de2452c962db0522c4f066b3bc4eca4970e3a3784d0b3120a803c72d801f475161ba871379e0959335a4a9ed09a45a5b2040251191b0c8f4c83172e234b912f8f2d242b8224d38ece4a1ad5ef2017902964907da694a1f04bafee2bbde1038a7af074076ee31a4d7cf76329c47a2c232686b0b85f92610e18cc091cf69af6e89f19125699ef1b3cefeb1be478a35106c37e5f64d01ee559f920b9ae38073fccf2652a1c9a6349b6e533479ad2447b57e1e3e5d2b36ea8f001220da477b44b6057d03ab1d98c142c6bbbe7b4d8fbf889092c98260043af69e7f41d45bebfbf2d689cf58caca26f12bc4ff890d0beef1cbf585e781a07435d550de6133a5fef962a8f55b7414d60cdc01b4bba0a5e2ba378ff1ee35f7c36cbb96240c6f349596dcc47aa2677a072b0807430a2acb5db47cc019fe8e2edcebb4659a48b49af39bf0efb99be653525c15a5ce4bf347a987b7168aec445e6fb057bc9c37a64699163f46a422b4934cc7368dffc4ae17f085bb2acc4321c37041faa8fad4c811a1be0401e6c0b63c54cc30a02e75347fdcbca62d0f797360bfc76722db8a4dc492f21cced03fad07f69742952c15818c4b74c1120bd95f1c7e25ed96064e52c11ae6cf5b5bad9cdc4bac246f850ca7197ebe1566673a108590406e3a475643305d23a9cfa29ef34891bb6b6cce357;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hc5b005cbbc2021df7c5c9d23713e12f59853c8529cdd578d1e3614a53d0dc06b1cdf13c7ee38556736c03a35378b5d687c8ecbe78386e73025637fbf849b3d7dbde46b001b3952d86a80608a7d9a0f4b1d77a1d16ae49dd04b58c2293cf6e3028b05e69e4a78fd6159a10dac316cd4ebb44d06751656a0a54b8ef9898b6e657bacde51ecefd26cf230e3267bb4a10d756354fc2f79c16da306da842ba675ac6014d6681eef7be168d5a1f08319327fd6ca99c0dbcd1bebbef667fc212323989389b6e005d61010e5278fe93c6bdeaefca20d4f416073c8095cb8165699a53a083f4359809bc428860bd7740834371450c27e3d20af5643abf7e96dada57a36c7c525bef4dad18a53ce01ca719724ba32a02c766b761b80ca74137d4c9bb50592a6b42ee5c5084bc26a25a43cddaa7fe59a262a4fdaa432fb63294edb50bd7cf721c0ce11f3eefb581e4cfc32aba56de010ca01d746c644468820c67439476e54f80793b93c3e683135170f51464da9742205a4bb3edcbe1e20cb058992278457bd00d7195d2961b539e5b855ebc71ebe67bbf0cfe315601f2b3f507988024f2fd647ba64aa3d95dace7fccdd6501fae33eb7959f82fc51196517bda58434f0bb4ac8bbbf87146d2086c2c506dc250515975532d23b772285aab9b9bdde7f3c1291f67e35ed053c243ecb1fb7f59996aec5b02efe579b7f0f27003b34d6f43f0be13667dbe58d2bfc607882a81ea3f09dd49a7f777273d9b98ad2fd4dab120a25a5d86351c6e1e735edb3ec813f8d2a1abf26759c31bdc82f213cbaf779c1df968fb2e26d19955e6df8419f30537f4f64a6dd20ad298ef9be741c1b25910facc6f993417cc59970ec5a5b6840b3218dcf51abde413288365c7033a903880b4199645309c07d9b6de64d1855b0f397322897f5e88552b127b8a95fda454c4868c5dfe13a2c1ba2d6c90ebdd2a5c9cded5854ccce2f7f7ebab4ccbea2e3d0cb08ca64ccd8041e88439c316c4594bf8f6393a6038bc71b4941c0812c2e2e400579696014b676bf9cc9e2a73a797b6d3a3368cc850886e4fad9e8b29b8518ac610644d14ce98447388c7929d29bdea415148dc94aa02ecaa09218110071a1c2ffb9678f1c91004931c5353375a991a416ca3412f4bb4d93968c2a597c81cefb2844baea5888b05a0356d999f858989e3855ffffbe9d9df54fca2a9ecc6d21e0d203f2b80597f0fa258adbddaa3111d87b341ec7c2ef2c81071dad101876255cbff3922e3c8c1a8c99be5f2fb4c30c6558e90c9882fe291a5855f5fa3356d6dbea2849fede50d4b93920879fa977c12413ec6464b8a0e7a1bfee4962148b2f3373af1e1de8a3d5c3da6a04d43eb55b530d4eed8169d64dcf9aef34f2ad1f2ed66f5026e9f5167a41b20589900c54f903845a2266affb3bfa41633e5db373c2bd605fe6ef0706096332fc7ff52fa539eb7b9d79953f09213c764b0e47742282a451e2695a8705b5b624b6fecd3715d7c50b62c29f5a1172daa6c12b8813d802de09d2f7e6b4443297b63b1a7307085211a3858ef3b5c689eabfc09ee9c61d65cfecc753ff49bdab87256fbc9d3fbc700ec89f660c573096993bd2c0790915c62dc62af64ef498279a20c574e51f120d588e3d630e9412e5ff3a04f54331d9e2e509ad68208cfac770266da1cac04b31c3aa3fd748e073422b3d46c9581162ad8dc973f613c8625e5b6ad1b96143e29118ff362fe739347fcad78c0f6d96f64aed2fe61a673f98e5655c0cee1d5c72f4b259f83cbdcb30dcd74461cf8f8cf0488e25333775571cce2bc563d40ca3378139806b2c7f7881e630a6938d189ead95a587450e0de4524599d60f5e9aa06acfe7e69304cbf502446451829c383af85371f7e473692948d075acbe57f7905cfe3dd73e1992df557e2a9e32725a529cf1c092d2785e044fdb222f4f016e5b36977377cc2ddac4afe16401b1e1123d5a3cdc42bacd7437e5d6f98609e269cc406eed7cbddbcb94ac8b2894a575e8e201295086a5a7ecc549287d2216426632749c0382037b4d9339f95107d01cd608ac43de097fa78522490e82a578d13bd999a714c76f50a34316a3951615cb4c6c790eafb5443c4e60d5ee96c10686a248145687f8e8c6206bb58519c22292cd0c3adf5f5d884be9e7aa167d53492966b7bcfe1c4cc7cf2974a0113539fea9a7cdee4d376d19be763c8ec3b991ee11b1aab25a10eef48c9cc6dfa631c5a625e79155d69f53593b8b4292939ca82b9f0deb2fbf2103a6d4637630a6bcb24ae367153f3c307cdd17d77c8e9166344d2adc3e30a04aeb0a9a6c4e7458b1816045cfc1ef3a5f05449797288067624842119ee7d9927434034b13a44e342c9bf26f0ffd1208342d3bc7d6a40fce95d4c660326ad66a5af897e61595b1f7938093c46336c2ab57c6989558fa1d5ad9b4477f5d3d1b8891b3e18cd63ff44f28a2193e8e6d5162b267026790cd19902851d0e98d492c57d0808f8ada5e327b6dea76cf95dea788d73b378360702b273a19d197462d7ff8bc8e6ce21c06493637ae9d8e17e3e5537619360aec9afc3a4a8559f5f8565b942662f465c98bce954a535936b90cbee2feabbd61e381d46c7f42f9b263f088691f7f000f2149f3c7eebfe47c9a45d4aa69ec43ab8ce35463a62acb8810d1d5aa84d8f6fd7d98481a194a136933f969a32a237922c1ab2229c0339115823eeaeb6e1ec9f402dbc56b6205b66359941f74718020d0b1aa8ed841bef0ac026a095b186bc8e34d5d2123c919dc9847a9ebc5aed68d859e0f417dc5ad83deafbee2e41895c44dfbaec7fe8389a31cc7ccd1470cc4b8a393d1b2053aa59c3af63473bb735199298aefd61b9971db973a299ae7fa15c4881e6417c6b7f9e15c9f49b6458e74fb6a0c346951769acdc5b3d36a5e34ea411dc799df549aa74ee2fdec9e5ad36749d36e60f5e04cbdd0621fc4c6e292eae13bcb237b88f2715c59b4d9aacfbe5ac3a98a62e57c15ebe1a4cf5381e1c4cc382f25112df8938167beddb1b4cfdbebb9274ff08c44ebc8297fda46fa39c5d0fbb9a855e8d10584410f9cabdec377213e6d487ab2921d256f84bbbce5fad429d24713b0a9e9b8e389cc14b72073e5b6d05eec7c6461a2b9aea8c06943bdc3e0bf091e5db838d6d6311ab1f4f2aed06d11bcdeeebe28c9b24f22d9f6831d1e78702e28fbb052ea7d12fd80e46e2bcdad47f9a3f70bc2c82fa69c67608449fdbadb9cc08f6972ac20959869d5895640f9fdc5608a4b37cec3adc4061eda85a27e11474d47514d6cb38c760d787bc5c0f054fe2d0a4388121124f1842cafeca7c8adacfb25ad85ea31d280f668e202bd05f868f7551594c9ebc185e938dc019c6bcbb6d78ba22b91c941f21822944bc060ce27d8b3ffdb89adf32c2ce841b844e45fd741f1f57fde8d7a4a5dfc9bb74f7be2c783c537876debd8e5a04b63a7e188f54f5583c97fc0f9804faab90bf025bc7887762d346c13e4aacb3ae39302eb49ca281ae81294317c1ee2532e398a9664d66079791bff758a47219ccf9ab40da9704a25458711981de641043fa7ce21dce4fa39b2b2112071a2a4fb818dfeab14c5ea7401d883204dbd62ebe5963bd416617482ba7fe09428d62d47960a7cee1b9e3f1bd394b86c6d9edceb323be341b11ccf2518a3a5d34711f100956d003ef4ae566ca68578381e82a77ba83aeea65b160a61c9f96e1841b2d73777a8929b007096cec29a0669a297baebe8c6503b9f4be49bb98fa13d697ac4c441f080f6643004b0cf1339ed2ee4167558c37bc92a1d8d848f8e69f615498caac81d1d2ca07d3350a5fcd2405be7f00e171c2453087433a1d26c2e61ca37b6be9b76131858557e08da19eaa829659eb7bed145a8a2972eccb1276fffcd9f2070b453d1085b806e6439b7689b93f00315e73c26173f9cd975b62291cac5625537d6d3550d9b1e84091ae7f0690b68678ab23772008b01cbfaccad1a4eeed22232c7e6ee0d2980fcd83d34bd7eacb93e3e19f20d2e75f2142f923a93f1810c4f6a9fc14977d5b6df62418a9fd74d8dd0c3dc351e037340c1b957bc8ad67ecb248d9f4ae4622a5a1b0f7e979533760fc8ca6ce3671e4b98f972610172c06ee7a31165cd803748bf821ebe55f72b9832b2ddb4dd0df3d26e51fa77b70bafb59b5e0487a72aa2e8e6d918578b7fc9e5a330b2e33dcf4a2bfd95fa1b28637a2d8476e7eeb32ca520eafefb1035b44c09f95cc970e907b16ceb6721055eb85480a854be84c5c2824f68792a76812fad38bc2ee0941b46554e4132c95968db82533514bff6b193f7db8a36b8f17ad92ee182e4ee48f2ce137a8248502654de606921a09b8cec72ed54140617516cfeb022a8e1f65214b1006a98f537882a521be3b21c91616149c76399c8f23426068340b860cdd0318197fd0e444e8068825c6e9454fa3396c34cb90a69ef0dbbbc6b39d5e082e2bc9911993c015e9776677842be70e26bc2728968de1c91af5ef2bb7f154d357fb25edaa7782409e4c1d2b9c53ae63e37f29189aefe5f0abb5ab3f26295393ccf0e6a03e0a09b046e70eddaec0a531a6830674886e710bed488f32e60b9df12ddc45a95fbdc9f8bcb445c5d1aa9bd5ed1faf7b47651233601c2c4d6011a435355d668f214c9ad11c00b350867cc1fdadce8d985076fde3e4276b1ae2763fbcf51d9d7f60ccf09aebc0789b9128689c33779d91d84d8d7b26e9475a509574c9f223e25bec0e400ca287c2472c217467a9ca2280796badfbf96a06aec340a05f6e66ddace20b610bef89fd26442550c7e1adbe2e4d0e59ad2fc895115783b4c059aabe4821454816f52e40164c43aa151e4a1566991a79a2dc5aa3ec963ed455686b719d3ad28e489e81f7b073ae2527adbd571292735d172d880053e9fe63610378222845739e0534ce2091270dfe18f34ef6a8e89c7556b1b5109dc70cabd8f4eaf2d3520f67515fa8a2fdf7e6b75afdc759cb5f69cb498a6943ca04df89b8a4c39de9d0996eb1a0f5c7b98be84494b5430a8cab53e4393b06abab5d5ea2e205bfba134f07c5190b83dae34d60628ae68a7b5f8d3d22f0f752777460f4ff94ee958dba37c5251a90bb2e09c50e8cad8882511793b3206468ec17156e74a6a9c7775da2d2a5284ea8f98b15fcdb4b8cf87b1e483cdd52f6e89f4025f87aaf83197ba39bfef1d0d679d32f9ced873ef8a4e167ad4a7330f2b256bd4368aaa9ce1999d2c6a855969c4286415979b88049a3a69eb58891b5e973ed3dee0a5bde7c22c028f8aa16bef2cce9f15a4662c806cff1a910b751fb24e54ca5539bfb5b4c4c1b482015203befa3b19dfc80b0b9d8eb0004f0fec9bf69bb01b4615e370badfb6bc4a815316c43959860ba8eb3d5f8b49557b04305676f9cd23bf601070ac61bc7be5f6d6c847a14714238e0a879f29d7186868cde8b003f39b853f8beece43aa6ba99dda7e32;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h87bfe5fcbc946f2639538df62a7a6b0aef4ec011c4ef4fbac72e2b5278973a8c377fe40adbf24e48e432dcc4be9cbbd31f6dc8786ea12a35d6d73755c32840c563102b54cd40542e396e622dbe2bd5bb14c2f887aa63820918ebcef161b0fdf1f5596bf20cbe64233d50bd00529efe1d024e23ff5a8fd3dd8b9275e20a554e8914d496b968b9e149fa3b019737a62a76771d901be04c151c20b6abc34209bf70adebd4998c18c9714c904e13dcefca567059660a65541da38e0f63370b1da591246761a0afdb22a91dd5d9563631799f48fe26b9dc46ca16c024717f2782387bd14cc826cd745020c4c8b5630f54b6a609ef48a65d2bd07e1956c1066e9f4f908b08adbac6edfad7a1e69f3d31c88044c3515b0f73d64b7d9d22bcc53bb2a508a065d170bed91a1d25cb34f76723d59a853fe06fc589cc9dc658892e8b3d444fcf2cb0dd7d0874e898c81be3f01b6578d604954f93752236148535efc155492fab4d6aa48b44a0d4d43bc8a8a840e1136a586af03740338cf65044ed356b0b5d058fccf383ffec69230f7323ef8c3cd097c3ae3a71a96fef3e2dae4d1bdd58fbce867f58013721c762b96858fccc356782adb13ddec337ff7a4e3fc7806fa9b6398eb86d86ec077ed63b673b12d538cda59cd33894be2ba730c09b2e0977cb17e4546bc6dba6fccef2fb6c1451344a6fae3798cc17b0588ffda942081dd21392782900da2f878bb55be01b86b884fb9e039a33ae168dad6cca4808aa3ac7a49339322b6704498575bf7a99868393bc2693385b4e4b8c1f74239dd22c8ab80dab35558e8dfd7edd5fc1a3d42dbebeef57bfd2f9ba7e599640c61ce132622bac53efda69860697b19131a22df458209e380c27fa02f0d3bb0e86e49782593a86a50807c6d15a5490ad23bdaca8aa264819567f80c49296fffae02d8e2135840a54839403b3bf01e00aa282b79da1a379c919f16a95ea9ee91ce41fed153596932a1bc80d7fda80d409659cccaad89fee4790c722eb9884305a46827aa0a301531ed6f8359b7c18f1a8b8967f6f7c1dffbf701068e37b01fddfde7a6c9aa0cfed3f962da835cc13ac49f66e8dbe95ff3273f1f6cbb8991c90f05f05310e05fe165f82a520dda5ae379f83651c6fa5b71cc79226fb811d40de5ac70c90e2ed449d84af13c46f4feccb545a39d70a11038c6e536dad7ee832b98bf3cc5e7f90f0292eeaef7a669509a2f1850630c0a8d5e04dd8947e010035ef26035774f062c979b029a48cff35e0f8efe5831b13f0128e3193d6106fcdfc24ed73bb5c4f7bd076d1f12ca37bf28cddf51ea37a22b822305d2885b1da2bef18c269baa6881c83e3bf3a7479593565125e53f8068ab95e36441fa589dda3bac2d4a1ff4c375b115aa3e02b0ba59bca425fc60d19b720a766d55c0f5f0218521a0e20772ca94ff1bb58257c57b7a4b2164c78a5090f0deff92e2cf21e22f6775e5241e3e929fa31cd9d2cb874e667a167987d3737316ca4ef6aded16c98ea92ee356bd3025c248d5d50effbec0fb528a1e7ed8cdb0a68ff108271f73643deaaad6dccff4888aa398bab5b66f50fe4adef41bc07ceca9613d1f4d7a048499d72cdae60e13326435633c838e58eeda4915456090f6f8d9eebe91bcbb0083efe431066646b712f83420adb4c0a76ed88f9077899f01671ed67d93daea64cdd9e75ffb6355a4ba0a61e9a381506e8f7a102efd4faa862f94eee541608f7a82c528fce3fcc661e6282032a425b712942adad0dfa5655dc59050c648041c7f6fc817f5b9c61dd25b1cc721ef4641c9f4e24506cca6f9b042769a95d2903479e773730bba2489dfc34f302d84b0935ea38bed80b0daa312b96258eadfc9f169390334155fca65d1778aaf0dc83620e6c0eaff1e39377f71d17e1a18b67b225127451462dc274c374b10b207b02c45467bf1f588e1221235dc411eb621f313976a323be6da6b55c6ad4a096ab50f63b418749b64fbe7eee92fd1cd4d6bb7b929faf57eda5ebf91a8144832f1df06c7668c5227e3e8ec378cce6b7abcf5bdd33b7c3ad2ac8e96c2a3ab44768ba87516c28a7fb1ab2eb756178fed5f60ddd1c99f89460c2e8d3fd05e94d3eb126d315656cf0ed43f0131f7eb1909db74465c8dab41c6bfa4182c0f765b675b37a17f087c8ef00b7200cf57f3e0ad30f56ac709e98213b0325ca0f4de7a4a950020af95fa8fcac4d575876bb69245c6465444841e973357021dab8292da410f1d70a5f69240415cc3be49568730e4fa174d8e4418558472e30314e4431ab2aec6b085e79e66940de74a251f926b6d3377ec50bd80a48931b08dba979bb9dcfb6f1034f89851e52c0f5ea1e269018d1e96ebc5398f840589bcaa44412f8ea3dd0115d4c4f9e28217048495c2c358f9897feafabce3dc48b5d07243a6550576ac04bdcd4f57398a5131c6c5ec0ba5e2dd1c550d4ce451cf3bf8cf61d0fcc9c8360d66cb5f3e0839f6d8b46f40aae9bd8a0cde36e44c8c4d5200206de5378c1ebf5d49541178126119ce8a708f046ff172d00aeddbf6a9c7e8a85c96dcf8b1112c0d3d3c64e51015a7989952fd44fd72ca3815ebcc129df917cf4694b0c87ceea3a1848d6641985717b2fbba6cdaf81bd78f05defd0c199e935681d5c49a962abf784a034406fa551c8ae3ed8c65b606502bd68af796b2f2428067c26c9f4a4f6374ff3ed5d4f64ee9522af7e47ed3b91e2077ee3555284d973acee934872066274bc7cb7a883a846cd3ae5afdec45e6a6d82875f4013d1da5ade97158e567b005d5539246357a02e6160499c7e3fe8ce55d44da694e26691d8b1633d2bc77f8305d4469be741c8b509aeada10ccab8888642b26f0bde603a7c9caae780f660560118fbd0c7df0d0636c3291eaef8d3e2649f502d2d33f0469a26412c5d7722003690f0f6b1ac2187f7a549a9a7803f9e2ab7e9092b14d5420f5fb000cded43238b495c798c6af04d2269a40561afad03a4c343371875353c0e9367e02b30582063a8b6efb09fc493dd846d3fb94ecf2dd6b0bd650a291b284a04da0e962ef6819497909145d7e69b75a0515e16190abf4ad1bc08fc98f051a75a40f4852a4f50ac996e20041ff77d528ba18688cc3b505f9232c74ac4d35c62a575bfe9dbdcbce4eaa9d0686f689e7dfca58a6016dcfee3e5391e9026f6259a92f4cb9637bb32f22b84babc83910dad2ff6ac7f76788707c9f69f9f9e2327fc301f0334e2c2af1ea69dd49c10883c3fa44967b7f7ff93294c8803bb9df40433e98ef2797d898757a7528fd6d33f98c65fc87179c9e9ca8e8fb7c2dbc64b7611afefb1fe580b80723033a9243b7f7f68a100f99f7b2531011a41bd6154c7b9316bb483a9e272613f24b48f32d794c125f978fe11e2c6d822d9b2fae51377ef3ed25a7b3bf25ba0995c74e275ea4749030b706539f1e3b4e03c8783bce1e2e5d8a14cd398a9324e2f12f01ce9a6f20bc811bddf72c819bf73e60eddf60fb967ff2fc35a9aa5a7d16cfa96cc2cc3b8dcec4c48fa95ae5d1cff43f1ea80ab507ebba3b13daa1eadebcf5572aa316712a21fb665c78991d587f04f84cc7266aed2a26c66600e2774159932732db59378914603dae761fcabe670e9ae0bdf0e0aa82510c5c414e0449b376d6e4c3da7064f6f0547613eed40f833e11d2902cc7f5972a490fa49d174bf3dc6ef4dd85597e93932701466119608e0b6a22cdd8eaade2516b5332789d5eb39ee1cdf8aed47abb0f832622af1924a52a5cbeb3a7c529730476c87b814901b10c24d78e8b9f8491d189c95c89a3ad1ee5faf982329b950ac410020ec9b09ef3eaa4467e0fcc11665984da4f3fce6f2f54caf273f059d2298be76593b7f2e02adb98be6720372ef19b8a2e35610c0e3766b7d8afdc6e3355d3bc178be236f6ed8a4ac9430db33ba174f58e104ee1a7cfce180742597885a9cc07ef16f79ee22a8d94ee7c6e215dbd0527d2f4e62d989637ec1e2f8bbd581dad7c87784ad1f9551bd2f74893f21eebab577ae38e41733b95e60fc09dea93bd6143a4845808e5bdf50d09930b22cca92402a41a481bb8c263c0aabde8e856cd48bdcf0de909a7bd4cfaba47e3a336429f32c873f10aa5d12f197adac006ee1c151062244ba8d757df5cff679567c263f9ed05043a570f90e4bfbbc21de5f0a7ae5ab011898d99def9f8521a6c0ee348b6676f6a74c790e32536549383a1b4529023b9c8ed7706946bdfecef4aa838a7132400bc0ee8aeb1bb6b2892507e61aa4b7fbe793ecc3df8e41c45a5b9455357add29e05b3a6fb279dca5642e905c47af3db55b20a00f763b137e11d88d9398d4adf87c95a15f57d439843197379b044ba76c1cb89083d3014d23a2a05e946a676c4a8192c380c33d7caedec8205a9ead119fa6c5b4cd15bb7310567d48715352a05d4a017c4e0d4c9bcbba2126f2def621ed3877b1f1ce7e1a89de2877d8344b51646ada35298f5c647a04e84362ee17ef0e226303ae872ac1b06016c4c714d35e5a93898a561ffe20acca93753d867c2f3462a29884c8e56cf167e5c5d9871b6bfadf362e3b89b5c77fd0a6bcef2c1b25ba6e5ea72c93c1f281870fce0675eb84a653bd0b2bf286646af7cac2ea90c033056977b206692b51b6115254536c578b8c9163f102719960ae2b167d09b3a78d7a8461ef7daedd003b5282a6b3c7e0cbc21e7f92ef6b79766ebc6da879bcd722177e2f291c54bd7103809c6b6a0f5166d80185a3bacdfb37671ecbd0311ae03561ff21565955c1619659df26bf09c809d0d7ffc1c32481b7d227f7846f062877cd6159a04b05bf0a719933d0bf542095e2e40177b0dcf3bcc7a6e2f4f255458857f870d2460f5c724a3941ae84583dd5d5262ec55e0a18ab54026b1a84f3dce36da12b3b35ba626185c2e94390628b7735fb93f3b10939ee2201f279af6a19b8e97a62a005b2e15e77f2ed44ca2be981d2345c360608b31a53a237ba16f39f1b68fa21dcebc0284c308c62267b89175bbf3b58f873b44e33965ad8c876f32f402a1cf21e34b5f0e4af8ad5a57a4467e073e7f5346cf19adb07da0a5cfc6991b255d8246bb5c541f6da6110f7557e2f616414568274f99b66c1ff8395ee2fc162056d35428776baca15bfe0ed6a4c416dd0991dd36f54548958465f9661cfcdebf13217d5befe295c13191838750784c59d7de77242d660b20ca83ca86c659a7bd35cf467282b9b2d4c518389ae623848725750f1abdaf61842235a45be321415545ce6e3ffebbe0350ee46de01d16bba52d934376d190dbfa02c656b70483f2e9b69cddcae4f1e40898b5a2ee7202443d9c6635bd13d444b1648f2aa9eb95b5a896c061b253607e2b3207b11eb9ef2d1c0a1f5d39ddde3f6e1cebb0e017012e53c220814e6bab37a35ad7f4025b5876391093cdc7fb86e5c91673d19147c33ee2769a1192131a80b433c090c112671dad60bf560290a5ebd6b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h26b44b2515998886a88f3aea13bc74f6e15cc2beb8dac766881d3ae1f946d7446512d2453677afa7885083a470e2af9daf5a4e650a387d051ccb441e04e98ffcf489c84bd9be0eb41274fda03c9f955bd30f3f004789512867088bfd8165b3f4977f10448e9729f29859aa17252da92b98da5957bfff6a8f49f3ad2ed0109c5ce99d83347026d0dbb805b5847bb8724ae8a3310612c31f76cd39db76e4f8d7edfd8099ebe06144c1adb520ca5b24c64fe0feff7e91afc18914d43855a35e9f6fdde61b3ca4b55958c1030f25bb10e7c21e31b2fc1579e5441157e788c84f3c163cd4eb2bfeb5467136e4b998494d7f3426d6aef23d813e23ed85734ae7ecf26eb2a483c9ba3539b071e13e61c0c7ed2f1f91e01b6f75f32d457051e4a13f26b1ecd0dc167a861b8a5685b63eb463b14b3de4526f02054389374ec6dd4b077a4118bbf5c7915a039f1f0b5eb47c7e0c8296745008113ceeeda54fd04ac6d55fcfcfb52e68f23cb710212d6a588a1d76210aa9c8673f9fd48f2a027b00c137970bfb5894572d1b80cb077d9396d4ef8e35926aae824d2aec02630083bd89e5b380b877f8fc04b4a63d51ce1a481cb45dcc31bb27141f315d0321f31a91a9cd8395a1ee90a39e6a4b6c1c3d1ae1849f609a81438743bad15b6225ad3d00ca558f2d1a4bbbaf577a625f540a31c47a1e4f6881a9e960a59c43357d026641c793dbca472cc6134550f988bc7944605069dce09cf51b4f7767c47384a451488d93a4461626ff66598e488d756c8884bae2764e8dfacf7fc5ae4b780d236ea3fb17f274f11c7176dc0dd4ff8cb4c7f375053f856792420c70288ea2d07f48ac9e2694031be7ead1af1d6a64b1e77a946037344629e215fc0c334df296841c81ffb9afa6041a98e87c542362db73d4bda947febe58656369c9bfbfc26bed4666938ce7714d24005f0bf6d3f5f6759e9fceaab4ed481722d743ab1c5f93d5760c06538a3321475f67f72679d75ac13ade609fe4d276949fc36dcb6eb6e68bda8f81d27a3c084e54d81aaead30828095aa928a877405f24f604b7bbce5878a4d9d2ebd4ba46ef917ea82871ffc0b3d9d80a2fa975c310f6c8dcade0376104f4402cf9ad7925d3ed5b9b5eef8fa1f786668786a9a85e5a56344f1f36ce307f5cd4524c3f1e6d851c655e4debc213c73ddbb4d4aa0460f50dc91b9e236b9f298dee0cae4ae427bb377334438773590de61f08876d6be720965475d2f0d4ac7ea3c9cd0e6cc413005725f530a9052f919f3ba14de38113674e1ca0e56e705902865fe82b05097dbdbd357bc4a3b4d9462e16abec9e122beb6050310c38d66b2b8d8e536a03b6302c4eebd7781e85721bbb7c7cd923ebf1954b0be642801ea523882c88bb1f695e6028edfe9d4ed4c0476128dd63fee4e71174abe68df8361f1232961bda93e2c88ff7ba75c57aa404658f63c43e0294e5f39c826e4eee804f5b9b440086d0b5855abe152515b49f75238af8a7c98c75eace95722e47c61fe9e5c339ebc99bd708c3f82b0d0af31e118f4bb64d89552bc98860cd0040604651df04d17cc59aba16459b24cb1bfa2cfc403b624edb8f1dbafb2a69866c60399e244534250a31bdc30c40b01b9bd5c8bf3e47335eecf263aca714253da1903118c1fcd911cdfb0133cfd0a714e042f5fc9f0fbaba43c090603c766d587e5c33ed296f64255dde01868ed8096681e3ff0fa1755f58de088d1fbfede904f8255b52907d03a561f0a73374b4e0c5a9cb7b2e01908e4d8527e58df1089edb3ab40de4d9c3c2699d0f89eb832516f2e8ecf8ee9a31721e5cfb1243a47e695185a4f4394a30765dfd6dfca8181a28b072513e6b27558ea88587361bc5e2382fb698b0030cebe3fe87ea69e54938aaf25b6ff7acaa6223a36feec4b8894737837067e85a04da8099356d680d103e00d076d856d71400517c1882edece413cfe19e866f677d72ecf1ade4bf00cd79b396e0f5b6182f50805d75c05c3a60b106a36e13257a460fb13b9e1c783df093de6a6305b36d9cfefb09e9dc1279f9ccdcb9a7ba3e0dd049cfd53f04bacd6699a86d30d232f755f9ea6e35f045c805fd08a769782a0ddaab99c19960d62011ba5bf02edf99bae2b7f752f438ae25822faa4459ac6ee150ed36afef175f36ea737857a9feb7ee11785c750e636da7c7b7b818836989ce5d61780a974b75dcd19c3ca6d20aac7fb5b751500d284de053c6f92077c148997deac59428e5dcd5ac4c38dda4d157002a81b1beff948bb21356fd51a11b8338b5207aa2b4123f27bf8b6e7545a70f3f2c899b9a99d6e3069fd2d61f17b21bf199f313bf549a3111be2dce6dd7082ed2530606daa17bb28e17667a781ed7ec2bda2e4685866b2563ba1cd37a207bd23911268c93d8214730461a755f84164ec539c5c8baacf36f2ae428ce2d9015458efe1fde5474ba780d785a4baf23c9c30db234f3e9f0fa68c8329eda4d625b43b719d505bb27b52f3641bc50b8552b61e71eb6b310e0d99493013d17ae84556813ed44ce2a0f4637cbb4d4f3d1b7d8a9ad6c70fd6b50dd634a10079060afaee619f02615c9669454efba1c1ca4aadc14b5c9ce8bcf5a366003eba51029247c7d1c027e2ab01556350ed2ea6c9713de5f59b4d140247693372f5bd77da0bf9017f5c65cfc3565dd7944affd1c6344f13acbae60897b220ebfcfec151cc113b6abae400abaf31bd5aa26fc38b6de2ff3cc3090c1211e51235eb8ee232127705432591b85ae79dd92e2a3f57b0144413a9d4d1424c16d6c360fe54ca07c58e031161ac69a7c234f728038a42da2797acbd4ce709cff0d0ef597afe828bd1ea170ecebbafe249207dd1a10fd58d6307fc628ee5144db167be2375561ccba1186b9eac0c51e6518c75098c28fefcbb696758869259a2294fa010a6663699da9ec8799ea02296fab6141f35a59da3e4a820a5150c9c9c90752d43ae2ad1f092ada1270da896a0ecc61a6ce3cda8407d8af441567ed336a4e853abc52ec1a7a53590256fd5d76149a8feb5b950462166aa3d9b03d6f932d6dd6480c8c1b7e8f27973beb0570ef28fbccb25d173d15e670fca2726898b3f81fe8ef80e85b6a7e85641463bd17e4df2dc1be984ab6c38d9dc22fdbb54163eb9bde8a4d9f46eaae225a229e744ef2f9e96a7e4898022e7b6bcb0201de8d5056882a8dbe013290f32feb01f1044377271c462fff35aa03e9d8318a310c6829d02f5c00c37b449432a1f732766ef4ba31df6ae0cf6c39f25cf7b0fee53ad91a47068adff865402b0fb4f406071f52010a0320fd10a70533994a6235f5ad0e00f36bf4f7c8f58395ffeaa2729b4ea92de82480996a591b6e2d984e991d0b9e8c2f956f81186295aa2ddf12730ede55040d5750121da6064b8e4a512e0443cf131316b329c6383a7546ff97dc0b039cec04fb924f9a91fa9a43c2786078de104b8aca066b1b89a643771c4f9b8fa7817cbfed81e85d01e63e4a80d60f0953f0db4d23b09380ce39fab9a1c5b36a413236d802edbcc1263867082eb261abb91ae9d24bc7235bf7434ffb75d44a41cedfe5ea381a8fe1b248c4abfef882ec731bde6a20eb223db2d66442ac8a2cb81ff041d344227157cd2f3ca96b2eea4b7615cc23e27fb8fcb2baf78a0362d9736d6f596ae84e73d64b0ff9e7d663dfd92c1865d0451cc172b48600eed556f593cfc297e1e0500ec9a634c5ebd2a2d7838fe06c72fb521c0bdb1c06cf281c0c47d8b9cc3ea46ff4b8259f847c4fc7f87d979d46a3647aa58520d3636c453aae169a5aaa522033618434640c710a7780aa57019afc529951fa1d78017a3c6ade4b9b7f1f3876eae1a5fec9bc7d3179e3b7960d9c905899c4da62f1955b08cba8632cb6bbed99112def2c82b5376058e9b2e1cb0436d7eb45969987c6b800a8cd892bc59416d9f28edaa49a6e330925980e520c79c433de6ff78b25f01db5dc48a376e4609cf6f762e9e6f245222c04deb18972763ea92e1a539a57ef0b2c4da8e78bb47d98dfc64b4d6e9169a40b5060c08b2e7b3a7595c817aaa54e487a5f4e4d7d95bc7515e2d13572547b28542ee338d9c1b661aac59b6bb75354bc666ef0ff85c09af5927711d2a3db6a677465641729367a73312dbfdfdb4a11eec100c73d6e02798c63a2ce607fc4b67a5dd9a6c4e78d12cca968000b1ac2fd247b0deeea338629a3351c0b6f96aa9a4163ee81f7ce78f2e4ec06e54117d10eebe2753d2e5d775122c7406dc81a5c3046cea0107a4ba9b91776decc8a5ff13944041be102dda14f983cc52e724fb051fdfedae4ce41084daa1dee86e4fe274ffde6ab8b69951de1d006131b1813992b14726f3111bad08773ac832f2388422930585dca1ae74e6e8eeb4eccd2c82fd5408d548b632f4c1cfb7db45c94a53124d1457da54168d4dcd6745e4d20bd15f0c06075aaae1927fe5bce7e5ee0103864dd9fb8061da3a607acbe20a7bfaa3e4f17900f99b193b125f7a528aafc5e6b39f323b9a11c66df2c079b8cb38ba9358a57f2e5cad95332452ddbafa9386f3730457cbbe6b2a6096d8a3b1b957d0dac67f7a68bb63b23764750c935566a667b798b07ef36e506d31731ad357bc56dec1c90ddff0cc89b9bd061c794eaf8a36222291f21c0013fc3bd569becccb6b24db8fec5dddeab629ee3c6cfde220df376eecc00bf2fecce2762ccb9ab4903847baf22224ed5d41cc71d1926061e66f5c2551e41772cad53e37e05d1fe74a669f5431b9336c3db629cbd7add1afa6467cf5af404af3cb5ccf019f513fe601b92b8bb34e721fed5022d246fa79068639689c56ce4bd8afd21054ed03caef702484f9744b1583c365a0406ad1eabba93d74be7cc4e6da26111533124bca0aba96564d032a0ba209f4a66e135c55d6a74c55027dc0a6a898f4ef59ab89b846651cb9b089aaf43bf0a7b02821cb34b7a1948df7d37f27ca7fcc5d5fc78c2e720d80f83ecdb7d8735309efc01e648e36dad772dedbe5c556e6fd7adb644b59761670603e9e23cd71f51ef6ba8ab2f3f2576c466312e37f7dcdb162e7166e79c6211123a9fb415e4da84199cf7c4afe683ad357214436e0ac4292c30aeed265d4ff3b48af90b60358648e1715e1a77cd6657789834a215967fc6c6a987dd91a12e007ad8ce371fbc1e584115fa6e84ff88602a67cffb7aafa6d2aa49c8f48d1d36764c2f860fd9c69381e86e07c751ae741a81538488ec7583be0cf5c6cb6f3c3069fe5e7ad7884e8d648613b244c84d4a2962c04225711b00fa31842b8d9ccf498ccd1937632c01706de4629a3545a611e8b5c12c3ea61f97157246af161ae8d3ee2f92a12f97e517dca4403a0244dfc42ad39e9c433ad9b96ee8985ffe42e7b37f2d0acd3ec971b0341fa135acc95a2b33ef7d47726977ab89a238f9cb1f78bfacc13d52e9e5b89f5aef5f8d5be7c80886c1b7d5c58f8211a2abf7b5163a00d9ec3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'he2878b8abd7554b3dc065f32802956274627c82bea1aab787af3690578b9f99b2a838572108c4cd4c98d9bb8bc5ccc566ce24c9f73ac7169c85450aa3d59bcfdac5c7b3c5ba62edf52e6d92448d778f19faab00a4de3649d4839b54d0355fc332a9426bd1ed24a3b0db92bc8906e7cace54fa6608861f44960679a125fad77e44828f8a1f4a5c3f55d4f91f6a0b070648bd0688635e5c92eed20eeda04bd100cf4a25b8a7fede71d442e70d4bab9b0191fa7d0c6f5e90e30b6e87a9250a7e4bd0d4c2239a1deacc1f3d67b5097ced17cb16b94b6393a57fbc537e50ee80a05f0574cbfe28a160cb6436c8aa626721ef767c424e4ca31f221d0d8e2f9fcf08a0d8b45c55af73026a3eb28d6342b3048a26338a7d80c2eac8466046720c71a9f35f7f98c762da5b9f716af7e125d2d0d6c221b33eb259e1719d73170b6dd3f5c015d3caa5226de355f7ff9bf7194f4f9bf364b84daca420aea7340ed6a0359c3d82d604f03804d8f02ffce8b9b3fcc752571e633eb0ab6fde5295a3ceb28e11591dd3b21f20e134a09674e036fe7697d05de3e06fc428e4dcf97e3438f4b42ca5ab9986c7da51af7fd94364939315da02a98af372e3a230490a0674856dbdd62dbb823d5f6f40a2ebcefee71f44208c3b91b5f7cbf62356f565fa2c88042efe0f6944eec53ba12223c1d58b22cb28669133f3229c3dc9d93cd1bf8c1570f97e0bff47d8e053b88f7541981f7ac4caa497480a39675cd77936463928450c693dde37c91a1ea8584a232d9e73d4a8eeede4b5c02b6eac9c5bdda043e6470af210e993eabe865dec54410579a2d7a4feb76e8c4766a40a3fed312e993d05bd93b707d44d9722a16e1637773340294a7061bda55e496e707eb328b41ba8db7379fc63ab356b7a795eec124b7e267efebfa08baf5f8f91d4daa70cd798f248196736dd0f46cc323de4e68679d27fe30697fb69be4f0d2334fe64cf25765dfb4eb7f5c8a343b675a68c13d862350be1518ca388e6b9d40f896a4356042f0cc2c90fb68559494eb53e7f2d6b2fd0d30be393b5af6e9963c16e756bc1de4fb7fc65e35894c2eac25ce42dcd2048852d4857bdd35ff996b9fee0ada6bcd07c8c37a861bcdddb9fa75d5ee133dc9b6351607ee9805d2b3fce5d94b34898391b1089aca260750e68456816b40a0dbe1e21620e1d88fd933f4de1e879b2e8f477200445aa69a2335cab38136151e5d70ba1d542952d4b37e9fd505dddab0425be84289e647b08100060aa522f7179eaeb36912cdba55eedeb744fd78d2ed193fd88a4ecc8182778a6190493fc56a1234ba41b5be9710f2338774d87ac42fad3924e3c02b70d59c61cd5c87d628d80569261fdb7e8052e0cf40b1029d60a2463dac92bc0fb6479cb2a64082c0b9d13cfd02f1ce1fe2405fda03bf9ab89f97189162ff4b475f45e887a4c04ddd9d7011e2e063548ea537a09a4f0fbe2a8530a5946ebc6a182975e1132cb2800ceaf18b7c060ac8adaceda40184952298e81c6e47c0b4af3c4d748b434c2006d64c04afa244bc200be7bf2841f728d46df30982693097a55182295e39df440d7906221201cfa4d6d6f4fe9950b139f89bbcaa7007d613adaea2e249afc79aae5f57829d111fad188f4e8519491c330d23ef596a5358cc7e6ce5c0a00b958e59c88b9cd543366e604956fb8fd5f311a09dcffcfa17b5f25a0025a27a302a0792415bf6356336bc3721db005802f19a530dfe437c6055428443b4df2e380aab62b850a77515b7726db030221e3d396cf847853769608f7c91d0f4a7c60e2fc487e386a6c9552ef95f1f0ebad21b1730caa2d19a5107083f9b8acb5b745b1c11f92e34bb07e91c5817e70dbc0baa67cd924d90b32c439cfab0b9f11d11f5b2bb81968d89dee60895a9bd28bbdc3d57a1607d6e95108ec1a4b1adffcfaf7e4f214970304d4926d0459e1f047c0cc9c8ed65d965414aee827d2573b0d9a29c4737195dc0042a1801398c2acc0b3d531453e1da350a7a3db0d0f085fbe89e59d55a2fe5b5ff0345c2e5a5173c07b9ee63783f4826e608b3d307d36d3c75508e36f32f574c1dc6b33ce9381d19108d49c8ca2df339a18f40f8e53b26b023dd420a650b2e2e94fe65e3eb6cd188d64ab65adddea98465b9884750d0e7a3728d2a24fc851ce90d2c3885ad9a58b8bff0df53d930c706f846536a5dc012a481e9385f689791f9ecc8cc4340037e96462d74d1dbd21d5ef8e4dcb78aa8f16cf9511e4922993a34131872b987b14d364e5452280567f61be51172d1ccfc362272e5e2025b0d748a2775b0d0432413b78fa4935d1a46fa0c8bc177d63698f9c170c1735d1f3867b72c6d9b01d5dc3ab91fce78d6fe9667b85828f4f98a474bba692879d5777131663d9285d83906937ad19c0b961a34ca3878adb6bcd4d8f054f2187024315aba5c287b44e256bd17b8bbeb9790a2a8b14a7d246f83de2e99506c43b799641bb72c676f52a4e96ffe90361376ab92d439740c53167621aa34e0af28ba0b0ec38e3fb0058480a00c234674009c90276223124e6d9b92cf59e50ff43f6f0ffcbfc429c016b308b439b6077521c40137fdce2dfde8cc9b1f5c6586305f62ca4e49457609a5730059a4de0a02d4eff2cdf7bda745ea59ac001d18dfe35f3318d25003c8b88808efcfd74b48c9db8a72a7bba74ccf8274c1fd1fe54251c3594f787af7c17363bfb207e348412191f546d6685bf144315780615fa211012914163d232a53feaec8d1f11790d580959d23626edcf475e9ee1bf8ec283c2435d8ba04e2fff5cfe0391c8fc824a771930d7c6d606cc6345d991c38ab3b7e401b7cf237014176ded3a9b158118d58a9b43ca138a05a42ddb15787e09fb77a49999a186a86aa767cf3461497aff5f59ffe820f8405487e4e41c4cf73f9425e58b56b3859040b170d38bed78c725c794173e74aac8f221a08a2e35a2a730875ec16a18c023c48ec1f8eea2b0d8d724317c41a408a7f90a4686455b537e5caab08c1e489cd4cbf31e97da1b0bab65bdd5b2f2ca083cc71138727ca9cb3b6026159d9f3b22bc08595af953d1e986e500742a66810ac244a2630aeb4c265936f64bf255d67c3e73128ed76af0ba8192262a100cd34829284d513e185261d1abdbc32823745194d815c234856d16ab734ddbc289e43dbc1eba62b6327c6d910388727b62a6a12e97f4a4c0a87e42df1ec5545531bd4feddcebde425bd62de1256958bcdc524f1408767b351c0664ba710a08c047085c67e3bbd5457d31715e38d61d18f76a6e5ddfe9be5fa7cbbde1a31e17cfa4fda104352044b04c0c5980b3f0871bafb9ee94cc4204d926c9aa8dd52bc009abe3b22ec1ac6c32e4f2241afc1ae59a2ed15f3db1b34f88cef24a15363835e603d985823b49b4d8bdf74fe04a74552b03d35d5f09ef7fd15d17e2dd33ab2a16be8162f4190889ec700b580d95d6ed4ea202ca225f0ea26a5b6a202c42279774405b55551d3945416ed1e3df7cab1b2faa06de074d84079becea4a6909f5be42fa858c7c91f851a46b46951c7968945a8be388412d851449a6c5fad94a04039cd8af002d1964a68e1d5b0830df6d58ff1f9edabb3b639dc1ab851533214b9b38da623b70771944146639214b54b42fe2fa8d0d10dd6766cbc6ebedf7568dae73d883e3c64bb7d5da462680c5cf7ca0124e711e7a759714e9f25c6519138e9071b5c59883d0872ef5a136ce70fd406ffc8d376ce1600e5df3c2f9e94b640d41948cbd42ecbe77ce57624726056b39d2e10bc0eaf2ee0d04903ee79c8412185d1449da328e5dd13f7648bfea4c3c3270071b37b2b8260a6d7ed0c79d9eaeea922423cde1e52b38ca86c4973231263c65b73840f975ae165a90687c3d67c13a7a5656584ec07495de07a3707f7fcc5ebb0cd4d0c1e5596a15549714557f075733560d43efc42c4de8d97b34703380f79da39a4e9e6b583c40a7bab72d668e524bf5f7b2c5dec238ea255b8a74cb45c8b29227bd8c72a23d7cdb401353f17be7addde1652351c3f194fec6cc4a65807d77fafdb7e4b5a609391961ea07025223aa8e4aed1ae826677cde6b534e1ea39bdd2c9e79afa861b55e62dcd8895b746275ecb30b76446e064f1ef03ae10f6257ebf0ea8b639282f51cbdd21989a93b109a932dc9347b433adb9309a3eded324ce06bb5e6b9bc447101f05df8a820d53f5137ff824d6deb5b7f70ad49c3d19ce03c6a882f8ac89eeb31a5b2133c1c81eafa24346a32a6ede005834f007fcb72e33cafc1adf77deb7f5e19944adef04caa9dcc1f83e099c21deb8a35e0974ce7da29c734e92dd4b60ef0a0066b5aa025b57bf9ec9ad4ea399e7e5feaa57e1dba1b31a047b5653c82f07cad0be9c74926cb692c836477e6b08da05bbb1f1fd222157a69f3de4210faf2edff8c4a9fe85833a018827cbc32e44cda59be38e95dcf576a1afc59a7251427ff4183b40edd3636ba6c3983ed20f214c3cb00250d39205e2a6632578bee80ea08d041113292d97af7e1c77cbd869e7a4d4f5880ffc676c2b49e65f368ce1b8fd60c00c99ce1ecafc613b4a66dec4b813d3e70267e130f979a2475e3443ad0c94dd19ee9df2c42f569ea32290f35a1aef23bc7f9a3fa35b4e4112baa5e803e741909157687bcf4e9ab6f0a62ebf23dd531a732903d5eb9e0e475b0606b80f963af1d2c74634132759c83e2ae77403d0e0ba402828a0928c366e17507b8fd337dc7b1f067924bfde8c54462c07b4eb2ec09ed04e7558771e8379d807bdbdb7d1c4afde6289bfd8e3be0f257a3ee72dacd6627d32d994fd127d21fcf8e6e205b223d1789ac4a9eb7e903eaa970dea1ea8b6525d86a1356109ac432f07a4b660c6411d20d7bdd290c3a3268f20fc372f70871de983d8495e6ceb577e7ec50549bd322573bd3fe85f777fd7cd70e7a0159e538c15c0eef8da6aac7c73b7faddf29515f59574286ee7141be794758358379cd03623fb3af4cc973c6b191bc2194cb12c1bf02aea20f00f9d8c94645ff3344c2cfb0efc01582e0b08791cc9416c4509a92c514eec8f53ac4d4dda345758803fe90927beb0722a2cf4719f81806cd6d47e6a963e7b4ab869049ae68cc7b98ed2f1ed42f0418b95c68fad89c339fa41eb6751db1667cd99b0b896fe4d978fc0c51b4e6dbbbde7c19f59c374815b9e117ab0eabe05006f2c3068a926a2527a2ba826bf9fe2ae01d16f8ed2fa59ed28f1e287da4e8b09b69dd23296160df0e1b58ecd3bf31e3747ac2e74017f0b20004328bf31e93e68f10eebe55f049d0ee40bed57ad503235b4bb85cf29253ff7347ffbd711122aff535af0c2094498d63102ba85716b3fca015a1bdbf93b0e67b3a182356296d2f95c88f9724a83828f990b2b1af345fbfdaf30d60fcbf52dc0832881e97a38faad2656e2e795fd3a55126478cfee00930b2df36edf611d95359e168b2cd698ed1f2dc858346f72;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h5fe43a0db32629a44bacb586f0b2b536200dd2591862ba79e8525317392d681d66835a3bbfae696bf324292411be344d513b21eabc667ef1c57657098fbd4609b50b4994bb653a32f56ebdeb97443a9f1b4af421270b59c215c15354a0cefe720b99e2c48176e25afc7d08d8356f95a44e3147f8674ed46282b5dd507071478917591594c3647220d1326580e1ce9190d3044d17947452a533689c8f1b2f162880c0887d927bab6aa6b1d6e3f31ac90f4d0480a82f984196fac9e54202792c05a4450f07b2672f8b6db34034d4f379491247b647b88eac6b8bc578b979b69e668431a4b1c06fb8fc66f89180ef3668119acef12cb96c212700335302edf80ca84f22309b75cd242b80d6942e49ecbbe73264c3c379b6c0d97dace5ac409cb792a83f238573aebb0bfed7bf433622be841d773d00647ee66cbc6c963315110b8473f13792b40327c5198a805b89160f9354f4cda7d669b8b11fea983ee53e9be14f91e57d8ce39bdbfe4a13ad7be9c4d3be1314e3cb8c771247e09ce33ba06234a7b650e50c0939c1f768464c5bfb59ac8ed9d0a23b86240d1bffda0e01dbd5879615d2ee49cf05c7d9d7506b6ddd8402501c5e870bde0681e45325465ba3ec1cae5f64009d8825a5923cbf278d2a1dee595f862fca75b965d8730750684d7a9193c486215ad12206d607bf30cfe66cf4154bebb9fc768cc36414774d1ac3c81209c22ddfd64639ce7d0856f5b5c95b2cc26dd2ad92aa2777c1a8144d2989b9887b4ae73cce1a77d78a498d34441109e27b5d20f38af04523d86e82c204b67499252768e334c7aea0f44d0c14041c0c630282a8153e22a86545ee20f1e216a234c78860abad613bbf20c56b173dc5f89fb31dc8cb06bbb736bb4cd4f00a9e5ff735f8b061309baac282db0a49f0bfc66148d81ab29d698db169851fb1155d666d3be48c8bd81b8dde42a6a59e64aef4bfd9b9f1863657791d5dead836ccf9c4a50181dea2c272b6203f8759ae0018fb809d34e859820dd27e9f02be9db861cf51e123a002dfb805d99eddeb8110f519c5f05afe2e202f76889aabf87e85461ea467a2be829c6105c310788276281561e57b3563cfc49ae3d01b08d70f07d4e31fe1e4e204351d51be80bc6b742ef9d839308502709a53de3a666a3b1a2d29de998c41def5461f2e5692b6271c77d3c3b05110e067f6213e684f0bfb68e628158ae6925ecdeac5d82a4eae3388bb9e89dbf0fa44f6e4bafa19dc078bed75c379b863f81b9787f41fa9cae224a66da28923a7b3938c7ca6b84351ee47b71089fca306671f28f8b681bf1e4c9eead797eb82005acd1d5d59f6cbb85f39e2d8abc91ad406700ffd234fb7096da47eb435ce540b7c57fa6210b867fa3f1a3e89dee2b1689b9921c2e94163a2bf36a4fd92966630fa42729d1bfc9e22ac24c58fdfb932e73df0c9fcbf0a299e1c65140f8326fd0b1c9692cfc388add27f33165c18eb75173d4f632d8cea36a0d2bc2155b4acbe48debc6ed3bafc587d3ca0baf403f34c2713aceeab81db1ce5ee039568731d86639a92a4af2dab07736d56818bcc49d1bf515cc0c836e6a23498b57eef464fe5c5b799f0f3497fc3e2a32d2600755c230dd5e6a01854c9862d41ffc620392cb703d60acd2496d977bb1a0de915267e0a95b57a4da5df2585b6c9d0d4d9da1fd39385406b5699f8a1f4a226aa5a54a8c7587edc4d2b0a91182b02c37249454b2af66c0ec428fb18c6ddae5ed371d3073a1d809dd99ca0f268201d2687152c0c376b90cd77f3ccc2abefdffb635b1ae113b88830feaf8f912b065d733df1d885cb275962fd4e8553232f37e9f5eafa614e7afaba15e6e999b588801f964ec31999121336ca81d5380b3f708353b51e970bad5ac91efc251ab87c349c9bb40fe36df13539755048c1b683e64e9d3fb58e9809532b9e683f5a901e7c735f65a584508d5b5da3e81b8dd8b3138e9b19c9d76b47efe96ae7b77dd815b9fc9cdb93acc1ccd415763d3868385eac30b92ec05b1071cfe001c5697bc439f71b010c7691583d95b48d6b8c0f65e759bf816815447d877ac9cbf781a64e2f247d140c82580b79261d2551c400ffbe3e4b9f9b39986789b78677d20232f1e5c7ebce1b08fe6f8a1ecaf2cffdc60a32331c7f1958f30b30618f8434a567eed056aa2b2bf443ca488c474b6cdada9722d74b13e36ba083fb0042fd2c6dd01375c219b8d8f0a7528c824fce998f8949bce8e2c2d74047ebb19f546b0c3a82ed0a9a1b3dbe94db83c139b5151b766fbe928d3043524e669534179bf54082d0a102c9daa7b264eb3e287baa9059b2d8552f26e991e758511275efc64babfaf9ae64a85f8d76c24c734e7cebb20fe41c6d9d2902cc15e830749d58cb6dc5ca1fa83e6b20d59b2c0cba390c1c45898b6a17fe408f982e8716d4e2b995138fb2faf364463552d74a0a1cb050c07cb74168c0d0a7cca0c77871f376f168196e397d58638219223b343a0705bc9aa77a2c043080169419e7ca874f11449f83d5374dca8c9be220f8470c598d4ffde0892aaeb79704200aab1e89a025372217db55ebb0664be967d3d4844a1dd91111a82ab57b64ae259e1e62dc5e66cd8c7d5d254261b2be4c6f64b48bb1907ff49296dab6dd1b1755c7c0cb76b4288677bb8f46433374c1e2282bdd3a6c4e3f742c593367cd2d964a1328b612f7ca2a4d6771332cd9c10570f55e36d50e159dd81d265ac6f12178c9bf5994e33cea183a229d6e5900a81a3f7c0bd648a6a41330b838e7b95e793f17759b924db91bdd8d63b7365a26bf54f40dd22e82250f3d574aa5261a5792bb0a9b31debf9ba2f7db97107bfa91bb4b5419b09cf52af8628eba6de86e8023fda42ee21cbc4e563c07ac31069f1a84718dc88264d37775f5aaf22996ca16fa8ad20409114dee9ed1144719d523b533e5f8d03f26e31ac0787507d7060ef2c0755b5ba56f97c787e22d4dd7159bd8fedf5c7ceb7a69465a24c04e990c01c780398e582bd2eae3fe12465dc97ac58e5af0781f96f25cb856a824cbdcf120eb63f509cc67ebccee7a3de24c0e556c441ecbe1de3e2ea011777c25dcb7086fa88f362ba74e1ea0f750aac8270930c3c1b67f5654936c54a2c01c0f2d04d824111d93e738b9db63e7b054a5e281d358cd6d33c476398e85f81535f18c44a193c3a7234706b013a252fce74b1306ee1da00f835c2e7f8491f42b59b09592d76f4108b900545d253705ebea451487a9df8b1129eb56915353a6420818cc5133702a1285d40742e8a5e5a74f10b71a1d9431f3d238ce4f8ec6df19927410b1573ca6dce54997f0270334c596e4b59b68a60a65368f41243fab704377ab9c08bfd5f5f2a7c56a031d1f75780560ad43a202fbf8ab3b501a11a45de45ceb5a0ff1d138d48114be58250b59918aec7c22d987f82bbae879a4f729dcb6dbd3b229c551fc5b847d520ab948afbb2b97cf1460aa0ddda76147515a3ef1163654de09ec02ab3fe5fd4bdf80108df024a8810d31e3d0b1fb4bd2ee0146a4d97ba37f37ead24a982973d532d6acdfd4d04a31419f88067b83615d553110642931a212ec303d5a8473e51ba7b72d72809b0a28ebe9ca4f64bf76c2f92f88b34604579c8cf81545aa1a9380c1b1e1bea2d3fba3898002cc96d43e0581598cb528703072793c97aa6c2f4895c05e8128680e7cc91813c22649ee473d125a4d4e31f666d409b8e06e11bdff02ff41e57e3841075971fe0a8d9c408be9497deb063ddae8500e4b3c1812aad940f6f79537a85c0b25dd2d10632011ccc84cf033c73283b61801961db849feb1d963f4917d08395b684f5a4d9b958b98d59ab7106e46788e5e83a06340a2d48d26947cc04af5e158ab0acf6032c48874d69c2dd6b8b917bdec63f42684f6dfb8838fc3ab3cea19d6d3fa289468426fcb87ce8db0bda8e4e17b61feaf9bf496a2d223887d49f6f0d4097337744f80dda1f80df83744cfc48e544033661724aa58e42c28f6524335ddbfeecf7c7d98f02a460cf24bca366371506e28272c69ac5487a00d98692c1b2344e21d3d3de8e30aec07c0d32b6b88a6fe2b560929dce247a50a8bba26d865e47f8620bd48d914eb3012292d93c094a5cb81e9532ef7fbcea8142d7f785d5700390c17f40e61d879f61558aecd012f76ae57ddc6c3fe933633d3dd41b7c06104858d75d1116b2ad1fc6622946c9b0b18cecaba9fd52e37563e7499fcb313ff2b55a62356196196f27caf39dce2fe9688e8843ac5fd4f7caf614fc6ef26fe109a6472ab48ea58f279cc84acb9937eb8e928158fcb1f9f0fab02480d0593ba88754be00d190272c3dd4b8a2e1632cb4f252e98c55155235bf1d9df718495162a053cc5002cf5db15617e014af3715dc07df964c3d8f8b428a2c5a021e8d98d434cc9722d9037fa0ac6c0cc1c28ae942239b757c970c38daf7d1d587428a491d2db0beb69f4723e0744cbafb27059eb73c0c7069dd46b23f3d47d97edf3a12cf30ce1d43d00c58f0d9f0f03640bee862b0383c3bb38c4498b5fc935e1b83076ec625b42409f0f08c35df14239bd7680d03bc00f51fbcfda49f5251229c0d856695276ed25f0b1c13ece02f6e6a5a1277c3d4548637fb7fafb8475654a92599c4fa27f3cc7407e0bccce6caea34ef388e5780c445ffd29c3183074f4c912e553538aa6cc7a9fdd68401e0bb7bb4f73d1b37a74c66d55e24e95e9b3249e8d61a8f768093f68e2ea67101f846612077d5b7cc615d94c3617137ce6d1409ed3659762e405ba43785629eec6e94b88a3ec3e77277c3abf3a7c41d4709da71d7f5ae9d87b0ec033578e864136b5a6f84da52029503ee09f870f853feeaf18d45802d56c64ac81e36376071cd9e32b1b6d12ed421bb12a24512f0244a5acd2e1cb802c513ef3949513220269a0f36fce245e4f6089201f532631eb657f3bf7962befde399ff7ba3ea6743e785df42dcba279541b1b754250313086f97a2d3bbf1702288392f29eff70c942ab18f9027ae9859e8c83e7bbfcc7d0e3ea83d2b79de9fc8f76f33ccdc0d011d26e4c44fd51851bc2c6357d502e4f3356825ff3d4d09b1504a72320dd406d072cf7dbf7e23230245c1fe470a23817375f807fa64fb8849866d9921c9ead4cf359e91d445bc80f577b2ff808e3e33d35697a0d994fc507176327838d2cbc351795ccc3b5f220f9b7e09549c0d385445efc38feaeb717d451802340a06d6bf536cc0174db8d21cd59ea852e71135633164ffe9125bcfeb2d7f64237402a7aab303a2ef711b0242a86bb6c30ed2d06f7d81a7e1c6cb2c86facbb3960589d6de549c06f003422a6008d0e22520469ae6c01775385b12e9c13911cc8fbea0687429062e65e40686abe25facf1420c561ebb5b49bf65802ede38f4a61c0f93eb6f457408e92708b035e1cb561e4c5d9ae2914f3b7ba9b69550eebfeb112148ec50eca0bafff6db893c945;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h827e5b2fcd58a901b2a3582819b4e727d3a0c91e88bbee73505c5e34cbbbbd4c202c30ae82e1b43fd9b9949d4e787df16859f12806e71239d72ee1677655ad15a23c8af727a6a445ee8a027c18c3ed029ff33bf968e743f8059fdf59d303c22ffbd370d990125c7ababff308016081e4b5bf7b7b377f0c2cc47e2bcd7c4a2bc93ce8faf4e39b3d98eb21667947c067f59ac063159b75c617e052605672f32af5586c8561e181f1d560b16a63b79132b2b0aabd5de0c2f79c14fc7c82b14f9316364abb0f2706979c3bc920ce1e10940070af5adf907224690b6285b5ce8becb76f9b39f4d45f3192b79978535d3effc353766d7528118d49e5a6cc18a7cc4334d2f08e623da8f3f2f1cb12397492308f8809c5dfc367dec467f833fd76b37645bee65d7cd7c3c29c91eb2e1a8f56de0e0c05fd92228e0d3908d5e14a652a4078079a307b4f335c0260cc0664efd705fc41b48c88213da18b4e2630d3d29092180133835dcc53dfc206960b353d9f312770f80bb8df37f10a05beb0051f6595e49c52a775b161ef20275587ffb8f98aa2d7ffe1bcc5b5959b5e7a6dfe5e565ec3ded84a38a0cc55237a5cb76d3e3067c8e27a8d3939b91507f19c246327a78e2678dc80b4f1401625a82aa84f15b9308038f293f10c25a224605ffc5132ece9f9ff5135ec2ccde12906b2e423db38093971db906e04509b41d6b72cfdcedd63ee739febab9c7047e191b4806ec1a19b4c1b9a2628e3a7f5e00f28f4eb329a561dcbd9732ce3fa8f7c3e7837d508aab917094c701108544e7ea3d88253150daef6b0646be4fa2c8ecd2a6416e5ae94dfb72d8a03bb8a575ec197fd9e9f48c43ddb05bae5245db01a86f735de745d6798afee0300054f4510d3cba7f53a827dc5eaed3f48c37ebd188826592aacc4998a8dc78ebd00f09a8ce7fcce888d35d923919ab63223c016d6db77cba85a4ba0f04ead09337d0094bb57afe55c1ab48392bf9de60bd3421bc5591c57bb5c8da1e9b5013d71edf14a832d6f2f7e28dea83518e0570d4cf7aa119af38b7bb4ebbdb5e921679efe7e63c4d6679d7aad8c403c50e9f4dc5c7d48b96c47d1a476449950f2e5268018d26e94df381a54d6bd7bca9ba7e67bfb52d0c7d3574d40d28631cee5ffbc513700a2e04d1b7b0aef44fb5041a041113e53d85179ec3bb72ea037d25b9c34cf6ea28735e7f048c92f14b4a77f28578a0f7b0a1a1793cf60a804a40259ff62469fbb5b08b6a5a2a884f7981773c086944cb6c8661aac5d0cc1033c3e51a3b765c90b4c21ccbb8ed3fdc4b049c0d1a5c9b650c4f5e8908bbb8d53a73286572fdb7e26a3de35651ca114de2b8324d3adaf3343598a69782c278b4c2f54bad30bd980d01fc2f8c5d49216748bd4057f5c512646bf4a39bb613d57710164885ebf10df12aa2c5c70623167912ff7a73036ebf5a2a0215205f8437d67dd2c6913be366b97c87a130fffc48db08a83bd4ed323700f6c3f96d7434c6123f423b309f016f6369bfb94f0d96bdb8ca18c4909d8826b3352c3d324f17585a511fa81c3e9f5ff6d0aad9f9bc524b7f73d9b495b59754935e0da5df4e21b8992501a23945d236de17bef0aeb2824258f4a89ab068d0b59ab0d60845253272dca1c863fcdd41c789f1f27b3ba0230516dfbea883e7e354f40c361e07980b780626cd171e172ac385bbebd4385a6675fd7fb0daf33617e09852d578efcd22f64afffd80463b19508534febb04841af63d95cdac5cadc60fd16ecdccf0ea3a5bec1f295b43419cc0799d75322e26ad3ba788c73bd6b06b2c40f71cd2042fa35a0cc46fb717f2d68a6b61ef778e3cb5b8980d75e5729573949bf81dc5373c4bd619624d25b54310bce71d294e1abead8fde9daf87350916afe35c6009987dc77df5f2372e202066bff97afcfdab09c3975b5eca19bec760d8420029fd9d034b53b0a0bfcaf78ba10721d21ee843cb4819c894a2a050d469136cd33cda9b4c9b05452f1ff7bec25a4d69d4b26a040b8bfa639e6021cb6a449377460051b39c8d2f5370fa1c0b9d6dfa09bd9eefa9b6b74150d4e7e9137e8ec4bf7e792c38698d9cee6b305c41b0a68e1a2429b60467a888980794e5e7c9bd6b90f7eddcf7ec3303f2494269954f912c4d4c88ac4ec57be445b24899e9f9343f729ea37536b174a206d0a9939abd6e65e2b0a5f0da5f9d7a735d52768d3ebc33b383dcd77085989949ad5b43ace873260e6c65f7283eda74514cb926cb30e2d0f9544509cda6ef269422cc85db3a49b86661d31ff064b9b79ab8879fad3d6533d23adb6d8e52353f5de278a4a04e7f3b9aa71bf5538370ce9999211cc01530c0d8807a6f1848c80151c385eac9100aa66b79814cdf5c79aa0214d7be4e72c11276ab096f3933fc89325f4ef1cb52ef5bd6c5385b9d2e312f5c280a790e09d6c3dd525fae548466f30ee54de67530a3100fc00cec54fded9548be2210afe8e587f24dd67ba077dc0abeb5430e6bcb2f2dd8262bbd13992452c348bdc61acadc7f3f42d00d5b76a8e944e0763e430e8e13fa7517882a9571ea30b9b057cb424a8e2d1ecad7b03882ed2a5261ce77cf66d78557dd875f9b7f7476936a26b06f42e8a633bb31c3457ead486852ae86edd8d2aeb74529a39bd1c138f49820cd1c0013e611ceac9759475200712485d6c40421ee8a9768342263b9e708b1c954b0cc133c96b08af6ee39ea97030ccfa21eb1f289267c77addcf871c398b04973c8fe51d973cf62fb993d38ea536260d5004b05768a1c05bec41af3934ab6f49bf71aa59234f6e3cc1676a4777ca98ef6b99a5a14abb0cf671c6665941cb2dc9f1364037b43243b8d46a0284ac10e9bdebce84f8cdc8984546c86e10f9d6341c28c7e43668c0aea7b947bdb254b37bdd29a64828743658bca9ebad35e7df804a05fb994e417088578de7d5eb74583b0628392969a0bc6619a87ab0f4fbd6da3683611cc08558f36f2627597b0dc0f92c1ae08e3d29a2414a0ac6f4a9ed92b8842e24947ea2ff9e992d29005b250bb185fe0b386a4b4cbe2aef1cef5db17945996a0245271c7695e00ab916bb298bc1a5e9746b5bdbdf1343c13c2529bdcad551219b3ac8d4dbdaa4e79cf6c7e10915cb7d5becdc513a06566303708d29e6d3a94e726d5ed4c212f152c6fd108ff56962c1b32e864226a95999fefa544537fe0e1f3ae62ce00571f05d55ca57a5b8b89967b1eb2fbbfa8557ee36556a2c3f1582693fc075a136c8c1c54ec144b2488bcec026f74f63d38db7095f929b8a2e3f85e3238d95182224552aa4db4b128e82ad56520594b47d0397d3697b05f37b99925501f5b86d65f74a14742dbef30c9474dcfd7114de757457b60440bee3fd4b870b111e4518a1f2b8b533b71198627482d26a9a99d6029e292fa07babd86862f3601705138f703d1b8166a5e0935d0d2b2a796050512b9f0989367c3f172fe34f9b174c579ee2f9b2c3e4ff66f59152f177c4eee21fbe7a00fae8aae0a39e883a09ae3c9e6f04afffd2973f1ea58c5a44650ef8c6e6b8f749e4fc90a4314cfb46109e82c24f5e938ac236c7e6905768260e2e28a942681fbcbb145f577d68fe5a2da303a73cff30fcd1ee75d9cfe7bb3c14721b7cccaef368d806ff5385002d0b2730fdd08d9f18446db3016b8969d12be48e1d26dbf0382d83eb76d8137bd47e3ec7f956f0d26a154e7ae163d3fbda8ab643870d1386477e05df05154911522ca49e4bcbc4cdc0c9a1e9e11fcc705db1f4f0935e3a80bac7ed96278e05ce93427a92f095925774575d5e95412ee0dacefe9f7160edbfb0ec2ba35921e4e542e1232d15a7a7454d92392c621f8cf9d59c54485eee09614e34f197978a3a9e706bf49ee81e9e02c07f840e3d76182e815d61fbf865f0e4d89ff5fb306c64ebc4644c4edd82f930d6c7ab1d341df8ab71ae5564304ecaaba3de9ef2d778fec9d97efa5b90c26e37e96460336479426203f70b4a1cddae4c96dcf8dff6f182dd5716f78556dd8a93fd390018a954a263a73a86b35d3b6de876d7edd9f63068b80b2c4a7debb5b1b5b7d417b3e9a3caa1c7ea2078aed9cd75737a9ce057a793a56851877f57e97005d6cc7477ea1ace767ed9794185a4d24b94d8f075fcd37c53c1c7abf54079d6ddf6cd2576f0a4eef0b0e6b354d0ae1ce398156f84a3091a517f3f263ee0917b17a65052dc5728b95e8e5b193e242b3b5a93af3d144d2871062ed670cdc077be1b1564e93a9b974502639706a5418773e7e0bd96ad11d35b5594e6738e434db9f10d73e1467aa66650869434f4ef9a8e03502c3a11932d3c0ee9a8902e1ad27835c9151bcf3eeaf2a98b8b72d45f309085fdd2a369aa82035f65ba1d35607e1fd717f945b227a3ac39b02b45ff2dcf9e124be2a256b0279c6ed4e6c7cb2eeaa9b5d5946931813a8e6af7f44d51fec6f18017ec19b5ada7c9f4dcedfd3e0962d69578f21db2d5dd3511f28630eca054d5fb7831ac9157ed8fedb3822ea91d588cf6d94c8e96b1c933e3901efc1cdefb6f457c7193f87f61b9ffa5ca178f48822a6bb4256ab4807a15e2aff407505fe9b40f587702af0ec6d8c829a6f65b16346d1b2b1404fe2fa7ce6227c684c998623628c887d4443fa2ff93b422e53c3fecb661124105a5b3a088b25aef14c596cf30719226a3400aede7735864c10839593f25f691ec622b73afba8e5ec46c5eaed28cd05125a0eda56b6cc49a1386f5ba39eac1ccf86096e910b354a5c7567fb61bde2f01049c2a82240ba993840e26cbea7c571e538a6832b1f16013bcb59244fdaeed57d46840238ec7425382defc1d958be27b18327a14ecd4c513bad17561b9396bde01912ea9902677b950e94dec3fd58ce9f95bbf5ef48c3c1b2c2fbde8d30cfe1986ea626d56c473619855d8b79271dbc3d837a921dbae7a65823fd48382088517e940ee2bbf8128ef7339ea0cc05f9356deb14dcf0f6de12ac8d26199c977ea6a69f24f96a659b50ce1e8f0deb4f7a8b9cf2acd96495e9604a0819f5d92b927b9c4c043dd7cc776a302e6a0b8fe649bda2003325b5bcc3e9cb11cf91ab73f6538db546f77c4b151601fc59c3f3de4f5e7e3b02bc6bf67c7eccaca9314211a47a5b6c3a797e13118c8290418cc79b2fa7cf9eb4906a5e4d70aa7d959ff15ffd2cb648b14786caf8139c281c5ddd50f28ef209bcdb4800d815e464cede85c37b413620aea45dacf2ea98eaf9f2b9d5580a2c80339d5b3f553e63ba65f40bdfce8d54eeabc2e5e43cb8aa2206e2209a71fa44049c3a54f44e34e0edaa6d74684bb1bde63ac1cc17835da16e6a3dffce3f7fe8d44f8cf0dd55368e44c5ba2c04e23d25e42540700782cb56f68a2a833c1e361da85121ed5e9a95e86107d39a51740c9b408dacbea9bf0bed60f72156ddd3c06dc0bc4814f0cc1aab35f0b621753fc81817061191ef72361a7ab9acd7e7251233435e618167d162e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h278783df7d702578f15122f0e1f6079ca45cdfff5e5168d9495db19f7f9121c21f30218537aeac4810d1e58467c5aa56f59668601b5316d5f753a2c37c0ef9ccd7152ac48773938e6cb489398781d6fd13b7cd3f90da77c36b91c8301df7cc63c11f8bcf9d667a31cd7e2d303d76719faf8a6da742c9cff3cff7b41d944ffe070c416ec9a1da3556b3d4b501ae34a7490c13d2d00ece6a181389b9fa2da63ab39a04240883f6c2964888b907d0efb750d7febc90686e730db98656513c018448d8af158346fc5d3fe58ce2bdf5d9a1562ac6b882566a4749753847d66ce4942f9c33cb19d54f4ac3ffda411b2f98eec3ac0fd3530facd19c8875f5321312ca56883b75e25e55e14d3cbddc47f4cce94de0f28b63ddb9bd13c4be197047911e1a3a8dd5a0e0367fbd7d5693210e49cbc0e8ca52f3589f67eae392e85db1ea9ce1a7a11cd8b2ebfae37a63256a89a75bf594556855a00385e543778f9cda9c3fa82bc0aa93614364396b0192c3911b4f127280f2ec4e06e6b6e93854ae0953f8a2231d236a0d7c12e7d5386818e0729297ad25620dcbedbb69186b0c873e83a2a71af3cb56d8373b9b4cfab5d6db501616234e11143e08310555a50ba14020d066ef92a83268cf486c52ca58bc58e7a2136825dd959a87c0d61db0538a049eb153977123130cf1167523c7bd1aa5df21a6b8d6585bfffdcac2afa56718a215cd444af533fcac20db6d1fa3f20eac0735b77e265e51f086a8b3a6048c936e83b92647e71bb481e64a0f42b43e1f85d8ec109e3427aea439751186a903885970f2896580b77766126718d8b709987ed111e85071a2159a54b743502f12a37ce4c166853c3dc390a2a29eebecd22ca9d89f2aa73fd17ced8feb79b62c224992bd57b967ac52b6f49c054eec7e3733173eeb4b180128b0de5365442032360793100c81208b0c3edd55ca42376e83b3fc97e198c2e8a17e415c8055862fde8f9202c83e80b5b2868e84730216d35b1603dba6fcd5d1aee24d863cb1732decd83b0ae7da4d63c29f8dcf7fa065f09eedef0cd38fe57093b9d159598bdf962eb07a109b2682e9e677032a2560ce1583a864157dacb4f5f75fd577a19fd12039f108574a5bfabe865511b2a5ee1dc5ca68c9edd20b094bf783cafadd536e19f043603338f9081c11296df1a0e2378d4dcb9a1e4be276cc7b3751134d9760d6d7b6b06e5d5c5e69c24443c56cf5230e21814ba7e00f5af03ad1305693d2a8ffa01c1a16a79b37e5f5b0423b1ad9e30f64471b379540fd233d980c8a1ea076e77a55031bcd5035f8c41fd76be6b220fc9693e5de911086f11e4ddddeee248afa6603f6227b5fc49d2427d49204f6ef3228add74cee6278badb975c30622649699a34110ee98c82c6e99838b250c074d0183f7e315782bebd7ee8b6a4408e96e3cea8ee04ee875693fd4b38278031b5d03b53ff11b9e0b6845f1cafeadfb31e0fb7b5ed160c5c06b1a34e2b179da2446ac3d9e061aa6cc0d30d2e9f1e4e25aa33a7bbd7b23ef796d1757227ae31cdb8d69d55799d7b9463d4248721eccc315f8013e8e2a22e2d0ca6fd4ccf4ca8d6e16ee87bb3e94e4e3108746318178e9f2cd1876d26d65f4c9132d18eea7f5106699d423e6ffe2cb9a5692e3e229f9d9f420871ad5af49e0dd46973b2297adae50a2825440dab3cfa658be87a26949463f0089723a0e204b1bcbeb17b171c9bbb930dad0ba536f3749d7db9172d761966c475b95fd51c193283ac1fd1b895f249489ef1810040ac4a1e789766608cc4df8efb1e4f7b3e5ffb348f95812f5273c09827ad1cba9794edafb09e2b97c7ebbf7bc1b0544dbcbf16a8bef18ef69be34455ad191639a9471e9f88a7d7839546261a7742f45477e893305c895653438099ce9fe43b47a1136a2d19f8dae6f70035c386883c15079600f2169bd6428b9e36d0eaf051464fe4592aef2e9d43e180ed7d28535acd037eb1a7b1713794c8609c391f336a9cd146e5d910ad85227aa61c614af0a0184c8afb85e70a81ea3cc6aca6d4ebde6ae8d49b07783edcacb3886ad7a10912a10f3c49c053df3994db3d4a4f4f029655db3e193ff6acfaeddcf01d5457ac72a5e5b1a52c100cf197fb9fe8da2858add296c16e2ae51715cfcd79788c2e3c44b0936d237730277d3a4b7cde6666571ba7c150a324fc087b60a151550a31eaa1243ba73c0ce62b86cbaec17e504b893ff9aaee237ffb6e872f45f1139983896bebda7903154b933187b598bf2761032aca51c47b2a8f06880ae48545f7fdbab071bbdd02c18b225cfae383ef6ea9863cb80a6b633cb0866f8aed824ff983773b34ec5a91b2228f1e080964e6eea1dee4a5f74043bbb1c8fa8c40a832b5721db4754df01b431f0be3c154bcb65f7ff2af9c7adeee24022b859bc8551968e4a5cdffd501e4fffa3754c77a67521c63498e59f8ec2faad037639bf2a11abce2faa5dc91653e3f345a6d8c2bb9d0a70fd1ac563fdceeadd97c74e042ac38c4ea85f08ee4539d732728b1a531567d906a6440ade5feb4f3614638c2a67f613e02f9f29d6994399243cee5294c84d338100332fbbcce9e2f09db4f01e0aa34ae24b82940b235aec9898b16920fda17bdb44210cca63f5748a2fe653a8a3c9a27281133e1df9f0f9ad8d5214560230b8dcb3df4b6ec213edd620eb8b4deb079eae88a0fa5ae8b3250b8a3df205a5c607944a6b6683f038a7e141bfcfc406074dbe753f8bed6fb2c0e1bbf48d614cf710ff9227f4aa559d397223b10e475c7b166dcef63057c88b1ea0939d51e0a6e6dfe8fa9b93c979cfb94c4502fd6c9d4dbad6c62a8b806b2229445999e1b38dcf1dd302a04835de9facf60f6d8e644b6edd0523384188453d59684be5c10a3e6bd4dff5e63d7c70e6ee6900b63a21d2fea6053576684c419874529cf21800e774680782bed16b2888592aa6060fabe65335b7c2b0a69c86ac62f78f901e2066aa039c9088987df7e1b892028201020456315ac006f390baa0ba2113cee3a9d0908bcc07545ea91fda30e719049519e88e201afe985d1f16a5d283cbc6569b9958b8409a9049313cbcd1bf36d88707a4640072c82a82fb1bfaa5b971f4da2f3599f7a5c6c6690b5533ef2582d9b5bd410519cfeca181d84957df4b8c660a9f7084182ec0e6590c82c88b8964051cbde6610967c778e9c32614a2739e9d34e53c0fd24c74fb7d045eef04acc151685d5b635def302adf78a45e62666c315ba26e608ca47d2c2cadf2565e86a5f91b38812b40423b3b74beb51a3b2752d4e51e03cd121e29a5aff77d99cf3d41b683c8775550e23246990f18d2158894d24049b70e0cd47188d05e987383544ac34e9ba5120df12e00b12519045818409bc95a2c71041ac7c41a90b5fed325e9b5f576ad5f7185afaad3cbbfe224c93824be3132cecae9bb59ebb01632097aa4de467a8e9b37e3ba638db0f0b26ca40d089e0fc10664b73c03d5160614987b6dd1a9e745a82c5d73aa3ccb233cb7dc69e1873b438a1f1ee05e0d6a039d5443b55d76a0c5b42daf5fd28548723fc5a0e1bb588fc30f966a28e8f7a7aeb3adbffdeeec0272c027ba43c27c3506a26cf78b7896e33ef71e03635eb668ac898f635d0358bb8610c317c6266a9882cfc2b3cb910c72ffc48818abad5d668b38e7329ba042bbcc15f835e6a23c00d9ef9a614ef3e9084c65bb4a7c55f6f54fcddd19408e49a25ea64bf75706eeb07623bd53819bfa0588d0ad7e071402ec97f5a2cf9cb8dbf02bdec307537df09ee554cb9c55e075473d9a641ff08ae77efe616f458b5697275862624f5e642dbc66921475a2f35139a789a2319c12db2ac3bea99d8589d9973ed30c97237d9295302922af232d71600d9a1139adc576db207331535cde70b4e70089e12476541ebcaddfe13fad4cc86a2c4bec77944b058ec86670cbce2e188e4e8976c847d64202d091dbc064da79633f6c03c6a216b850a98513609e01def4b32a84eb552b93fecaf5b64bd690367b1b527f3e6243be24b9afaf6f497f490e04d3f5a8f108bc5603baa6399e7b84473327d0bdf0f203c18661434126b8e7b70e1792326bc2d18fbe8af4e7086f84115462ca4e97f07cb00e167cbacffaf0d3f40eb28e7af41676270045f019134fb0721381464ebc07ba3b7f2329e450865c4fd7f026c7f742a1992b992a7ba856690a59c9d8c37d15458ea5108ce9d16a3af84ca096bdb4abf601da6a73d73e4e2ef712718c65dc876fbefd45e4251eca038cbb512859e5f47f788139fbd1c151beeae7fcf64cba709cb8353b74008932d69647b5b65f6cbef400ba8b4e908fa7d8c210aa7d75e618c1448194f89155624b567d3124fa6c850400866c13505e99845cd2ab8ae9b5539d62697c1db2740a461b43cd2e41c96e44ba5566cce40749d25173d862b333990ee7357840a3f9e94458a15df07a7e99743cfc6e020f6ea2c795ebd1a7e2aa2125e74650d97920222de24e3ffbc67991bcd5c1da955698296ab8ba65bc90f153d29a860c7ea7f1398de6ef32c5f5630c587fc15fb3e5eb339e017eb0a887ef2646e14807d7708b67d80eec9bb7aa1c72c7ebfb2dc705ddce3a935f51a54c418ad21ed41308e12ada773dda93b4ab360d69021a214ce98fe8ad35597e1796205ca35e1ab0044dc857f92cd37a151bc402739f7cfebb6689e52019a9595ac14082792a73e88e4c58462522b8bdf18a7813622337dbd28709fe3372cb335eb07da572414804d4c6d8cfbdb1a92d9a63e7a74c5957b16cc2a500e7a9b4e67c074f1800f158f25bf27323bb6d737a04fbbae0f2ab070547a5e34bbe7fd2a563e9ad244f3f64ebb13f34857cfc65ee589fe8e9f08482fababd4e39ca3d4cc95fd34376a8958adbe7c874558bf3fe68075a0880d01dac988f4fbd26aa6823d4dc52524ee9614b5cc29ccd305280d0224ba4be027b05ce9408cc1f4450f8487aa2532ba6621434d3081427e64481d1a86b391f85575a4d0527f79a8d4996ac84e5b53dc8ccd59e139bfb6015b116783ef9b787076e13eea2bfbe989456cd12cc653315fe2e5c8fce28fb276f712d35ba848f1a6796c9c72cc21b9b24cca2b6e52f15dd1ac3e40c7539788967b5394c9c2643b44c43719ab37a1e32154863da69d8adc919bea50864907a619d163b378cbdb35a237be0e2735d02f5a1abc22686edf10736cd490d320737bb48abcb01ec342c617cf3e83026d38b38c3ef25a3dbd081538bb983ffbbd80df71fe0937cfdcdff78b7008b56510bf36c7e66c3e6eca20da12dbc085d6127229f4122a3f743dbd6bd02593cd784258512425601e0dd8daa181822262f100321ead44f4cd138931733e61e4fc0d5df708992e6af9ac19b0a0f8c4b363d7346445ada43642b667dbb86a5419702ee02550c0baaecb959ff4d3b86d9faf331dae6cfa2d3af0f807d68f32d04551730fbf205cf01a6a1600bca4207bf1c8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hc164e6047da47b0fcef2487ae38d3c1a49f8da37682edf2a38650e5cab976c3fd6f201980644029eed15cd2a10747ac984a0068afc3f5be149c8e342f72f1615f16fc1b1c2617ca4ca8cc4a23a673e2e8e43b4915116938b372dcabaa814663fd88efeedf33611b688a1e0115589916c975d74734ce4a690ec280094314a0dbecaee901acbad8d43a3bafa91809a8f71066e45dfa654414db10d5db3c145327f46620738e3db6d9c0b22075ec59c8945aed185d4bdba79d3dd4bdd5907cd192e633d19ba04ee6e29da24e453c3607e926c719283112b1777e4cedad82df3b59c95cdb2d8a0dc4be807ca90f3db5fe0b9bdfcc830259ed294f275cdf83eadcb2ba198b62f4a9a6a88ea8dbecb75aa863beae81c8fb08cfe1ae95e9d0e0cf98b6dd7b615809082817661558ece03989402b6809d616b90de7f0b93cde23882e021e7f3a658b99ffc266da4d841c66b6bcbedb17f54e60bed11ed62761fbdd88524640f2be985a77e6057ae2b77e05b14e086c76d7f783b6151daddd337147f13216aa0aef3ef5a48eef254f8c54d70ee9c7d845d47e71fc328d73e048e50fd2abeec78e33cdbbbd37d5137e9e9e535792669907c29325026fe88db8d57fe7110fc86974003f5992e3c8ee84fba38307b5c1f0404ed31f3ce3a1e0b0cbefb1b60a73ddd22df8ebd61bca993de4e68e8b8a56cbabff02fac39002188551591baed70cb2e665bb9142524174f00b487173a287fa31ec0e199869d8ce14723e2f2fdd0fa2737187c195662d7feb6c397b7516888beddbd5712ef4a78d0d5a350a0e1b053ef5ace004ebd9663a5552cc76cdbac4eab0351400f9f5bc777c795154add339c74c5be8ebb502815ae4f5f758139b00a6509b3c4aa91ddedaed495fea5359c2ec56073a3d7e28d5a1966cb262eb9d5b6b86e07ab481cf237786ca9c6cb72a8b823e1caa7179d311121ad78bf35ad0defdf189bd1581d1ccbbe10f89a4c18b4f1b34207067b5ebb1ef914aada69b9295f10a672fe312e8082a32bd4ef1f546071a697901971cb0b2f0bd1899cc364748594f00c1274a2d65d50d7878c8643124034da4dc6f54538fb509c1b12d168160def18c9b8ea01e416652e4468706daac6307bf3728f1799e8d6479b629c36c314b4cdd0dadece355295e3710fbafcf2f3f04e13c93b43f85aadcaa3e8cf54dc7daf66f773af1d99f54dae65da2fdfb8490f4ca5fb1eb0e669af0620b231b45e6d944b11e5a8452b4f09e4b7defb1475d23c5668527dcab75110e8ce26da35a1f92d4f2c09eda0a6936300a2c2d4d8c66fc403e4c51e8645063205bf0003352994f391701f05e05b0d3af09ef7bf66ad7611b69cb37d969b26cf3ec8741d951fb984de376d0129d33941a79c85aaff6466f11618e2704a4b5a853f0f6ebf842e943842e39d62c68032f62cc3b9f4d068e634cbe7141dcbceb7b1595784c1a9a69a3d9ed2e389357587510e88a437670fb4cea8f0b94b8d45d9d92fdfd30020568de34fa773527f3da4c12b9ea00985f34e075903e758cda577c99ae7062b4b164b0d1eaa564906217888088b85c0f43d58f5f0461beb5275887e53a9e21ca8417bcebcc445473a62ea6164eb4e2565ff45cc26896562eab25e1f69f5ceb0cba5f461f25b88fc8db6ce02b95cc62f41b43413691ad96179bba779dee9ec5eb2c610cd64252b8308b2d6a2617f4353ec11d26ff8c5e6c75563acd4dfdd17ab918d8b2700319cc36a9623cdd10f8fb96dbc387165cc11ecebd70f8b0fff0cd5de9f382d2e0ef761c48fe88594a1616249e8e89254b59e70d579fa05de7881530f39f31b29e8f1fbd3e59754e0e13dd007424fda9a70529670d9e728b5f6a18a28fe72fba26a2af2298bf9b6a44d98a35653e3a7b3d4ab7d7e4c8f98d74bfffe16ba7ffbe029fbc992ceb097f15a3fcb7bd736d589014dd37f1fc9d867056ea8770e552bebe999daea7148b1df90892731108ee20c28ba090e17ca1402703637265622e844f70b548571f5cc05665e33dec142e7942187e93b2c606a7491cf9e70417d71dbbe28a53c68ecb3947ee90e8d08e85a02745fa9956e9d07a981ee3c500ead00edd31a90d3d55daf36ffb2e0d78673e846fe92843a477fbd96288298c9d25e2c6f381237ba89484a16dc91837e6a26504b29bd1c9027d2561fe5c8467f74b252bf57b7676662f9b575a892ecb5b140eecb5f9b8ee9c58de8056b9eade643db0137d4d9614f994bb040960ea793d5a37b1c76c7949494a7d8193fecc2ea5d2576770c049dd1ca7150c64906e8953eed7f1afcc27c66c87fc03df0f4006df0c386c26fe1a429ff640da8034ee93c6cb60b4395e1ffde8fe656906218a40e2fc335084ff8579cc62ae19a6a97bdc523a928de9e4a3755b98757de73513f4f4c996fe91c6de564bd642def7b9f33f27c5b4d5d1e0a1935d6a68e50a93042eae0a75bb31ce2af8bebd82f1f331a0261ee33783057e0c4158c9916f8419ec7661a1d22de5a853f4b88ac969e70ec418f0761dcb90e5aef2deb9ecf0297e0e66c93b72613dcb82ebc7e97c494cc610d11642682826e9fc80b989458f59ac4f04fcec3818ad74baa4ca16ef5e22e779e9df4d677d0e499a062cbc16c24960f187be0a870d7f59be76e79ad99f54ba1f4b0ad6b580759de760ad304f831eaadca6e36a6e5b56ec833a65c68848f0ceed7fdff99396d4727b21becbe820811c260c3c6fd4c4f23a00460c0314afda4c7ab6c0510d535616508e1d5a9b10cb702851d3a8d79abab184780645404be324c12aeba7eefbc33c69afd13e85f223fcf3f1166111aa5eb759ede4efb52fe70d1abf15e6de87317c8a318bd0517cfa298599c4b9e8a8482c66f236ae20a028028b8032c8fa2618b4ed1204e08a205bdfcc1c4141167ddef32a8677191f71c1da8d0e538955676b126894a8d0d7e4fcf1c7e86e38ff7523a4183f2e4ea9e1da192862bf1520a384699dd42b579559d80a21515fb91f3b20a2c124d62e3a0d0af30f769654f9a2b67f25920ffabe23d6e493b53290d80289d17269aeaf0ea235732137404c086274f0e226c86d9a8d225eaff325fe12777df8ccd16473a875f36b7b13bd0fabc848fd854fb6b2e5b097dbe3e130e8035e8ec76665cbdc10d634c6d1f7fcfce451b5c4510671ea025fb2d5d9b37fad91568478c2fe4b41953e01ffe2655545dd35fdf7d2668bbec44e223b0046bb506a065032350d0a4ade9db6babdf3471b2b3129452dae92d46632652e47e542ddfe215a356764d7e79fda57c29f8e2447ad419c7cc8ad41d742fa1ef88a8dd005d72f6f855f9e33697e052b9350852942608888bedc1885c56fe85104511448f1ec70abefdfbed6aa1ca3058ac5bef5a38dc3b94045bae30b9b8da0f566928d33568a8aaea13df387d0c1331877a7061fc505296eb8fcfa13da6293d23ca41f132845dff7061609a3a6843a1d32c646800defcef49409c8fda0768a738dbd29c802f901058504a030c8950f4c403af1578c6b53354e13c8f649938b293765ea91176eda7a211858bfe96d3f6ecc9d3ba7399b1e15ee04552306e75813fad75b9dd0b5aaede7ad1769ff35ca5f325463e47e103ad81fa58c8fd83f61773fb66f3ef36220af4cdf47f8ce11b8236e868a50f0e04efa0660edb6b3c413cd8f7585fdc36fb8b842a7bb7750024ee7cbcf84103031db855c82130effed3faeae06c344838302b8ff886a2aaba1ea0892177b6403731f59b5a11a919d7fb6d9f8752d0b5a0ae1649c93591bae6babb4a178f44f53800b8dd075c934a42c0560d930bd3a42ce294c3985d3d43babf51ac7acc45569e1de53d39492a2856e0bd9cd8df572cba392f2ae004271e47807556249988a6e8cd7361522e17476b58d36523dccedf7e9b822a4161e4e934a48591fdcf860d2caad821d20bf54b1042304c45e80af0d90f2e34c99a1b90971b65cd6267deddddef842a959db965665410e3a925ac69a4c47df414704106eae5b67f818160e59baceccf45f7c636581869d540752d51ab9e64fc3993564513bf4beba53e04b853932b25b015fa66789876221fef3506816de0fb2f4e23d2e00b50644c717ca5525cdac5eafc4fcd3e2f4bda6028f4edeac9c73ec869c45c1fe91c5e50e552ba9a9dafe3f8e31479e1e5a734810921cbad2e1ceeb1459069237d7f2341e15a6feeb188377ed485a44454d6777a124213e1a69ce9934032a4b3b17ba6d81c20b9b0883418522381043dddeca5f158b69d4eb095aa5ffd9f8ad3127a0db024834dc78afc05f8f116e76cbee76d0bb0621c8d6a7a2a200b2f8295ed8730759466491995f8239cea9cbb45da965fd0e2ecd2c7c609e7c942aea30b4a1cbe4a6bbdca19f67e9657fdf55be84c47ab3bcb9dcc2cde0dd06a0f261ae1e6216f57160993d4ac830179e6a1a36ea7fe7f8cfa375f398dc791aeca5bde1b1502461627d184bec9fc02f6b3cd354516a4d03621bf9a10ffc113b40b32bad5bafb34d55139cbcd63089ab2bbcc2c280ad7b861356f11d52db95b24079f89789a10f1c103628e5605a6b63480a545edb57226a6acc4e9a3f25117f8ea3939563ece3263ca95cc46289e0b421a69e415b164898bae9e9e6cf89c14ebd67a7d1f1fe619a53f0397ee3793828f2d641a23a6a044718114fb89937c75be7f74f57f2373d6af869552bdbad65cdbe2344a06ceae35bba1189b442627151e10427cd4c2daf948c94931fe1119a1af2e603f4f34cec5ba793a1a16e7e641ee4a2287f247a397ebe3f229fc1097d961f3b56b9049a326d7da263e8bad97b6162d2434116468d98e982cee5df3ee8f2cef3b34104de21070b7a29176421ad824c8fcc13ca4d0485d8e6b918282bb6d4dfcb6e5dc249c75252dd7292d2f6098798d9bc5df36c35bd100a6805ffc177ee0fd57c17a8d877b9a1d3a05f066cd370170aefc0a4fd8c41f607cef0b7fb0974027a55c76855cd45b4cf37f1e25c056ce92b7b1a0a4da512c1f692746bc1551d2905e34fd53f4d0c4146156fb74fd889a460384e2709947ce6aa5177917712b11d92ed7ef198b7f263760812c0df77d3e5fb673e081ac9a4ebc5e329eabead4775380eafacca4c60dd6e914fa879e6f2faaca33fc8cb8185145a86991754eeea6397adbb43cadd3bcfff0454a631add62b42c281858583e1a455197ff1a25f67225fa82272ea6a217d71ab564e275e30ec9e96668f7bad822975b36be3b755ce3f82475c5a62235534186dc447ede8f4adaeb37511d4f473677a3741d44a585e25e17de5a920b04acb1212c276efa215101486ad8695be13e05ad8ebec95a55bed4e724756dfa2a061e24aaa3d94cb9a9176c883d0d271ec88d2e28af4a908a32c32e752bcafe0f228ce2a330c5b9f2779e699614db28fc8949e142a77719910c50e6cf11a7d815064646cf648ae41e683893654eb36e2e04ee137b51ac47b270d68999472eba3b196f0d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h5ec8bd86666cba1f090948c4c91dff02092d2e567e4bc83c2e4a08c62e2d1f6e96d30fcc45d4bbd34a5659d05937ec287047e5717115e29cb941bf3feb05d974bccc3b2241a561e0ebf51118853f338e891e7203c15140cfe21bd937e50977b5f1105e35b6290f361502c960e16bc362d6cbdee03475f783bba5e9ac0d9a6d7038acfca079bb4837f6ffee527b834c3b631242119a3858b499ef1ae2933b6e2a9fa73ef9ef7aae977ac3d77f7e0e71fbc9bfd84ce6642c7bf1eb5adcdf3029022baaa09852e7bd97e08545c907b3e23942b76991b939169e44316d2e28ad11408d9c9ba60f8910caf0431722db5072b04cba01f0f663412793c9ef103c0772696c14024929687c7d65e10f7955489ffde274348005d869f0c42503dfbb906dcb2f49651af626dc5d54547b1973fbc6271241410b60966cf2b4578abc96df7d228f41bd0a8744eb291c653b5f23f8560889bcbabbbfc3c3e2e1e2f7d717a2529cad7cc0e0f89f44fdffb91c13fd4473ef36b462468d6f4643fb6024f25fe0fa2882093d29ecec9c75432528559efbae5e762dda352cb0bccee9d4b5c8162744c10a155308bb0c8247cb7a8fd052711f8eec8f6aa6fcf086896f0cf36648badab89f7d71894d9dbc2043b6a2453622589245c2e5330b2443c5bc23eac93cb894669c450d087fb17c2c52ba7831a003bbd60597933a728e716b8386cef37316b601ebafee1e5c4a781daaf216bd012f921699ae2b1730fcbd19e03e7a3afae15922a2c2686cd32bbe3e411ce61c355ea6c5b6dc39e17bb7af223763b57baf15c8a4f6fa5e3265667dd8d1cea036f5df8750dce4fe687f1de8214957560481e3e167bc48f46264a9ce537c46c70efe6bc63245c78da3a5d8f53864fa7404db4e5a6e0af34dcbc2695ed246c5b9a573fa283cf8eccf0197a91ff7ef7ea99b6469f67072dd77fa40e26994301b4f82ea9dadf62338a0f091f2a6455b2705cd59b697ee873b18d0d69f3e66e411c6eedfde98d877410e2d21993579e86ddf57762491518057019ceb01df848afa0d76d61eab326b3c5ad761b89098dd776d42eebf55429761e794fb459f7229159645b2716ac3f6f3d2dfcc15792af52589ea430bdd9b5aabd5ad9484a197c10adcc4f9ebbb17c800c6314cdd2c0ef155bc554bb74f5a675854ae4bfdba7b19d034d1b52e29c4ef21709ced7a647936eb9e24db3f090763750cde4e2ac37f949b824f0f91e91f7a97ab2d515ffc0009ede080519b1bdd1d8ddd634448bae97b426be36f39ebc0ee695f8fdc7325e1f48afa2df357700209a35b364a5ed8c20cfb0e06ee1f0c6f23717a42191b22060970efcc3eb92aa7b322e8f52bf025cfd2a8a1807b997f0b6dafafbcdc3569b1f1d09795f4f32a28094b7df1a3550d08d5ad8d7f88e7d4e8042ef53cb2bf8fc5708a04f95e528aba1b061b0f1037e3b97e4b8e0cff93dc2c66c3ad387f893a06302ed4a45ec766ffb79cacc4782d74b013b50505234cbe2a7d52a373a1b46ec7a8207dc4e0436829e08ed903076c51a7b8378664cac10f389fb552cc9c49495cfa037b74e2061b09590489f34f78531ff4df2725f97fe3d5533dcdc11ea40eea263d6b197e20da2f66a776358884ed4c1cc8f093f4a1470e40ca43cd1a5d11841cf51456cdf072639d63879c4852a1dd43520f4d05c5c5ce5590e791dcb69462b7f3756eb6a80939937100f61c05811efd36c7bb950dac35496f662e94f371e8e9bc170945c3815fc4b85646f3ed8da5269dabd725966c67e85b3ce94c47a8fe24ce4dde87c6a61c5af94258b8630d94581b04f2654654b8aa349e70fc7d2d3954cf24c6f6ac7a6551242b06f7babe4a271e4ac59bbdfa3afeb1b7ea20624192800b1deaf1e486074d5ce7d280febab44ce7da6b2271f084ab0bb3e19be4368ec89280d1052a663889c431d3232f678239de659656a81813d0a08011af5bb2d5da7f49335d430e3eb433c18341567a0f490b8b41c7dc5d7a6c39209ae43928c6351be92e8f9ae9a118120b72cbf5afcfaf75a582071a994b729ed73c7af677e945f7e2c1df2abd6afd1b68eab802e103f84e1a54fcde38d732230ce974190d78ef3a81027fe6205e07b02a96202785912c1a31ffac5015e733b234ca474d7e6ae647c7c08ed0152577455d7ec336a6827cf9054a3656898b208a07b5d37096e7dea5902f52272e3ca7f11739d58c2e34b51c17cebee5555bd8ce02987dadcce5c7cc7270fb8c41651c378fc02f7c573021bf0e131917cd5d1659b4fbef48078fe1e8b5ef44eb4ef2a04340b63f2a32eb405692ac2764932e98436001e8e958289c0dfe05dc149c40f31513d5442102210e1f711a6a32e2fde586e33157c222b727b1f6f3ac4f9d0558151151860f419f5ff526783a1e504b10c38e649ca7357125478a52605c32d44a1e7abf6aa6b658ac4231de1a65c2b0d397ddc10237a038ab854b2383a3c74bab0323f321030ceecd9e158b4367224e6a85df5dafbdf776b0092e6565b1cf4693d63a4d052310d7ded23cbd32f303a9173c535493682595a0825fc16918aea12b1ad4b5ba8a1f19732e5835be4bc9201b5c861d98591de34a1a00c82f7283e962188f2e7485ddb9825c87db582d40a2bbb6b58aef863322fd04afd8470f6134766bffe5a621acda19d0a0b54b1e1f63d3bfa06616647b6875995084955e8af2f956543ba15b1faeab7f38d9ad3694d0df004e485a5257463558499dd5ce2030ea407413ab71f8de011a5a0bd4aa4c254c57f77444ac2de94bd713768754b5ffce2c0d02254c82f0427a8613f04b9e81606d94fa25ad8fc3591f5d5d94deeb566eb94b24c78852c3642fba5cdca84ac78948e7a22ac8dcc56cd8f314f4ac274598ad0d248be0d2d62a7253f3d0ab1c9ef1d73f7271837fa5677b1564b20de894ebb39c7f9cb774a656bedcaf27ca82cd12c2b108a301c20db1a4502458949dcc320d7ee306df76fe1f6a514395cac4236ecabda571c9f93a7f78fe07477cb046d46a3b674af03d35e1e35b16a04a79004438c412d5dcdc98356ee45d7b66a556e0810b585d2897ff2283c478a7df00ec6f084fa0155f0922390657f594682802b80cb0805e5ef4769af7db98569642525f1916ccfb3a3d1a570d5e58e51b9a611aee9ae24807c9bbaf3d5049ed1d11970a9122a6a288102f7a06ea504cdc10f885800312478215094da5f58e4f7673f2485dd43a4198f0f986a9e98d43e58938b988a44a4170054b7bb3a4a5b6b6b75246522ca30bfcaef4eee947ca9a58b9ec42aac69c8bd0626919f35f3b3be5845d45292b8f87ce4be2517eb4f133219636cc3dc770d1da4c8ce2d621defa2cadc7eb93cb470c3a0f859a530b632203fb36e3519349fdfd4700962a7e6544bbcbbe7e904fc49476320e478f201e3e6cff0ed90af1f441fbc8d83d1773775187e11628e95af0a475d928af88fdf6b05d8e4416f76fe02b2356e7b86778b67aeedd55629939442d17d2031020cdcffd4bd2b4bf68d2eb7f8d370651304a591f8a0c768b95cf8408a911287d30757701dcab5756e0fe5acd6e6cd01d0a59294dd22134d7e9c3219a5b02af45b0e752d9d2258cd15fe46a35df5dd6fabf6c6ed439883c949b60458462a252f608d0d6264ce341da859036c740a544ab618e1e224a9ceb5d938945df73642d182c1208f0fcddb93651993644157496945b417fd9f319d88ba1455b70c29274a940b448d67f03cc0b3e3a13573bea85569bb5ddcac75c85741455921374b3e8f84e13cfb26a9a7dcf3f00d1068a846f1972888cbe222a61eeba747902341acada28cdf98b6c23ccb22b9ac69a6e9379b6ac92ce1ffd500ddc1ab2c1baa74fa4e0b4072d37b3c2aa117c97ef588d6595e2cca828f4f9c62995d294e3d461aca7a6754163beeb88d599bca12dde136e02418fdff568fed0ae58a5ad419b31b4321761a61ec290b77d0318174efa0e7da7e0a84f0a18970fc0f0b950da950dcab25f5bfd5fbd0d0bb8d1cb0eaade087634f6619dac4787c3edd202ad7c5224c544b06491c3d8ccd4361e8570d43169803dee99da8c204378f0f1e504a2fca3dd09e88b17a5a7496be34f1c98c2a6e22322fd79cbb9b429817de35c92366c6db6d547ead2f3f1632ac459081a0b311b1279746cdad653a6e0987c7973517cd2a1373c61c7cb7a599244c7ebe78928ab7993fdc39d84538ed013614ebaceaf5e0854687f5d82ef9b3316f22c8ebd126e1609bedc72ddc3146621611e53f489f67ce101d9927d3f716e7e8da44ab7aa1f9f99775c870aa2bbe7c360bf37e947f65ebd8456ee4a98c7e5fa63ae31aaa5359abab3b325291d847b1f8213013dfc9a86262f767d83a1d7e073607a7eb3a4d6876abe673af97e7aeb8a14bf5d6c9d6920b0da71f11db08753f3cd28ab75eb53e61867ff7f77fbeec1f6a0e8f90b3880ec15148aae76a3ee20a55bce0ffd2c732108aaa5518c453106bd5a6d90e16ccb8c76586e01f6098c877cd9f1eb243431b9e39b42d92501774a24b38bdd0255b42f250a30ffcf7a19127a8675b6b6a27c692bb447f26480bd2f95632db58613aea4065fa33c1ba74ae4a801c3e7049d4db25cb7e11f78654f392bc77d333a7528ec2749d5334cd35627d14a98ed62416137653ce50a7729bf450a5cf55bad98120ee60a6275eb9bebe558d2841760008f34825e59779e54b33f439541faea17d51b959212364d82f79e861e86a4b306db65c493fa0e54fb99383037f98ba12f5aee8c7463c56fa0ce700a342af458cadbc15d17fd61a054462567008913bfe6656470456ea888b1e9bba28fcaadcc11ec206004cb8b6d0c4ebe568d3bac9e72924e359e4be218231fbd6e3e1e54bde8d56866b8ecdf41d5559d94470b2bc5a9e3270d6150496cf0bf383251f526548eb0ac75011fc521550553f71a24f7926f44e697c3130615add3bcd22f370f34d33fdc575f61dadee01253006fc74d2c37623103fdbf89fbf4e686f38fefe44f1a1856d2c9fa4599b6479798a025185cc3e400b52f6736b1850895a57b2cdd63bd903367d8ca499729f73c7cb923f052f015433d043a38a3e4b726934652c964ddbb4e255c26d459c663d7d9872e2dd22ee796c9fc5aad14c80094d17e4a8ed4eb9372ad553b0365b2c7ebe01f1a87d562d47975d743beee5b0b59277f138135f18386c8bcf1acd80864e821adf9222041457775c0fade2acffd428842f2582dc9a4b315f4f3a4f067d8393d34fe916de916541a30e12b3b72ce0ac6c92bdbdd4aebfd970d42784b15a86c995ab87793d5d5e5c50bad4692eaf4b8475efc12e28a5c1e1468ef881364ee68e227673193ac94fc9fccbe4e6bc158592693fee831f74a6eff88dc2539fb53ea05e09fc081352f93ef5e180fe4b70740ea07637dcac8318a333b765ece96b3f8744a38f784ac095f3a9e3856b735c8e3e970724d46d3243ba7e0be4a004545d133;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hff2ae566d9b0784b9f3ef28c0dc598888d1ceb84eac929863d270682e83c688b10c1b1a6e18045c51c517c32be6fd57c554026dc8085caffd5bdbed598f69020d12832ee89a05c0b660bebe5539bcce42bebc0b2e45dadb94ce55aed799bf9fec92238ead0231125ec2bdac44d6f301650b648fc6eecbb65b18808d8733043fbd1c2ac1150e16ca13b358709fdc2a877d5c2931ead892c0735ec6a80e798fc5407fc02aea0638e2c353c4cf654588b663dbd68c176f565c2db5d23c16f0f8ab94e7e814b36877c0713d7eb51c02067787d3faec4681aaf1606b47e81ef3e6a5ba5393cb4f56b54b26ac26783415ca3ba910d78ab64bf236e9ca5fb0b2d1a302e20ca8f678100cd00c78cf6fb518df5e13a051348b17405247774f8a0290cff3b1097fc609af8dda69c16a52b99b9bc70d3c55e1d70bd2c3714339357003badb35816c2e935daf45d27f2c76df236fb3d46b9436b29603b2e1f40f7880a397872caa6551d8ba0c23536095e1fe0ee62007f2ab661d54051a873a0c56cc4964775d32a1bfee949d9c6455b9ec101b883f9fc4ec874e9b8e3f88fafa68207e2473ec5d8e323b890d41560d5c84dbed72b30a102c6526b2bb0966c28529c58ef9f0b12c9499bda406348108ce09dfcd7778b57fdb705784ae65274e4014d6e3f4e14e9d69879dc96e07c88db1ee88bb85ef87b0525f2a2230185d6934b24159b9a7c0dff52eb85e62182773f5a07d31b840f6b7364a3719e98484d67b51762de870f1dd2d2f6b59135bbaa449d2dc375ad7504d60da84ec542a0a9b4d134c246f18d98eb8cadaf14fc4004bd50f682e93d976c93522d82477d64fd922bc29620ed0424f476d5bb5375833b09099733004ed65da37b28d8394e5e289157e90e005827fc33f573e5606eb0bb03b28badf1aa87fa816c1a5fd6e9402a7188040eda2d80665d316dfb218565ecd3b2300b5348b9cc5315fa23681a58149d94c0349a5d6a8438a0e5fe6661cb6b04c9790774ac974731f42aae017167c426c9649c8c23053d247ff94f399092f5538fe285cef96e58b53cbd578bbcc500530791d52c9a50eb4daea1f648d440344b42ad2860ac3986d667d4bffdaaba0c5012f906d3c6c320c9b00c2e06e2f6550ee99fb099cefd07e2bad090329b67eeb896256d284e3b8277722a3c1963e94f212acd2ead8790c78f15ceb69eb57fbeebd1918346bacc7a1b1564546be496879773482d97e6741eceae6260ae4d3ee122dd4dcb85377d764bef3a606319db97623d25900a4f50c768ee516aca0b820c15c173a14bce78dd361f5679111ed586c2a9c4f52200b8b3aa805dae566c4df58cb51f056f61e0426c82e4ffac9ca4c8a301be291ee6b5bb2e3641641b7926438f8427a92b98ce929486e3037e1f8f01098d7eadccb01934c31c7cfaa9e1988ea01bc644ab0a97fcbce2c48e27655bed1502dacf9b83a5d1364e4c230eb2e7ac68ad89f0472ddec9363aa70364b35e5ad3ba77387fc864bbffaf37edeb35202a613fb1dddd08c6a8e97b74cd0a11826aa7e5ed20a26053a75e2aa545f523fc23bb3756ec7fb119c9b7fba34485bd39330e30055331706f0f1ffd7bc9518fbe12505ad8b43ce518b63220ac0b38cd539bfc26df48284b62407595159c0fa85c44c1c110608b2ea50813beaa8dd01aabad140b53c05028c50dbaba7bed52b83971c6ac7eb78c3e8e8f363f5cbf5724de365d03e51d3eb5bfe20dae7f055e9a08af33861ff03d2dca693998b1813ee91aa11d29322010cb2ced02f18ecc58ef05703910526fe984241f94ced768be4589989a28c1bc93d57c308ab182428b3929a3570ad3707590d8639410b4865d6f98d98735d885f936ebd3f64c0dd9a28ff63b05514f470687c6ab2223b38ac8d690ac6621677555fff283b78c16b133444110fa4f948814cfe6ced76ab06961962e97f4339bd8a5fbeb17020d944b1bfea983856a27778861e4a3f1e4dd071476ca10c836f771215a321d551ed1f1e16a161b7cb7a56d56593bdc52dd4cd7d28b2636112cad4562e034bf7fa58f22c90a0525b20bcc79aefb5334c89dd0ee0970b0196026c98cfe89dd30f22e40d9c08ff2e91bcfac03d73b8a5c9ebf7dfa4f17c16a6ad54b9a6281273c1df29e81dd9c82eb7f685c93d06553c32cd01ee070e376c3af1d99c6594c2abf727aee8373d3b3670760d72613cf5196baa8af4915f4a06d877019a55e716848aba6cf7cf63b5a011b1154d81c8ba9cd19b850681c71e7a1b5e7e83ae03d526f30068f854964e59339a757087f87b22ef09ba795593eb441f88ce87d86b26ee26d3e05041631caff264bf1a9b79693a2569e8dfcdd98e5607084b7a661968a30c32ced34ce86137696eb727a1a9742ab7bd00104f02434b1992eeb1df895f477a868dfa7f61dca1e1ca02c8017190967dcf328f57dcca28ce10c756acdc716090a32812e2f2da52d09bee3337ca58ba3fcf06ee41f5216d91768e8276343cc8c020049a69fd9c3687e8b3064d1d101d4e9592c481281baf111242cf350d7b221fd56667580796041e7d3cbafb3379d734b9ed6d1296d440b9031e9ce2b3f4ac33b9626a704ae54c6822ecccf9ef2a3f992a0719c55a6af630e5949fceb35c29781ddb7aeeeefe3f41235655440ecec67ee84221cef7b5d52a62dbfff23dae14a41f3512359d34a22b56c29b01f9fe0285e028a4c8c268e3c062338583824b203568d7145ddead46ac6e2c2f15938d0a4223a18b38fe953ead50915f507469f5f2ee026d45bbc03ffc163c49bce6d2438e9983def1236807b58835bad955ba12938729e9247e7750c233a362267aa8abd3f2c92efd91d259e2873e31b26b77e3614841b3ee6b614f43d276f783feec8eef444a71d39bb94755797cfc5de3d994ae6cd9a4aaac0afb6d67d1964c114dbed9024e34aef81c88a41cce5ebb6babe7d5c180bfcc0df4f443de96e016f17817a4c9a7276923fb7b1a2857a9ff9d0854e5bc4192ee4c244f9835856ba6bc64101f844dc0d3a43bb84b06249baf5fefb9036cc21f84860e9aee5716ad57f411f08912ef71eeae72b8153b3dfff821367a6129caafbb187c77e290d79b364c7ffe09a80292377cc6a55a35964054f9a86a21c2fa00a010d128b241c51445b6af0cbaa0058ecd94d7e0639c3b4166227f7b06e39833d3736b24610b3d47cd62fca7e5e6f513f6fc9226fd83eb056f7052f4dc15f3accdfdda33197fd4cb0ea29831c81699fe75e9271ccc0881d0cff9ad3666f448ccb6b9085bf745b79fe9bc8c208e6a00303abec94b9942b53507eb4e4845d84ea455ce217f476c87002063cfc97329f9597d80c1cb98aeb927c96ea5586baa9a0f6119b9f4a8a0d8398cd5ca3f800310148b54aaeb5c0e0bf887e932fe7eb79715dd1fd9b819e4ee3f216d071b6ef94f2daddef7ac9a4306f875521e809d6fc8c8defd88394158c196953786969ec864eff2ffcb649a5ff7189ca4b58ad9dd39def90d49a87cd0bd98d3fba324d5afb1dae2f506d347eb501d1e163b995e79bb501852bc68fed669ac5622006b5b0fe5b1c648464a568d7ed5c9c02c83032dc4ed3c2141aae9648a0f94fb8ffc3e494aadfe3d0f74189287cd3bc0df694eaa06bc4d57faf9fa331b3bd26a74b1b83ecb0d3cbd298f7bbcb3aadc5ae3bda447d7af8229259f3853a23923735da6655e7b669e1feabf9a3ee53f45810c6e9b42ef27deeac113d762cbf5fbad4285be7c2933b28f20cb98fa150374e26edfe3fbf7f5888ab8e2e9d8ec84e57cdcb72754a2658c10d7a880a3b131c6c7980b9600d659594d01e37a1e6debe1b77a6681a07bd44bbc99c244a9043524e25ff5a09fa5333537338d50768c2a7ba4f068121db4a53c4477ffd1d9d91b69552ab64ae029606e879ed136bc487c4bf6007e4ff57b725edab6fbb1eebe5d795a47558be463dce9d590743947f682a8fbd888708ad6c10e50637f85f6ac2c118b6c7314f62c046f789356c438690b3b29ec7aab6ed8b9ab9b3335f9f3bbbd822abe27e74ed9b33cc4125290dabbfeedc9a7c86d2addc2f3e3ce4c0880192460444442bdbea7836f7f971f8e72c5543a0387b5afa31ae186b54445c7a2a893ea86e80cab1d763b3e5e710cb1d7eda06a4b7276bba283a61f93218771a0b6fd21a3335806cc003af1909c2fa0ac078846b5714c5b106763f019f234d0eae62dc796be6013a8184297771d1864d212d2641afdec5b8f811f209de5c3cbb5cda77599766902e0b6464c1d39a98dc298770fddcf02af447b045a1f0ff568723b15c01e54af27eafeb5b959db212e1ce2367fae89523c2f911d0b25c89d8f0c7a1e34dcdadadbe88a3fe29d771b84cf9280e48032fe140dc5e2589dea38d2e13e0381036caaf0c78dabb45009f8eba9f85c7231d4eff2ae07e5ec4e9788fb6d8a5e25898dac4a866c3a8701b67ca47919f3d41cc48c94c64c368ada36c630e55bc996833c90114c07e8506355cbb603bd8ad01cec3643c0e2daa018d1faa8b479651221f5fcebf5e5704f6aeb1e2a9b9ca9c8fa75d17bfcc6b2707f43399d2bcac59f833b19397c2091658f5aa3c2fbbf9b2781adf41c909ed27919b5b60ee4b56d9eaeb23523671b92913619d8768333d9d02c228200b7286ca98abe2501eeee7aa1c6d5d93d83f9eaf2b82355e59b8fdfcd450025f2e87123331fa087cd195920cc883d36808539088a332dd77404722f9f24f110b53e65ecaad3eb8bf0f8eacbbf96e25b89bbcb2e13d8d2aa59b819d549f8fa8fac13817d3dbd71f604ccac0311e1221a0133e6c209225c78d612a97a2c03a063c4ad9f363bf05bf07dbbf5cf98e96043505f7db975797cbaf85bb90ed9d09694946bce01846409eb7fff7d953efa4179653a766f9142e939f19a2639d53211821dbe4d59e534946ea7e4cd1ac4745c6b382cbad07393a5b0cd98fac88184c3a3e46886e717ac335610ddbb17068e295868e2059d10c11845e2ddb4649b5a716b969af1cfe26a625f414a1092c4a673f7e89f618ddadcd23e2774464ed7191dad493f2178f539906a2c24b3ac964f288631f41ed6f0ac2951c7550c3f09e3554a744e0ddf0fcbefa7d09c2d70bcae50408ec144954b14281835aac4d8096e938f445c57ef48a5b7b9f5b974dc8fb40793e849502d3de61d02ad74951f4f23d4750ee6abc45921b24cdbb428f11f671f0c893d6ae12525b3edf04dbade9166403b2ea7620311eeb4a1d8a0ffde3cd04aebb728b3548d2896b3c1a0a4691e3db19c80beae3e8a00f34052549bf8836b602d0f315bcf2f8cfb63317a6fd4e7e8ae65d754a4d9dd8e3fd22cbf265787d5200b594edff28f5f6decd21fbda34b7aaa46769c0994631c148d646ee8b8baf55552a5d344e466de385ffb62e165cb0510438d414521b0260c2e2efa9c7c9d70a7d8ca33aad17adcc4d6faec833bf82afcec1faeb94cad252c2e769489e4bef03b3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'ha6b08297a839319cb5a6b93a082787b05045c3dc46637a4449552007102bbe33f40cd3315eada022e9b4416838ce20838ee4534fda44c0263a79b7f32a69e38f9e8863953f786cbcd64d7e91c07302b97d1e97246f5df14d4378adb4d23946ed432163d9f08b3d7227db87624c418329a392b01d33f676769194ead87142572e327d02b970cf5de8b7c201b367cc609e4f46eaf3b2f70da3dd228ec232713a21bbc64393326ad624273c4934b6aff33eb6b2929ceff7711c2a87d7776f788f5489ac98b37b525419b5716a5e8275971d2524a071985f4e9de45c9b0e9511fdf95290c1f8e00cf6343220c7ca3b2d5aadec22d81664575164010985e0aac4ecc1c13a0660938172954a61ba0f721b1266ec2b755a6eab9e24b387f497719a2ac06c36b4a37a682c44755a4864ec258b6c5c63d542861fde873ac4690ce36adb91df669cde93d45f7a5fc40796615f92f6e69cb4cfddaabb9e0cf53116cd426f03e65c85698a64f0abda0274061c537c8cb3914f961355de8dc6fd4a0404c94b52042ee7955530790de984c464dfe3e9c7aa73f892ed4ce1e09b960f57b998c4bc60c090b2cb7399bacf8458a963826bfaf30cea38b24cad438c48475317a3c8afbfe38e1277177e9c1618c51c5a47f15b5684945c1c752b6f6eb98c434c0cf1a9d989eb9264165405b4d85652b9ce6b995b6f70c09e755b71c6a2ecd26dd6b0db8d48370d76c98a9ff6452cb47e596a1f6289368baa7de79dbcd06c64c4fd26b6093ff044e48557a388de3c24904e389a5355f355495726ff92ec564d8ea028142cf5ab770852ade1645177a314d045e8916884e8b1ffbfd8328c7acfc1e205c096771dad5131a407531e0c1d9766a7302c2d551374a6e3677df04844ac3255a9cf623fbb3b0a7a34d2fbd4325ffcf2d46ab218e1351ce1df6f468d54a1c46add283dfe62654712170b75a64ed96238549c7f008aa4b3e414dc2a8eaf500366fe5ec63404d896012cf8da1972d43a78a96fc3ec5b14618ef44d73ba6f212cea4402db0838043c0f0a0206a69767a5341cdd1cc84fd142fc5077290301dcad38143e6793f1cfa7364f78e2a38a101865a081c047fe759b4a26a65b275e313438424c660d46b6d87ccecd215db16c27ef98dbdf26bf9cf7732dc2d6e4bbaee3109a1f47deff5efd445dab3d95b90693e6525ca0100abdb736aae4434e5244d24f4904c84b37256cca5969ceff8b451391eda10dafa72e5f5cc06cca35b2a765954fa9499d20b617d40ce1ae17ab0ee2eaef17a7bf5bf44b0f999bf6fa1422e700e50438f86e7ad341144217eca1de3872d3eb37a84114d8fbcb11f0209740e2cd1d0cb1fabb1c50ecf2e599bb78a6299dbe897edb503fb26a6c001da6a3504f4eeece0e7701f62dfdac2c2ecb32b61f2850f0f247ccdac023b7cc6e57c327505989fd9ad6c530883faef049df8e96341901459afe7c2000317a4c4bcfdf82003f8a718afd4ed809810a3282e2f160f44efdaeffbbd41f0f095ae1a564307ce4df2f21b86714911ff4374baab157678c5c1e555cf9f69e394ec6afc4810507b1f2b39e730f27073d41a47726290abc826fcbd63e34ce8bc706423a4de09107a5642d29e6900987274f766ef5b903fc98f2ee4c60397c6c83bd0c766bffa0ae60126410dd64f1417ae3ff2cfe00adc49b287fe47b074f67f9f131105854400d9d164bd25403516b90483636f1f592080a9f9df5e34a98a2ccdb1eed557445afc0856bd943eaa9a560b5cbd44e5dd295b226f804e5b7fae61ddfaa74f5c03b6075f9d5957db93c653aaf9983f416d2b777a1f94035ee1926761d824789bca744854fa53094a426fd1f30f6920711a1f57c1ca3fca153e4fa73f7b5bf6cc4b05763747d104972b4c398a23e12a3270dcec14621be64ebf7d63d228efb524efcc472fae34c6893fb6a9ed4dfb0cf23f33b8d1333a1ccd1729621791b94a6b7e829e3650f5a85b28813702688430b163cc07d84e4bbf9e7c8994be21c7260a738581d8a52c7a001e472d2908d4f0d84e08b7198e3dfa46b5e64b6db0d49a290d6ebcf795bbdff4e7940913e933db0fbc02f2bddde0e769125045e2bc5738cf0c1251f69167bd1af48ea683bfbe31a5ff3e4937729dec7275b3ab13ba5d2995b609a1d58c83311cec7c6c6dd488efe5ac15f950bfd34d3667cd3717f6799c96537da018394305e25e3c017d7f079e102f460c9d93af9395b80a76cc7f4f9f19b9fe4d586b67ed4f9c232f7c3afaddb275dab9707f549ef6780777ac5b2f18c4785b655986086d6affd506d37c959013ec485b196b7d5f45d4b4dd42ab7d2e37df73e2162d73c3be788c3f520da0f426a11279413a206f632f5617e527418db34693757cb7e870325081bcc18383e6de0f4871b75182d4392defcb49e11275278c1e0f92f64739d0506bd781afcab5927551e9099dd610b5b7911028581accd0aef71437cb39377f52f6fc676efe938385ccb44f38f3b77581d9403072fc86c80dc9297368854dcb7ddb5b060298a921d992f44cf2d2866ccd72380cf643d6f305d21590c764e7122c78237ebf1a05e976e363ab9cde654b7e129f8ea48a4c706005d794ab2b2b158dd4f9cd80db356c9a041c5ef1c1a71d8a227336627428ea197a2ec18d5c8b60d09c2ced0b60e733896d03cd8035456a7639af249e35459d19129102aec76c16ecbedddf8fc42203ccdac99acde9e6e53ad91b1de71a3976df29b50084bd1ec3f9d39108b9bf128fedd299cc572a809f2ff397f70eb0da9521b2d8bf506ffe2bcf8d04a1362d3a5a10151f039b67ce7d8a587e38edaeb98262691a195efa416660326d3b327281a89970f7c52ed8aed5e4ae1f01ed13cdfc0aef1fcf88d24a90696a4b6a792df35210cec7f6a6caa2b052d60c6577c4dbe82bac567d46075bb5141419d6b4e6d5a4984783c8367b2e154284547526ae7cca15b0e1dd66e1c4592a4dcfa5fcfbc368408f64d635ffb80888008a548c8126dab62f2c7d8d402be1d675183576a888eca63c912d5a40f4235b1b6d2e58ca43caeb140e52e21a3e29df1ffa40bdeec8ea81fcaed525371dfd9f2ee73b9252edd0d9efa05178f0d93d1e8631e879abe3d4ab9746aac481ee462368e02d0633bc3d4c47aa2e918220b41b1d0f1fdad6b52090ddfea78894d9c18415cc9f994e183929dd986237983d372f30ba02fd8a1ba0da90d20f5d3300e87de2f93cebbbb361a589e351112beef889d5bc3f47b8faaaac9995542b426d2b81292d7b72abb4979521d0c0c531b0a1f369e5c83bf05538130faec073dfa644d626200196cb239a89b285041baf596cdc4331c00785c91981f324702d997bfeea5faed655e29ec6903ab269cc3891bcea0fa7be02dd38860e7a8758755f2c677f60cf5e9dd777a21136b743549ac0d3469f216c960baf3748d6904f9dac59d007a7e9b67ab8983c906b90722aef07f965f98633ed9c84834138a7d396c33b0a46cae91f54390bb8854d8a8daf25baa17b94c54e5b6b045ad23fbd19057fdfba2062c3a226b42a00513979798baa3c0e3fa16c1f640b30580e517ab0dcd8e597ec5d4dc9ba0d8e9083f2b060a553c81d2fabb6f924d5e59be1588ed1d86e7381eed31423fcae21106b19dad6bf4dd8262a1ee127cb1151cee1747224393a0c5266132cd47506465aa5c1a5baad169a8657a57abe50a12dc8ce414a5e1f8001ed1704c508c91d60c0f484106c5053afaca95dc87aa77ee19f61e8ddaff3ab8831d0512c1deef9af598c080521c4d5ac2517bdbea206ece911a5f3d5f3b8a608829c1cef18558cc5591e9cf544829c394bf9bf28cf1d3be5658cf1be2b2dee0047e914ce15c0260ff78310e6716d4e8c130016a0e3c74eddb384375be5a377862ff9b474815fd20ec4253efbd2501b0bc3e311a4867fa3c197ce19ebbfbc347602343dd52b60bfef6e8f6581780262643995d399860603ad1b4d61f4a3334725e358d1203e1716dc983455e4060d6b4b695cfd69557f33e80bb8fe060e4fe658a2e9544708056f4d00e2b0acc6d46fdcbca59b8dbe083210df7251ea794bd4137263e0df4cc7b2d754ea98ab06943a6086fc5ac5f8ed5cb4df331f6426abefa2da2678f09d771c7270e8c31df5f007a51e37b9626f2ac1e3dca4ba409dc15026a292e1b29c7f3554ac6146aaed979d3f6beece5b36691230b0d154db30a26b761dd523438bac056387cbcffbcbdb4e51d7de3a1c769a7f5bb08bdeb0526b8cb26a147f06a28db5eefbc6e2e2bc8700da2d6022fe0638d685f95f85b1d76979b18251ff52e44c970e2910b32d6ba885447c598a72d23932dd3a8094cda92e37145a0f56d871fe95f7cbb44b330793713aa073a730f77764315611a27c29a5ed6c6842bc4dd07346af52d185597ad0161b89d93c6b7d44222412ecdb2cf9b01006a8150e565c82ba3e9d7284dbbfb367833288e176e2822cd890f3dc41713a87687e3ad435cceb94504bdeb67c14628e2f04fd9298ebf209f3fe9df3c85b28ee86a91d31a4a114378c580a6d086f819c0d12cc04ba1fd408f0133a7325e982a3080cf2ca947bc1bc3f40780798ada2f6a7ffed12f81fd5308adbfcaa08fcbe8b56c02ca05aca2ec89549707973ab1cc51d2148b60afc6a15348fc4853fd6bc872a795d9b9c6263a13672b88e59f075be13040fee66f14e67100d986d032ba0f91b66614aeb124868e5e70c85c20b9ad6631f008f7ba82532e900578ddfd55edee088a6a30f3e9a57d71330a72747100ea14878a0ecaf0299828383a96cbca179cd39387285634befec7f07aa1757289cc4f40bbe77f70e87482a179643e84dc0bdf9f6e7eda23a7d74815f3f7f2ca08d7dde5540316c9bdeced522831f57fbfbc083a4a2672a5deb97dfda2594bcdcfb75618f66c284454c2dde2960588ef53fb6a8aa38191bd437c2f9c28ecec3c8d30315aeaf5876cf1575f9e7317a2e47095f4d8c4de13f432f0999e1c7284f9524eb4bd470acc21ebddd96a86cd1264dbe81338b73072534ea4c878ceaa277cfaa9f8eda61caf66064af41946995bdd88d8643004cc5b934aaf280056b1e2d66ac69ad21398a26875aa0a25f46453a172bdd591f9944adde9c137345447a104ee7ce3e61b1a81aec79284051a73d75b4f77934a63343fac29a9fdb5b10fb952330210c474defe8f6c63c809031c560b76ecf5d8da861110581e08b1c3cff98afd4bf00a0a6b1734da88fc2472ba3e6b17241134ce7ab61c99cbe187dcfd5ed06519d0c283c19508166c1739512d9f41509c19c25d71a41c18e2714ee6a02cb98f35f8b9da0779faf2f57ec3d7ed3b8f7a51fae9caf4f5229f0002c56479db9ec76bc8f40f3c8dc1a566132614b3ac01819b585ff131a3d08f61a9e700a051692cc707f83d79f4646842ddc6eef4608ee7ac7dc081ffbc9ddfcfb9d71f33ea9a8f1d43ce0915778b63ccc6a0bb99a923d7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h68a230d4eb5be8bfefb71f9f9bfb219ea770ad6cc8cbbf853d1d786fcd5db574905a00d19cfe54f4b279689663b326a981d5ae9a5d3df3350b230e850b13e80b29d74d099fcbb07c7fde8e068ed7d0101a016396c64125e780f8786f06024c5a5b57313448c7fac892a37d59dd79a80731dbe1eb588097aaf3bf8b4cbf4e63eeb8fb44c5e68a1f02310372ed7ed3bc48daba3b498cb2d21533155159c8128d11a0b820c0e2176267fcaee3e33e9eb1ecd47770af3fd5e5b6d6149b7c3455465da506a0daef5d7a50a8b0ce5232211b82a5e1bcae5feb789d0a5c6f5daf1bddc629aaec744fb6f6adea048b61d1f47ac772aad7083b2c6c857c1aba21eaf99a74c4ee4ae65b9fe251cb5d64bb019572fed1fb6748995712117ad0f22c2669ab1e6bb791f595ca9ae4c6bdf4c657df345f39110ef2c3e29a054ed37b2a16dcab91b412fe8afe276975edd6434ea1b5cdfffb1f8f373c9dc28b996a5783f94dc0c5453d6678ee4380334a845b36775f2916f947327b3f73b2e394c966925992efcca87c97087425ac1bfef0bf40872b49e5da345ab9ba4e0ce56e6b638268701fe9bbe3ce560694f1e2381e1481cf3008d183b51e171e062a1a5dc0ce45d72d80e791a539905268497cfd4b1d5658649f37bfeb4659f9caf025eb0c48e74ea6ea3c5bf4b893019a279eb6fc6d0cb1ba3ad39e72287c840e44497923623a5a959a686d6af7f6e8181c45c6626b8de0c6782a66d85ffdcd1a07a93a0c7c3de1220a84be552c3afabc20857cc8fdc952228e7e2874e7553e194019b113356ad907d3afbe313d29c1e9590c59e4303d7171baeca8d1453ea68d900b314e0da0e41ebebf5fff5b9a43798362aab5ed85dc9be563cd67820c17aa04b326e17292aa6fa6121c367b593b4914ff3fe1d635caf5df633b26666151efcf8e23f44566f0d43484fb5054581ed66a0ced7aaf4decb55142d978a45175ebaa1ad66a0fbfc9d0b668e7000e3b4ae45038feb5be7c6c4fa54a0809e0d489b09817b5bdb2a634e18d61a1df71eeb90de125bcfaffd34587159fa63f9e622d062b934f829e935b16a739362397c2b0c6eacbcf796cf8731c65d5de8e8e81b517da55a056a77b21c3fc10f05ca73b10252719bec269726543e6c0a824bc11d8d96168c5c29499498c48c6ac08a71d38f70cbf1a485d41330ced0891891cfd209114cc9c73a4e4cb240d8bfb5842f51845618d39bc254351f89250ad1694a1ad085e4b00c5860e053a8842fc4a686747408efbaf773c1c5e88082d51721f48e988aedbf60f05eee21756523d7728df2f8ff97cbc86ae8ef978242eab2e0393b3270dd0fda47ea8ba95f9ba8c3e196e92dbbc48423e9175086e11908efb6441d1f74050778c118db1a6715b6b2bb74be04b06188aa2a2e3f39e514c3f325944ac6d3ec9c5e737ae7023c87b9f8101cfaf4947739de6b42f3e7f1d697e9c4cf8967b73cebee926839de41803141ac6ec82e131adbf95ba65afe0de4614877e6725c21a6006a6117e32982ea90cdd8befb3d02bcf6785809307fa49040d98ca8c62b032d57e3327744ec1840a52184f8946215732159f0eac76979cc54de7c0520b1a08db178fae37d883a14fc911931cba48cb61b32012e5b23da412717cc007a6db9f88f892a600f442a640e8643087e12b6c872f2c3c8355af13a0c314451030e554ca3f65fe2832bf5688dd50e6a96083a9962a4ac541b8eaf122f07969d89bbfe945beefbeb74c4e73ed303be340856fd0efb0db7430bffa710df3465dfb1bfd33bbc16e1b2f9603e224df5347a2d7de7037f5272a58557d3db1827e806e40898d5d92ecb9b04a1a5ab6214f904d1debceb975eaddea267cc44b186e067867b448a9f926885da69ac3bc8ceba06327f33e5a2da1a8f1ad754a3246b32f376d060966171e929993464cde53eac76e259a77aefe02eb9be2dc401d24cb36bded77501b7173e46237791e71daacdeb4c29aed88fc5fb2c16b0e8745d71213a9b01b01a6ac62816996d88f62894201cd7d66b64fa0d328d8d7bc9f66351de9f340b9988045175c65c7352120eab619a45d56d357c0da464124df9b3f9f090798791a3f42dccfce3475f93adb496c060e2404138903838db2f50cdf78f68171548bc4c47c5fcff6a20134ae7a35f6a1e9245cabf9a8b09b417c756e6777c578d9c9da191b39a8848f9ae0ae9fa6e9458503f1e5913d3b3752bad974040081613fdfd475d9294149aa86bd8180a8ad483f2bab544025c8fc482553ac52e5f0025e2c2299f83c256b04218c5e221e82c73bb0e5dbaf0f8b2d8b59903cbef150fa30da8faea2d298561b6bb08edb66eefbeaef50054874670f5c656186e6ea90a3d1a01321eeb93548cef63aa87d7078361362ec2158b5e5b999175e595a282cd8475124e640876c8b3896444d9d08e34f70b0d7d70207d35a1bf54b6111361875e07ae832d330909eb0ead84f5e7dee5f98ebf6e84e89c03d5f9e7340c4d9c6c73c0fce240a6d3de4554098bba2faf50c2779e06aacd1852fceacb499b04175dcf8e4d2ff8e1f83db009a970a4ac13213282224e1a8939161e27d1775e2d444f263693d55620c4639414d61ed83df11379f21b72cbc37b7d2ead5103ff759eacceb52b6cfb71ade56e93d10a62cfa4c9d102f1ba7b3c18e3dfefd42df043f710016304dd9f828964be8416ca2a25ade5f79eae5b2b08ad9743828a2121a921d176fb9a1efa4d8ec9090e1dea1dc7b569edbc3f30ef83988f1e3527721291d7732472fb440e6b8f103d6575dd525098893e23e7a06a1faf01941d8af6b2972031e424ac8a426235caed99165e975a5d53b4b94ae5540a7f9fa0f3a4cca85e30a82a94137cc6d72cc34cc61e0e53920aa72b508b703ed5d8c60061dba843e62a0ea6b90048c2b40e943fc49ba7b5878128dc82db3c6418d0a3a397632fb6f52e71cb7208e105b69a82e41e6dc4a7cdbd063a0466094b40ad818a94a915cc9b2d6527bffa2b649a4f43f8b3c2854e48b99ae27900271df40070b06c5d308d4829f2102786a2d8f49318af826f8d85812513a482691a7c54624ed2bc569352e5472121f7d02644dc2c6decff47feac2ba890c923369835b999b18028745a24b9f3eca4e81578acfdd57d7831606a186cd0dae2f4c7ced386a79f2e21a6225bb59ad11ed082e1d63e5c09c97c4eee4cbc67e18301b9014186630b4a837f813587cc4c250eaf0c4f900e9d589146ceb6ded3745118a5de3f41013fee233144f7af6056e3354f3f705000f88221c63799570b8c0d2f68d3902c186013107937ebb9128634df4c438269f5c2e8ca08dbc28c235fca022819f12c64e9d0663c2def8cb59b38f36af072d74a88ba6c8df145838d97b8abbc4df77e538ca43a5810a361510fb90b25b24b1f305e37f05cbf2d1dbbaa85c96ba4a6c7b38919d45524e68ce2601d8a3e9ad86255c786ba38e718ea158406cc291d470a98537d07b034e42e4a6e307375bf31b9390c3663d05f535a93802a73a81243623a79ce0e8da6e6a0189e508a4e311d70809e688cfe27d965a22b02fec5860b547ed0d61007720ee762a59af02671aff59aa7181fb1387b878462c613dcc7f5946eac6be4c9920fc0fe78215a17b5c7a9f72ce6cd73b8849bcb8c15e34fd55ebc8738b00d49eac7a2f50060caabf9eab127c32db77e464620771f2b0eabb7147a4d53d3e3a50722f00f2361be320a8da4409363b2832c3bfaf10c80d78763a3f9609e0ba6a918fcde7eee7cd205cfa011eef99cf03ce00a304b09be559706ac0ff029224d41c59dfaa6949d8b9da0817ce44e0953040b8ecfc58b841d02659610ccda3efe97da9d66a398ea2e6430b2b8d257d065460d00a1b0fde8d746f8f3efaf1d0c2efc6aa2ebc5c88a360f0da854f6493d3d1b77c4ac66f661d9b1ce461811e3ae6073bc6ff0b14f4c560fd826fddcc85185c41ffae93e2180d7567637bcd39236154edbd27566eb25ff787d43b5feea9c81cfe94368160ff59be0485a65bf6189797705b528e7e139f292a660b7a2499e8416c21ba5cd334e14074281bb6fbe7f626df22acab3f369efc18642259061e19b9540ea10585c12972e12aae0412f18497ac0f386f0ae7d4d8669bad697b65a6847129a2600a27797438dec982170f7696568e4c4b21095d5fd385be8a32f390a815478d16c7a5cdb8416be907d2bce18c7bb312d181ff4bd40f2fbbae4ab2a4b9e6e6acf5fd74b155f1a8841a90dbe2efabf955331133b27a7e62dc102523dbd706261fcbca3edd9df54145782d63a7c177ea17e96871766924eb832cc056901bf64db4316bd590cfa87d6ac84dddefbf69f616786b3c617fadb10e8734de19737a79f0d55ea0d4c3b53135b898580ea6b075e94ce662b0566b6693763de554463b42c1ebec457037074800821055f2c663fb869167814ca2698bf784c50a78b3cb151c5e5fcfc89a3052600bbf2357801d0754ae99f14ef138fed14b12d209bf8c108bcf8ae3255abe916c9e62a023ef5a226ad0542154451e1a787a4611e2266c2c1d9a0f55948fb65a356a3f769bf797c3429e03a186d81b3a595de80a1be427a1f28f81f46c8ecc46aaa37165ed719c14c5f9b07ec4158d61f86e2c5a0a6cd1b576433faa776ad05bb0183f3cfa42f5fc149d2601e4907043a03ab046b9238bf05aecfe2e769a8d10455a2148a41a930cd8429340209b944ff2c983f8283498c0513a3411bd602050a262aada436fbf30bd29cbf5c6e402d4441fbd01284d72531e70c3523fcb856b17e83e3443336038afe37a6df6911bce5feb4b5f63ece363616cc97afb4fd66fe2eeab3878f25990907de97c6cb9f5974e36ef6698657eaafb5e0b1b4fd7f7032e0fe0d5524361de77ad8a4dacf7d1e6c2f179d59281b189546ee3db2b007d684cb38175beb0ae765bf82e9e33134fc3eef53941b413bee1d58a70550e9c677bbf34dfbc0c507212e7e6e6ac16aa8cfd58efb0a2889046f1befa86fd3e363ed88abbc4adcb5385d308ba85bb00a9a4f1b97b2184befbef4fce206e7ae930bcb1e3a39e661cdd1b9f585468a6947db89dc993fa67e92a96ce05ddb39f4f9a7c815ac6fe9b9258d343f30ca503bf32b62b170c71c9082a7a468e89d43c159b68ea461427683eecf73be1d5a48c8dd12d74cb1b5fa98176f25f557e1ee5019bc72b8285d9c7244a2d67a4fcec07754745c2f9f7c28501dac799912f548eb700219d7ef9630785170d52806f827636f3ba85da2d2e85b938db496bd5b627dd3737aaf80fb62ff17f01b6d95b54996408ccfa8b329b1b3805e588ef286daf8eb1958f4ec6d44f86f59d98ad015cd65bb75482c11e91d81f3014bb8c818c2a664bf3af7a70704418b41266dfd02b845a278149951b730382a52d133e402b33595a0c7df376847f23c6a26feca06bb4987cecd56c0f904120edc4f0069ef62a7d0e3d6e202d83c852d693efd7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hc9ec86cc2c0e68ffc3c75ed0bb062747538b4102f9ba918f588c4da8187a2e46ecefb24a51cb4623759f069dc8c48a04b1d5af955a28b38a9e17969f2004452b43403b8f3add3dd485efb194102247d31180541feecac49747e78790cbb530f54dc0dae101774a54df724a3c595f5293da1b9dfad87621e59ac17674305ab634544e95865a5619b812cf674362941224f7961edd8ad132d8846768131611296400102c364febf8cbeab75418f6820fe775fdb15aad9faa0341756b6185d8a0eebc87b0e9b366ac0bcd36d82eebd2bc4f1c125d2c18759f89656215f97b88326b3df772a5285a8c26d060b01acbfb94d076e04cb55bde716724dd5584980966688dd7b8077afc00d0b9b359a00a39d5e87d3044c76f40e7c6a9e0f089c6c9af5318e6706a746295bc0417b2419a1a5c47273876dc7c5f025bc49ec364cd603abf035e9e919728b1003ccc27c7e65b7d761f09187abffe946cfa94163e4077ff2fa3362bc6ad1f96951c097048294f6f8ea06c2cca2819cfa33d417d67319050a73acf7834877f826a5ab670380fdcacedd849fafaad9f80f9d92dad84cffa4796f119dcf80b2c7cc1ed1d30da6f4d350c16253e861f542af143ff3a2d27ff9e03e61088ca2d756e94dde9c00364d51b2c7e9efb5f44e88b8376732859a8d68e148267ef3ecb5f03cbf15bf250b14581ca4a54f5070d93793680a340b76569d6f50e01363509c2c3916c924935e7463d8fb8c1117a8979820879c9a27a8550a9bc222bb539df38d55319a69751c3b9e1ff3fe4630772ba48cddd5bb5c28a27e7aa6e9da285af8f81b1eaee81c97d61239fbb154c0b5d6d065cec571a97405bf83cc0313d0058e7f6c283f6580d72b554f504154978d712677c44f36e3b7343a3f3833c129951f92835ee439a294d0f90c70a2e81d042e2aa1aebb4bfd7a5657557b55413279dfdf86d783ab56283fbfcff2829e76cd087fca036d61b16e30a5f0e4ef62df67962b206c08d19f3be25a3f1a68f4cae185dfbd54dbfc750ce07c4f7cd84fdd047121e8acf0f65ed27200ac7139ff6ed1819740f4593e749f4018ac2bde0bab04054bbca6ad65f1854c9fb919518d58d8cbf11b723199324b1d0c64462e0ced0938e7d48da661228525de20e3612109d7277b1890a99b2a9423193ffdf2fe0c664999b01e1bfc1f5e70f9f86758cf73de0deaf07a52e9165cc432168bb994b553cbd87ab446bef325f268b59e53546cfe5d5a543d8738f2431ec60e452e9d47218aaec20b98a90245ad950f2ef1139d512b498b824055e0f882895bd70ffe4a4857feaa355a8df75b4036a97b3c25a85aad97f114c372f9e4dbc82cc17446904bd5bf06f10898a1e1ad4b1282b8728b4cc60c4b430c6a710dac1fe40259fff7955f28037610e59d762afbdfcd83aa04996018bb18653a90cd87601cf8111403e9c3299eff1939b5a6ea9605797a610577ca72ac87bf9d670f9eceb6686635af143555f47f640ffcadb603f0de94e59317d88ef4d1433093fd6b9fa307d1ed4962de438990f233a12c10862e7620d8e7e3c4b1c58b0afc880390d0f5bfa4f18b73791bb4b87ba88a60e1f24175fa99e6f7766366094e7e1d099501815e35775c1227e28f21e474216518ec958d28db8d595f34153e747e7393b9cef7b18c9a6c1d0058b7ca93d646dfb6400b2ad52268447d25e91298f04f0658e79eb1e4d058b8b4359295c62cf8e478632020cd8bf5ec76a33931faa27fb4cd06132fd159a062d45a73a3bf405dbdca1400372ba9d884ad7bec50039bc21a9393e58df292dd4e75c6518a56b5554f22da444af6bb17e5049fd1a6c401962baf77e8e580602a4a4bd378470c7bb91fcc654c80b3955d4b209d38c84b823e2f038de4898a63d2998eaf305d353207aaf7cffb97d862e0bb941db72b2f9c388fbb5c6fa0847bd84a18b01d12380642dcca2363c13d8b63cf71bc15f677ec1ec0d7b128aec2a077fbd762331423b9dd53538bfc23b18a180be1a28e674cc2b087361be751c9c238f1463a36f6df1d942dddd437969cb32200b6fcea7babf27a9f2886eb2c408070600ead1566b468ec3dcf3cb8428179f25b7be160ee639e108a38964469b2f9dda031036c4483b082c69e9fc0c6e390ad07f47955be91a35cd04a5fd72642d8dfb6b2d2764f05e16042ed619b829d43af444b80182802211afc330f3005d1a25db08a03e1a135bd3301b8c3b1db4755f73b045bb11b695b800145301058dcd6430560f410a08d5d373921d495045c723ed272c28214bddc63409c888622fdf6f5b3c777badc596cbb493e4962dd79671c7f79612e68351e7e0302f0a51b0cdc7d9ed86e03c07b80e9c5b26f1acb2c93ee4cf2ae260d486da47a545c74a0c56de626df5ef55269ea3cb9807214ed834a56ba43be7ab95ff0a96ebab9038f24fe09810d53cceae790e71dd2ff20d50ed10f84c811fdd32ceab7b0b8b4e31750c4775fda74c0776c7a70210af90fe9371abcb31b5998db2df653d746783fd9acbc6c1c1e7102cbd08d9001f8ceda6ce663377a95d20e071c0962ee2033be48c2ea5b95381ec090073da8735ced63990d541b5bfa461faa943bcede1d92f9e8db91fcc8619c3e89b42f5df869903ad85026b3abfa99df5bdfd141e6dabdf4df4902731480f9689957fefe44b7840f2aed15a7b9facf92126d7f4caa7f12ca7dd08a30b40b9088da9a835266f3d31b87e5785d0d66e70272b7c80cb29db50d028ad56c91915668abbaef37f8225dbd159f3eca95590717b226fc8111f6b98c66a8b9070242dbf727d3d2fdd345fb3649550cf6ccd175fd7a5e28bf5b665ec51ae44b0a51a90d60771447d047884e30b8869f181529f2dd11ebc95f4782972788762063ee1a8eaababf6d19e8ed9c22ec2536f7afd1a49c9feca93a1d6206dd514fd9510e3cf0880d1937dc305e2c3b383162c386b1a3a75f58068ea9f91aed22d9ae649239686639f94309cde877faf455554004f96e7a1e9ae6f4127e7c96bca59809d66eda19f5f2cd764d469694e30abf12f9dd6b3a800d64606ed9125fd72a8b2206753edf6d0d80b553d7324e78416cc78eb9d380734b27a4e85e29fc0e1ca32bafe4580064b34a87b89a07aef1c4fb4cf962b4776a653b57fd4e34b8831d5fb6406d4763ef79978fb48992f7ac14f5e1541363dbc9766805045f4cb2e993d6a35d2e9db9b0092dfa0b5083ad3ecd0953596efc55d61fd3b386f634f010c9d1ab073a924951c379912c25ae57e070d724bb70a5721b1da1f1d22ca44afe6bb55b946b33734557375a2114bce83d41c1caa17038c8b411454ab66cc2238c6506b4e3bf2fc431103163cc83a8a4685da6b98bad5d9dbe390e11a1ab3e3b15903742fa227633e3ab05b17c87e4dad75897dd52b76820d0876b13aa124a8361f755c9ff42d322e9e1cb46e5d5a0647d46ad53785b8623b12bf0216b7cd83617fe763aa10ecc8fd41eb908ce15e964b4f054047d64b32584fde2e413ac99854a935e3841397d08de3a96ee95fe500d68ec0f7c5c9d282895a47111f728f636fe5c132aa5cf33195c9f199b102f78428b849ecb8276e761c4dbee4d1609880b131017f3f5da81a6da8b701d9084d388c7cd3d55128282e4ebecd43b83eb81422a0c1da2d2977fcff3ee6ac93de81a4fc64f8743ac9514d1a9c8a051aec14c6478ca5269d2ef3558d54551a0bc6e61fe05f2323504c3c863fae3e2fe817b14e31a5c9ead4fe92fb837a061269c9d1ad118682854b362e44b229725b4a12d7776f7a0c99ddb1f0163d993d917c792e98aab0e680cb31d9726a7aa1542ad38cc8f2c0d57d4ce5b75d1b136de1c7d948a0ca3e22da017bcb5edc22f30975dbdd107683c8fe52ebe51d2c93e2bd65febbd8807a31a5553e152f0f68dc9ba26bffd19c3a92175f766f445851abcddd5626b0bdf287319b7ff5b689da620669bdf216a4d292c7e07d57103cf0a1e758433f12a0f035b23f641083f77e63c7b06aedb1e8642e90621ee38bcc01ff411a26df082af91cd922dfe5f19b000a08989d5ad0d58898c185b4272bb2c5e660bad4503430b799e811d9355c042337675dd1ca826eabad0bd82968936f3deba7ceb5b7567e15772a068f74d695e45b6d3334078c423360861faa2996aee7b34833946b14569e81266aba01077f76b164f5bd0989a577faabc0377e73607db93fac988eeb3d2343448d5b0cbc2526f47c55bd0cfb22e2e5a5e4df330fbcd553d30c0a3039514dc1e08c269ac6d91f4040fd7f61b523cb8e8fefba96d42d2128487741e287a404c6267e6a3e457fb1b55c9d0386115498a1495e39947f50fe053682b2e5797ea1a76e452a7fc488aa4aa510f438f2e9791ddc8c63aae58c932f9bff90e00d67cbc095739b47681399d85f84929ddc8392f7943a2c07f82b66a9deec37ae9f44f06f97e4fe4545008c86bf633d5be35dd57917a6a1d6382c882b72d01d57263a7f34a15ae9fc942b0322844ec26d6cb0891ddd42e9eb731d767e9768b7276af3d0bc0f61c86f78849b437d0cc88348f921b395a706de5a6ca82919fd55a2ce5aeadc0962510e3e2290a4865ad170f8065cd76da69ec8ef2e2d4e49d939aee3cb8f79970076456b97aa80f218810d218c33b9d0f57d2cb8f13bf2af0f8bc906e5dbce4fcd7c6e9d61901e92addf29bb4f86adcce2af9b2228a84e208851b7507786f3b9b03c43d911f6004484c34fb01f50f96b8aab3756cfc10ee3640bc7a2bc243f531761a5c3b309a20dc199667a436d4e4d88361b15e57a399c3bd053a46ca8b63c63660846de958ed7ba21657d69876d05a25a0116988968c91da76d90f200305387acd5efcfc1f01d24cb57167aa282a235a3f6f33aa95bcbae8388fd94d509d730d528411cf2059085dbe94c9e3dd4256ee05f5c2a14ec9deae46c64b189994d04de4bac652875a23234637311284b82cc012e24dd361787575f25b2ea4d1121518d69b2d880ef5bbbecaae9da60bbb121a505a4cb18362c217cd6feda991dc9aefb1300d14531e7d562e4517ca3822043bac7af32795eb59550f368450c01697d41a113ea5b2e1fd0bb7ef1d057638c2294453f6d9bed06ec64b7a1c3abc2e9cffd963b35e8ecf1ed1992b4ee724b830673c6726042f4daedff365f099edeaca40e0ca6279c46af74116af8ab7517fac427fac55d1fdfd226a736a112d71858c0f7a3ac43c427ccf82c968d88cc04e6d8ec29d33c4ce8b7a8a6e349de2af24baa031f812c3b454283890b43ed0c35a843d168133ead65327a829d24581c079b67a8ff5036bc7288f6fea31ef195a7f48c6e616fd68e20b640fe3a6fb622c06c233d18761eee37ef0622fdd169b6a4e7d56bc1c848a95dd673fa6da4dceed1d399f32e1545454ee7f607e176d2e800d6607483d70cc19ab8b8364962e0f88514912115f8f9f25f03a2d1080759f8f18358a0159b5336bff11ab966126c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hf86664c75653cdff252cffd89128b1bbe7fc2d90221da076407d6d3e173b836954b63ada5998d5e0fdd34c42a8f45a9ebbdcbda6fbce7296e43063a1be2606174c99af7e2f47d30207f5d0532fd96bafb17d356e38fd4d30bc49f35d8c1b30326f596fae5fd3a04a016036767660e33fc6f301094bf965c26a0534afc958f12c5d5ffd4d3416718c8929295fef491a04025c3d470bb8bcc9958f3c65c087fcf140b1463822b9a809f7f06a951808b46d7af2fb4eb0c802b896ef236919ea071b75e22b9fbae2da9382493aee3e67a856fa186a84ba3dae2a2e9de83ac248fa24545e09e9c39940b2ef09aabdb1d2d5ff9a8a23cd41e4892998775fca7d5367ebdd52ece0096eb979abcea1c45657bb3c256bee0bdf9c79e291069e1086b7ec265fed748c7934282aeecc777343eb9366e98ea333ff135292e3501f6fec26dd74efe433ba19ce64a52ee8da48c16c8a158c26cf22491c18a7499181df01ed21cde6c8b5484269f9ad2e872c8cad729a43d430fabf277194323b53dd8488bbca45ab2b2b4d5976df0edc6eaef6a6e99fba41ee10aa35a1107747e63e8f38d49d955a874e2440bf5a03a6f375ce2d312328dbc2eff7a1212e01fe64776bcca3f169fcd55e78a6217640f18a29bea53efac57505384f4f2a0ac9e65abee34c539d55d842cc3e5ec386aac8a4be5e6916eefc001f64f703242557c2be4f61fd8758fd8b5aa65ffc35c0f4cd77b8cc6c38d639de1686f3c83a06faecb1d580cf72f95005b0070739f671760f011300b4ac21504b63190973bae500bf2eba4d14db678e2d3ae9c7556e8367179e281f8cd773a434cbead2fe620021dc6b4a16265dff5a3451008ec924eea7485571584005b66f4db56c5128910527825ffcaf27c7c64df58040e5565c8f85b1e5dcff00a5f96ea8867c7f73a24d856a00b74b94a05b413641233bfc876bffb9350df6faa03e20887560cd01d27e0bf497a211559f91a6d5a1d1ef362a6b87dcb3f882b57e11381a6aeb35b879589e5ede9b8a99f795a81c3d3196d37864b709fbc87d725b2e2da102c3e397f8914e03f9d892c309e7a8e301b3e8376bb44cb48bcc8d2626a81b1f168d2b1e10ed770c743885ee196493aff7f958ee3001e72d44c44a99954e87662ee99c884920d67edde8f80614b99a5f0a1746fb473fba8469858182976e47388237de1c4a78a4b1f3f4708d39684793630473b401b4794e995298c2f85f04b7236714643221b3dede5333f65c1626940100e8bb26e32407bae81aba3a9cf91626237c2c02cfbad50e60b989eaa4e00147ee79e510a9f6b0616b8265ae7e127bb498c04ef40b25f81210b67bd403efd77af3803bf0fbf25c95fb817a8a89cd77d68f8e8a3c920ca2cfe160e5895f53a2bd206b9882a6ce32c8ff56379a4d49d9bbba00202769b7f380f4d18f292f2caf2ba19c91acded4b2445653b60a8e63be0d619d9ed8a1e4fd844e4103780fa8aab038b3983a2c2ccc36c644ad37f3bef0052335a5c9ffc994ff3391b0641ffbe50de2041be2a272de741cc476ca97f62683956945593e34e36aa53e2e5d31b661b07d61bb6669861941a7129ce811bfde8c81a16e9efcc914234dcf8dbb48aff5be0c9f7c45d8c9fb12a36b325df964b95429ed3d5800c536170e669d2c973657773250568df2eefd764f783b4ee1ad39afd624e01acad388705afc8a001055b39fb96e2f125c3b0a2d6ec38acf51bc5b23537a35cc51e22e362a726a74d7ce4d870b60774be12604c3a9bddb9d6fa29572465d1e5f07144454d84db77c75841a5f1bfb79c0694ad395c8a8fc102b5704a6f7b04ac206f0f7cde47d2f00f6be41bfe2f29a557543b2bde99af9feeef8df67b39a232e8164f3b8dd2de76bafe44cff89217038cdce98ea0afb8508d392e1ab0df8f765583c8e98bfc0e09ada764c81396de4c6f2bb684355970c1525eb757ad983efb4e2cfb8291f1e9545b27b4127da87c5b0e8c5b59989fa7f7d40e44c99af6f5560481d1eaae88b2ce0b4b87e2535f4fd9dc01525cc62246ae3d17f9b5d76e8736719f064fce4230446f51831f74d0d4bbca59b7a1cc8de7b39df62739a77dfdddfe9d74d143f2def2a76e06490c1507e7153b0002691e366ed85334e343237e666001b61598aa2bb40031e0b609fb06a3dbe4a0f8d284c44f165d849137eec1a9c69002c07332bafe2fe856c93cde8c9eafca251114e5f2c5c349c4be01a3473de3c95cf9e22c3731b002afa2b040288710fe884d67adc94d3624cdc75229058fb752533ba6e176b5eada40f04431e50dbd70cc0a1663a91c9a0dd62845fd7e932bf280c7bf9fc875e786e5684979cc67b5f3b1c2f27054eb71a95e861121c309e7cb79065145133c34b46c1b8136a80f74801762d687b234e7f1651a30325a3f860f052cef00cfb93c2a4d9536e3849b4e86ddb80d3f5ff502ffce89fe2bff402ea3f091a04fdd8fdf7c7d68201b64841e1fffcaae07a555dd2340da5aee7bdc5f7dc8db45f88bc59b993602532d7ee0428cf6f309bf4d8cdc287bb67abd36ed73264f72b2bec56dcd5e3dd3e55551454767b51ce1f2abc56aaa76526f267646d4cd153afd797d5ee120284e9430cf83ba341b7fd7760c57cc28dad80a499c363dd4af01e1c2d07b687d258eba6b31bfc5d5fb03df85c8aa098b016216d0d6efef873a40564cf8cc3c8ab96d2c7c42ba8efdd58cbaf9a6395a1f0aa58077ed818b95730c6aebc0d6f445a74bedee29c68fd9fbf4fd3b1dcff99d87d12002782becaa26832698f022b22e425bed8083680df8607260d2718b153c4bbcdaf2470b49766aee7cb4ddb16dcedbd48dd901af888755811ec0d975da843db420361185189ab58b143f5556d19ae4b5f8f3f9a061c85d72154807bf89cf9c8a22627fafa1a253c58778405906b249bb2c226174cf369384bdba6ac639cd03619debbe5bb992041a2f4fe6ce76da95cc218b55b152da20e57fc27fc687c84531a3508d22b9fca34a8923b0e8e8103d89ad09316bb5b9c51c639822da04f26a451c9c0a72d4ffa9af8c1f9371b8d9a06f020764a636b9375d03791ea3c3fc436f58869e764897ae8c80143419f319d6d47e476f437bb0cbd00aee4f65896a83777b182fb5e019366ded9fb153b530e100a3909dfe14d829108c403dee7bc9f4076f19037e2e72861b2b8c7349200ac84b43152e221a8af7f1d6506371e588dfd849303ee1f6f08d0198c89f805dae2992ab30b2f05b8071b78084354d195e32cc8b7d88863813dccb5b6efff3a3bcb89d37f1d2cf489adce811148b91cf547b95775345236c62a29d7d332f8b2f21e6ea8a5df8d9c6b5daa783fe6875e6459e859f84f130e122c9d60256f8cd9bb7b7e09442e5cea1bda948c3804041c4acacd77ec137513d1592462e26c1d7dbf8761a1747bf0643eae1f6f918a35ab5dfa31ca78fe5cc26103a20f1818eaf2b21142a6d17e5fd6e00f5d268ea5efe88265caed01c989435250533ab2f78445d943502610a7ee479551657471586a5a2d6fc6cb8692e0da938286691a61ad6e30c6c1829036a67054c0d34819f04dcbc4659250e87098d039e0458ac205a094cdcafc6e02caf07e57c4dbe48cfe136b9948391ed2d1fe52a7d6b4605faba38771dd58f0b19c9dda18d7f0f6c390e41292a276df8de2e470e2aca4e2815b5c939cc12e231eb54b82a8fc53c8471eff9d9bb8e63959fea43a2fc78e692abbf02c2157bccf4315c6c68306bcac44ba29ded54416c4c4b99f273bf8254065a199401f05d4e0067d37bd1ec0eaf4e5eb42cb0c66d084346261819365f3d5780ed025f86d342dd3a7fe7d212ff08f16bbe0084fdfa695d864358ffa7d0df7d95dbeb8b0201f0fe4f743cedaa8cdfb23ea4f31f606dc4d0f10b0a9ed80a30e9a0d0e8f92b18cb8b4ecc7febfc6220b867ae7bd6fe5a810e3a9aa53e98ea320ee305d8dca69281947dd5d288d1ec825346bce8809d3b85109c5b2e95a3749d3bb834e96e0492a352ce1228aed7f2bee39f49ac1e1e1b50fae478f4d010781fd49205722eee1ceda86a30f81313beb950c6b6427c9570b5b5f53e452605487569d7e60166993d86b41c41463f7239926f595148a22d1022beb24871c42b045e74cf8ec6705a2229de5005a624fea1754728caf65ffe4358f42ec04558079a9c408eed91c2c55ef13b0d8b4b45606ad10ea0d799b23532984e7d2e3bb9720be2da90a120d01660d0834a34f9c0dddc6b104930cbaec43f7b609ffdd06ce7cfa9326121bbf35b7c2d53dce6ce33a78fb533f1aedc47f53dee5dc8500f1d44ac23b38cde5a6dea295ea3d632f18d665b47ead6cfbbda1fabd5da9cd7e045dc18c404e5e982b16afb2b2e5176a1f878b9535b5eb334f38a53d9aa322469ffacfb1c414c585d5b1a4c8a5655d8377bf1e19996dbccb1b978015404801842674ae21b3519ba39d49b474d8b793160a5b30bcd7c7ffec33dc675d24ed26a7ed8c7b179b93372b1b3638ab9e4de726656172d4357122ba93200f32e7d814547b6b829dbcccf20c9b55cbb43298322f14768a389d47957360017e9400419b91ed00e9a09ec57d7d3d0bee47a0c35ef442c77d3c2e95acda5497b79264a764c2b154f7986f7143b01706c559f70da3515ae8eed9d8945ed1bcff40f6df43758aff90320222b01d325fe6dc38d4ad4131b64ba4fc31152cf08dce2f59902124d4d601723a589cb6e0e25c3a4619687b7f2b3fec43a18e45486d73285d49b10232ce2927b0d211358522b8e30650f3db3fbc4d37f387a5432341e4130cfa8decc8778c263328375f964c6826d850592c1c5873b62fe7c2f35e626623e6546648310871ab1bd6887e7824fd90b9f5cb8012be3442613ad4d778231593a95743d382529461965b23d32da0d5c3710e448604d76a76ecbac0ec22a3d5d00ba5cff4377655d116ef25a6cc69f58fa288361fc15fc8712b8460b8ab4aa36d5ba1e5c5c38e253bc7b8a4d51fe78688b294c7a6ab0454c88b6b043ad77615e8ef418f7b21106ac6d81b230d58a320f78df6b0c7f6040cb6739d1a154e8e9f61ad77309c804dce5e40d5b8654477d9ae3f3600110e7f4476ab8eb45b23d66d8935a07a64824fe506bbe83269816f34b5dfeaa0471db1458557288d1b33574c36219e64c613f8545f457693cf2a4e888bd51c2d264fa23bac1f339b8ea7dc4c5a4722d87baabfcdb2e839434161de444a82531e6414a2e0aadcb5f511a5fad6c8603a2f55c855e71d3d056e801a6316943ac7756325324fa6905a3901272f1671fea2b4bbcacd8115d0c1085fb404be4f601517d9aff858a386713e4ad0021ad585e914b49a3e9291f3cd7c547d0c8f0574bdcb3de4773c7e2f9e6171c12b174c987defd6c57f3fac946c3264bedb56541420ac9214727bac980d1ae63cfb06199f9856d2b6019790a49f09050d7f1dc3f25b78559ce419a8e89de7e59c773e72;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'ha3acd8041c4a4e1817720b050783f3e882066928f92867fe5172ebb2724285a0b72d7355c94f3496899ef6f78d2efc1d3e529c15691830b20434b07e588f27ffd579c34e1e2637d5f82712fb2ba53414e384a31c3d541fe1d14c49bac98c6df6cf09e2d2889ff965d079228fb1e4c10e98aa5b5724d235d540c52d866ec3012dff6ea8def38239d28c0465016faa54da025926e82850f3a8c3358bd6991e399cb1f253d3f2bd20e454249394e95f10536c623b523ac586401df088e6604a906414171df79639a23702e5dbc34031c4123655a0b8977f9c37cc0059e5ad96b0db49ce7617e25dfb941b9bc453cd9859aed74dbca14d36cbecc02068242440948911b3d4ee2aecc21cf3627dce3a7d355a5af8afc7403cb5c84c418dac801c428a622b5f002576ba71f9c3dff56d507bb95b658c1c17e2400978b27bf75f4d19295ad9768a72b1359ea8a62db4dd23e9616886f8303c74fbb3d36fbaa790742c8a63fd5b7162c60491183548fd44685d60d0fda736d0d749b211f8c198a2834a9e23334d9ac18ab4f731136794b03d99c612e6b8174c55cde14b5205ecfd80bbd31ddc22914d28a1ac800e20e3938cf24135a65842f63c41549c129c0c6f32abec180fe81e8247097422617ebc07a13e19b5ef836c6b732a3b36a9ed6936807c804bf48537d05906015e7c2d09a4143b4d68ac5dcb1d39ea1bf6e4e9d978e4ae56fa63461e84576e6883c90d9826465b9924b02a0b0919869c4fa5d75e00ad6fc57b06a9986750edb54679ca2e53298beeacd527d017ec3eb7831864e1920ca6a95b86d5b7e506b6beabd4b79f584676a6c867629273bad4e57b0847ab6a7e43eb2febfb3d70f87d592a5b8cd00127582fa095766800cfb8ab0162fa2d7b35641a74f25c8b9df5258e1c849dc6bd84a12890f0d7063ccbf7b398a6ea2e815743fec10f2b33ec91cec9143d6b85ae3219359f55516c2c67e7d6646f89e3325ea1b023ef542dafa031b95598633c99a6040d8b8643202b01391c3fe85258b921c482aff281ab3089b013bb888ae3d609a93fabcaac55deb27608945a358acabff03d693b08d694d8eb58be73c788d87993981377c90a902e90c737834f094ad338e6b8f2480ecab1bc1864f5b4e2c83dfb6d4f5e17b8e2f6f52f56552000586ee1407557f9f212aa8e6e236f7867d7678c1fc5c0b327cc7de787c5c7ea218183c9ff4a6a1590cfba5452a42116ff8afe8ea36815d71640915cc18e297c39b9c57cf5c46fff7652d617caa4e7251c2dacff958750621929378a5f3f28d80451a2e2ed5349237a15ee6f36b3d7d6326aab307bcdfa05d003dd3f53eacc38b90cc3a63c71229cea7351d1ffdd0208d3f2856a7f157bc553fb213c4d5c86c3cf1e62fc9dec99a0f34a7205d8f72e04f81708ece2c2d212e960a3b86ac141992b759bd357f4e9a1a442259a6211cb7064c944c0e3c3201e660511438c1a4af8e17a8966f5809bc8af7325b4ce3b514d429d17094e4c860037c675ab6c90c94aba2ebb91fa7427d344151ee9c2364f3b0ebf50687770b2a879a559eb55a882a4f33383cfcd7e2aeb221d613724b2b7eea812d1122ec9248f9c582fcbfd4efb361f82f5bfa3086429efa778018d437a800fc56e9241413fdd9a6bcd387fe8368f579fdbd9f0f04d875feef4d701ba32d01082fea3c6fb9f0d28396b46cd83bd029bbed4481a8cd0f19732a70e0ab0cb310dbd559f9b6ae2734b7e1d98723268e40a91ad73107eb84aa7a0578fb211d742cdf81625055f17f0f915362a6b08386346d900abc7f89ac686af9fbd2a0649b15c080963381de855a09e3ab2f52b0929e9cb17c0ae938a0238123152203e5ac2c637bcc88c1a1703d4a96af419bc8a7054e3bfe225a510457621506ee6c60c869c29f725f02c0f3b1eccb008b40c78124f0932ff01048b7b4b76838497911f37b34881b9734fed63f65c615b0adb0feb284f5c5b0f73450d92b8ed4cc72c0f5105dd89c38cf44a7df99f93aceccedf84989278ba3722c6a09d8f3d04947a8be33a454d507eb8bc6f181e97f22a0f25190d0ab5c83ec4ada2ede4b26e323af088e8f03938e851dde8275f6e1562a15856475425a6e459a83b4bdd6db0d63d9d75e2eac7cd26c5c4fcbf3d5309fe01ce6b0e9fdf735b09679fa6625ff607b6ee9a4db3f952a65451a457523698d194082d19ae57d3b093e3026d207b900bab7d5b51088c1af2c25e521586478e575c3abd7c1ae63a0c08e4af2be0747620aaabb04912276e0c4e28f93f21ad2ec595d10fab9b67240ab0779b8aa37ea8dea6eb8196d6b210abf8a7bb2dcaa1ca4c282391027af03996dce1da4824500c6e13b1f6eb9aea485dafe3adbd398c792913a73e94f9bca777a69b08a29a4fef213c25aa888cf31ec80a50ba16aaaaaf52bd0f4f8788b099e144c5dcd99ba2b968d3702d380a3d23805aa6515979996e3406abcf52fad9568c1ebe424a23f7358b3ced54ae82e6fc3481b33e7774163238d1b5c75d3584c67f11688b8ef7fa1b4726fec50a535bea00c954316ddf81a198baa4443a68168e06d274895a207720fb953c96ec04f2139f05628d6d280d0ed01a0f6f809c7a3c279df7eb1624e8532850fef5ed38cf6cec6aeb5aca6431a57c82cc0c8ccea523ad1794fdf3eb8e872ceb47a0bc23bf1aac55f6e890dc0abc0d296454ae90fa205dbad5de92799907665415c803e0d1c760638e3c2f43a5961b737b6f662e915da03ada958a25c0cf0e8868b77cf676153fc5c11864085e49879631424d606afed9b8589758f2f8b3ee3e31d460c5d5d12caf97d4daec232c5cec250745a6726298b4ec826384494d115f75096a32ffb018e8c5072e15dcde0038e2b57911692e698c91ef95fdd8b1fea9683bf70e99c17a4772a5db7cf333a5c09a4ec5912964bfc3326fef90eba18b5dc8f1061b2acb1c975473009d290c5bc55ad358ecb000af5d850a05b6eefe61b7019bbb6f79036aa1ad4a23e0bf8fce508cbd6994487657764aa6193fcb972217a74f20bb3bd9a7b740c4159fcfda21550afb15d18e1966e78d799b0195fad0fb5f1e57e8cc9d07f47e060b1a97a39634285841b19e7506425870053dc459ec25f8983b7c031399d4ea07a6c81528041d94be038fdbc46dc3c50c4c46897b2f7012666659bd3acb75a159582c6bda635d9280cb4d1203e07d152fa9e3ba0ae9b65f35f1302d854c2802fa6e02e12ae99eca577d808a6218e19d57203c2c3b05fddc61d4b70b50b6aa31e25b544761702ac34f8d1c3e1f4b1b8fe76ac1b6afef1465865d3390e2a2936a246e2cf59c116b954fe9a297f42b126f124f2a54b53e8908e641f3585265031984f96e8650bd07ff05f23504847dfe7c1badc90b5539a5c637b2af15cd6bb6a2d3e6df6067e31c9d37357c9724098f4c6548eb85cebc45d92a329a98f876b985c982bfdbc1d21237c9a06c41558f05c41bc439c7a338580be915bf32738084009cb998e832b2b247e709fe73c5ad994113cdd45163823397e6fbb5217b917baadad29cff2ff8af7ffca36ef63823df23df8c9b10a33ef17abdf55c2d10021ff062c2f7f29d4ccb7786d100878b3c4b4b2370e7aa9604a0a56f8e17175f266a5bedd59c77b8d536c501ee0532412ce6755022f8a4631d660299986bb85765e889815db7e91bc3fbbae8794df2eb9387df8d5dddd5957730c4cea4278f7fa2a006bbea70cb419835467ccb2e8a086b1b49a27b995d159c35836f6b396a03f4773b4b245ed52998bce139ee27ad05dbbe9dc36cbfa4e49a661d868f8b6f9dc85109add1bf5e83642adc8240e8b74643a09407897eaee2acc3f924be3bdf29bddb47037f1d0e1c3c487c400e5e710b3e770706b7f76060ec22aa6d87cacc47cc569f40237aad99b82c6ec1abc52dcbad3d416d170684221752f1eb1cddeec4bc252375ec3952b825616b1dc3ba4b7d763366ccdaa49c22e4e7990e87c86d324e289c097a493979eb6f8c2c3c497f4a50eccfd50b5a740731bdc6479459a081743e5da6d902500dc2b1721aaf74eb5e70e95f5d48e2a9eefcc9989e309e9198bc2d76b212d396274c0ad191e0fc969c3c307e3362cb5fac101cfaa7040b001f90b03307cd2f3869a99d01f12d091672f7823b886d901d646cd061aa4bef13a4633a5972997c741c740a4e173b1f12677738d1f392f9f930e458e1aa7e63b83e1f6d7892e04d9c85cdc49c6fe641dd602680cbce0d3b8320a5b1622684b2bbdd333798a60a49ba5e2463f82d80cda3af8082087b3d5a8192cdf41dd6c765308432e04a8015977fd93f56f267c13acc52c07bffb1b27c1410b081dddc2899f782305da894ac1f8f5a2b8476177e8cab1e996a816a736c0df2dbf17cc1e8d2f3236d50a6bd66d3191f1f54732edf92ec3065ed8e8f10aebe3d58fe1f61a2bdd0a2cbc8559ebc45fcab5b8e23c5d1923161dd0955c70a0e0eaa89d3282dce8e6abf03ca3d8b261f049858ee8e94aa9a26992f9bc6442a3f7a5eb7ba6004ee09a0d64c53c0b4750aeb9afc56d672795e8559806a1bbaff5f21ac9055c2291eaac960a86b24f072b3b5863206bc718539480dac124f5cd69ff543c024674defcd5cd14892c4a43298a0888d6e3b572814e713a693f47a91dc0cc4cc0db09133fcfbe2fbcc8f2ac4720fd9a91d2082a4949d06f6b0fae545d8a2dd75bcb2fbd1398f3338741bc6fc65e094a6e5f35768a02cff9782a0f0675c879f278929d78058aa93b1c88466d1e77fa2d8eb44d421bbd67483f6c6febe8e11cebff0c9e96929700cd36995535dad97fdb426ddc2e8472bb3cf07d6d6972176876626fd3f898ce66b96adab87750ee3c81af6706ea1f43700f7d4eff48d7a4219c4d572a11f63c65271eb2ebffe8aa051ea6d91d226df1fb6eb37e5f1abc2d20fdfc32f0c65af2a5d376adb38ee02a8f84fb68eb84c43a97e6da546b58dd25a52ccd0d65f3285fb193902d7435da94fb05aa877417f83f268b922acfa9eee0c298fd5026cd4458ac85af85321792fa87349e1ff609d6577366687ebdf9d12936d253404915e7925316a4bc013c7905052a7a0106aa2d3742f428a9edbe058c4565472dd1c80ee8df66fde49b50f0b4c9e13555a58a2a772b21afea63493627b280eb9d68f94aa69105b6114c81b67b370a830d32dc302031426afbdb6bc77bfbf74e0fa0951a7027158f4bd865b9ac96f6fe64c29282b366e718f1dea02eb87b5dc24b2baa50036c7610a63637702c1c323f352b5b082c067632c38f5ca010f1c160f3859f25a58587663ebff5508974cdf1efe9da2fa5f722d9a6b24a9057453a7ab11d0b479c551144aed11ea53fc4d12fb47b11f3bf099fb8c75b86e9b1b59e58853380dec105702b13113b06c4b68f748d098f69daf57d54980d5645a0fdbddfa0e0f5567d661066afd1fc5d44142af30960ee1d6d49a7b7a1976a6bf0c7d08fb7c72756a3ccde1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h7f2ec5b1e6b997db46d0dd2dc663b924ee9ea8483a036c7420b7815e83fa097eb202846748729b4e3b37c133f9f5f7d9303e145d2b3490ab98d8be6a39272303fa3dbce755dc03f3bc7b63dc8329d978a4130441b792f1491eea08c03bb7c742472293a1e9f0650fed0ea52f0a796fb2c58c4b56c29bf5f1abdf1fec40bae60172e379986caa3582256c38437a06cabd0af59ff3919d63a92c456b3abcbc502c96b78288a5888b271da58fdb911caffdca9674c65bfb18358c1802d12574f4d44cabcc24325a92e1899f70cc6451a8199f3ec4de2671965f9a8c3ef4467156b0846519409192ae7b78dcaa763ad93fc7ac22b6a29386ac704bd50276c7b8bb6f2df4c1e1bbb7587648b0f50a03ea120cad5930be03c8ba81ccc33f9c356452a68ace654e05cd17cf1b53bd9fa55fe879513d6f140a7e5a0c9223a3bf4d742be4a4c3d0fbcdadad8d33f1ad4df76a818436e9ceaecc00277c5735c5c9065d0a7fa788659abfbb5b047d1fcf41aa6bb2f67ed9a06c165204bc033fa723c37db51d452dc1729fd5ca53dbe195c4521012c30bfdf6bd9e3c5a0cc9c4d65cbb2ce427a546467973340c9d25ee1caf8e6e6ec72b536c0c128a120d787d2d1f46f336b56e509ca180e9e226691becc5cc52b7c1ad08a7e90696f53f6f842f8896027d5ceab80b4cd4defdd33c8c2abe3678b4b4de0663725070f1f5a416de74123bcbbc0ce4b3e7766a4b11bf7e885e51fbf721423aff46a6b671646ee75b4b1e472eaa305c02c4631c462bb148d5ca7cf87acac45972cf30df8714fa0b20c4a096095fdd53805f43f7bed9813893b2b70545c635b2910803ec6b6efd4010a1374c3afc01b2f65f67551881632b0648c8359d754c62f32d500b9424bab05b5a1f796537799586276c7b269c4b6f004ae7544f78dc10f3735bc7c6fe7f571cc3892a28f7679b574bfb862a9fb8827f2851d4a14d6df41b916d59b2dc09bd90ff21f6576023d76d78c229d1eb94abeeeeada1064bac065554e0302d182b6f6d6523c7ccfa89deaad6e5ba4c0f9d3885113e26fc6a89887daed1ea5eeda0bfcf8caac0d3feff1f91a83b5b7c1936b3fd6d53673c30899a12b04d38c1d2adb6bae195011afc7d3791962a7abd6409c85de1ccf8ae5e022d8c970aaccd254746d6ccf53aa719cbe3a54666ed9db0831557da313d99d0111614f6eee416f369324231dd5321f86d37f5c1f117e4da8c170510d4ff480d267152e79a2fb6ab9f612b6f3e34e2bc4c3aadecd8533e40493f212bb26f0098ef22b3b147fdef84db0ccff7876aa816682fe8e64d3ea93a4e6ab684fae44768df67b76582a72ff765df23db24d83d3a4cf9764825edcaee454a37c2597b50a29399af16b16ab944b63d21fc95c64d8f7bdb4306043ff7f4489c24d95f1867d6ff965b62135dc15ebb4ef30c9eb0fd3b8e1df81f86ea9806bc0ee7fedd5631ca990279cb15077c4d2c93806ec19ceb4d9c6af0623be6352420d4963bf857712e2e0d46c7b8edd52d7e574d53780de79f9409c57e28edca9d9488f359d67ebe2dd59feb918d9a76b640fcd54f79090a064965eabbeb4da1d1aec81bcca5d83ddc584c6308e01807d5cccb0c95a34cb476972a9f05e44148d77e5564c0b866e8d4c521f2511267cf3ba23ab1238e970021b71de0224faf4618a938772949634271d9c157ededb995c22e695962d55ba458baff3a7fa67534a132c8e76e3188b14515f6add787d313fc74a8b561293843ad26d8df13a41dc8f209bb86316e57fdd76ec593a546bce0c266bd4c2a2bb3a8a24d4fd1669201eeb5fc18c9bdf9cdffdf2af86a59421d2b6a5860aad12c8dd95d23c26529b1a2e8cd336fa07d40038fa20f5e34ae52bd3f007f22424fbdc2758baefc81dd185f56459c0635a520d9d69e95c9edc4a3aee7e7b57e46739daa57f6a0acc77a5421ce198541ec58843213ba715ae4c54a112db98dabf61e6c0d0fa90a5c5363b152ba658b90a806c769ca95e92456c92239babbc6327a7582dcda5b09e008274a58a576539b1435c57cb7d69df1a3ab67420b6accc25dc4cb891765b31b303ac90e7c15c062788053961e0eff029115d168f6b53bf27e8b7950b68adcb39e0eb36662b8a438559e145c9f9cb0de42712fb6dfb169ccfe44a3dfbe415b1ae27c7d55e14597cff4724d2d7d3747d9c9a469af4050f96077fa5bcde73c2b8a2c5d0afa19ed434a4b93eb9a74671942e5a6176b7b6a4c3a47201f45804e643e3f7401b856527bb6107ea036b91e93234ddf8d28fac924c8d6099290286783aececc38be86781a7e60b5c41a4d6a405df9e1c3061337931631675107b043e6db3903a0b55c260561657dc2e41c381c292def3c7cdbe243abb3bec840e5a86f4bff4e7577f4af95fba0012dc40fa52cd6f2f4a8ed0548b7dfa69b9b02846fddcffea7b9967a5d6493bf5b741605c80658720674a2432037378ac268c5b5cabb46d244d89e8166f00da6a4fafd074b10a06d30a0397701278c0bbf06b257dd400b8d535adaf3d19e64522c0d19db430b2ebaf8a3fafb7cbf04c117eb7040cafedd3802423fb8ab67736fda020ccc4eb93b4c321bdddcf0a3c540a427186ad1b6a931bb99bd4d336b2e37e41f3bce0427ad7570eba405ba790f0efb93b90e9abbbbc64759964466b4821c8f94ed828949acb7d90f6a25a6043b34e5267bbf0368c7b2ea3a092e7d94769a64511c1b8d99e1c405feeaf2b09ca717c8a8fd9a1c5cca8b1985cf6d133a2a7019736c2c9c2c42e721045ef09279574a5d1604356a6eb71a72e554c820981bf148d5cbf7a2b3cc70810b94940dedff80e2473b228ac08fec8fe82509fb002f0ac91ddb0bbb5b4729d8643cdb387568be054ff8fdfc1c6dcd8f4af57a5ca5470ce67c6418b1a3535aacf689e182e6bca89f8e3261140051adf14cab941fef56b892bbf292fbc82940d53e311a80bcf299e5fb7ff47ac2e7764f4a434e9d559dea71af11caa0bd16f6e997308c4c9b0104b49df1a0b6931e76e0f1d75e9c7cb930551fa5aa37613faec1e666597a8cb42a0e825e7d52f0877d4c585013b867ef9a624777030df1dde4b295700bc29ba8e0147fc4cb26b2e941128d4e58005818bb2e588cace0ee8be71d33fa1833572300c7595c972b513731f1ae080e49a2f8ceccfebeaa1b93acd68921300b1a1ec0768ce6f70115da45dc844ddb2e9a9577864c388d2ed6014c45be022389353860813b32498c5cb8ce4017da24824a80fa50918f4b610ae92b557f17be36d05ad2ac21cfc98c4c6cbea9821acbc784d7458856b03cbd510ca75babd4ade93162c7b64202087565c3271ad4d2d57000001f28aedffe81faf564247830308163ca091d33609ed0466d06666dea4ae66d3f72cf6a883cd16c316c9c085ce2285607979d5efed382e99c787b4c27cac7073ad2d61b8800f5ba43815021ff39b5b91d95ad8e8f3d42d0e459ed49596a29ef2bc145da139d645620d687645a2498243ef699044b7b072c38a92921dccfd3e4675511d68a3ab5c870d5a58661307c40768cfd0d8c8fb34fec34c2d13b212f8800de8db508f600005c589a25cbb6ccfe9884eb140ac91b1b35282430e79831cc542adc9bc720813fd9a88ec326bc983f91b30bcec2892d50f64bd9696bc1afa85ccd0554d1acb43c2a711f11f24a65cf201ea7227373833032a24d6f6f31f8f7b58b829d3f318096c7ada28771e33a06726d57817048b5bcfeff603c30a04b60c92c9ba07b7a793330f481c1ac4b1871286dccec60156a6e68adf9bb4cc0e647b6f23cc7bb2c7272b2cc43702053df3fcba3edde639c3201097e9f44d09bb183a122e7e4d9f5dcf1b6261335f3ffdde584fb1217e707937020ec822c766da78084988f83d5174e0f17dc785a57b11f4154f4880dfaa9a2904cfc5cfc76a5367461c88ecd606d1d3005944a4293639bceab5e0e8fc1793295a3696f51587e6b7e7740a4fa196160b6d52de9f9d6e027db365b21f83b66033fdbd73588bf0fe5879b75d48e7467d5a3f1e723c22263e93909917e854310226f89389a5eab694af963dfe76a463f06656e15022294478f93bafca8aa34420596923cc3dd904ca364df064df671d4c7334af241b44b66867d28b52be5a2ce8289e74e860685733a51f2f19a4e34f34652d90d29c67cd4dad6ff93c44c7fe32a43b64dddef942ab0cbd96bd774852d1b6b4016822c045fe005781245a4368a8b01e572c64a4d7deb2461b1eba13f7f66840119547975ee82cd7133c48f6f1f51738fe24f9da190bfb24c8366b23e7dfab1b04358aed30a846328ca3b776caf80eb7c6a6f79d1024566804903606009a8651a3db060508b24902566a5a6e1a45998a3d787c27192304a8f8b1d6fe3dcd6706fbd09c4676e8f0425a664aad21be2fa3d2114e808ce39e6cf92c6fad82586eb9dff7a9e1a6d94024e8c485b19f94db4b1b14b7c32aaebda1418b63905a5fc0e110b6aa05713349ced6971d4ddb944d38de0228769639e44a3ffd44e82b9349136282bff00fcd57f1834805ca5618943f1fe754218464f5038226099e38666efc0a7a57e7a4991c2a17e9a9a111e8809d1faaeab32111fefa355062e2adfaeeadd65384a0d0beaadb6471b96ed79a4c16e355f69bddd4d25c1b177e63a4f03e6a66b1cbc8d86c7b93c8d3ce19f2dcaac7581e956852b8377fe148a24e4df0fa7182c9d27c131d63439379dda35dddb06d53a36d269d591d3fadcaa6bcf9c23f35e3b9ffe6c471830bea19e210807cf5d78499ddc994e668c31f0bbc5d3bc58a30f88596d2126ba699efe7138c1c50f2231c735e278867992eba5faf2de51db4337358340aad479d4cc2ea24d691a98ac3bab7af6c65e419076bcf1a6e086983a8354e8bb62b5b7dfb8ff2e8ecd5f85d360aa773958beb52b966bb67fa7d5974050029ca491ebfe3ad8e617e52ca2929fa9c6dc7288b939d339c8180f20877ff0f7ca372ef504fa87fb322f2cb900382d7be63ab3c6aee53c7535fbb9e6b8e97110bedbae9e1230f121bde4d843f8fda64917fb6c9baab44d2f5ba39b6ed811c13390058ea362244ea35a975bf4877efeabafe97ce90517d3113279b5ffe5904a0cba49b3b92ac2473a356ea9af2bb2048fea1f05f5bae1972fcbbe9a170064d1cb3d5e52229dce05cb71305a6ffc1abaa1832d2bc03b284a221735e4c7515fa4759397d04e371c74890385e27d5e370cd7744fee69acc6520b228c7d1b2a388bcf6458066a0a4e54c89d040488b34cc9d9de6300b8935f5ca233174e48148bb47da01cfa8af148fd15fd76c2ac4688c81bf8d39f2c011acbc09c6c83b4fa164d359b03ffcd0726f4d1bbfbd14b20c56e0a5c28a37b32e609826a7fd3fe56b18c6265f4ac3e38b797288d7ab0d705fb7e1620127a87c99305b1f08047d9e4afd79a999687aea92539acd0e63dd7570a9d59c3d3880650b97fc6f63805db9a1fdd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h1e34d11719720916901d04768a39248ff36ee0c2ad04647a856c20583677113f5a62f092de6be2cd5376f12708b3953573490f4c895b28c43af13a933ac9747cbaa0940d18e75be458ead1f7eec7254870637cf2f7790a6f16066504083c133cb5d4f7df8ee13262af78b70a28826e62df7e91ed44a6588d8ace446054f8802edf251fd15b9a1489b391ac860d82d81058ca19865956198e8da50e053a20ae0fe1a288487b611bf16c82877f1d746bdaede57230c635d839a1d06c1a70ac4c16508562d6beb4955ee99a76ad453b64abb206cfe8e4eb8840cd6ba1a70520af8ed7ca32049be2bd645f40060906eed99c5fbad452ddb78bb48aef42aa718faa77dcec1a6a978b3505fdf8f4dc19dddf24a943eb7c1d6231cd95a15475115627b43f5368303092653633ad9d1feb06fc71cb118d9c1bcbc2d752a23f4f16cb091272199d9cfb8238e136c5c9b76c672259c85beb94f923aa150031215a198d4d76840851087f01528a3bee50fd1b67aa0cdb359edc1ac9d2b08176b70a019bd054c85bc9387a0a7260e0cc72f10640e6b414e4af0b727cdc07a24562773182e717da5e60a5b72047ece7ad7aa263e1c31d2aa7579bf955d9f623880858fe5640db0bfcc4e4048e86ae7e4cc37aa5619a55b845242799d73d2b3b78cb83ffc333291e069ec56bd0f45646c2498aa01ce83dd5c1309b1220b8eaa56c3efdc94aca607f94f06cf43ed5f4b96acbcb8d8363f46e89675a9620fadfea2a291b73568db4d76a0e2d5f358d171c7ac9a691ec8ca2a671dff46fdbc041c0bdee5f4230b77bd62aeebb584b3b32a34060701ea01fa60cbe5ffe4a8e59f7748a3103a231877daa3927d3461432a993c5a5830d9fccab12d1d654acb840eb6fbb2f79d249c1b837e13baff22dcaf870d4847aebd045986303510904779f2df520db72ca5625b84ff3c226d7edd8f06f1dca8a98d43f60058a82dbc8c53361b4e68f4deced7fc94548d6442e7accdabfbc2076ea4647c80bf10b86f454a9a2829f387e5343b3e170f69e7353fb48e5d61ea91435448afa61c0afdc86f99861cae46a63d42af0c7a329000fd792692c7919a0e525cbc5381eb2aa9e346dcb3f7352e0d0c60422078ceb8cec31768244628b7cde54e1f7000b6a2e4f8097c26d84a4826b6fd4ac0529e791206df734d1bb64c08437a01e2d7c59e8e1220794d076e04b91dab50ef04990436b2688ed2fb79b43359c8dff21877b63d4d41f71c4392c56c87a3244a5370736838325e3cd09d7e671e4a65e3d033c4ac421c4cb0fb1c206812d74a34b84125a8ee2e1c932344a22d59198d0c501a7f0ec471c9bef41a0d7fc9681c5b8ec5f53bcfd2dd912799f8da1572847cbed756bd37347aac055cb371a7a6bc52375bd457f2a71c7b69b52b9a297d22fba261cdce76c89f7b3cc914974912765cec9ce9fff3d60e40148e56f88b194a660d491c9fd90ef721aade210f12a2bcf6cffe213a69742670d23324eceb20513a8b150bf3dc22fb904b73f7f33c12c1dc23572a3cadf056fabe804ab968a64ef174934491bf9a8984948d45433f42a76691c38e97f0ededde2e2697941d5b7f76eac301298521edd6389edb829c7471c36758eea80cfe4ac2401edaa0cf2b0bbf3a94d4c2bacbb79e634472108fff1e5551e835734cee52c321a614a2377974b82df86ef070e0c5eb838bbe608b97bd8c5eb56ed57ef2cf8e57c8480e652a93550cc045f289eb572170c112b6dcf58ff8c8e7fbd95575c30543963648899d0b6ed787618fe8b1e8239ccf4b4c3e0f5a3acec792e8fbd2a1a480c69952eca7608daa3fc8b0dea94b96a749de5bd07de060d818816ffc3664b165be0ab7e516881ac248ea36e14cb2f37c916f7a713861002b511c1eb1feb046821f5618c8db2813b6aed5fa7310bf616e6836ce4761ed14e3a6d8e52d504f047648a58cc24688b0827b5a0ef9ca7651ffe8b81528938c7f82ca411e40189d77953361f6650cc1e2c174ab4eb72fc30289e66a2b5bf4fc74a04b36f706e65b7ca02b803f58fcc6758a677a0f2bfddc89a4a43d145910a8ec14e90f258659f5d7b9f47ea10ed6720f5e0d8e070e015cec52fabd3d1162b380f3d6c17ab6a8c6340db8cdc253c7d4d9caef1a05de75e1f9a7271addf0c6469b62acb1356c4bccac7911c537fd3b459a3a408246a30e63a2bca7e09463abc65ee18c71bbb13fcc80ababc04fdf81e7b7729d1f099d873492f3d123d1c243a28aaf7476777e968e0281999d2ded30cc6a1684b034d39ed2a9ce0c501a37da3a373725ee9a2ca7c19002cc7d1d098857992e67ebe5ba36377ffd87ad3fa5da49617617d61bcf5764496dd844695c7b6e33b05cd4ecb275dc38bc8b4affa6e43313a865c88f6394adb54259017a3a54e30281701deaf02b5e8b88f19401ee3ce181ae5cea394506901a748c260eaab2827fe2f4ee3b638598a06a34a1a0e31ba016dd4cae2e5e23a8f352c5babcc20013f38affe63efb622461b0b272d71dbb62258152e02a1fbb7ace8b2fc2dd966bc6dc4b10a4d8ed0b3dc272ff5a1ab736a651b98d22c1f3e5ce8296e500312c522eb8870e2d8f4950defe71b155f52b50c114266aef1de35bff9de253ffd229a8306af9686660dea7544e36f437df73338c882f93afdd66f1d0742c1b20ea79e41fe9146c6fd411071de2cdec0790f16c76000421b48c6817b1586525a47a8326f46bfba9fc388b170ee252904929e16bfbc8de1319a98ac103a64d63d177a6eafe06d974a24867e402a639f472c9b4eab3d0e505fff7965fbfa854da66d3db07fa225bb892fd4056bdb78419c409b6dd95d1dae8824721d3e75e2fd009053fa2d90f078b15ed02006b464f7be3dc656d0d51ac5ba9d05d4d569c0d6579eaae2509726fa2a4c9695c088bd1aea11f58f33ffd538060c7f508e29edad07533ec59aededc2eda48d988a26bcab443ae2b1046938b505a2d1607503b6c49529541fc2020d92adb0571756b5e5c9dc7e8a05f1bc4d8826d61ce54e2f9b135048289b8635005300fb5f46db87e43131068bf0f0ba2a05151ba3281f31ae115377b48770549b9daf29015b037aa5b65dbe37e226b7d26ec8535e6e2d1419439d5f22f8d7d5287003974c0a9c1532408f9de20125c62a64892d7776cc76a85a2d0f1cf300abad216273ab43159091b8c3c09c2b6193a95f57da42112a16b36c721b8de414d0c0cfa785b1e42ef0795792a4158eab03fa039742b8eb2b8027c62c7a7a9f248c63348af1c009428168a063815f7ee3cfbe9d1f4f7b8d293d6efb2f3a73eb5f45c7e6ea0e17e883f12ba32b498dce9067451f9fc93b55be379b6bdfa6633a845f406628e653acd5f6d9c35fb9dcb99e6687ecd8c5ae23e7e38b7060b41d585ed8f26585cfd1e672b07b0c287b03166c1f7ae71e66c96d6c3955b586030dd6d63d21a8d6a539d448f2a67d0ac859537b69cde319a5b80cd20877d8c326055e4e5f661d1d431904c4680cf700fb632eec81b458af3e3b03fa2e72ba25e4fbcf2933c7e4d861d55ae7feab596df282ad682708d2bead0b4fa21e4c2beaa2e030b369202ee4764a98ebf05704c1db20b7963fbea60583342a81520b4eec7b18eb44fce58d6cdd19fab22d60ccae8d33304d4ddbbda11c9d74523c1fd6701b3915e09801b2b9ccfea6a0dbafb33cbf1f3468b3b2ea6175759b9c2a72c28aebc2c1d1f6d0c13f15d794cda8c3bad1e2be6c978c370f800c73200ef3222a7c8de812016e92427fdfc86efe2336daf87cf9ea88d6c267069819ce090e52a56c2d1c8d7779492f2c3eddec8569e3239c2cce233ff2a4477e3e5dc8c658d9ffc64a1bdbf652d9decbf854d5d861fd95a59d3d7fd74168e291ad089e3e1cc9e05f980213035158c4c11f21df491b6c145481a12c2a6b0c22eef8c1df6e8656c7eb9d44c9e181edf7b839a05306ef40884de75c0941a390efd7a4b602fd9b469cd7cff5d7f9a5dca7dd8dcb2ba93153ed6c3950b0b49d990562bf8b15d90007636f869eafa0cc696e14e8b09e49b2b912f28a31c320380931f982dfd0da4cbe1507e3afe05dab87b94d4359334da413ee00e7e358da322c6b36100c66a083b187dffd6bdfc2f55292d43a2cd97d7b1c8f9c35182a53e99e5db0e05db1913b0d67ca7ff21eda92da780059bc3b81b6c4705435fa67791ee0f5ce123387d61dede5e36dffda0f2f3952a372f64ce0c8d08845dca2b5d774d817fa74fb3e3f9f02c283035177aeb73a757e975afaa9832e5e746afaabd3ef5fe0b34d556c497a2a1e62d9015adba7733428b29c5cae28e0929cc2cbd3e0cfd14101988c95285a18a397198f925ab6bf1794022cc9bd38799f4b7dafc56517f6f89045ada18ddd9cc636c793ef9580fad716700636c5684f880e573413d14854fce5520f467af737457fcaa7dc42fa81fac8e054c4a14c24bc7eaee13126ec0e81898e3ccd50763a09c7be78ab6a94728a56677928899bbc77a7777db2ac36c2f0b91b99829c0cda97cce7e494b6cdfcef367ac929e42e742d8b4350e57ffba5733293618dbb1487bd3543c02719d5f0ebe2e1933584dec265a5c81b312a087f93ee721b09d5f319cdd5eadd20bb9f1e83863f6bb9027e4487acfa69c4a375f3f20f87fd285298d5d7e1d638d34054a956ebacf7bf6139266127b89c5ae0b0f02cebcda8ef2145414378cb6dec505d6e27881cee429741815ea84636b1c4539e1a05463a8a266809fc2f6afe8da7d68563fe37ad439264fb6812671bc4ae06f8a984c4637bb5eee098b1fea89f828a749aed65117ef74e23f89eac14a9b841e9b43005010c292a4db4d824cc8c533a1c2398155cb58eeaa813a8dd812d0f591876b327466b0a1a20625731cae88dd1a7a102ca526ff36c355d22ccbf132997e81f109ef1b4a7863710a0fccafa470e334d264879772b6948bb7632af3e2b685b83a85e0682539785e83ec5bba3d6d8035dbeec962faf542a9d7c19eb77932ad4a27bc59f22e3fd49a132a38a40f841362450add6f23bdd010188fed84d66fa01d1a3bdc3530eb2a902a7484d121287fe89446125b02e6edc1821be69e864b00dddb040ac5cb556d0ec5d9543ca489974821583883350c108e279edafd7cb3743c129aac8e6a7efcecaa50289964db051d59f45997b506e7a6a68ee25d8b9b5911edd294c6852235e3205b33a488f321dcecdbde5a7c6a4f8925070d29c101b6881b33e5ada121aeb7c5c46190440d8b20f7e08136bed252b5313b709a779598922f5848528e0122f478d7f5f376a1e23236b646b9d318c63834a62a29ed7570ad836285c5ad25084d65266c8ad1c5b15c92b070c8faea6e84eef5b57234c5041509e9532430bd7e4fb0cbdadef2cc99756807981f14d18a19e024d6858502390aa55584469868b384678f36871d14dae4ba95dfe6e3dcee61cd1c78491699dd0a52895774355996c5ee170ec73c83f45;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hf481eed3e8bbf5cb4cf4f8bf353062c362703449e054522d88688995ebee28b09b8f70c62586593fa11abcae89d4b918823b0a348d27bbcf5608f74513f0184bbd9f0df374785de65ab9eae6836daa8c70d0b76db90b693a96523bbf5030218f9181d95040387249f5590cf33bfb1c9f982263d93adbfd127fdb3befc38d5913663a6862760a9a57e35e57bb3653dc2f7e2fb7b313ab8103b11819553b9ddc58c5fe52a55c6f9d79568e18a80612dcd3c749f3a334f826d1c975c5b0b7770db9ae1306b202c16b43e85f5ca489ac2f8f87dd35dcaa43dff1663a1686cb4346c0932a4602efeed5789389a58db165195293d86d6793e594628d6c2e0948281e0995961f88953bd9fbaa380a638df27f6813c3458784796d647dac4525fa7f9ccf45e26e6843f123ed1cfbe23605c0a68bcbb400c06c79f57d8dad551a2996bc9c7ef0af87d87eb8f263d107f9d4895d663e69f78f43d232e602966f9337970c0667c022dafd023c099fa64e2bf3112148b841c02c8104a8a0698fa2ebbea45e01ac78ab56c0431c630811a310da93ad6e6998a8353e1140890b0b5e0399e26a90b68ffbeef158856341341b665c5f0815a1c75976167ee4e5135b62a0abbb6ad7e9255e1cf6ca93cc838a080697c0e6d8552d46181a6a34b86eeb34f3e7cfabefbed5bfba240e3de191ffde31c500bc6aca1251872b8cc26a69d3b60e50f511606db10c887b12147c1e9434e2ca77287f9fed2a1776d40e77b27c06fed6520c9e21ed7a46e9d8b1f977af34442afe2929a2dd0ca23ca0e6c42587282ddde739b6433572be2d4e2abdbddc76045ff867ca3a24df3f3dba323c93f5e62a4ff4072b3659e7bbd0791293df141fb8b5416c09add994f2f16ea72b8fce3c72a3645b173b1f4d92561185d138435ce3348685cff77e79f406a78d1c14f7aacf14c74b0122db6110abe6ee53b4307435b51439787190667f91ff2cd315bfb75449f226e01eb7f36a6ee49542d2b3a6a02f20fd2384a3591a3f749e799bb3c971af6e15ed56c8bbec34c43b59faa1c9e77ce67b38f8ad69c87c1644dd876d4fb2176c0eab7c372eb5559254ace32ecca56bfc1702df7ea0dbc7a3f52c064ec318afd2cbdbbdb5225f100061a13bd8e7daa8841002548af0b26e0e313a74dc1038377923c03709fa76217aeb0330fef81e137eaebb8e2cc048376ff7f5479a10bce0b9f96f4af43cffe1863a15b32ced379b9f275eb40abc2b51179d6f754106b837c0cb6315205f98b68c64046b81e89d9fc1496038e9784948f30d066256086ae27491a067e6de3e5dda2b3892a9dc8dd37e83bd3b352fd77d07cc1739d8c5da7dd5b05e711fed67063ed9bd877174de5ba247c7fd346d27fbb3ded969b15db3eaee471e8cf43e4574324bc102d830c2484ce38c04838217461e0a925c6c7e9327a42e876fc35518222001470600a092816049d65d0360a58692041133bc70da2d8fbc6d89bb881467cfa515dd288994a594fae062aaa631d7d8d13adaaf512fa6ba33dc6247214c838a51633fad71af00c99e9d06be549af0b0a352e2442999dc6a1a4d4f2ffecac8c2fc31d4f09ebd5f18e84893b02a9f2c2d694ab8b5fd7f7fba674fab56b1c8fc04d677cc9a964a6ebf365e79688ee3b1e01024e92ce98e6ec8806daf2461d433f8ffd560ac6a88da89e527338aec7697f9000f5da6c0cecc3d97887ec53bc3f2c4795d45ec6ec70f19f060b2c30894896f094076277f53497c92726af81641a8e12966a0e045cabecaf445eaf0982857c2a3d85edd85507900b760a7fe3364e4d3ec52df6b8ebb6e5418ca0a5f472ee58846887f921d1b858c14655152f78f95f99dfe62bfdefec790a2f809019d4bd0e1e83b3b14f86c08f584dc35bfbc230c73b88391605e1afb399bacb782c8f2af8c5952ffc3cf671b319fc1564800d315975a70ffd6a426009a3e02db4be6000e833d7122d235c8ac4ecd748c1b88615c08cab588707409d3bbc98286c2a7838596c86bb6500e2985dba00c8dff3d09291163cf25ad760afb40b1aabc2a7483cae6cd90b5027b3538b4c9d261f36f06bbce7fdc3c74d77f3b0624788e9ba29a191f4275ebcf5051a615f5c92da232e1177a21af55f8eeadf53a751448a1db3092161deace46c076ca0f0dd55f78d50ddb7a0b194b4bf816bc7423ce70299c5f5dc99ae21ecc3f90179e87b1cbc51f5532aec2f36ed22c515ab7081f08be1604e5e46bd09400d2cb8d945ae78a46413fa2f3eb71a09d9a18640297bf22ee08c3f52a9a32bb2065cf659e67f027f5f929cc11d25364b4a7c2c1ffeee27e88340ede473d2d3e2379528a22c33811448930aca9d20a824d2f015c3ac7b0784224c91bc328e98e096f82699221f66e09e65c72d9b43fc4b1e6e464a2c2ad9f748f703b7ba5269f746f6228732d09367554289167a45eef070023ab353928f36e42cfd21c87ac340ba588ba2b48d2a2a656be1aafb0773f539bc5dec4f72a9ca004e344a14abc2852670b9d3ff8665a91dcf4cd5e8ccda5de18ef89c9c89dbe427db5555c4fdf82033e8d2155f4bc75e54b35d1f755c3ddf7e8e43751b9c0bb9282dac17e8ee1e841162d57f75958c96759bcfdad68633c8b57e1d8ee5f600d5d3f800c70373a450942483c8d3d821019c05d01740a705a7167da6688d9511181f88851d4787ea2aad358031c328ee5e812cb040f655bee0b6a3d973d76869900f37245bd58360789148cea20552145117afb9b4b380a33f2684e489e09bdc7dbe1ba86ec55863d652a6e6c3c467428176fa50125532be56fdfb854309c1c78c218500009288fefa04ed703c5c322ebb51d4216636280191e66f6c6476c9f843cecf936f0f72badde8325321542ca46a177ba0659ca670f209a1c0a31998b15d18d3ea4ead09f2da9662a20cc7993552a50bf05f28082eb439dd607408db26187bf905b219a2774cf9362291c2780a90c372bdbcf61ac832a9523a433bf9a657c0ea721157682b46fe46bb3aafb299154f552c22b22e931893d72539c19133cbb991ea4f2eaace495f1df5be0cca38929c16611eda068f3eeff75376d6d0b3477c5f1931634f6582b510c1d5c0d3d623f6494327db40d8e483695b0159626c9ea2e576cd61c4c61fe4a8eefe6387d2dfc8a309b63ce4b96955c115a774ede309cf1da1e6c0e76e6be2200dfb1121554687d49f51cb398c5b7375e5f01e834026d75223e5814451d77664f22d23b6f5c9c7e35931b833e9c3d964d7996cc33a59382da8cf6ea2d7477ab2cb724cbbba4c8b3a4ec0ebe72c00b2e135480052bb6633e963b749df3c484cadb3803e65e397ea8d80bced5dd8d701f0d0c8893b7430bd2d1d3ad647c92010ce80c21b33682cad5901ef8fd800c1923270f9e944d17eb032a1b3c77ccb5c228f826a53251b0d1ce9ad04582b3d08ce6cbc8d02856dc9aee107e0e4ad4bf317032ab6fb0711890da37a6bd419c5d3e7fcd75734b176067e1c28fb515a555a29200a990d0b1f720bf76ff376ebdbe1fc2f54ee693fb22df28c831a162ea5904c98af3413ddfa6e1e823fe300af0766f9e8b5bee6fcab7125c09127b63e60435c0f57273a3786d2dcffd1edcc6cc1f0677c2e0656d6070bea82f0bc271bd24b112d131003e1e0a57b075a709af30749283f6f055a1783c493d8a7f8096cd69ee0aacfb510f034f33c32d4314dc776bb5cbf112f16bc311d648d2847f43f5a48e10e1113bbf716ad569542b5f9ad8036e45efbf827f74119b719098f742642d47f40265ee04dbd0988b2b2284d1a921d8d9ae8e022978dad866f7b7ca45f320f3a69f0f94187a3c7a5dedd067d8c4db49236042a442489d14f249c0e5d8f04e3cc9c3c7bd6445dd8ee7faa9d34184e33976edad5b3687102cebc5f4eeed63adc29a04b9c40548f93798471e3e9c6eacb0931575aef9ad470e7773656e676194657612604e86a8fc8723b34aed0b8404428ead7f56d7a5fefc0be4dd61e49b654a50709ab9be1405ae78c2c9d3672118e4907da33ddd65d6bb6b5adb656416caa48928c12cc67657b16fea27de2d183d938c8f140ab9bbb2a1a70457111c467777312e0f1d3bf7da8840de16a383794ace89f6a1a446b6ff27ce37887e93de89bfce8ae90c683e8e3bbe45227b0e27e0f864c11f27c975d3a299afe88482181eac5fb4b635da5af158a7253394fdc8dec7051de01a315c0b102f995a0abc18a6b1a42f90ce1ab1f63b2f98c8894f31aa07e0ad7d6b94f7b1f5e4877a94737123c30cb4c50a6bdfb000ed1f2a624606a20ea0c4d60a7b45c456fd2a6c7018da72af98703e38541a217ef8691cb59fbcba8bea9dd478d4ea09fa50c8efce372dd6fd6a344665a6773df2a24501163061a8c6965e00efd31eefaeab2c865a279b60e6433eead027b87c203f89362433ddcc391b1509fe1417fa928e95267b0358c7ca93d94eeced127621bd0bcba8b54b07ec570474c4038211b7b37a3b4d7c2c7efe52eae416b57417c31b77dea14ed2567986c76f59548f1ad5d7c74ae9a63d3f9e34c738dcacb1442b8991d89cdd5339147072190edaf66a9aed468b41c5c348b39a7a4e29d307af004ce22b594db96c26e17286ffea124ecd189469abaffcec9754f806f99fd09e06d68a4056453c3f6b11f1f084db3889daccef642f0b9a4e53a37fde2a4d3b76568d95c429d60da0a4c7746e950b9348bcc0cfc44ddc9e8727b8fb24c98d80fd45243cd60769d085ec5ab6d9d9c9e492a5bb4e7cae465d5930104949caaa9eea9e8f227e5b3f7ca1dfb35e7267932cf1d9bf089c45670104d52fefbd7bf8ebf6760e6e8036b4be04168f29d43ed5f0ff941e11d948cc88de62535bad8a83061733ad871d22e581fc869a6b013be94a766e3fc6332b06bcc10f2917cf94e0e0a420bf5155c2568e3510f01f13111cb93b9ccfafd792fec5861dfeb7c3782a9cc27e9376ef852077f8b627edf1ad27e023abfd6cd6b5fae5c1504c3f55ccf5a0aba53aae365bfbd1eb6206af5b5d3117d8243f43ce22b844964fcdb15bb45d64cc83def143c0f46213b3434d7816b25b2ffb2b5cd77ac97fc3092a1debd8b27a1ed910ca7f12af6999d451cd4446a9e8908eff85cebd427ba9c5199b6cc0010454c6ef49e478c98ca8bc9accfd4207715768cf888cc55fd51cfe278d1df41311fae44d8cc4638501a63f21b55c0c3d37e6f1329ded9fc2162a2042d5e9ddbfbfb5209960a38bb2862d79cfe1186182d60d4befeb7653a6f58e47f86a3df1e5f89b5805190f133d814162bf425739cc4324d2a3bd4eb3edd65cf26860f79802f1f2b5eeaa327e6fa9237659eea080e4868a4937e2c084ce69599fb4f7b19267159b3825879f68ee1862b691e5f5050fdee172ca45f2b43a58c0927c9d306f5584553f981989f6ee23a8507d9d7aa9f4fd046db5cca461fe1aa4072d7d9533c1a743d8ed2f8faa40f921dc849a92df6b24;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h6604e1ab5fc62437297eef45e24ee07a117c9376fbcd03560b4578a517cec672b179556fa452e5e32956d62e4e37dc2dd89e0c77620a2608f84e158a685ba7e0ae8ed0cab225d4459c491b1e32d817e6f1ed592b53dcff85a357a7ec08587cf5226df56ba89d3b9234419b9dc4e988fddc33405e1b07fb67c86abbd1509fcabc59ca693066f34f2fea9853ef53d1d6b217ea776e3be39d0d4d24ba68dc0a0868fca242af41364dc912f2cc49a094a524aeebc7bf07266452204222b3dca65f71b838fbad7c11128a4b36e627a1ee9df1ec3541300a17b1fb45c70683d86e537a74273c0d7e5b0fe33c9db1380a6d7cacd19988f5eee82e8e01fe44e2718b1a18f95fc4d303f530d7bea3e8dd05bd5dd25170b59ad1469c2dca95ba85ae349baaa7cacf609c5f072e818f22ead8a77303cdcee0351d718d014911849ebf64f3cb7e9a1150dddefda449c70146db4fb49ad56f640b0a6fdff59716f5aa447d251110ef9454fd9a512fe355eab7e985bb5c27680c7e2b989a63f70d1c70c24007c9341a024f4b38a7f5a497bcb96f3b9eeaa18a1f9eae77ae2627c3f32377ef4ab02e3114674181318a4d362491b79ba6f15cf4031c52484bcbf9cdada753a4a0953f9c03fe11f64148be27905a2159c9e7aeae7acf5a0c3e10734d059eba03fe0954c4fe8c4bd88a425b55b4c0f5dc9fd880eebb9358335a744bf8a1ac6c2a9de100dadf6274b506b30f13e216365659a43bcfc3265c1c9408bb52d7d4810ac7cde5544b6900d4a0680ba7bceda46befabf1a2e07d06a5e9288e6a37080099517a09a9ab736d62197801c570a8f6fdd3526d56e46c9ef8f2544bdfdba0e930936cc9dfcb4f208c3b68ef4e505abaf32a054aeaa10a93c8690db6dc4685d2ed49e91757f4ac5080044519f5462ff568835bcd9d56535f20d70fb0d70f1491c44a54caa94337a9a778b04de8edc0c01fe33656d9f9eb281e71abcee90e6b21794e62633257300a35b585ef8cd64441d072d70525a2390d11205dfd9b77cfe47655d968c3c2874687c8f65d5b28717d433bed0b47f83594d220681ae5d8e4a56d809d69dd805eecd0fec9374a3f97afad1b1a3165533fb2e379d3b37c1aa0eb78295a31c44c46751545c78ad1b213223f77f137010ea301a2208fe93530ebe1103153d5e181e4ca7b81dc7e02fec9230c8e3a2d7dd2f3b4e393572bc6d1f7be8567c3d7bab28fc842f81d9ffa44bc288ace8d4d427f0fbf2c13d37214a2b47c1ba60222bb6a0dbcce414519465179f0700c2553b8972995940f2a7552ba4cd0418c8a2a6f8487bc63670331957bd2070a67a09eafa2ef9ab7141ac1f4900f6702672910caf86869d3e3d9d7d7c8a6b7c23ef5ab5ce6f8144792ff301bb8c1af7d55cd5f639a49a4beef1089ef19c9e17d3422b4d7a4e2431121bb58e6ab7bbc643ff241ad22db3a997a0f2f4670bf739b617fa6ef3851e48b1b2d30250970cfd411488724a0c45e94d04d0de2abd76228164b3f539f1296d52d932000f5ec5474a6af274c33385fb89de0ba7033d4a93bf090198724f403d70f5753a9abf5397b487d503e4396c6ecb4a037dd6f6b799ac383d7983357928bc4bbe861ca92dc1758bddecb6d12e049f0e73d87c3843df4f69ffbf8d9cac61a9711e74a6662846690077ec85143f1cd2aec8ecc811ea75460e248db1cfb3bdcc4fc99f476adbe94d9aa74ab1fa97c436ead6c7c89fa566c8acd82b2ceaa420482c2a21af5f65de36aff59ccba428106560d2dd1bc99958f5f5156460beb5fd8bb030599e0792f64d39416dc65266403a970a66aa52b6c9ba35d15876ad756773f0311ef38cec5c631acfb5acafb0a26b46f0a94acc9dd3563bd83d4ffa1680bf41e126af0aa7ecf492af46f1d40acf8d4a80a555da851306b451a67a71bd5ac42adf7eee0008f2b49974f2daee43a205a8449d6f5031caeb7933dc4617931e90f676a5ec6868fbc1cd2afb40e064ade1ccbd68c7cc0b8b3f61a6a7eb504f9dc8962b881e1b9097218f8b33f9a1c1b89993c3060ec7f1a266caec1001188b6f7e4a5d445cc01037c1bfd7c511de3fdbcfb9ec356f9f94eeb74fa62fea64abac7e9a23ac79f527f69270b8839ef92fda78baa4750a762ceaee40aa8a9013bcc563c415f4cb997df14748ce7f9cbb8ef3bbf0498921727a5e4b7dc7b572b486e60aec5083631adf21aa644dcdcafdec1549289db774d6c04d81d86a9b83d25d217eaefb1406da860251cc153901252491c33c7a4ab67b383f79bf3752862a0e435913976e6bf9efe2a263d0d8adfaf6194d493624e8fe1e00ef21f2645e360694a3655503f132614fc6fc302f01e1d1a41e0ce660337e4c4c8d02dc370503bdb7c1769c4e8f756e036cd4ed6e3c795e3cf0d39ae6235d173715f1c1569095ce2bf0861b0708ccc8338281437843f3c2d52a6cf4d4c8bc234b7a3678f652886b6194ea1abc0ce50121a28f1e46e9207bd3b0ee9a5e1d82f75600d12402468258fcc00cabf2414b560c900bb7d83e8d6692e0d619b13b1a579f5aec0f83fcd25a6460f24900b95213b3aad340db400fc1bbfc6c67b5db7c520837f6a3e0c732f7adff31f0aef12ce275fafe0aef19c6d43454b8448c17f7d3b2b06941c1e28729256f329b509b4922d3b4e904d587ce222617b6b8055895281e57fdae91510abc253dfd0cea166fb8ca26e15c02a870fc0f6693bbf3a8924cac92f949f8ed26033e903993f1775b549029791fc72e511983ba2ec930b901d2a7a9839fb2fa3888ffb09c2bab60a19f34f3786d2e41dd867e1eb15723186e7a999e4c985516e129c165f92bee355a6c6694888cf4844cfcfdc1b9ea774d85350f5719544cacb8170b1cd368c12238de4710039200bc493b234a111ac617a4f9ab44f133e81250814f4fb5d834462db8baa4c5058f86d5a03ac325b7d1e35442a6106058e9f0ce40380b5b7ff3d59f114d7c1d8d64fa277db0985dcac6b3a65ba67e89b7e04b0e280fe439d1f9bb3f08e1dabb854dd77f60920b6e4c7418127ab7233d0d2d14828b82d5f98bb4faa5350f0658d4ebe745ac5012812124db07098aeeebe66dd8adbd41c06646cdb945dc4bb67448661e76ea18b5b4020a1ecd8c51cb4b0f94be87671925e891a38471087c67ccf365131ba0b45b72d2add51ed1e912b89dba4720cb68b71ae85eeb77aa8655a3008b269a2974d09faf3b34341feca56a4b1a017b0694adb561c4286dfc928e88af2871b187e4a76bae8e56eff0f13e627c6aa9c986093526dc18fd149c0098b9ed4fbbbce58588e94436437d246bd00415cc769502b8b53584a6e957fe85d7b7c3868c4996da0837b626c1fc5bfa016721aeae7e97797206c6dfa8382079a4d8f6cbf863d37a6fbdb33abe191a22be1cdbeca2a0161f5d86369425d230ed89eeb0fb6c441716726a29c9472c6f7c5a1017d51eaca52b428fb55b9117f3710935937fb5c3cde2d414640cf57405041eabcfbba875936f7ab74fec76f36478c7157e4babb3f351142ee943bc8ff82dc4cd131f9520cb115c009767624631a20ebaff79ffe92824c569953077af7d3a0841b8776176e9e9cd05ddb2ff51398b59ef58a042847f1c8ea24296146f702c517269d2fea1f8327d3d64caa48889e6aae930d70328b8f879e053dda07fd4db1868cbaf4c1037936e51b7eb046d47c2c413ce4f04ece1074d01022845e4d4ee01aea2e92d654a3c8bc60b10542cb0c66a714d63a8e98246ab8af3f94873fcf5fdcaa7680d3c1f5fe3636d17fad6ced79bf368221862c0cafbd3aefa95cd393a646d53eb5a5e2173c2a0ed6fe43c48a9fbae40a82ef286d7aa552443656644e747d5905520e7c4077604cb3d7a2cb8be325a6c611853993e766af0ad5ee3d7e8785025102b3c8e38c5d8e9249e814236e1503c98bfc99b8125e13d25b86f0045c82041c1cafa82303258fa9a6c4878d1ac315903c3ca53ed77d5da1954c0412ae0e8457a82c54e760b58d5edb73f1ec3d36b5220a5be4e3ecd6d5dfadb63d80d1f26764b9e9871b78054b9629badb89657ebc2ce3b7a3f0f74039c51953641edbabe7fe9f2d19b2f966c72e155a4a2d6165fc76915ad8137b77df1fe339a5a5dd7714fe78c31b221c9282d4e44129e38fadd017629ca59287258b3dd31e721841aa71f3accc80531e4f4573f76b10eeb36f341a0153f8d1557e454899364934e63681e5acf9cc199035aa9db253eef223335feec4b1a8f3bfb1726ee384e838bf51cd8dc9f3d98b7b567180ccc7e3a3dde0538f8e52dae098ce9ffae860f8207b35f17edbb95a106f47dd3cdf4fd76afa3c1f0d9d2b4c857f844a2d0eff5f69d01e361bd04418b2c447990961cce689bd05cf081468b16cd88b0d6283345ab7b6d68dfd9b7995d8f7114c572a5c680ae96690b261fcfa132606c4f2de6567258e671d9651dc5aca9b48ddced5eb0fd1ad24a34668083ff0dead97d523595bc5be9256ec26dbbcf499b7168f3413871dad1c0e9e69545e1ff49f5a088a60b86efd2d31d4131a2d74d5ce0a59a4309787f34c389201825e71321a0c3e2fbbb086cc7a90389840dcf0bacf2841cbbdb74abfb551548c2685cd5904224123e4f3e717cc0e4b271ec400a636c2a44b189b014f172f3c5b450d9486ef61f6324bc3c7497cb353420aa4ef80af8927bba8631149806cd066be303a9e03e9dd342a7ee2d2eb11772ba73f16acb2facc29f060bc88c9e6ec9a9d776d1503a0bcbb83090b3039e16ff645b251cbddc5a8a497e303d3bec896fb47876e4b82bb6af9028a91e8dd00773e94f2187e797d2a74a18d0c4cc0ac90687e74eb4b95ecc57c4e71b0e5facc458b792f5381412f2c21efd2e650b20e146413ba85ac1f34a8576ebf0de8020a8aa6eb0eae46f66b0e321f3500a8f5dc9e04ccb1483f49e36cf6836136560dd386da34d012058c09dafeb8ae75fed0d2446139cdee013908bf672a1801b6f0088726b0dedff32f4b0d1e2e11adf2a628574fe8170e1676b059ccb31889bb0648c2d0b13a40f1ecacc78158c0a838e1951ccbc5a2c166a0e7cd76d14f24b9de3301d0ca0aa6ad754703002589d89180d47cb36beef31cbad877eeacb118e6e9902b9fb865a6ccc19f5bf163b014c0790c759a634ec9a135f0a11db7168dfbba628a13eae3ebe8e07ba47d86a408a98d60882feaa0c575873bdd2ae0589aaef179cd4b801ee13256c3282cd7793bfae5eff4c55a8d8a50600938de1836d40123e0df2637de3208073a9301cea19b3296a5e4fefc1e84e3d7c42a50266286d6b523a22add99df9d0efcb69f3d691a2235122b7737773f9ba2c3324311227aa3d6820a45b2c061f9f7c2058003a829055067805f40017cf9c73cb0406ccc2b3b649b0fa7950cf712765c0d053855d61d3c789f4ba2b59d9bf396abd1f0e45fdb9fa002d3133733653dfc2924d1a99c0736f2d1343b6446b94cd8d4cdc7ceb756ef56;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h8b855fd6c594edbfe1982392787fe5f09f1f699be2ef2f676825b2e6a05986ef646e0646f12b8e5a212649ed10c91ce3be6aa18a5e762f1f732aa19d218e549a7e26ca9ffdf4ff1dc31ff8339ffd4b84913c8b8a27c7a54c8057000f9c3a3d6517eed0d22c988a313b65ff6f414c4bc046e9c21ccb0793aad0aa5c928dacddbf257079c43c84dc525144f5ed24b6c27a81e9b0253bd9223c1f350c23b6acc85d27e17297f0fb602166996888e314d52289ad05100c8f2f6f3a83c238ddf18b1a879be2c6f1536dabbec1e3933c057449dfc8fcf3e4b0c8ee16b49ac588b50dc8ef2d5e3b33da5cd45668f73baf2dd3f93067d80072ae7386c84cd0779cba7bc9bfd8fcc341ccb552336fc597c50b3055a34a536d9f647ea3dcd63c067904c74c24300d3e1498d4960eed1c8f04b1c6975c5902bb3b6d91a15a6a8659b3471f49bdf9c6cbe796a0a7ba5a6c6a9ea387a82121a5b856068a4d46ed8f0cb08727dd812c9f0d8e8b306663ec46de4a7b3cc2bb174f5f764e14a65d0560b5adc3ad6458db278ae6aa3ee1c6f6d927cbd4f076a8189238713315f985199530091ce70b774df7428d835d4de70d4938ddb9f21327c92b0b7af07a18d6c56e2cdb279e8c5eef26609e85409fe1e28e828a9869c67d281e153133ac2a69a17feb1868cdc9ee2d4c9b1165f776fb20ccfbd066d01d4aa4a8f7161fcb05dd56f2267484fd78db168b105a29a4bef44bdf7d70e21b7c069e028a0101921c94bc12e06d454a1d06c5bba949a983e520960fc80b5e3da1e4ae357cb1980d8341f1b7e0f201f338b94bf7aa1f0eef29fd9c5928d488d4b622054f193d9b7ebdeddaa2aecc8330ed0d0f5c3da2356ca14588f49dce93ec3a2df8fb497d68cc4b1e9447522c2da3d75ab1e8e6c67fbf470ecd963e0f243075bfc3349957b62f136185e66e5de1d18926ecbd9ba6d2efc71477dc2eef7ffcc5385e77a4f21f5b4b55004e698bd2c6bf41fbd5903a467a40c3707841dc89d7c440636f4310e2c0ddfba99c6886c67c8f0316678d2b59cd4183b069c1d7486c189a3314a3f54347b51025555ce6abc24fc98397e584d3971934e0fa287380d6426b44151fbf3da410848e7f91545940a7091103f3f60fa5c5a01c96f14f69a3c5c62d13b70b561ed8ab8006a98f4ebafc91f6c1f7fa0e54acd716ce13cce9783391463485b68d242b8b3acc5f7951e59354ae479c77dd4b1f5a9b65a0e9eae90b7d083b9a85012d0d79b2eb8997b3051401c85632ed32b8271a7ddddc4b2f527fcfe5c7e5545c483dd181790517943b4b2c713a154e5bbe114869a0389c5c19a5976fa1b9a6928f9644a627287c033fc9c6c284fe2d1e456d346a6cc4a9b1a91a4e15b193c09c63631215c9eee41e064ab88b76aa239e1ad7f222accd4b20ff91d15d1bf14fc623615b04a366d38ad8518112589bd8ad432b34b46a1ac9019895fea5ba685c977702573e31ca31847e1d85e9a0c7e8d634aa9d811efa4d6ec2a8c100987d1d0b3d0847c752163c94c942ee5ffa9d6aa40838e14527effeaa087ce5d5a3b65494aceb31f0e116b109f265aa4131a878e9152903668f2a405e7c6290f46489ea5f3d8d41f7a3dc808f67c86e5a8e8fffbee8a63bed0d531c350ae703630f703c91fbbe4e4ef75fa2fc59d13ec8b3c7b3e8a5b04b3393f1569dd29e5e12c365dc21d9521916011475b11919cf2738bcca5b179f5d17d2bd6cc7f56119ed52d1c76cd2d79387cb97b821067e8ec6287c0f6a93acd7dffe2a6dea758a1698048b78f7532a1f98ba271d19c6609e1171ed701cc6be590678c190444457d2ed98dc44c5c4d7e39ca7fcf92d660950a6951fbaa2572ee507ea19ac92ca433632a987a14f7e78e4a3d51e76ff114a6643bdccf6d4412c4bf24aec01dfceed5da175654240b902fec360ce7e00f27ea7411925e53f5ad881f1e031d434a692f8679c7ed02261cb533c5a48413cee0cad2215f0982798d1a051f2d08147d8924ca70b45ccd04a517e3143a3a2e762c6abf7c2f568e4a9c62d9bbff5229da90e96a94dd8f90631b46d88cc35ed0b2bb69a0757256e0433a7794270c80c4b93a0b9c46973588479f1e6dd1826f85ea331f8a8af889561163755cc5175746f19446a7316c340dd0eb5740cfbf4971d38e7e528848b5455a477a94d11527bf40902160a46c72820e8c6a57a3ef203d4165309b27880f672ac6e35863515e04c273e092967dddd8251893a867b0c62ec18e8d21fd3cca5af0f05215699492cbb8e35963a993a16ae322d53d5985bcab569e5beedb254ac9fbf2dc38820d86180537c5058498298566c576aa49443749c0a5aed2ad968ffac7344f70d5275e6634e7b3ca475833e9bc7dfac83bfb6224658a5cd055dee55a8fc171e8f693821f37d9d006c5725a52f3fb5bf6c6e84b016d10835b8ede1c0886829ffaeed69812824b6fd9e76e1139ee3ffa1fa2fc0c2846b44c312ce8544f7f126eea506fb7667a8b94a40b67613caa6759d62b1f4d725bb8ad38d46a9eeb99fc811290799b442477bbbbeb6dec8395a4741df816ed1aeeee37062725b79b37a4fe2c9baab03c1fbcb2c1d3240efa343d792e5cccb11b0b8929a015fd0da336dd11ec8e86070d959967ff73a4487ae715e8dda933421dab4a25fbc7b871f804ab225335845ea8dd9164d08c6fb56955e52df87beabb0844b100832b933db55fa9cddead8d3ba6699c6782b50f5acfe556baa1cdfb4cabb0ae9b721bce87967a122da128dc631db0f0468560eba32aa8fdd19bcb4dad626cae089e98075e1d4c4451d06c9275fc11a3fcc7392538eb31f2a6bf937c2d70b10786201399dd07916bbac0033424f673a5f77b55b76ccee60f5f45befbbacc59e255563ef684e268b2744bbf21df00aa38e197a3d1176d95f2e38ef2f46f978d574118593cf63cef184e52790aa2dfa33135abe442b0e0f74e5f0e0394042b5b56d85f20b8249d35a045decc1313b5cbe6d1e671bb5961d1e4594cacc18b61ea6bd88251b5563ca50347aa9c9f6baccce1459d4c1c66338bca65e1a4c375ed1fc49256a4dd62769b4104d6c8387ce5a46e703f331c0eed330904ca0118838d57a35867c1f782aeb30edc574efce4e356484e1651572be53aff65ac1c478959221ad2cd28e075290d93df16cca3ed56efa6ed64aa519a950e4643a3b458361b3bc9f1251c0ae1ca80da0cf59dcfe2ca9fd402f7488eef358055689abfecd6a70a0364cee7ec003d3efafcd26a5696ff6c601b692e7481edffea7528a3bf34b12aa924a309f20b51474fb29113b800a256d35e97d067079c57683cf6aadb64320293696635c5f0d65d1faf712e0568c28cda88c6e52955a374bf4c7d3887fe34e01448bd26a953d72797c59354ef11f1e892a5256aad90b09a9ed15279645a08c305995d305323933879aca0755616666e0bccb5ba65e7c1d384c36175b895ea2683d9e78572c8e479e7785e4781dd95435834202a7b297cf1f8c49237b6896e25dbedad0a53884c2768c2c97ec31c9d3428399883a49c8433352cf5d32f3db2d7d065b196bb0404f4d3f690df471abdc4dd7db71e544ca952d5f586ecfd43a8da170ef57ee2af017bbe413b1564d3049a58342da2a4e7fec512edb6f0806215b6ba5da6f5a7863a2dbb7b2f5c0d55f62f8734f2b10a2eb06b9304fe3433e072f7c51fee343cf9bde5d5342279c2d268e0d77b397858a8412da67efe488329463e820d3769d0bf374ca94eec36731c15feaee6a978229592040c837a2f1ca8aa25a5703f6cd96e9f5db35255a6401cfc43b3cf98d11970ac6b2d5bd221e77f9814ff81b0eb5efd432a6697881f99418d3d3d08389e48a1daba723be745a03ffe6ba5404543e14cc3df931b8c6dd158b4b05e206142309b206b2e17f2e9fab81d52d63dd378ffc1aa78e75ffb6372a292b926813b8c4627849bf86649595e5240f04da39481e10345dbef73ba98194d3e0dee743f2daedb89a72258c8661700e3871f103aa4cb9ac343f6918ec5b1202c69adac351b5fe376cfdd3000c2238ed970103c9f34ca5315e0e2e8c88001227a0d2824bb900e8ba9426566bf50547ffecda966b96efbae6a0a4081d8a9ef42a145e1cf23b457ee1e115e2fcfc6d86c2850f23c3ce8914d95c6006f20b6dada852b1c41737376a1d681bf3d7cbdbddfe89fd3dcaafbb283686d15221175e4355a8045048f2abdab4fb92fa1256682e1ee49f95a73125fdedde64f1698f2427e4f0f998cddc97df7a524566ac57bb2a5e8772d08a1acb6fb77c256e2dba193fa3cc32b52a5908071516c322b5b74f2d671ec153294ade10c7595a7aab3b2bc4ea5e5679e19b01947d85798e3ee3a8bc8e103447fb5e5d31d1073b3a0435f9cc3dca254ff4b4300c8e33d127180d78b9438c911b2984eb48392c23cd7ad84617d8e466a7191a94e3ae468d6be17bc4d5615aa4de96d7827d43c1b544bba61b15c1e3402ac934535091a81de482ae19845840e67b1a6977d1d0065137b6c0bda1da4aedb464f7c23adab3b0afa06fd1004d081b6b8036f4995212f9db6d7af68c798f65d426417b9f09efa01ddc9bcc016674bc4270698695c1f9c4bf0b528ebce7f91f19e41583649d40605c2ed2576140a2aa0543dff6070fec38f8dd6b955b99444a20ac4c33046d91d2f3e75c870c0ccfb35ea7cc4720d65ac68bf6f097d263a35c9954d7b326f780aa75a16db4f0c5c28e4ded45d54dab23884be17f8977d64218b55eee68341494a5a2c47dbf5a3609bd4696a12a8e99e74aec05cae8baf9e2f3509e90a8f77ff16ce2d05d7ef85a23b0ec903eae9c81fe4ed7cc275e895cd2fe0c6d86a4b614e5e41301aa664fb409265f8930e66a9a36af5bd1b662848598dee220385ed77ee7a6cb0b89fdf87e46b3f8fba5b87abb3d2b2ae54f01666f97fa59aed074f95c3b6d403f7970f91efd18bfd0b23853e756e892bc2c7246b94bd75e0a8f632ce01a17687663b5e4e1bb76f015100124e3ab24300271e7821a08f8abdff2a5655a2659b52db49aee6ba9c260bb26f0665b670bba7e0fa3449745a2a25f4e1666c77e86d3d197592e3dd5b39bdc174706cb2e50a213d4c2d723f020afcf13e390d15ce9494ef6e11eb897491c4eefc9b7149fd4546c4251bf1ce62faf5eaf8251dc2d746e3a6bb680843d31be2114164bf7c30ac70bdc24e7e6be7a6c72f33575684e25d084c25ddc5eae4826d288e7e8012fc6be5ee7005eaa4466a28164a76ba758b5a5903bf0db473bad1a030faddb42dd9d4fbda3e778ddf332dc3be4064eb3cbc4767e032567814d1df1c498843f08de69fe5c5d53490be351b74a242619bd704e56d9276a6ac58d661d0206805a0be69e8dd6ff1a738663a21c2667b7a964c8716cf2b03a9f0fb63c3fc8fc9b0875e6722ad05f2c399bc8321dcfad23a81d925c8c2a57beab140b933c7db77e25f2af86b01836a0fc9da25f73;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h89c7998a94a4b8050e919722521f8387fe28995edd7cd41981e20d496da516bee627c32e2ac1b22e6773ec2d71a96d3e8b71d8a1b94c24dd578d1a3735963787a5bc7a63e4f641701dc0e663a6fb1cd857f3faa07a595d83a60bb5f5eb6496dff6fe0d8fee69ecd66879c2034c6726608c59f25ee38d2db2b3c888c9bad46a65e53cdd614cf8ea326be35d0d8a15db3a594e24debb6c1b86e72e291441cbf23c0473fa1710bf14f27093c1d05dfc3a13a65a66c4650add688cc42c78c1911f7ba7f71206c368a5b5f0be9cd67380f872e469bf07b185454e335055cf9db8315e386205814843677aac9237f5eca0ad027738132ad11ff7fd14a5708676f7a63abcb0b4f1524844634d2a9fd489a0b7d6afe48ae8dafb47176c7043e867d6cf07bfa2733cc76f0e1aedb2c814b0dbf8b8378f78bc0a2679305eed77ca349b37da0de389757043f74e850497521fa2907efd615c42355b45c1dcd4c3e74f0dea97c2ec32764ba7cdbe4efce3c952ccda087e13afd5371f064a5d05db3c1fc7a9146f85285344ea578550e66016b7d32b1b6d24d3a7215a20f1c9c1e3c6727f00e6da1be01d02ddeef5190448e449079a405aee4ad126d2f9dfb1450424d2b576cb9dc1b1ebb3c8414cd1a6bf9eed481b3d02de296fe46e88f6cd2d3f8b7ccebfe00e66e7d34668ccaf749166c2d9c146b837dfa4ea9ed8f7890a0e396c3cd92b535a65e7aed89cffa284d23091446b3ddd46b4c75137d72beede105d09b8f1f8bf5c7672afcf42bb059728c67d0d8b0644f99a72946dbfc54824caf6386c7252069e7577db28cb486fb4041c490950ac7e867a529527cea676b165ba3850247f8d29a7babe79cad007b69a6ad962f249deeaef4afc77a85a91907fff3bb078bd23039f8752800f12bef29e3a184ba3220910cf0cfbd47c3cf6dc3e8f7cb677eb90cbe0fd5dfd0b9251e4743ae1e8a4a8fb5657019a29e62406d905316f510885fa2e6d6998dee9bc89132ef4fec109ea5c66b2d4521da4dd537b668f2be91b7bbffff10a0a64c74d6ad43605a0925ddffb4684bb894f5b42cce9f62a56630809837b03c17c0345818b3bb6668fa256ef1e3fc4d327c68778d8b437922c5236904e1b89b22a999bee3f8bcae16deeddfe3442ee3397a62fd535dbe07240b1170e8f046f0c7d7536ebce264111461cc8bce1229f7fa132a4f59e5d66212bcd63107bb71b8d91819f0d7f6ac56f24d67dd2f70f688d157c1034b6ea02f9e8e08575f427558b24193a40ba7013d3c0fe0b30191d991a88d43dc1afa113c47f223ad060659718970c256e887a8af5e910fa1f7a949d34e4a4d210b689f38f80bb632d13fb6e48b21d053cf49f1840eba2fd6ecab689e435d55f6fad64ceae8eae3d4d6142894a89bcc2741994c4cca09e7a6cdb0cae908ef73b7b51b44532e73d9b0bea55b2a76993e95bcaf731e5748b49e18931dd799f7969ff325ce652e2a3b30bc5cd68318f79a4b7b5603dba4206a7bc2d18fc82490467cf04fd1d50aa83d9f04c6b2822bc31ef8496617f0161f68e99697c310110156f868a289a45d439138afc0bd381316c531714274ea0b044de093046bca18d86932061cb86625397ff8bc63e1e23e275547b5e3ebcdeca95798b8f472611d0e9256bac9ee968bc4219321aa56fc37485ecac6b1f3d15afe115cd6718f338619508e6c18d5fd2a2361fef4a5929a1f7d51186e6d91431b7e3bfedccaefcb08bef8aedf9670caccef25a567f7ad503ce53f50a3db3f102c570f5fde27ccdc293bec124582f23ecfff126b369447e6058a770f75510f65ff185332df7d11299aad9626e1fb303b275cf28101ee4c20506fe8910cec7a8037ba5064fb1af8e6b5d3575cf9984e3e0a05847a5f1b9ebe3e1020b13015a7952942a569274d2a91706bcf1cb438e6c651cb933f722a58e7c181cef3a3cd90d8acb05520d8e8e732fd9e84a104d876d0eb41af47a1b597ccc982f8954ccd071eab44e3e03f3ab0f94cea1d969a3e2692c1d8d71bc58ab4d2c00aa29e39eb4556b873c998ad7bd9de67bff0206415374b9ea1a47c58abdc442d10eb82d30745a03f64ea63bc9a8068bc58cb79136cf373cb31a3c3b32e0b1749a3ee594207f2efaa06020bf2020729833722ae763bbdb949691685ced8aa0ec7b452450ddd9620e076ca5820bf957518c1c8638c78f38a0e13806c49ce44025017b24b2f89d2b973b9815e10d39068c65f68d7d3c818d03137157b2ceaf97aff42d66dbc6b55ca6f3700dffed787a1bdfb9f6ccb99bd678f4be403235ae1a21b08e57576bee6bf27caf4858ae6072f7db7aae3d251ca9359dff1fa78b69acab27da20dcdf4503aaccee10810693bc19818df924c02e098b616ab5ad74399bb3eb2b649cbee21c92d19ed251f0c08bd505e5b5418320ff6aad9f5f35de2c26e991dc5a43b43f64d75429e7507c9aad2e39a43a70a9ce4df3873314a32e0fe5ce759da355d709acfe24144978e13ee92724fde14f8fc5892eb399adf46f4c0cd0b61f7dc3ccd0eb472bd0752dfffca57a85a83d7965ccaa9935396bc65a6e9ff85ffa64afab12deac2f04c99ec49f7cbe6263281709ca66af1dfb0255d7f8943f2316462fc3af0839358705a0d5ad3cbf05e36988fb422067cbb2db182459c5866c8b7e908a357d71ffac47bfa9005520ebf675cac22f10c775ee5b3df68b65acff39563ef39963f79b459165a8dbcc2d99dfdc7fca9a4b09d210ee0bf8af0bdab6700aab52eedf5ef319c4406b8678ef41b3560d755b531ed9c027bc3629d6cfffc4e346395c5090f3aa8b7b73b2ef78c433aa3139b1abe912c03da0f1da61060098e42bd1833f245a6ed2ef855921cd12f05360b2503da83a3edc27726de3f622a1772a1dae6de4eb4f60105bbb0303634c30eed9c979357f4e05d9c45dbea4e95848ec06981c5ee45029225b77b955e9ec352f634ddb7a05eb69afd2a3ac4572fb843dc807fba4e96a981fdb3745d07a7320346ac4ceb5064cfbb42244f776f19e830835f4ca790a8242b237c7c130c0100290aefb5fcc7aabfcabe34429e4ffadc84514632f2a7fca0c6e91092b0080944f4c7dfffa6bfefa38f401a697e731c37a16ecc65b7cae89be448f6444a0acf7172f93354821579077bcbef6185b11cb9aad9845313103820963a6805132a71391eb91b8330fa62c8fa0ca0ebfad92c3989a426e6e4eef421f7cf4c00cdfac8a46f5af925ab033f58b9f9e690ab0bf5b6e0a927c8abb4d01fc73b8970cd66e8ce285f09c43d663dedf04fdef54d68a4c90e6e97d16cad2e3549a2ee1fc2c9a0bcb84e7862ebb5e4d555cba2ff78384f49a167aeda3b30dd6c0882be3c567e59ff9f23cf79bf7d5594a165c86426bef4089985b3d226df2ef84cc481a842abef5845bd18ee05999bfb61666c5f4f2de6a4f4e3028b99fa540ae8e02804e88d441fabb23418e5d9d010b1f78912d60bc6d477e4d46c7f793cc4f0f2ba423e47c49e17b89b535216d791a751474debda0122ae6c695410bb42db9ae8832101a7e5c8e264361902ece4159b0111e058c3b49321ab9a6bd38ff1517442991a2be2765b490af46618294d74ae6a17a81a79582933ef702123d211238c678e45952f83d7eb871f4c6a59e8be82510c8e1b17849d3ad70f5ea636413916fed4bac6f50b4dd102182d370e511b9d8169bb8bcb48f1a14ef90933ceca01dc85cb287a8236aa7eb2e2c3e0888a222ae178a1d20d177933025c2a5d7b8945ff246007da0a7bb438119b5df83a7f5c0d1803a71ebfbeade546632e2596b988361f8bd24730fee2b69afa4ace71fa66694243af7cc2d43463a7822a27e0ac4332937fa5ed9bb18b281645c5343c3620d19887c9056f4b0720ef9f96850b8fed052bd068cd73d2f8a23b81bd11dd07feadd05d3d3ccdfc02d49ee1455d771f26781bd0f4b9bda28cc9d8661930b6be505ce8fa1a7c12fd9c79d727ef2418a924327e4e9f31ab73221caacadd60f3deeb68c1bef564dba3a4563ad12e2df214f9e9c84901b78818beaf712cf8b70312d239f49cde657491b6036083caf651ecd67df2d13e43c5a33eb2b4e8a71f4de8a95a973bfcf8a8ab780b7b09344ae62413945dbe1b1d01e1549e32c3d7708964fc31617cc63deae39865971a2700dcda9b97983c0f76b113a662e171d4ce4645cae359909d0b30688cddb5226ce957c4a2ae1efeda3b50aee0dd012c51aee4e62091195941e421753f1a78e5a74261dfc31376e53089d5261df46454d89a240af6d28dc6a22d01acfb0d693561fd4a5e6634f4abab2293024a53a80ebfd0c99bd94fda886c09c91915292e1a9ff385671da339bcaba245a5358f7a7f3df4a2925733eb10e6ae52efe47d43c1631d1883ef98dcc965d9ec75f00f132554725956bf234d264b4c3e5aa3be22ffbaef064b8f418841460d6e8f79534f3e267cff306d15afd42ecfdd5ed705e1b2231c9c81296821f2a9d347bfb53a037d0537bbe3cba06e70b21ed2c65604dbad382c44c6a3b61387b71b645c11bf25ec97fb9e0413817dbf8e0b292a4a2acef3680a6846a461e59c36ac165df81bb1849bb0e75a0bbbbc0bc700467a7514d7f9fe6c1a8e45c6409a2ba52d430737f836cf05716c3eb3d633d5a2faa05f8e58ffc5683a54092d36e8a443c5c944a5f266af24ea0a28665e6aa74242d45d101041fe8b3f5b69bf57cca3860f804e5a2319a7093d61af11d7533fa8573ab1e42039de28c983540ff47013c30528ed3b551320fd299b924e87ce6950487e3b0c8a38e77e81418ef47666dfb0e5c67b1096cfc4dceecd2e90833b58bfd9bf12d7ddaf92df3cb04e94781e8bccba6f386faae937d5db4017f172446d935c9691cdf4cfd3f0c30fc51449f9ce7d176bf78cc0e898e5c7efcecd20ecb6bf5e631df98f800369c77d0983dbf58d6dd541fb56adf927b4581897885df16d7f412e60b19094daf505d9cd87860967f7eb466d0943056f713f50ed2c12a10e92aaeaf1b451c25a608e9749da7a6fdb03bc30907b80bc66d25322d03981d5b573d702252284e4238616b390ff187e0b197bee545c4f7bad5876e11261b205b488175919f8eed2be1709ce5e4082573bcbdc285f07619b9982575ab9a97ab5ff2282d2d6ce23bdc6194793daca041abc50d371d657f7d46945eda7bd7dc88a0da528a6d0a1d5e8309c9608972c664e6841c07bc9b121f2ec25e85b4f4ebaea4007c12741c13a75e07c4bef5810e23e8490a3d0ae4cc9a0b336dfc32d0a89ed02cfb6a5305726e84467574593a17b7298e0ccb68f0ba8d71d0944fd2a7dc9128861235fbb79aba4bfbfb9bb6076150e98a27d7f6014f0ffd696910834d24ed02b81f9ec77b50c2284cee7882c86a9bc89aca1240a44fe58f632f86da1f107806b433cd5698dbca7c25a61e9e6a9503ed698e4cd0e82c6f2c066a26f8f927bcc2db3de64803147ffb289627f3195835;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h7af2ee487430a2ba407e7f2ba0667e1b68c138b9bf9a1cd165ff9070a39204c00195701687f2a8cdd0a9a7d07d18316c6328dd1648f396422aa6d4f19d3d0875d4f6b3e46ac261e7fcec9da245d0d29b0b70223897d492a5b25065e66a3904d1d77c52533a8db6e8af0395c343e0c1cf5769b2d4a96457e6a5eb16e0b795197b47fe583d6ff4baf4c17f93803abe23790fec40e97a2b114b3ee39aa2b309ae694439eb9d1e69c23651127a059cb6787e97c6115015bdccdff85f9e59a325915d4ec3ac0e53ec17c791bc03b673d54bf3eabe1063e7123688cc537abbee54acaf4d9ba859c21f1f69021e1f92712a7ea58aa46eedd32b12202aadb43e760ed0c81f82d0b5cc0dad6be3b4ee3d973a0a6b1401a52787b7dc015e7be2254931906e44b39cff1e5c0324069dc2b3d2c2edf909537cd2146e3b442eb545f17b5408ee42b71df9f1032f2a4ff3f8495de6ae2f49cc95991b965ac7a9a6396fc472510fc2fe432faf547ea3e98cf898d206bf7ccd2499d482cd36475758c6dbaa2214246fc2622c5f20eaafd44487cecaf6d99fb240e38cea295297681e58c30218733dcc88660cb9ef4b1dd7eb849d99f1bc2ef97b8c2c543f6f0b0ee2f30d7277726f0c674ff5e3431a19c3958a60d38c271e3451641b900fa4908ec6d09b2f95852fd7e2985365d241678c27351eb7c2e2a8e6d46944f30500307ccf5e77846b2838a693a71301f07b58afed4a32d51f3ed9761b060dcc9b6983abb66debc92e144de8d5bb2fa866e4792c14ff4211e3f666d98e88117465616898145f3a6e78adff92529e48816c3f5796d1745ff36887a8b27aac86100e13c26050add21be1f6c62bf6d53c6f3d0093c84d3fdc0110425e29e149c308fcd564a005cc71b9888dbb2d781c80ac519ea0e31ec818e49c707b3fbe047fa281076870eadd6e123a775c401ac58feb3edb679ca2207f4931a4a7923c0ef2ce6c28a0373ae241f8b41ec089d8bcea114e27d07f7c4d3a3b1aa77790660b447e8b381dce788d6e42889b2b783fbaae5eeb58a6c9e56bfaff61453accc0c432544836500cb2af4c697752077dc96a033fe243c8c6ef877e4fc89bc362280df1d41110d0e1dbf900e38cd8cef46d4a7cf0869c9f6cd623c70d0be5104c21798752809c377ea1eec5ca60698a55fe43ba5d2c60a462050639b209ee87666a082af660eb1c76328f66f1c0ed53d942e9ef1ea4d6a90a3771b4d9828da35f7d854b1097f4e6c37d4e0f320cb6389296e45c2765f9cffe5326c433fc60e8b9e3acd05e519d621b2b867896f0e4a45707c2856ab7ed0f65530fa7de698289795c1c3947c341b57c6caf95f19cc76e2fceaaa499303160cb67c0f1b692dd76d4b3eb4dbdb04b97495e15ff6d65a885e09c1ff8ac2cfead3f0dbaf9c9860b9d96c2dc57f458f1b82966a6142fce53cd329de5dc26b00186288f4120e1b34354f28f5c67cea6831ff831281a00b3f3291da5b4278c2c4905ccc526e2293008885d9ab8fbecc5a8e7e5656abc4b49cbc998a64589197ba621400d267624c6450f7afb9fb4c35b7ce7db540beca05bd554c2ed85e11e31baeedf5832ee02c45641ff2f21c0f60fa43e4761bc512a2f66da780e305f2953aa8fd24285661845b438c120097a2bd8435374af6b83f7ac7094e46b811813aec340972e88f4f30df6dd5027c53bbf3d96ee39837f7c3d5bd0d4af9ae543c9454d1465aee68a40895aa34158b599fdffa66eb94fddba1073808bdede2a599c976c49ff07d78e16ab36ffa66e5e4d278821633c3b9ddf70eb5b1e2009fa04906e270fca6985bc4575b1701d6a37a40db4a9792ab2dfe50bc9b76e3dd9663d4e5c31d38dfe151f7b06505a1741dd3a3ce00f143f23c10c14bb29626049f347dd7ece61bc1d643de6bfb4b972ca493e9d8b6632d65deb09329639d6654b65375e3263340cb30fac6018798c738c620d0b98aaed1c148f8c87502084381d264abac323051f088971231319e5eb97483787ed8a04fac9a836101b30c231aed2b987424de9fd790b3f5d0e84b7e559124b74240de05b38bc2ab8feaa74ca458a6a896ebead4a7da0882999f6e3c099f53eccd0dc8f0006c47104a9e004181991ab847e925e30c678a5214f966f7b392b22129d8632e98a7fed692d90637a56249638381ef04cac77a3d69a3ce0d2de2be197f4ef42e95c53d86a0205ad6ef1cdc7ee86525a66e0a3d6dd376859b3c57d114b16c48f78148da8b860915f257c91e96e9241af1b89b328af8c8afc73d8c4438f273a0454d017608bf968527ae02e64eaaa45518f7bd3daa053d151b00e2a12bd471881872a5d9d1a79e78f26937a3cfccc5450badb668198273213999a9c9636bb4e74c10bf2a904ee99e163f22e0bf3d15108ba4c57014870067669d71f7a9f824d8ec5e2045b1913e8adf0454419baaefe48cf8a6cefaba2569b1de50970f20e5893d7d1fc31b18f02f1ca4a877f3b1d8a6d6e8cd6975589d7240683191d46203ac3e1e1b6458fc958ec8fa552fa7744f79662bb75a69c30ac3f10508e4b144c8fc05af41f0e6ba60e91f6c7a8250eb0d188fca4f3f80e79f035997d69ce60ffa4a160e01de1df6d348b04cd0348928e9ee98d0933af2f02a9ee171bce5114bcf86e88f476a20692fd2b871430457a4aa49d1ee2a0f128813eaf1aef85dc362751b8cd533ad5d576ab9488ffb750912e366e2daaf96c32ee51ca4e644581862a12c45c35b3e2252f794bf592d6336d653f000553966c5408c907f01f216c683e6d56b27e254df8f5af631e106b6f0a0b244f537a47193cd67d6aefac01ab50d0c86d56e9712090d639b740befe2d8b57983ec579d1d7b4f32f3603cb9148935c5f9d621669eb6862f37e591a7457db6abc1b4a3a6e272c45c344560ab8ab060f8b56217e4a42807a199596baa8e78acc17b83ec8be9c6942cc8c3f6d1ce0cac2b0e0c7b79b5e96ec0943438a93f8be6fbe9777a2ec6f6a981577b1e008a7c00caabf8b7990f97cf63db8383f13e9889eacf315643983e7a79220dbb7ee079c3306be1dd261ef54b9660ea9fd3ccb41b80a40d413d4960bcbc6be277806081ae6f8143bbc38a29f45a478b470be087faadb78c2058d7b972cfa74207d48edd897deb221659707d5d5efeb1a55630162c25f1aaaa94f9d5147d0947b23696321aefc8c544d3095d9b800773566a1606ed47ad9fe8260216aa096755349d18ce411ab5de645d21330b6a2f1ffad34218dd18cc0a4b8c760845b3878f61dcf4aa184d24c83f0e1236f89f61edae7834ae0f77fc46373588e87cb01f55ae6c99b8154e7595a89cf7ecb05b7ca212f4c29ecc1faa2c38cc7858366b00b584a225e0ad4c57deb3d179c71321d3c4113dd0dd860629de727e391c44c94f6a21c8b53a78a1e2e8c3a0da17c0d42aa950e7b1a74bb86a76b1fecab59305208e2e566748fd209a7995a0c5d8ec63d349bcdcb74e4bc945423b4edd05a98a13d71f680d94ae06c30ec2be34e298b5025a53b2a61da393f0a2bdf17165724a0f81d8d3c04828f976b9b60007613bdeeae9493e81ba5ecf697da5ac84c9d3b68f7a392cbb66f7df9b61144cf66939520617c6204670fbfed2b748b562dd97728acfd4f15cc440a9b386a7ece4683b0ec8d9dc20ca9a5fd863664d1fa52c8cc9fc14cb7fa24df758bae283b8fa6ba03d267999c8f6f4c99bfe77e7ea89e420de32c7c000e0d7e4c92a84bc144000e564328c00655e2e9eeb1461ff0ac90d182360737b02adf8e9892c440220dd9213b6f4e5c9a42594c054fc237ec620469265cc7d12a31f4b6daee3fff1b19c2b645bd8ec8c0307b038cc6216091e4e800a6d1821c18a46a96e653a45230d47722f6bac4b4d65a1368bab6561ce63ca2ccd4d29628f26be0ac2d3c38ff219b604953b7dd0f63a95bada06e83b963af73c896133e8a873955b75cd664d82c5cacaa1f97bf53f43b25109f227ccfdc9d085415896de22b1080d63cefda7f00346b25ddaa6f72a39afbb53783b96dd1623f7027fefa020858f4f25666b426d990a2e6fffb5d28baeb8eae2e511db162bb0f0e32768ca6451aaf2c032913baf19d19fd2b5a332f829bebacb982b81e455f2f448b175e94dab587a6f6312a5efc942fbe0835e4fa11729c8e7ae6a6e725408e966186f23b1866b8ecefa69e43a43d6e03d65aa422e35f511e17633cd138eaecf52fdc9b668feb490e3b887f17f478cc7457b0393cdceedb7f13b92944b731192bea9fe51cadfc443256e16a3c6cc854bbb8e13277c72e8a79ac1ea5e3a8739fbe4ce26097bc4569a05daa85ee0c41ee16e9331b18bba206a937066cddfacbfbed84cb8c379406afedda35789aa2e6efb6bed7d4eacbb4c198eb628e51e00ad3200b88a561caf9d164a619a7242a35bba18c8d531dcad324d7e421b890c555849da0379327a4aa9cb77757832df9208713706bf58a9b0a365b424ef94e9b783941a3001cdcfd39a4c165dbd010fd8df077e9026e56b8b250cffa8dae53752217923dfd7e70a7b27d08cc68b7ae5ad50d629c436f34f1753506a20e0ef94202bbff53e3601fa87cdf05dc6f6243239a80269543603c8522a1970354fef38873d745ee48abb7b3cbb96198a8e0245f01e89fd6686e99f03f8cb8f41384caf406cd218401bed9d2af594c70da00c0b9c003b52da9b5d7f02430df6a6a0b07e0d6f9bfec73bf12b82b7c051a6dc647e9d9c7ace90adbbb74e735826ce2feaa4bd87d6af020bbd6c28503d8526f29bd4ed0a75e024a1495217bc942ad34adb87445d4fb38a07de89d057179934a5bfc706d8e1df146303a90ae50cb02ec888d2d88dfe4db6259334292ac39c4dbf9b8fc7ae4c7b3ad0d003ae16b72d988f638658f83e63c96d280f2314b5ddf4fb87ada261da7dd3c447602f1025deb4e6c7e16867fa2b5afe2cadec03564f90dee86422ef3129d6632e259d5e1ac11718d603c97b2d7e7b7624ef8c57c5d16b8dbc13841b5f1574a5109820daa03c84fe635296a75f29f61329e0360fa6a13bbc75d2bda735b3e4e319fd6cb98a060b7530f9991bd0d13b2546329efac68a6a49ed5ce4564fa1900a7f5dcbcc7a389c5150239b62073c4783827f03536336e0a4b9f819d03c9981467bab4c749f28f8a774b17c2ad88681ae93add6fee7e14bbc3622d3129fecf5b9d0ac33b1172d5ca7841d8f8ad515a46d18bd0ed03a3b9f8cef8e180a08a45d0f801442d65abfc39c4ca3402537ef038ba22b011d096bd05c6f383857a0055cfda5fb4d1f26cb5f1564e5f1199a1a8d386ef5ef63c57997f99a060b4e6c6597411a79d91708177db58c4877d60da4ae02fcba840ea11091f66ba7d3f408a8fbfca1c8713df1c05c96e8fe0a26129df1d8c02b5104f372a160593ba4d9922cfa480cf6f3f7006df278c8b85e3c1fca38a11b8731d4f8782cf17d15a13b24e4c29f0cad5b3794d7a147e0f507c561527972d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h5594347e2f099ed975ab27254367bb2525a0aec11874df23f8f4bda121028841e785b8d710a566ced34da3a1ee688a84b7bc76f3dcec073649834a5a6dcffeed8124f1355e7cc5bdc70f8d5e670690cae6a097dd7d505f9f905b5084b9ca699676193821652bc02e8f128c63a675323c0f1f2486a9805a85b36c34a9605840275332835b022bd6fef66eb3233ba85957e4639892d589d7d8a6af2f1aa25a82a4d83fd8925ddb5c1b0fade02b05840cd05974cce74c70f3ec50b2c37127f0b4e86f8f6f0257942b642772d7719ece4f77d9e9d5b16bbade0ae678173cfd0dc39bdf34c66fc0eea17e0dee4ae0e397d39703300861e23a40c656fb3068f82b8620b69053155191a6c682a7fa49b2083717b79d91f94afd74ce0b22ff24cfc7913c8ee91159620b522c03552ae2d43f77ca0da4cd7a3db03376204dc133937a14edaa8fd5a7dcf17022dcc719aa608f202e07591291d0333d71cb7d39ac2689854e0e9c65b25ec9ed47d83512779d6d2acb2d424b7e836cb4c74675031e64f79f34bb81e493070d53ff72335c31b57c890349c6861ec581f4f6aa92376ff86df1d95388fee19d7ec35882b20b580a598e2068b0c407ddaa4e61b32d28b932f2cdc7862f304649778f04375cdee023e3f34bb15591a8066dd17bdde5098f9ab7dc1cbc284c77ebd8def46f5482c82f99b058822018c6a5ada9ee98a9242cc564641150afb0cb3a87dc5ae5e9d3e87ca3ca7d80eec0a8feed3976d5f00606d9bb11fbf6f1035000ef4ad1d764400c58bd98b65a0db0ef24191277b87f0a66de3fae4f51a883abfd7518336612cef063cc043eae250bda06a650fb544a411de9630782382cfa8c32ab0ebeb7159db02e2f6eb18cfe8c7db10d6d95da8e822b662e335a429ea5e867d74050de6aecad17a926b85a3166607a84ad2182251ff1e2fe206a82b5577c3071dbe7cbe15e5e36aff70e06a27daa00035db607056c70b003883718b3195087d312147851c083966612fbb8f3230c83d0a26fa5c6332c94fbdf4312d890cf0f1681dd756320dca4d7568f165a49938e23333cd339d3a5971e90de701573fb3163465ecb28d56df8a35c18d296c315aa6e2e9c1a834c1d201fded872ac1e08e23d5822380cf0c9c7f7573178394795f6417fa5344dd734b0c6186212d68e5239c47d9e5c7832c45eeb876df26a725bdd1b595769331609122bd53ab1aa669f7e2f23ecff562a71427ee97dbc86ffcb0ba66a14c8622384d1cfa7bb3bc948392a510195cc44554ca20753d700e26b492978332ca4e0748f78943b9799e0e0bd34abc046ce45ed3a9adf341e3c039fdaade6ef24bc194688dafadc20ec9d2dafaede8da6eab3b27a2ea05b0250a870ff7d2d39cde18c6220c65ea2e579ebc3643d8e65fbafeb36502f780d14505ceb8e5fa4ee4206519c81bffcfc2161fa8fb4fa584a10075247c5d653cc2502522519864cb78132f9987ad390736a8c4bdd01b8639a8fa8cb0f5de46228f4fe2d0c7b4d38eca2b3d5468922f5d6f69f4284ffed00cd26d1d7a4b38474b7cfde0a5f4482f258d2c6c876ecbbcbd205d7f4fa431fb1939ae240a2f1f95ee33b5f30a83458d0456faa1dae3a65dddba09eb55af395c57abdf45f3ef2d702a7467bf2dc769347f4017e1b077ced86812b1ef3bdcf64af0d2950aeb57e469adf69235b78bb016c01b6ab2713c374b98388a5ee6ecf779f4efc9bb6e3dbe393a2ecef57adaefcfdc3365e09deae71358f2efe07634b727ca401726be4948d900386ae5d13020e707814f49233e1a0da23c4c141858f67c71d1f6e8860ea8899f65100a1ea70f138c9841ed4169ce5ab0b0e1fed3bc225637272d2e60bd415bd7f2b460398387b09ab5f80a646cf33975e8ad77dee27c24a449e6df42bdccc7c5a344ffc0fbbf86c360d53551658f4c33e05711b7f40af9aa1404fe0f24acb6313678d5d0f33badb98583f9b792b98a8b2dcaec9e5b1ca59df7d91fd7cc60127cff977116737e59f867a8df58aa19c47b79e9a742bb655efd2ee2bc121f12fb26cee6ce509a911dae23aea24c5011ada09cbb28ac67c67500b0aae29b145edcdf887df356adccba71fac660a111e955cb898ae2d3e44b22a7c986fdce2d4b5e22691bf54c993fcc04a52db368efa002ee248f7b4dcd6a27c0fec9222365478dc91ea1abb12c99fcb0b6b4c27800f3067bce776508ef35d1fb63b8092346003f20ed362a9b9f7fb164cc2e119187f35ec588252da1bb7f3d7fe892b769fdbfeaf6def35286ce94c8c584cb6775b05fbc1af22de45ecd24b6a6ce6d2033ae3963a6f1f16bd2cc9a3dbb875b2e3a3370c3beaa882fc796d61cf5b5a9ec818d2a9d5fd97b6855f5a7b73ce94ac102cc605ed89b8647ab80ad602fd405857c315ba85f67a0a2825314f2ed2028c8b2a19346bbbb0997cdd5d15cf2fe58b0011927e08763ae2065b279e54472a3a10a51291e32a990268a34e9f415711aa3e6ad379b2b7a740149e0df2db810eda61ff401af2c8bfbf6b2a93f2887af4ed528a2486f19f6fa95cca89be4ab7115996e1b9cf0643f3f1d60cca12d5b0364638171f6a90df0d7e25e938859b6d688c93da6fece5c6c1c75f4ae83ddd3666940253a77798bab156294707a60c54097cd8c16691b51d8cffa287ec0e6fe78f010b2e9bf54ec0bc8e3b4d461b243ba93afc8d53d084bfe87fadd1f7fe85ea92a1bb8bec57dcc2c1020ca79cd46ed93d503b0aa229f80e19cd1e1afbd8f4ef7c38162ac197289fcc7c1eddceca5022601eb03295d8b036f997d13de5b1fbde32798da7d1dbcacd899452993dfe59390cb3427c2097981bb857ab051b86b801f283faf8f73e4a932c4a601b2dd14c709e9494389cc16d3cb9a9f6be4fa124eea03957035238fb1d7ee3c1a6f3534b87317ea9cc5247297253aaa0b0ed121c64fd850cd97ce9f2699faf61ff70048ad67bf0b4fa2ab132de7e5c2df94b1052d1844ee864b2619365ef4010171c53295ce5ec2101c776a831981a072b2d52a2f05f038fa68c605af112dc6d1fce93a5499519822f9b55089bf92abd9d43fe7a2fc9c356ef606f85869aaaf6f9ac8197d8d07287c1fe01c99c0ef6514dd4e2f74ebd24337bee8cb81b1212e8d5a36533703faa7a2e0d032efcad8d624fc152d959656f550994899a54bc366968564146ecc6fca0351699fc0281ebfb4655fb01e20decfb30764c1ebc5234b3e55a342930e5f56395f2b31580ea790016a8ac6148d7f45ada35e8250b89c0b8a44ea2234595babdf67e4659ec1fd6dcf119dc079d10dd05c84249a7f3da9aa392f573bef9b43c057d5602a148a9d9c3af291bfd2bdcdb32acb78b39f3e6cd3b45f7f5a9d7d0b6d514235529e14749c8e92e4ab37ca5df306e3c696adc41a3a5658bdc95beeb35829f6333748ef021dfcfd2db72e0c769f83a7725ece666c57e6ed004d0047832fc6c9d38c5cab4610120be07578417f532825da92b8ca70ed9d1f75a86a12c7a2b01721aba7bb5c9fda4abd07a8b641b524251f7e7a24eb0550bf07bba738f063375cbeb7b066187461fb88dd82e28db1474770dbfe2eae9f11565be1178d28ed0b12412ecb685820f3eeca16ce4ff95bea8ecb85ad79916040c3843a026fc90abb924f92e911045f14614bd248b5184eaffc0d93dc471d91f5398700c35eb52e76b6b2e53964a110f9a303dfdf7b9718800024474be87250c19118abb64e2d05c903fa11f27247740f56b9e3237d4475a97cdd6864dc2851d9e6b127d9e7b248fe3151fa2131c6c1d171bc8005f147b26db7cf2bb5944d1351b6b8654e7afb995b98509fe91e31db30005dacba021b6feb9a0ed95d510f7ff4641bd42c1e5ab17165b2c7403e167ead12b8f9007055a1f984a9d327b6599ecff6c17925faaf7dea246a58ff93b1f423156400c9d364b29cd47470de23b49c24faddadcdad265ca11ea1410c79db97a0e063b27396c811a0017c82e71d14959e9aae308558ad0155cd2819ede896579fd1f562b3bfc34c9b98bfd2c7072225f6b833bfccb256f1b204472c3432a35691d137406e7fc8702d9b8b68689a48f67fb069e168bc6c75e989a72e9ff349410c57a0658b75716cf81133f1b574e99fa738bfea0a5d5e923037dc2634047ee6cc3b268066ed1d843feedf3e2eafa3bcf8b3fdb8b0e425a9bc0328cd464b1c749c39fa30f67b745241b3df929dfbb776961c5a3599e0c860128f08f70a5fdb15174c595368553f2b3af2c0a7efa268dc7b52f34d58f6a2247e22bcc3f09414dadba8cb14671701c827402ca0ff120b5d9e528aaf864f08f55cdd805e97b031b2e09b40a9b47455d08eee08b2ca2e0708e8c980e1892bc285099f5a040df5e9599bf43dbca4c4e3dab3c70d7d34d642e8f2379ea2b667c32f4f5a7a3a6cf4c393934d959395393a1da7bcd7118edf014ed44e600d65f2e644c1131d8075c6fdec6787cd0cd4b62ddc6795aed22133f1d97f299655d0fcd41bda01e6687d8433f7468da3654bdf7aa9b30c0f123e70d4a2679b8b31b6617342c9c24dd6a0118959e6a8842c7c93e702e2ef33ec204e51b4b958c4a9b182253869a000f5a087cb72025327aeb79774b002b24daa7585c5368aeef529fe95dd30e68fcafb8848cf67ca1b39345ba4597b9ea92fe415073ae2e89f651b5c48e13efe8ea1ea4798567bf936e428c7b6914f1d1ad6602b9411984bf79ba7734862d90a3af19e89915a489a67d3ac0251a0cf73adb5c60434b88592aec26ce6ca6b446d061ce5ddb262602e62dbfc06b5f999ed6e1ecfdadaa3b2737404dac92101a0d80d6ecac55f307174ced8b2d2681ef4c6d0482fad87b6905068536e1d4954139913c20a53016a48758980ef0d217435c9430b16ea633f74982d68b218de7b4b61e68b4fa1d5d609923950507e9c6a44f01debb23f57b704323ecdaaa84670315db6e201071fc4c75ad2fcd8bd40cc49e058f9c3a8e5b438fc53e7579e447f022b09cd7522cfe1ed0b108ff8c4fd5f7b746d5183da2d7be6b99603cba6cdc3e48b9609df7a447972a7ad5e3454c69e3ccf525c38b66c1a45ce329ab71854ab2489f6e4d3cb54f17257dce36b67be651f2a74482623f3eacc54c623d72dbf4d7117ae545b6d7d0e13093c15b9c57f879af8505bb05ff66f8a9d913232e79cbb3733a2501842052da747e5b1620e1908600f891c60deebcb52bdb913c262faf92dd5d6af254f36abb6f664f7000fca0bc604e046ab4c4addf92d6bd37fc0dc87d1c7dde4076d2130cbde8b9fe3c04f9c6e8ba884a3637c262bfa067ca61fe2e308f672c9fb8d627aa5e9d7a73a36293fe70054d3253a34e468990b63bbe693cca8552bec97ebb5529b5ed8ad317e16bc7389f6076c74f9ff1978e6d4fa9979318daac6a37e975be19f186efd4739ff1870876e8f3c994953296dc5ec8adceab5c0b9d6a9a9d6d80d76220f982fc22169026c4b13d1fc4d1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h7643511dc04fabdce250eab4ca5f1d6e6f0cc0ab98c2f4826194e1b924a4833f01b246bb7ba292203173600952d13e8ca73ea9480338d1265cfb92e92cc8c15ed3a01e15a74cc6e86e515fac13c058de6b6f42f640ef0432b98fb3eabcd292022c2fbf46d06a51b10566c5fb0ff8c13dd9487d808ec6836417eb543d3606a404b5774b2d69786a97a8f7558b422345e193434b9e781f25bda8ce664a6799c3aadc8ec03b27158bb30a873010869893f33395f8f232bd414a37d70475b77021db4c177912761313d395346b8c3b8c038b08380b106c20c16398195b50f77e6cdb2a3781bba8bc27f8a1038f77d3ef4223c41604d6969323fd211416b3bb25925cd9ca71020e1fa6a37f8a8c67b2439980f4e1cbb5cb726a892c3d4333c0101f8180e3e80c90f0068760715dacc719f1d05a24bdddc105ef22f4217aac63f6960ca73ce17f58db1a7bb743795d3ebfb559ae95545827c3bc6c0386bd6c8e4163b9f6181f04afcc4a27736bde49b5399f7d1d81a8862bc5b052f097ffecbd828fc37cece4c83c6dd6b966d09735e56b88bd1c58954b2b9e5b1136eea80367172daedd1e0f1eae7759e82c42d855c2abc8b6f6af1fb6540fc17f23d1405b3b06c9e0b5a932d4c10eec4f8f23b9d9484312b4c84d50ac2aa7567928166ff28f6dc195f3f2463ef750fc0125b74a883661461c831f3091b05f759f4c3c5e679bc12373a82523ee1bfb1a0d46e962d2a8bfe5f66764efa6cbcf977aeb1dc204988ac0cfad5018399efc49aae34c42fae63078fbf55237a6be8eb9fbf6a3d130d65b317a2a2ff22393c20204469416ef41762a4bbdb883f4e178f35fcb40742e098781d4c671c777fb1e1afa7bd67329378ca0d0c67ee528dc49554ca9baf55a7189c44d84f327776c023108cf9ea6b872380c5d6c840e4448c7554ceea4e8f655facdfc79a4fb3c747565a7a163a3c737206082c5b7c41dec8abf14fcdc5c792d5760aa1e553cfb3658b6c24fec3029a4a87400b7f7380a21c6df22b7fc0270aab8071207273e13d5e324a645b759ef66eb421401b2523579827956c8db1d2059d7cf02b47b3e1e760b3977a1eff19746a2cf946740f34144623a899382245c289350ec798028cbf0a19a773cf59940a902848468603910c3a916effbd81e9c1741104cbe08f0ad449e994e4197d952509146d6518c747982caa9787494a687ca81a16ac3544980ae846f8515587ad070d1c40eefd77fa9d361781cbdee776cc7115a4f2338b363cb42c763a80c6f7a91dab46def7fd544cd35781fe47eb17fc70de1301b9d9e7d09cfa08412ab9348b96fd67a28275fcf943ba5f1310322435f49abbc7ea2cca5a0b82bbf0f1420365556574cbdc883801db0ac8cd6b0e6f0d77a30d1ecd5e55763c858e8a4a796df47c8fee528acd3f791186756b07d928129fa1aa77d8a1a1a3d6def673964261d6cc941b9cb9feaf40117ad011601a6b32e9695396c1283f4c6f74ab24fc70c67ea0dfca45183b4d0cf4e63f79f8efcff7c1821a8ba76c011e17955ccb93298eb25cfee385b99ff64200dba1665253818dde65924f3e731f706174c52e4e53d7d870e293ed8179223b111d6bd3106bb23e72d6e667eb8f23e97cbe61ecf0b7d35a3860be4fe2e133218d345ce3b9142c8373cdbccc6190851a64f5a086e86bacb082698d37fc727205d7e8d48aef189a9d791eee0e8debf7dbc2901b8d237d08bf142ddde373709e50f20f79bc9b976b645272073e541b2a1e4e25a8e8300e9ae6c19ae0985c081f81cac623a55ef9b9d049ab1b46c90f863b09a3854fcbcf897d26adfc1e7031daddab813b6f6b37d8e3f44c327ba7cfdff7b6e58d6fe6d53ec04eaef21ef282e773cdad2c92177af343d5976fa714c14a5b11b6db492d9318f080eadf1609d71756faec0132175b8b0e7e79bc31a45f6cef082238b908466a056ab166b0b5e4f1047c29d83da7d38c50ecf3bed905d00b2053b6862f7baafb4af403f1a4080d7b827c69b01d5fbbabd7f82d2d7f561914ed23b627f10a1f316406f06bf269f91de7ccb6d7d2007b93c68e8daf45ea6383cb7580a2b9cca127d1d435eb7aa90dd41a42a94037209e219abd18963e9ed347ddd12d63aa0d46d88db59533f79c59018f69d6a986f7827615a7f50099c993a035627d5c09c8fe4c0b0dc25e0a58e17eec767e471a8779f84cf4dbbab7379a7ef76d4d2a3cfe60053cd9d5cbef216dc8f2acbab11baaeccfe1adc9a4d9d492ee0c8063d69e1ec32d3747e3bdf875444a16e720aff9ff691b131f08669baf83df3e44e21a9330af9835f5f2684e4fb8c0fb3538089aeb5a9de030f2bacc1b57d59cdb0b26a22c8cd417390561c4092fbe75779e84cdecfbdbdd9049b2c73372f5a2720b8a398b81e83b444a0d6b675e0695077c8e297177a7888d5a7c704fbc004d1e1852b975ea24b71ced72a123092d1c5be2a07ae595f2d06e3fa91102e45d7aa2cb2d8ad9d0d1c23a9476c2f2c15bb9d625ab6d5a1c539c986141e50b6b434fe0fe2af3ea61c5c0087dbb04799d61c7a1c7ecc67d03da9289b60917059a9822f5fab56b538a93da170f2ddae59ef577ddd6a238134c1876443bccd7b17d182b43cbe80baabf9dbe8d19c9afd86078e37dd146113e86210d331d4837cf73009efe99676e05943460e0007fe63c7f00e4b7d4cf8fff99bfaaa1f6af4a12091d44d87cc99d298f182912ed13840b0a64284d24e155425ab3238bd0dabed85acf8388a28bc59a648a87423da5429f32d5074e21146a8b17fbee32585bcf6169de850e5ff20fdc7db291067d08927ec8f2a23163071dfca8897ecfcf05e2f0cbd923be9a0e05b22b940e130e74d0fcce7750cc484ff3ba71a15cbd97e77ed7f0d540bbf9559530d8f572f478ed5642c1deb088311afc034b19aa6991a6e33d01effdbff44fe3926ed88a226fef2c69eee3f4a5265d0df850835f230245ba6dffdac54be8b695223d367b458aee64025ff3d5f15e539cdab54c91181886a9a53c3f56daf27e5bae9e8e9881471434f5cc4f4b791f543090d1ca9b64d090a6070d6067b38aa59d6913835f9f6fa3cbc6276ca9cb2be38e2e544fd50656585d2609dad61a7fcea8ab0bb80bb8a3e330fdc95554adc77c6f4d8936bea46ec687b53db0236d5d6dca4588cb74f5e7ecfd2751e660e3eb06db889af290df4422226ea337ce3b972dec4de4ec7473ffc97cf2fac4a589d509043304151017a849aba26f5232074a743c0a07372aa53a2d63b881a791e6a8e54440d24d6dae7d5ef496035a1c754330db4a148ac5f34f9ab20f5968ac6ff7b46b20803602e17e628f6e9d8badea0b32b7e316b9adc3116dee1213bf06aa5459c840c9d08b85147380066e7e2b56c08d35c68d4766f38de922e022f6efe5c4c834fa85731fc35a1dd3d208d6676242f3d43d7a0599eaf849baec68d66436e637d2bc30bb32575b8c889a4ae58f360ae0633b48d2a2930e5d43aaf5e6c0a8da59dbba10d4999750df0c4148b2c4ed953d3d5ab63d9de6b583eaf55f49604df7ff3b7bd8514038d8f0f97f2fef3a7bb5aba2c3eb8f849f1613c5be47233da261b97c447f92fef7b6984bb33834d005c64358d002cb7c86caa5f1d0c1b860cfec80a55ead0fa6580f5550a8cea5ee54ce7a52ce22a82945d7b12428611e8480469659c456512826141fc0516e9630074346b3b6fb86f257e5be8ac352718eca344d735403ff7374fb7be0ae9e6a48a85951978900537bc70e07dfa3b915c027ada3b4aa5c76875e95fc2fba1a04215072ce9da1db4e6ec1a36014a0b5dc982bc40adbe95a63652ad583d46f733ded57e44c3adcd1207c4bfec4157bb8bfd5502d6e6776f9b1fb88b745a4d487a7b3e8a37ce87d9eb8e41d4db69da1314128106748e74e76be76f9454b8ce870e66406eef461232430b84fdf28c847a3ccd1d95a4dbcfd7f689add243083d48fe9838a99517fd808aae7005a11d71ec8920b5a4498ddee685a5a79b0ffc50a2ad8311f9c97a5bbf5dd78d950e1f7f4d2f08b481b9d74f312568235081842767b9477c6d51291541a75bffa2a93fe820ce379316b13d2ee8a3038c08ae14cdc634e1ce8df745352c42208d2ca529962a758d6bbfb246ee44e4b244845aaad1ea67d5c486dbf30c81aa33dd32d455e42f6b9481a3efc3178a6c6fbca73d3cf35b3673a45a4729bf627e6437dc5566b4ac7e711f3a0fc741c8055257b5e5a4603945d887c419d2d561cc7f8ba01c7854d21d0a7bdc13808863312cf5c63f62eb58dd1d9dfb36a110a6cd2fb5cee299febd05354cd0076ca7270a9ca937a352a835192f1468d18feb27bad3e9bdce66dffd3e70eec1f4b0fb18d9448b030645026067230ed376616d42d3da4b24f41956fd735a2e45aff980a7bca229068d79076b4a423370fe32b8424d97b01b8fbd6df2c8f746df83363c55f1452f7f9646d930d43f117c68277030faa078f8472a0ed398bcecc2c17c79c40f5e8aabd0e5d8eac969ff3b08bf5fdfa3bade09ea463b379cf1dfc0e81b8fa9eb911e8f702361cb3aacea73a8228296a90c3f18cfaa720c4a068de36f58876a98d2d09a7fd6c9d2fd0beae16b57a4ccb3d6186712f2f60f6c9c525047a80341468889a53c308ef1bcf91e0610852b3072ac0ff6d71aeda82d078f58db36172f21cb228a52cf9fef4880528d6b1d1d78824dfc0dba65269b8b8a95c01313707a25ee7fab425f3550e9fc989f29e40f1eb8902c106c42ace0c8104709a0b469a7f3076252e06dea0a97100ff1180aff8476ffa3266b0381bf1fe339455d011bc94ce19bf35ad948ed8f44939f530ac63869d9c5774a6b34a749cb71b08c670cdd2d1a9ce78ced8b022e3c84d5d76d202d51fe522ab4f0079bd84ea531677e984b623e7ef7b3850348530bf7f2cccc16176331b9f93620364d708bfac69e7dc65de36d86402995650b84f53d1f039e35fd741f7930d971cd881f59d63874c72cbd52954d9d67ad07de1a3081a18c2abbb93805ff2f265220aa422a65919b7dfbfd7913e34e546a477e674af5dfb2d04cf3ea73c26816ddb7b106f676e4abbd8b59f0fdf17113c3f6e0dd8812eaea3cacc692b2a488b8fef12c34bcbe52be3c063e436f6a9e5b0e6a979cbd1b48c4a32ea0bf9fc80d9e73cf6182a83824db53eda5f1fe090775988ff29be976b39b71ad8a08ec153b24d072adeba0049fc9929e4916d6de068074b70b2cce614ecfa7b8ace862648848f418b416c8fbe9ffc4a9752d8f6a9efb5b43d968dc5a191f86c26e654202cf9991baf090b92cf9ed4ef856a400255d26487de4243992b352e71d85b2ded2af8ddbf58eefab0add6a74bee25e8d0f9ad697f0fbb6e1c59742fbc3c1916faedded3f7ade87e51160fcd9ed8b0a78354e2c8f06d73db4976533ee62e63c4bbfd9957e95e7dd05b592e2cd1a79778be5d5e3e9db451c8510d35dcab08db3887d9b0ee1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hb672b7c5dbd0bf761afbc2d655063a1b85d2282be8975b37f581777c5c0f74ce7d507619ee0d977c9864098cf84c52504940f49e5d72b119eb98a7a4abd812b305cae2940b75a565457111b0d1d371c4d7fbe8a62d83780dc838ba762680a404610ba8d7e47cfab587e04d67f8fd51b588e62d0834cfc414aaec19d5d10a4f144b996f73df8c58376be5a638bb2cba3ddb82441978de65e291fcacb4b699b9eea642faa242f526980b9780ff3dec919e5c87bdf282f3add9a84b0c834d1f26b5dea3462f672a98706f3a00a9ea99e9665c4863b9479a8cc13e4ca94a98b2a081659764ef6994570efc29cef7da7a42df862eb72e2dee61a98742cd7cecb837cf350a3d75e74a062004e26b159fab15356782c2eb4d39581b9a8bfae932e35a71127135f35333658b8f333accfccd2c041452a385f9fe0ca8fe6395bda3a01aa5ae66b2175edd44225bb34f03c306701c26664210d89158583535bb21ea1b7401a6e206a771fbfce7dbcb194fe24dbf9655f101bb3cc07ceafab96263c00e7a97a490416506fe56a92d926835ab96b93f1156c5ea074903e8eee901b40b7f4427ef5a8d7e47ee791bfbcaa2d5cb544e1798cdac7d3a0b825804fb878f783a867f64e1f140323e3b230e5901e9c5c4c722c97387c6acf860e54c44d3705bb8a946807da889f45d07e6ce7d372a2a308a53993f692dfe3231a404e7358af615a6f29f8c93ccc44944fe3b2e3e846c84c8617de572dcf657e3fad6aae878f452a0941060130f66f8b621531c5c7ad2be90caee5c37058c70c77a3eca104209b8c48c0c3450fa6bd5b6cf82458c8337aff81b669e148f2191485c11d3e7e9027bc4686afdb5cd04281c87fd65326765a57b726ad0b493fe48833838205c410f3efcc258cd1e3287df2b7bb9b96d2ae4258f4170fbaf4548160cd6f6ba255dc80e5b9a5f094ada571338a6bf3f38db6f3cb265cc7e862d121e8421988f8028333495434a64b1d09cfa4bfc824aa6b26566505bc49ecfc6de8fc5d229ade4f19d66a7978771203cd51d54db52c9d15bd2fbe966e1708591a9a2b85958081c269d92a6d57d3af4915b30c4f271278a86bc58cfcf38cc4ee83ec60772996bdfa4051aa6fd8cf4da8ae993c1d7df47796fcfd74fdcf447a8f347c539b6b052db3f4e5c119cf8196f8f9c2ea4a9ccf33dbd8a6b50b00dab4b711c0bb27345152139d3d43fc508ab43df9efad2f1eea2be5ddee3f34d333f975bb2f65adc8fda638ce1c54af74cba459bcc06342fe67821b1a25075186677a088f9f9ef1b82e864926f27f280f4d9530cbdad75187c3602b3b1b600a6484f6aec014e81aea4ab437b70ba6da7b0b800d238711902922babe0ca4236b07f63037010d55962f03dedc894bc66c9f17217baf5bc097e2606c98678848243fcef950e26e9acd2798e50a072d21d1de9b5361e8567e268b3c965d8202faaa46d12efc92c03977704e3251073200b603c4d3852273dafb266b457d73d286729328184e4a8db1e7d8db65cc31a752f85dec77c05bedc2df01e5cf89332b2c25b3a3c7389b9338ac66665fdb847bd7a10773c0d4f4b7155a0c0f31b6e6d8ba006070694428b13bc477592dfb97c3bbd73cfdb57779ed76155bdc87884e1ba9bfcc133af11b835031ce2387db368ba0636e8fa836780ecea257d2d7c381dc7466a0a52f8747b72352200f8923501f068adc0a0609e2566abbae12b556d1d53f21e453fa1b47a9648ec24b88597cb0d87e953733194585ed5d1b6d2af79e272795b9160f1e3902d9011c78d44207a8fc57bc6828779de51fd78a86dbe5a5ec2e5553733f0e22f19a6922e86d88b8f16a8ef6f24d0f8001a69a381466df8f02c2574fdb3b23bfea62f34a0e389a0885f7154c61784354106dd2ff1a630d87414b3798dff93f08ef9aaeea0269e012669de681d4908fe9601b82c038684a2e132d4d1eb46111ca5042cbbf17d77cdd14f40f33bfb14de183f9293d79294e6b8ba52af42116081cacb5e8f076970c17d5680ec81f0cb0e85105fcb4ec29f09dd45fa310d0b1c627f4f306557aa8394a40d8c1f6db93c053da3a9bdb7d4b0a12744c56a9afdadb900bbee99f02497e2dee8724e2bf16396e443941e1068df40629d4561b0a64821ed1e15e355a9f3d04cf3a12091f351ef6f0f2d4b47c7b4381448923afe520d83f630e9fc2670bc0b62ebff0d5b3359ed6f5c4a40ae698112cf7d6008cff8bf4f956fc66dc24803c2903832014511421234d7b098fffd03f5def66dae7ba14a951a6812511b066fc24fd1e8a144c0972d220aab1db1cf4df17be8da925ed228426917722608cb4ba65a02356e376ee1b7be7edec99ea8faa552f443cbc03e663754c33dd601170930f6917e63f42476e1e95805f4fe13d158804aab1a282ef2f78473f6853999d641417faadf013f65a28d45a9102506d1da0cda598fa0a24545728a6aa6236132e181d86c8b91cd5825b66db23b762c4b479dc2f61e5b63ca0e88bb58d471d32b97fbff61255ed43e1d662875be9e3ddab838c4aefd0a985ba6604a55ec064f8d03351f7c05b1da85a5676e99a8fd5a42486137a9cf9e9defe8d2e9807d3cba389b2abbbda4f1d0c81abc636a52c5c6a58c95536ec9741581c5ab412bf18a3065d8eafa8336b2cc6b13e26f6fc1f61273220af9ac75ac8d99566dbca07a5caaa29dab3a403e5c3d9e265675b603bbcc4aca4a8ee46848a44d62f03b7deec9a64650a3b2ab70f304f9634e999213963227ecb0e09f3f75725ad9aedc9f23de46fe4ea73c765597b591708296422b85f2df66125470ade3d62aa441bc078845cbe7e9665f70274d3abe72961964996d4165bd92cbbcd4bbb436a47dea77eb97c148d940168bfe0fa5451fc6d456f2c43906bd8f7ce1f7db2bdfe96ac299c183fb5851c87b4b82710b4ada4168e0356197369048e9bbd90f74eefc8d9bca98274264913191f8eaf2c9a5628827626fad00b609ba54c99dfaeb4cc1e42a18aa86deecdfde6556d3b4fc70e275e160ee90565c69412908af1bf4c1fcd4b307e7591eaec47e83d4bfebe450ed769baad4ecffa702d0a1f279e45a94e8a1e82486e1c795422d6f103e9ad353bcff4611d218b269f1dd07465072a8568569619f21e52021f609c1223b00f38bec26fb186b274ecf9638909bb8efc53bac7955014dbefd79586d4b9c26fb8629826f41acada2e4bc005e44fda17cac6b1d09820bc0383ce215b9ca0c20edf868b0daefda2f9ca3cfaf7074b264dabe698fe5b97891261730ddd3d44d1ea469d0e58d4564e1d815dfd8a45194457076fb8e8a94ef9fcd4e3b8e312c5109e5186ac6d0ca7f3b2652629ce51a6578b010ad46bb77e39657a373174d27c382e13dc5e3dc15a2c135b2e7c43e822c1bc370393abb3d71b51cecca9ebd35672ff409d36db419b1cdd7e07a8981f852ff4d0922776ab55943d1b152191b24fbeb2750f4cb368387bb780c250f41dcca4ed0badc9a9451851e808f590f0a36bfb5e51b28fabe8c8c38a4ee8ddf792eaf74ba8418f1e5319100b48422c7fe6d55847ed1b7b4146d314a9d7f5a680223ed87dd591ba5a228072101aaa62754271804521d72a7b025cf6c34acb557fc22dbe6a56c93cc0156f215005d9b42bba80485b77f86f244d1f15b491a99553430883c9aa1fc810fb938d15caa0b53ce80d4c73d0683e0e809aa7d0916daeab3b0374e46c57b0b2be4e59532aee9dc6075bfbfb2aad2fa388ad093a31b21d1063b4d181e1ab8b64bbfea50406214e7cfb05e9e48b230473bfb18242d1c05852cbe6587c8cb0a7c4f2c92923e792f60ff735800298e3021eb5e9e2ba5a9dc5289529365261ba5b2b0073018d785735d99064399c65d5bc95611c06e21100501f7f720dbdafbdaa6c10acd6948a6c3dc81ebd381141131cb1abc995355d04c1f8fa69cfb36eb4b6b7c58cc1b19ebb13c8d1e3acfbeab83f7084cbfde6f29e38366c6a4659123e1330a1b20403f7ebed947ef775879e735af2e1f1f489a54620ab7372872bf5326539bf2c82c6503f56b80a5b5e0c8403df2c0d32dbfea604b7898b7c195bae254bd47789d09fb559a641f1b0b6870fa8743c934f22aefd2b853fde904e1e3a143aea134e472c72dd84ba449c68897458897cc68edd6000a5bb4fc0893d221a4738725f5987503921c322e832ba52f6a1123369ba7aa57b029e44775c74a903d670c70f89473b849c86a2dd4533aaecf2a72592bbf3c1992fa40304bf0ab92b6d797678986d9875bd9b74a7e36e34f4949ac30bb2a2bdd61ab7d52cdcdaf0ae86e32f3948cbc853d47b1c25e259d68286cf3093ca605532b50ef3a07242ab9e22e5d4441fc25593e8196c2b165457b0b8f5a406faebdecdd13f49a9ca5d13a5c46f6ab1dc1d7cc55250f60938ff7c3f45a4a0c471df8a23474b254df17bcfa486ff713dcf63fa9b85edea9d51f7919d2754045c7db35a910862276d681dc515f43b72505ff9f5040bc0b9e0b8f3678ef37d7a93c078a9c20e60af96de62001f6802476ca06b8d22fbe92302b0f1a0f63b69ebc87feb42e696b83a973b59be5c77fd8dd78d0a9f1895c8c6525491b335b065bbb21fb9a11541c9f13f61a447ced517e417fc4e798d057faa6759471e71397c8edbbaa20430031cf45b14ebbe80968c4cae3c1fe021246b76e863dc1daf3a0a349a58170972145fd78b0f561d20f05cda0c9af8a9f4f07b910ea5d1f2c6922ba382e18066d03ef6c9adbe4ab6c7b8e9f76ce0fae5b7538bf965530e6b426bbd43ea0f58b7d73a56461435b7fce83135e2660393d588a8e1e51951394f6da42ddbcb4e7cc2906463cef3dd5a476dae5907e9db903e62ae0f0a03207ce7387d1dc17f8b17ba243bd6b80f029eef2e07a562e8a7c8b4daf2af89428e5c2b1374085aaa1ad9f68ec1810a2dc8baf9d1cbec5325f0facf6ef050993ec0a98addd6983e8bae13b0be25e464de46c5bad69aa62940d77b81adb86b415aa2cf5e3b3039d6d08678d2ae1f14177c60bdf996896e5a8e3536b0bfecde846a9852029b15b5338d4dfe0db394d056a77e2638cb7e1d3e793491968ee221fa14ab88d325e037c72e0d8bf844d44892a686e6a5b5a34ae2310ba622be888f4041006c4aa1f36019fc38dfe91f84896ba25a20b20c0f6a3df970fc0ada627b3b0dfd450548ae0dd41e10c6277d77c52596b03950b494c8e6e8435e98b2e32690293d5d8e8f0609ea673d0810d8f32348e92d2545094930d52fa3e723ab1c600901c765d043528905ea17525e64ee8080ac29f79c99984fbc4ad85c88c93ae7c7f7a76ce74c7a2068a60497086bb2f9073f47878f789d55a5f39449ca218f1fa73274808864aec0799e80448046f208aee3a1a242f37f457f69d943dcc751b9058727ec599e66c8daa7a24cc296de0ec74d20943386981fd71f98c876f3335c8e38408ca9d756e693d8f7724b79e2fe9246162b4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'he3689f86a65f9510be3d63c33da202df79cb2eb8d52a711a25ac5fbc50af233093b598a2a0779e83e512e9ac9efc0d125fb6287de6489b023832fdd174db1c5ceee0f406c6eeb2c89b2fcbc8cd9a6ac754baff79b346e70decd9c04a6a2c68bc9716539e859535dc87495c75d253c5dee72140c1135cb38b56d2d055d04d8ff002f10b6f36ce677745becbfc3e3198c1dc0e775894e601b73f99bf195ed5ff5a8eee0c591cf7f2e4ea271facb529c348af8b0bd18125ef8c3f58fa1b78ee348dc62af44731a76504b37cd22f0d6f2aff48ba8f9709704fe0573796d0087097b1864e0f500e301cbc9d8e77eb1c9c4e4b9a409a12645e1a6156cb041e948740eb7556f9e6e996c56b37fc456e7c1ab609741b9c171fa73b288bc25ade708a2f295fdea4a66f233460acb7209339602c883d5859d3ab70dd9cfd924f38e44a575ae946b0b5725b79929bffe9d22a69021d06e17ce16999ba272cb219aad05145a752ead1a5f4e782944f5761d31c33d5ce2361e0d1c4c6d42d96cbbd73f0816690e9e9e1dbe28f87693d1faeacb1a091f97bdc27582174ea8a0a29e0dae39ac4bd38b053ca8b2eb007940d29b7a4c5cf8b0bcba04d00863feae668bb2395145c3b1eab4a832ea96990948a5d74f8c26741ab2b60954b02988df38e468f52efeeedf4e17cb78cc8ea96ab31db6c0c3c9334e2bc5498e487bb699d296911924855e039d240ac33ddb2187583e2c33a8bfee767df35c77f1183560c22fed4b6fef2df704f63519e4f14f12348e9a3c404be9ab4d01e72b474a1737b8dde8173dbb9c5208074c25f84ea8e3274b550e2470dbf81cbb92e0e78b39e052a2793bca2a9499f02f4dc0ffd40db907bf8f771f8f92d5aab71501e0a8b1ebd7ce91fcedf05a9e3c9a2e2531215b8cfa6588c8d8c7a1661c0287eeb5b99476f2d7a1932e6dbe4f5c6ba1dd9af7b9466240c332ed8d7d0a87255a31e0409f5ccabc1a785a3c5bdce1ef324a3d80ecd669c45bdc70e4b4e675917818749224a1f45f4a283c2ac582855b581710f48a613c786586a2a97fed2562cad4fd85fcee75f572431d9f272ed26af899247174e2ea03466aac8d95c51f1df4e81fb9dd1fb92bc4cebaed89b21d3dd20fbe532440591c15ae89990cbe90e791a046683d344ae57bbf8b8b6662aa32124c43bb227a29c57f93b395a8f459dbe44ec76f7c550a9e16ff11e20bc542986915e5d1ea73a522bb0f100c5b14725b020aae299fe04d88ed5acdb48fd16fc17b3d92bbce49c177d70697c7b642ba1af4d0d1e902c5447dd1d97c00d3608294470bbc3dab1ff31e4224188864dd8c6097ff37d04c44cb0a13d11dfbb06c5d032ffe5912da4e0bb7749e168906cba3b55ec6f5db607f16537210735dfb410eca90d85567eabda9b22132dde4c6acc3a28a692b04052e11b2d87e054987f59c0c81a55aa988091c183e9003f11d26586b193c3f8f346bbe2efd233b30eb00f77dd066cecd37083db904059f17f9cc932030ac911533d6a5786ed224b1bf16db38a776963a49a6297d2aa82d6151554d4adef77f09f8cfd3cc528704cc344a0e1fa2813c2df91e6a79e697a8efbead52d4e1b9b5f56c77c1f0e46ecdcb00be3602592b9cc3ebc2372e2fc2f9f3d6905953815568da929d5bbd06dd18e2942fe715f48b862b0022e0be66e6d6fd07d86c247500f06278d4ac5b48ee07b24d2bd6d7b0f53efa262fe1eebb4bfaf5932407606458584b3b82f688b64b46617a58c798ae5b18828b1dd1226e8b1ecf6498c1a82fe92fd97774a9c7732594f189b3edffec00568ed634345c78e99405d152f350355840a36618f0dccb1c62f5871cc4d19a89d0f92e05767da905fa4e74cf993a5d8bc0240036a11a14096c67c000f96a80578baa051250388c3fff6af8ea44895d6ae32390098e018787034463f204c6001ef65ae8985feaa99d54f2cd02a563bc52579d51396ee14350875c060810d4eb055ad50ab461321430520efb1ef27c011b393e4043282fe2d3d7543ccdba660153b35e4fb6ac1dd644bd9f2509dbf3da40ab8df79eb44202cec8b9f0fd9874537bfedefad724c2a8269ebc6b2362bf593fb1ca729e7d3f72e543f3b49f03a638bb680334b8b757c647aab82fc77c5bb1950e7fd4974562ede8db9660d56bad8d80976a7ca03e3dd4505fe98e1965296fc8fcbfa8eb187f26eb42d6c94e3eca44eb53b413b714f8829be0f93e0746f57a1121b441b0798c26a9cec9bb4f4f61a4a936b536942c67b1ee156abe5e77a2bb86b38b726a7e7d5ad67abc443901e91acbe25195759fab182a88f9ec0bb6a0938c15963b6ac41a2c2462e3d2e94acc127dada43f7aae99a0cb8df25280582af160df147dab598f05085a23a0b1dc3de0e321e4b572bb84ae3184469435cb1487cb3daf2930181907313180ba45ec21d60e298641191d5fe5a90f5fe35a79574921b6fc4500e2b00ee101a77ffa39138a90c27646a81ed3ac78a1795d811f8ba3d18054703645e9e4fa4c425ec4cbef7addd8104a9e52e8b48ebbacc8a3448b289839ca8fc617d083cb57987770f4118cf544cf135a7e39d8d8333bc99514f7fcff7bdf46f87510612f2d88830919eebbcc1f7dd72dd540536625829781f7ebe894086eb7e8d9e14ba61f88d96077c296eb54c8e5e699b3bc157790eb13041159edbb6f76a0d91fc4060851e62bdef0561fe6487ac82a9beb6bbff673879e2ff10fa2098d27c9e650d5817cad3b76fe2f6aaae8289b58cd01d9543e008a71810891aa5dcc219f20f1c28c643d8b8fefc714be052a9be3664568858fc8e8ff537092d06c9b1a46277b81624623e1abf3ab6d324b08d82f51b954e1da8720a77621e9e492cfb745783277e446a78115a7468b16896fbd61e19489f528c059e3fa1fb8d280c91d45d9c9dd24ba251dfb79b5430784a244412e269581036bbe63e75bcc17911dcb13c30d898806b73e09d8e843fc275a0c72d808049a30e74d550511b41e7f411053c99c229eb4d2b04d3490b23e14e8944dd84f619883bdef0ac6929d61f777b06c348319eee176826108774feb82a844a52706d7181021551b94dbc69f2c120b253e24adc90f6d2c8de44a700664f1aacbff84543cee36cf7bc5e0396ac2f52ea25feb34c01355a58027e2d6e942b85c1b52aaebd0d007eb26429b2a7fc6d001289d909ba1be0cfa04275e55608a3f5de44a10937e4af23e7e302dbbc3a0a0e1911741fb2714aceb7eb2776ca22d346b84e40715024a3e8d3f173049ab348e3bc4136286b418eddc119f3e784c95e5d1fa2113a7dcabb93fb440df0bf6176a66c81343252516a88c6a630721b6489283a07c0819b2d9e2d8602c1c3fe809c923889e499e775656fe1b381ae19701ae10928a2417ec1d84e2c1df5244a7eb14de9d95c57a9726f467d9d896856fe22ea4a7b649e7dbbae886a219f112aab412b543cd395e2d888bd85aefe03ff19136218cb8e5f8c889e57e083beb49852a7c15073b088f908321e2a1979501ad11bfa5701a5b6415a28cf32ef417dda0a82bdf78995080ffd54ad9ec48702ae7d897956c59cc917f406ad0c78b93b7abf4914c4bf47a77f3858de8aac209a4b76c07bc485ae019b2464952c7e2c4a9fce8fe4a74866d666e2393450ca9b91de3edcbc659cb8e3de6966dd14bd86d161d9607338f52fda966578170734d433ff42a686fb2071873b1f6a5b62645e20773d3f354a3718ad02cfeda48d11b1fbe0d38b9f29829415015755e6a8664da548f80f2097f8be1e7db275a5522584e77bcb0460fa65da9e3e05034e268cfd6932a6c4d0a2b5c66434df10a291a9efb9c6698bb9166d7f53b212f97934936ace90ccc5740ff1f6286cf865d65aea83d49a195531d40aa51ad0c85fc01b782f7547c28e0a2922b7959bc0259ff429840883048da4eb663b95ff2d014a09ac37507b3fd2c4c7b0dd09fa2b7f717191c14e6b05323aefcf9281623d95560eceaa4640078e39726847253423f9c08099ae1e720b551ef1a98145f2b9b0ad2ce8c86d547e046e46f40270aa738b54a00314a4af03ce5141c8d6b428c11808fd2fc712918af805ff3f2879a538d3dbeecd3ac154bce1c00ef2c3c122d297bbe51cd983ca35ea12d193bc9e5846953743d9578b9ab94a0982e05fda6905b08813231bf79cbfc157ddb5071ed1e7eff397fa4705127836441fb21695535e615044aff3dc10d608820126b2a211a286395ad54cc87d96b2e3d90efbd315038611638685af3074c948692e9b232729d60201fb193fa4c6f2fc6597512860dabe72e48fff532a803a49152d010f924e2dd457186d2af322df8edbfe5204b4343aab7861c01272813d5696142fa7ef58ef4210fe6435bf273ee87fb2494e84c87d81d03e5ddb49e68656b13cbb1a0ac7ec3f38a17a00fd67c2ead0ea23dd1c9d9616885a7c5e375d560be5801cafc16ccd459114ebcf1e5f6dca0fdad6a3cf3d852eb206fd873c8b3f5e06d165c1870214e6d9ec87c1ecdc4941c04b64215a0c286c7049c3744aaed3e290e74103c476d472ca2857055bb17dff44d0baf9ba185e3d362e0e7189bfc499d1c17807b56949653ca47e68f129c18952c8918359c004c1ba23d5b89f41d5a1ec9186dec1ba25715034dad7324ceba4250e86bfbfb60c9b94572f211dae90250c48445d0a2a0291f657db294cb45a9432f00377dbe2365f065ba93da6a84cf58930ed4373adf4f5c10ace36ca6fbbc43814dad6c8f75855380b0218843e1048c6b75a3d5642d6d221c5b08925aea4a4ab99f345d10fc0c92f480829ae3c59dbd6d13fd2c94c4e9fed663ef0a61667d89c1f2d541e21d818b4146196a2948c181de66ccfbdf0aa379df9eed3d50365b1427744cadb1a02c1bb20a698c7e390122ed04d9af864e839ef8da410164d9d761b73cfae49532110b51d331d7f9bb48ff52b50b57310790c3df654f85f5057d37d47d8aceae191e3624d732ba05391173649d1570daa37ed2b2e8bd0b0a7c3016b365bcdfaf187709d9a911bb2005e40c9e63b09cff7cc69ec0f5d6f331b05aa6fafaef8d3696381a977bf0ea361140c857e71335758a71ce9fecca871820fa0411c1d307b0a3a3198e36ff6d368e009f62301ef6b8f6c547d3d09b8d76fc5ace17665c7844b4df5c301c0b50acc9ed201419449840c4ad562c27670fbffcc2303639eba933640ab6fb955b19ac5756fedec00e76b90c2745bda02c8a5abf14edaa4d91286e60a2a72ed4b77116ea157ae68ef735125ff46b46fbcaa89edb749d23a437a706795cef8a27cd957e6cf064fce7a10976c9acc33fe6f3a97e8be7dee3a28ab4d05eb1c3c4abf755567a4bb0bb6845f28a0fbf28ded4464c8c309d1d1b846509613bc48c1ad7724c0eca46104f4f5d9ccff638505dd27dfa0f7dac511f6474ca54ac5485acf12d35203b7ee3b1c5e01eb1d6757fabb91481a08da5dd8275a2b2e48a717;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hc6b409e7f02bf4aaa7d76b40a6675f5efec56becc81c2cf1c343f8fd5dcdf202b906f7ad252de7d2be8f0cd82da44989644988f9f7a69d4e02816a93297aa94a55f8a51993d4099d338d2679b633a4c2730a9c05a9155eca5345a0936787d7aa8f0f4df23131bd684c689312121eadb6c4cef4343d767906f3f44345ad878fd0613efd3c90b0afe3940ed43ef2207d7b39d48e5d62362b833f0d65113f3285e3faeedc960dee5fe3799ae83fdb35a915163c5bb45faea8e8198d4f472005cd1b15448fd14c61725be9c30da8a2b5b9b7da81b3f110f42861e017a8bb4d9f519b8f141da05fc211e3ffb98e6b84ad8d4dea162556d30b657cf0a1cdbc9135aa2a4378183488127de81a92ccb80d6bb90d0a58b4155cccb21cfd5639be4f7399a0cea5191a6de028b84ed559ca8703968171717c04ee596933c1d75be38b03e2317fdb77afb25252574a9b18eaaf2d19ab0834dfe251c8789d3904f656abe665108435d28f2143fbfba34b2e0483684f936719a467206c63fa95bc430bf960de6a51b66d7f8f50afccc528eeb43b0c2ef06c77b5aadd301f035efdc53fd274729f63fc5957b368a471be1c77ae7f6a3f901c3198a52ea88b5769b8c25660b605c6084e0d5cd71b0ee7c7932632cffb5e51fc88093f0e558888b662ab7eafe11029e0cc1270a35a76eff79ea286b0978e56469f0fea5a7b29fcb7c413f559218e58915d339958f15fc0229dc96ff36bcdca2f39e2d533e232b6295778cb800ad24c6c87698abbd000ad54621fd77391df44a01f36dcc9825c3f628f25d36735ae5bf68338e01919b95a7e331e6097f5b1e36d6422e08945beea5bce42c2dea7b5161d9a243b8fb636e6cd2f8259b2de68f1dfecbf251b156e650785cbaf6b19d654def4b232858857a751cb5219f1483134be8b19acd5afe7ba16f064fead1476fd4352d4b69ed9504906edb7b0e4c5aba25047c04635ef0672ab837ea10cd6ab1f331f09b54565e405925c2b75f0ac22f6c3de844208c5a9ae7ab7a50eb4bc5cd031f13b88406882e97dcf75be15d04764aebebf82be65eafefad3c1720319f0ae52a704a73168ab844f01d1f25c43d1fbdc1bbdbdd96107cf6b252b3cb17055ffc22a8e6563e6b268689367b0a00c915681f2d19dc7eb5872e103b50b7f6cee77efce2ef971c8ea75763d207db5729bf4eddb9131024dfeed32f8461c883b3e71af0873057d3f72f13088995f98566bfcfc38967a5a2a0f37b573822b4713d635757946dfce134fd75167ca3461bb71831681a04e2bcdab3356c5cbc8798a462b6a7cccb0833820031c95d4396ac755040b7ed53853aa081ba571acdfd7893a4d836e934705f67ba39c6ae6da5b65706394198a7a8777ba561145c89a8ca8d2dde58db5db5aeedb5a4acb9857936732118e4a1877ce3f848de2cd4b6347606ce7e7f6141a24d17c7707d03bf919ac941a1bf9ed426ac053179f63ba0b2a4399c18a9fe3ec273af364167f2da83fdd2780dbcef05cd393b41ea49a9120f9007e77e3c6370afd4542e45cc04dbe92a84d2147ee9f077b9cfa8e5e8baf4e6ff722f6abc0051e4a18eeedb79dcd3e7d7714c5e414c6ac0a1b08c6b4507ddd8e7fa888963f8322c143d0441479107a9efb496efef88c8d336c1ea180d2d72b923fc6c334667394663c477735e5da197c6233e43af3557bb6ce6aa700ba6b0a981aa57c838295515e007d6b1f049cefaa63ac5e7a1c7947067de9da46ed05252e9b7880cc8de7c81fcfc1331a0e47aa169f6cab8b152daeacc36f9d78eb7d85b9dc4c3c4d798dfbcf0e6ec0ab568336e1ee19901a84f94fc62758d00902cff0253f3d187c841876d6e7ac1a2e67b277224f383168a13cfdd5fefeaab740aa104fbf4c7cfc9a552977ef346a4971f62ce43d58e7cb4bd25878240ce6bcade8c1ed9844bd49c7176e57cd1d1448ad3caffed3125f6e9f0c5e9aa6eb2d69c5a6410b8214e3b5a0901c3a7e6111e9ea93e35e81a4f582b03f5db85f35c83a6d2628e6941beb274a351fe8ef57ba5937dc264f0aa44cd6dcaa6ce23c740cea6f0346a5707b0ae9284d935bba28dd2b80e76619089ae78028b62517516d2cd2103d42da5868e0fa5c2984e60b00600194cff96d30d760a5debf9d98c099784f9bf6329b9ba956b84186bedc4c54699e51d4437ecfcc41734f718c7be43bc363b5354dc51c4f7dacb95dd5f7c11940828dcdf348b759329a124b3c209032ac95ead8cfc59d7e527660f6a98532695188249fa58599c4d51928dbb84f2cbcd48f279ff71d158c8989838e37c7645160c590882c6471d38529fa62a0e9a365a3c935bd6fcb25f4053a2a9473b24041a1a6d8a2e2dd6b99b1dee3d6021956531cbf29266956773d1e8772ec586fd4fb2834035448e1c362a6d1e40896250a03f13867bc8d7768100c4ec5858ab3ed18538867b18ab3141359711d80449d533e214b73eb6c8b5b1c034562b1fa451a02375a7a0e547be4248a85a7256e5125df93bd0e9804d5b311e596540e65442ba3507a7ebf6bf4ad8f5e2c64827e650fcddfd309cd54507c26828b0db6f9d2ce7f5e66079ecbf10b5db6ca90cb90fb890902c7dd7d4ccd73f819ad62b5df9e8092dfa1cc779ed4ffe84de686dbfa8765f373a1cf276f53d7458e387080fa27537f824be1248d85c16dbd132c060ce92d975ff2805af04032869690d15c374c3261beb088681061c49047078df32990845f82c610464e42d2c7faf525651f5195d2b9b69254ee8248e16840fb9acc9eaa2cfeed6da83acc8097456e9c253ae34aaa39ddc0e2f7c273fbc484b2b9f782ab56f6c69dd78574924785bdfd8d64e582ba177b693edf62ad8772ccd7a0f227ed93e17ea875419060e36bad590ed3dbc9c4605c48f6c99e76593abc891a7ea126dd39d9ba3578991f7da911e8edaf878d06e905904398bffb33db138b2487b78d334e54f43018ae664d17b767973a6fdfb32a5481780cfe9fbb37f7e4390cebe5591b5f68125a09b3fdb299644bbfceb79ea76148e63252fba069bf20c79e02fc8ae6e9ff3bfb9f6deb2742fec063040879270de31156d09446389aeab8bc8fb4ee87cf2ad15d3fd9ad309aa060ae54dc33f96fcb82f8cadf6b4032e009680660015fc7fce321e518790e5894711feb08d12d22400669ce7ec00ac8ba4749bf861d0fa9fe2bb3813b9f995ca22c5a669e07e85b8935082b5e7f6ffbea4c64dc508888efc096f0e62da819e04c806a89296000f54f93641c075c8d6067d2ba3832e9c47e930e701882b366391f75d0d0f1e2f168f9948b3ea260bbcdbf9f836fe22d19bc0e0c0f4e1e86bb311d570f306204a72dc3ceb1de73e450a531caea90a5071392b5a27aa511f4887b9e2f3ecf9d106fd4334abb7721bbeba26f07b8983b25d93c7d7d421330edb93e89e3f2aef45cf1ee26668751aa30ce372a94495b9dff7f566ffa159bd2105fb87a1056f29ff285c219f0e7ed6924160053c82ebae8daea69532ff3d8bdf564e16cdbfc5d29d09d70910c7d049a49048c03a2af2c6a4bed259205a262be1d21b5c3af9893f4e2def58e9bba868e9d271bcee9bb4b48d31753ab895de4b64c99eae057ba17bd77ccd15b867dc62aabf2fd234607a4be3a60a30eb0b94d42ab90a97c3fdd3a9b9981844af4d8fd3df73dc797c7b334ae60d4303fb840642777012ef9b349721f3da7e5d8d8152272675b9615091a16742c5675a470669261a03e1163882582f2adf5f4d02a866b3526c9a17a31a16a2b92971f7ad1daabdaecf9e7cc27a78365ce9c9cebf5eb72af3400b0b6226512aab42c632774973e6894705738ef88c0bd7e8669667a33481773913021ba3d6d77c17722e1cf86206974748f23534d7aa27f540d7a11c79d3ef7e949897c0374e64c20475b0ac8aab89f007f69c7c0b82ca5ffcc5aebde0884d555e88b9538baf225722bff94743e8773bdd7d6cfe03f8fcbedaa6d97784894cfa07b826ee026126c368c2b87a92eeec796cc54f3b7094fc78265d089b1cd27649dec28199c9d7ac8bed7dd0f720b168320af32c507bfcf938726939ab68d0c07b59419120e396881359acbb971b72387dd65c30cbd655df798f392fbf4d702b4996c81bec479085d0adb0addf07d4d6a0a543b337b12067eedd0a628b6b8de8498375e20e14f247ef3e590cbdc7ad9b9e9bc46f48a74e621db02ed7c32ee71230646f80d83a9f5c97b26572289ef441bdbf3c050f83983225805e59a2e1f1a016f65e0655b1247539697137d9d7b0ecdaf75ae0f5335ccf0c57adb1249862749b18ce8e100cb190d644d588647aab9f96f5f033dbfd0b7873aaa7c300950cba29526d9f6e7d509b6f8737e9fb5d6022a5ea902b4a7a39c6446f203efada1fdf78fb9dddf4e468242f064ea5e99a42f4cc4c87b2401195018e6363e441bd07ee5401b3fdfb18988d984fcd5fef4e69c267440e91d9e7c768e0e533462948fd9b5347602dcd50222e829fb23ddd5498913e56c73a246b14ed5a322c39458e885c5ff260dce1a48d48525728944efd9692c95387e2379ca9b98a9ac9c786704a67dcd0259efbcd2fe187ef9d5c92682064c7f03065d326df5bcba28e92d93e8f286458d55325e68c2987b4c063ad0befc57db5b684224f325cbaed82898afe517b931e9bab5069e47456c5d0dda0b60329d2555e1896335588453734352fca9bcaa6545d87cdfcf73614a3e29b6e67e4753d43ed7e4c2b0b3397de36814b32bf6690ca6ccfc01e79c6bbd5cda132ce80c51fc45b77228b274097b477c781aebe31526901c4ed02aa980b89023ab3e03554e45a1841ab3c8a23aff8f716dc63085245fc4f84dc4947fcdd10ccaeba1cbcd87231f5a4ff3ac0f54ef45ba2a3c0ad6feb14d29598134e9a00aa7649ffc57849c2341e96e327256524d8037201391940e8c1ed111acd8d914fc8d9cd97216ebde135538da4e837bb2a1bae7a4e029b0cb94e426aaefc7d676c4ce97ceaa98039764a7c9d140728d727e9862c8240b1a47440a74d645443f9decfd5d1d1126cf68ecb28ec66cb7506c6dcb83c5b57bb6e64290ad10d496a3f3b616060eac06c2e8f55d36201ab72f58402a9070539f5c374aec0ae4868c0c4e8534a398a5119a7c7af0a02f8037f2d5c9aa4cb90eab39da5f3ad5a0dad7f205d03ec0cfe4feaae3ce39da526580597397aaafe11d345406a85cf25cd66f511d004807e78bd06f8f747b8cd2c1ad089ac38816e482895d8273fe94dcf88b3441e96ca941a91687b5c8ae5a6eab12b4d376994ff75e3a0fa0849312bc24ff75a1d48468d0ee4479f06ccbc83ceb0632b9bccad73d768c90b96ed14d7af77dae08b2a0de5bb4af19368f5d5de693e951992e2c7c4ecc0d896761e70e392f6cbdab781bdb0c2b4948f1747938ae803856820523d0198962d1c722e9fbc075d1c967384d762210c5d0f03ae918c78cba872db4abf33a041105a09;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'he9ab14aa35dba047733deab68ac9d0debaa86ed7e29c139a763f290c5e6b72c1378b9a6492e7badcc42f730601af59c0b8566e845394a597622a63250b42c948e5ce23d809bffbf82a2ed8ab6a7f7ee869a858d471cc3860d8610d372722bb3e36a5ad99214f3cbc10f0e8386281a3678e842486989ff1b9fd3c516392d534362b2d45192623eec16a4393138b1797772b3d6a7c5a1a4eadd31e489c3a607c084ce0a6b18600c2374e778509938c584380a874e9faac5425a25c75844b1557dd542a10b7d05d811c308405d14a50e00fd710b94be7b1e94b95d2de72c7a8d41c8e4118fff894048d494fe51fe56f2b0edd5802d0b2b69d8afd437930a1bb6d2e8394ac5d29b3f660f7ba994868a4515e923bc0e067edc21e5294a28406986ae07337d5ddc1d87d56967ba85beed17aa6427148afb650577ce26787f02b62984fd2d32e1416e67e74c9179bac43245511dc961300c17c49feadf0d6da43cf7cc28c0a4a92288729cd5c38d8083d0f0ff9723087c74753ee09bfa1d24e50d3db2c9fe550bcf009ad44b727d4af9feb7e07614e3ce82d421639582d9afa023bba740613a9ddd7254e68f0e6f8ccbbbe2c1627417ec4dab5647475e39a3a617862f311623df99d3bbb92ffdc9ef167320aa2effa6fb8d938d51a2eda356c879a7a75de9c0002f3fb871a60fe02f552f6b40d323c516250b77820704e9911c5a162ddbd3c3f198262f1f7e52c4c241fb9e057f05ef380181e8d6a848f6f3bfdf8317c120149242183513d17b05a253b40f7ce84208c2c514adae5f5fd3134cb0d7efe875c1066e6601626a0bb6698ad798c68055dc306b22158a0df6166bb6566bc86ab30b6eb5e2bd52572022b6412c580841934217c5e8c083598995097b15b6824f2d762edec59383c66b0c1581a8cebf9cc1a76473b370f9b9abd9081066f51a0010451ef5dab64442f572fca9fe4bd536e9ec79150a411e65364ec5efb6908573d12c29b435bacb83ee73b3df78b5ededf444dafa6eb011ad67983bb7d868d3aad9e14e4c0565fbf3db95b499dfca8adcc380758efa3d7a91b5eaf58aa70c632c097f41cf2d1238426d64557ba6d1ce7aaf82e4692eb297851c47127b2bca8692ad8097c731c3dcf0c9c09889753e61cff33e878ad2024ad9d8f0bc8bab95b4023f524516b58f2673629ed323991aa21c119a14aba1cb395e7d05e8d440464960a5c36363a58b835b304f782e67962a8dd2c1ed464128db5729bec23d876a96382baad1335ba119ed842033fc13aec52e1c59a53a273421b0e6218fd68c7b141d73fac784c147ab62ea4672ad118e2d5e838402bce1bda40ce290f17704baa6aa29dc570a294c096afcd0e8a84f40d7846a93811822973f4594129e4c3e2c6f3e41c80aa5edf97a85f312f2ff643f3de133fbf56f608e6208cea404cefa3b7175fc239b9e580ddd23af6228da26dce1d415582a5400d3dfaee8f76c6396ca112d6ef8e8f5aaee34c5cc89304c18a203e09ed90e0deba8f0b7f6693925a0e623995190da370f29e13ddd44e92bbc17860216e1d8cc537a06a15942d9b517a47f7739043f1f6b28c5c0a34cca7f5f4eae983f6d2194346c0b47111061785443232d07f26e14e9f1062201989f8250128b3639d34adea46ba0e042c72543f46f7a14154f07dd24a6e6018e429d4086ea31b2cb4eac4e0827d6de4f74112a518310ffb4bc3531c7779b06785aab42df5e6a07113077bbe1df232a5805f98b7ace7b63305c2f4359ae9dedbfd33ecd160c6f57a8aab3d55016db1af0fd94b09de9b0514f5ce4937239812df1bc2298d1d1e442fa8d11c43ffeef4cf25eff20135780eceec41f46aa332ef1f78d288587c292c66751add5be9be1c20d00658c1331bbc964475921f061021d79e480b2c6eefb411d5b30dbe1e76e5c2f94b4557c7a4334a8d8b3fe0ec465f94ae33d0920215e5bc568ecbb45977debc6ae1030a2692a960cfbde16af776d87f602cd1b9b372bb6b86681212405929cb54dae76c0f9e8334904b690f8243d39df1bd24d3dd98b72b8b620699baa919087369cb28446122c3b78db8c9a37b85d808dcbf0bf8c7e17d564809755302ca98bcd8c14e4307b7e971143063ec7fb3dd7b76905c7cbe3b5905ab67a81926475f6459c6f827c4551cd62466ac60d039e1546960f952d0a60f82431b4c7b26ccd6eae427d12cbe435d9a21d09bce9459dcac6041fced874b6da3681aa1aa166917dce96a9cd661bfc53fa293a19a16f32a1285a2153adb33b5ca30a07305e932c1bc1f2f31af3ad17608ef2758a8e90de49c0da984d5d42ba4417917fe28b1b4300dad6a8438d61b6db87dfcf76ef6ebc74af5cd6e92ae14338a9957b077e26e38baf7ea1ac29b81c9c2983af6a9d8f4acba4d9613cc505d0a3fcfc8caa2b2488ed77ce87eabf8bfea50af79b33c11d69689200fde7493d97f9f6d693893955eb060af2b0530f92d3f0af4a20c5d14e30c09f4f525fbd5ce7f5e110df3c90f23211bdc73c61a7cc15b93a318f37ed9374e6e879052e4c0a9f1d6d21017c342ef82552ad5ffdb79f8525437ab85280ef80d1e8c71f34b7701d02269003f98ce5d8942142f37096694d158f565b9c5cadbb4df1e8cabb5ab41a33880fecef0a38e528a2579d613a45add925c697433bbfb7667acf095d094836e6ccf795383f377d2e4a6e455e006bbf5106da47a78b9a89c3510855407230046a910b9e12e2d7f94631dd8e8f4c667f1cfea389d17ee721b31ff2a57d2bf3388c35fb0955931c7f53ffc4cce47592be654d97819fa0c9df9cf9c8194587694273c851e5614a98433119df8e47c6244dc60e4b60aa3682df444571e2ff291662eb598b0bb53214e1bd1d6117100f9a28acd6b2b6d89a502097760b0b7df122d4c3a5b57f16a7412de1cd57dbe99faa27120a8bbf25e925a4fb2fe8abe2995509fca0baa0c563e2a9e334d19a68eaa563e707a1610ec31669ea23a5870e2bd7d198ab1180a05aad7d0209ad86e6ccf73aeadb7045b109cdcd07ada99dbe25b1721a767cde9a517c5d4c8fd6d581e1e63ee17c943631d14226fb1b604c4ae3bf7f8266f63726f08bedaaa03734df827064b1279c9756e9db850202ee9ca2dc22a0c1112221e85faf78ecdccc6d0ea3ee81366734e5fb4122fd734d366c4137b7d55b5097491786191c205681df50e0c44fe07706e9f9f3f8ff8c51bde9b56e8afd3c5cd175a8a9829dee6041a14ac23462198a79fc63ea17dfb2f1ff10a422d4e57b15eadd24b730ec8684fb76d5d77da090c3b92731b642cb76eb402581bfc9dc4c03792a340dd3c7d8ceede6d744073e69e89298a5c0c6925feb6d57f5bc39fc94dd833719b28880bd90136b0d731bc37be6ba18d2701f0cd67147f9b1ca03d4da81cc2d3e3c7414204c07f34a8f0a6515fb2ffdf59bc112cc7d6a087af18881d94093ef80fe71279df742713cecbb315f0750630f7008670b7c0be629d981415c4331076c79c8c7e2cc6a088b87c04c94ddc6673c7df8c4c5c2b1667d425fc1169ebcf634292312282c31084a63203da8bbe22b720524d927adcf2a774ce9d5dc68f3b5571aae562bba46c935ea30ba8c6c17a74114539d749a2476ed6204dde1cd5699daa029815b780c680e686c5ebb756013461a3c6c1b0d31d2903c5713449ad3d726793244c473a649e46462a7004ce73d15065b3fcd39d1b40e975ce574548efd7cafd1896676ad53a211422a0e6e2e062d996c74a3b98d9f3a0859b9103288535058b3939df6f9a264a06c8a9acd041fd423e6cc7fe072611c398bd6ee2d54e036504a7f114b3fdf7c19f06583ead05d5aad2b98309515c3e9c23ec442f0f38cbdbfbaf620f2b7e2dc19a67295fe8db5db7850ce56c618ae8b01891f0396187220b8224b1328e1a7382dc4172610c8b82485a91ece0f0c3e42ba06cd1ffd32c1e61441057fc947b00427478abc819975cdbc41cd928708bdaeaf1591fc7f858077d4af09716d5816659966df89de1c1208514cf3d23d9adb3f7f21d31a44cbabf9fe40c807226f282f2f6305a02316121df8c3f6c8bd2ae17ee448a6cdd84e9a86bd176dd19230da0620f5e564085d33cf844991e580fbc9a071c5a71acc35e032ee09c81bf8c7f4113a0d9f1bccb27bd52dc0e4c81b098b5f805655e062a11f3d5649a84d7b0f6d728f84aade3461fa5bbc8795d80e3b3f4fdef244588ba4e53c125bf9c593dfcaadab2b4bde5f0c0a75dc96803a7776dfe3038a279eec728fe90887372fe0d184f7e5304acfc71cc47fc691175bb71fcbdf85343537f7289bdea06b761c8b661ce23705547e961ac33cc86229a864d908b3bfc22a257bf8faf178f0195cf7cd03b6ee7ddbe03ba81033135951dfadab8bd581f9f18103e0fae40c322fe3fb512c365fb8d46c1a480db56ad8a238d517e72522894983ea94ecbf2bb757612c2261dad0ed7c0ab0b00a6e60581c1610c25106aea71d346e8e4685ce7a1345955400ba5e4be2ce8935158e00444cfc1b01b90827da856b0433439a09eed38367135f5ecd2527986483bd2ef1908d7185331fb741848a2e56e1f796983b6d48455c241e6fa6b873735c7862456394ef33c4df6a94738559cb1646970715f9b84fb0ee68b947996ed36a4edb3e47321cd20d83b804ea2bafd12af072490ad29d22973b4a8b7e95951992ae2560d90b32373376d09438bad0a95a6c8f6da273d5b6b969608073278b197dee30e18f449438fd7584407209619cd0f7442deca68579e6d12d7fdfcb48eba1a8e32f76db960b9f3b015ccdce165f1b987321be34b337bd27ee9db72af967912a8a62bcb7899377f4447a3e4bb660e33141b06e926182292f55d7d336c2d7b9f16c1a4267701dfef7f62ed01eb63da2dad77dadbe70cd50748313b2ada49857b2786a49b3bc825d407910bd12b635e5ce731f14c9ecfa2dca69651b4e540b0800b3713d6f7bca0701f28701f94b760494c902a12f887dbed144f36674cfe83e201a10226bfa556575b1224144937894fa396ee275ecbf3a35c7002d2eed6dcc8fe2035d6d90e7208449b672d9d72ab4e70b063dabb1eff8b390f8e5db715628d8d9f1086bb29b2bad0fa1832ac3c026778d7e5534048790e41646a116ce17713c40273fe33f7036e8380fb6f02e400e013f32dd8dc596c29a6f86edb6a2a5dde5a66e13d0f2b8561b448f1ab0ef142a0ec97b0d2d5bc079cc006498923deab4aae929e2336d1613c1c8ea81fa07eb0aaa3b252bea8d6b90017b198d981d04d5f49e91b96d672b278d4d335c29508e1be44dd04ed3ab4fd99614c509159e84c8837970471cf979bc32b9b5dfaafdd03fb096900f9e49f7d70412a9c851173f48d0a8a522395c6a4ee8d8bc1d4602c347b3f71d112c6c5700714172863100d09e2f4998d73a0d680c18bdab69a910d634a9f9990d32e8d8a78d3b079a12ce2e5ae86ee02c9f6dafa3af0d46340;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h759052c95c44a81259ba70da30c17d91bc1781ffbb894072cb33aeeaca934589a397522132a15c9f5ad85693cd4874ec04c54d0890d06f7f53729ccd833e34c99b0af98b57faac871619e04d1de3b867fda45000b8700c9c9d95e56f8df48a65248d5ef4edc69580fc068d3306a3123d743a37a0ade3c3e2c8d7506808b8d3b46fdfd14e958417c9d6c5fa6049a4e13194ac8d7b489eee127aeef2fa252030b0b809eff846a435110993ed8c43598835e51215b9e3f2208782efdfa9c2af63d3dac0cf4d1bc2040a868d640a95aa4c69f0b92471df5c6fb2ede2c184f72630a68d0827247c26e555d08c8d297dc3727bf0c0e7ed3bf6993d22e3cd223eaf718729c9dde113a1398f07d0cc0f6637ca5638d1aadfd8a92d92aefb5215a1fd3de7aa62d6bd0739608095047a9362eaa0af2dde00e9c4b9399da8e881ad0860f17d210a9574d6c8575d6df7587df17abfca01f88c310eca72bc2bda669ec94db21b6f39846d62fd6ada72a837e060c902064e042d26431ed33bd5bdf6038fc6a281584fdd9351e61e63cc3d59560e9da08d6a408f12554df9ca5a4bb77f0960127b08bd4c9067eaa3def15438f1c20902af66c8fddd0bfccc1c05c1d56db3f6e910cbf37719fa08463ddad2a27e8cad3b3df65824859755766c2c9d7e15d27f1f7693ef1f0935d25ec7ee6272b04e8b4bc89d0c9ba855f09ce4427d8f8411fe67010863f3f3c20b2fa6a15d07052239a7bc4037e9e85ceea2eee408c5160195ea5591c5ffa0d013590e9c67919051143332936d064ca64c9708fef947dcef2479263aa80a853a93ecadbe595543215964e05a89efc6a8d89da3bbd8fa7070b4c68a413ade80a7f0e6fbf0b132c720a080767f060fb439ecd89987d6d28b0343d519567217b690ce116e72fda7e6cd84d728f3a59f5d684402b620e18703bac5365cedb630e388680046fbed73c047394e55a8f7cc23233ef0d16fc4220daa608efab7a4e38e485c4c278f4ad34638b40f3285f4b96f0a0072e8bc9b8848f539997ad0952890c82140e0a1737a36db69ca51f8dc1ac08b8387b127f3de59e74a9bf228da7e8e13dee0a6c10b2f706e149e0ba3bef7c71dc5b2aa55f501380ee57dd3c83e9966e795dc245d9af786ef8e9e9e4ee4f55ce95c33da6eb06329f1444d0df68a393b5bf021ef7ed92810bee9ee2c00ec48fdd23f5d378f80cfcfb0f56f690dcf00c3fa96b997a425fb147dfe4cfb6236804c61adfb504eb6b89d4707f133de7c63fc562852e84b0b6f7618b2f0ecf4c0639d6929a0fa8ddc628e6ecc5ce052317deca843ec6b8525edb5f6a4ee4fc39c65330e89d8dae9bd9b9737ed3c6e93df6b366f8bce14eb81134efdfbb07bf03e961f4f2a963533c9cda54a7dc6d554eeee83a5eab6a8aeb55f50443d6e607e4f13d754305ab8116da8a9b48bbbace6426025414afea425d15d5347d8fe2281c3cf376c816055cb9aa4b4df1620ec665102598dd919788deb0581a9810d9f38b70a88a5dd1cd39404326a75a7a0afd1a50b072fd493881868faa04b655fd86d76aba93b00861b68e3210a50b619893af0a40ba0fd8535bb4b7a8257f81337643e5806803547957b5b8f5c4d0afd93dfbe518d28e7f6c646acdb7c782123626fabf5cca15f01d7013c97dbe59f21f40fe722ab5a23ff019ade90a30f13b8eb2d3cc5bb7b5512e326abdb84aa9ce55ebf301028b6abaef747f3ac1daa2e1efc5ee72bac316189f15e147725b13528a00c31c3fc8ba9fd252d8c5b4018b81edbfc32728a59563cd077df101576300c8832d52db1e6ed50548d7c1cf95b55f4e6052cf7a8a5b7e7e42e55b65375f131018bb91689f89eed2c4cc139a563de0e968216b40af666cb6a9d5b342f103e508b293630b2a93a05dd8c3b8c5762167ff2546d26a40569e1a1cc69448a2181659790b1c415b4ccf40656a73f8c93b0ecc743f83a1d226fd2bcda2ad3fbd8b04265c07194382efe4dd41109d060ba7020092abdec1eade39c257f6f421d304142e26da20c0a843a836fe831c55ad95e3056ff920a2a519bfe531b5e3fcd209b4d3393bfa3f45df5eede5b13dacad0884b9ae470de6d445c607e6bf755911346183296ceb734c64dd5dba24d1851fd037e0c4bcbe6b25e23fcbf32cd98bdf0cf619fa63e103509255569430118265d1bdd81d11940b0f7186facccf37f21bb7f7c4058bf9df74911bda0600c34a54a76554bbadf9a992141c2e4ce4485ee0f51295db57e63ccaea5010f87c3887c31052f78be8dcfb41c87145af8cc983c6edf906fbe6aea800c0ba9f7e36bcff2a0839a792e5b098b6d9029424e6afb9b217a86b953d0092568639d4ce3e0f0dfdd454eeb1e2f0112a19a744de25a7b9728a9992d8b72363186f9b81dba731310e78adde94c762c159532653e5de2e37c7d96f04b3dee004026f9f2b1dbdfb12a1cca1671284adc730f8b9f721ec85d9e5c182be1bca5869e3779dce887737d52901985aef5576c154b88b44c94599cf08e185dc7d5811af497bd4e5e557bdcff668ccbf5a1919a25dbb64861bc4ff8bd7f2ae96e58c0dc43e408c88c777d6a9da6f8d2561a4e501c92149b3a3ea60045085e9b6829c41f5e11fd53beafb335dbc09238cb2e74b9684679aff556228c50eee469602fa82fbc5f5c6a7d488b2f212d68870933747d3fe443b764f88018d33002cdc0f4f2047a769ddf01b22b6aea11ba15ed78910811fa0008b08bb169efe9d1944829714779c46e75a0ba7acee115b6db5684aaa6cd9fb496322ea25bafdfa62674b9d71293da910608b98ac8feefa38e2903d61d2d09a1c6bd5b528b42546db69582bfe3a97ea6672e09bfffbe0703e841087dda1489a4e200d292cb63f3eba1033093ebd201a0b82bc2988de06c68deb917cba9caa97261b161f4674f9e24b0f4f750aac4069bd7352fa9d0206dd9a4d589bffa7077f48d15c7405947967676b2333538137a720b9a5aa06a17ae61e5bbfd32efa3a0a737ffe7e3178d7b352568aa14fb97d9f8a91c37dd4e1ff2e7ca27cc64e6c9c5806ca51f0aa7c820debd432944d99a1bb1faad70327db7652499378eb6134725d83e7cb52cd48dc899e0d5cc2cfcb1ed62470982d9b1bc3b1438c3e0638c6a35734ee4f61602923b648df25d0a8f95a3fc82dc1be05cb5849fa0637584310b9ebc55e371769b690634d073585eb5d1842b3620e8333f38620e5ba7ce188d38c015a0a8000e00c034fd13c914bada04699dd116fa8c44eaf8818707ffc88297d5292d3ee0061fbee1c3ef3e330c6789b4b9f6232c90bea0d6199555275a832c6a71cf2a3b550cea4f0514d59e7eb7b413e1c96b190cdc39a41ab9af1a52a96436e16a68e0764bca447c63654fa1e7c6b361db476f5c55214622020d01957b7a1098d14ee589acabb0bce62fd509bffa3be8ee437f3aa6ffc480fc61ffa5a4ef41b00db506102e1bb4850edb1041666c1a27af4f1d0ef50c2f34ec0af396f2b646f93f2c69d74269841ed94fbe6746445ec4ccaa65a1424a28fc937eb983b212128b0a0ba77a6ceea6a23a7e640b12d7759891cfcd2ade5438285dd3eaa3da2e4f34cb822a06d9d17ebef7b619a3aaa91306f4a9c27c840fb301f9076b6190a8abe649c8d3a08d312d5ce2a6061416fc0bec18e45e3b8a409c577f556f5ab11a910675047bbc4f07b751ed9cbae29df422edc1f32b06cad5436af43b104050f332e56ba62740b4d6c3521e4c3f7db5f64881eeb8c7a3a679f5f5a48a215ad77cbacc0becd7a9a86e74738ce4f247528d71aa979da3123da6fc730cf9bcdc7b01649f2759625411eb9cc96a7fcec1949bd5751a7911d5fc77c3bc52f7b3040e966c5feb4feaed284d2f2da7b80ac56533814270b5aedc6829a2524b7755a28abc7a147fd295cc89f942b894ba1421e0fd2fe24c30e47c56e86f13708b8da49ec7d2b8af3a58c568abd6e9a638c24477e41fb5a33ef00aa979818993a7d72ecfa55ab23170b11d6710c5056d6c2f381789d8851dacf33ac1627b69018f28ab375bcb1364c252b4d893219668039dcac412393197ec97d8f0af032a6b27eeb7705193c8233efd30f8208a98491ac0b525e977d72adabc735ea758a47fec55bde5d6877e3fd01cba6246bfa8f8ce573de0dcecc26252e2ee65367c96166c7bb9f9eefcf28721c3acfb73bda4f2c8f8d3ff87e6d594abdda9d65c688c4af5643afaf7c647f3f0b4c71b0852faf3d0eb3abbf740f3aba36edd0e5f97ecbb474f8c069e16172b7c4eb93871663372ad22e51a2263177a2f4aeba4f2a8da67329621b59b6ac958306bbb662ce105bf7c3c691e781f56a8adda32abb91f69cfd459fd2dc90fb3cb63ca5307dfbed2d1228673f7019ffa57553f29047998ed871b99dda046b5cd3f4edd1f261933a897a22fc7c0b4c98e30972bcf0adae0fc12fb9129f935780e04bd4568b24d4bd8d2c7f98e03949034438179db2d3fc6cbbb1d948e222a1a9c7a13b74cdc0f01cee3dcb355f39b0382cf2d80c57e1126af87add3b32c086e0d78a61e4fdab80ae2d4f2d6f3c64518aa8e33d00c9796392d4aea6d2089da0547b221ce110718616800df7038728d88ee3d883d1789da54134549a90d5aae67a883350c7e66d37e3ee3cae2bca7af7a94ae9232a33449e12a60dce86285f5f8cdb327c464be08876db3fd6457a9f14f9777899eeac95c6d4c521194eb2ea50c0ae030bee1a99e1dd15bc50d32bebbe94b83a653dac12114ce2b20e3938aba198786e2ed5abaf0b9d2f08cbd72050986d17cd7e5337283f3de86777b70bc5a2c4b987dca92c3869278ea9d39fcbc05dc777109a71f9b52baa8ff6eac0d642c0039557c797d8008889086f9c5587c5049257cc3eecd2c1a89aef9eae15e319742c3104a65a661e84e51f4d02dfe840caf41d74388d16a1f5fdf0c7e101578734323fff254b83de1ea15fbfa4ff2c2e8dfb703d0b0925599391d142333943045ab25e69a5708cafcab99530aa7e858bab1fb22b7f7c94990558d64009df114eb992b4956aab3a58af7646015d8d11cffd79bcd2b3e1adebb40284c7f5ab2d89709add79363446a28f903e93fab43224032079df3bfebd7675c183d746ea41266d21a2e142411deb8e95d3cd5c1dad2f85a544d733411b2a731b0255bf5ccb3406b8c1b6cd01608a4deb97b4cfaadac1518dbd0ddc3fb2f0fcbe8315fc4aca87a10bba2ffddfc706192f6e7a145876716090bf5ad092f575c2357d4a6a097d9407c0841956df37765e0d63ee96554966b130efd0f383c67e2425c70e1551baddae5889a3715eadf04879d1913078151f91b44bf08cb6274b39cf91c0d3313de30080af13fbb00c4bc0e7d854e5c422063b57f351626454a6e2857e6cf74ece1f2cf211b7cb7d31a75cfed7f8d3d1712a4f66c7523cdd453616d431ed25555493c714d04b59e71d6098a749e35f2a59b2d51ee8af96f9601263b4994eb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h5338e6a10fb177af1aa479d930a342c96e10739e9e8c5d2eba0d21df1b033c6ddbceaad9c58006bdac4f74094e70a01bf8eccb2de48efc38b25e049cae3cc99e530eb00ce5b61d19cad02403d8e08488ada69d36a2ba2a5f524cc18c703c21c3834b3a778e763c93ae7fbd28d6573c8c654f9f3b9c79bdced0501458861e4b0e206a0d4535d53c4bbd5d936457aea38e093ace59d8c0a30b68b90a04ed1cfbcfe57f74e19f0a223ba0e28b6df923bfc6e803e1fcf0efdf3932c16889a3cdf383853eb057978a781abbd467649eb8d5bae4033f3daeed6836fd0eb0cd295c120acdca2150fd0b746239bbb239506ff76aece2788bf64e198a1fa51f403eb513d1a9c44a8ebd7ccaf46d1527584c28ad67b0c1dfe024a73778a2a398ac3fe858280a03b80b5e9104534d7cd875e425243ccee7b46698114d9cdfbeb87f48c0100b63416753ace0a443834e6c403460acd30d6383b82ea3c05dc3d9785fe190fe3c1dc5cf7d4bdfe375680265d47c4c193163a0fc07152ceaf1ec66b0381521d22d005cd0f4253b96342e8bc46451c3f4a1a9da45389a7ff2cf35f9025f6771b0f82f3e7be53b89af1192b4dc142a39f686683d3d187e9299301cdc690f52ab1dbba0ad3b97917c7d6b89f07e6ae0e040b057727a059c1e0f450357a09a23e4e6d363789012a27ba0c997df01c27346da0380d1867b561ec8449d05def8cc239b5e689a92ae9d55b43bd25251981a05853ef6099dd6ab7921341cb0a593c9b41c358941faef30a10562f1ea72c4756b4a4894317db4d6b0d32b252e34161bf0acdbc6ae58ca1b305d661196094dfafe36f7e4627e2d3f1c81d8ff3dc7a70461e2783cd215e6a17c1a93a50f3862e7b9ce84319b0d7a4261c6f230d41ed2830a978f83f88ebb866041d65aa3cf1944c59c65f086bcb334fd5b171fd27cb33098664f66db69ab142319abd62bd9d700fd72ed489ac779d508151eb06e51d2ffc4323a9c5459826829222ed5b7c85225a6c3b9cfad326f8f681795d428d013b573de3dc491a9a3473694a86e38a13e0f7f71bc95895607d519a5578bb895ae5f52594841727a677880026436e13054114b4fecff8b3ea306deac193871dd2f27df36d57be4d964b89b2a874976b85c102e237bf9efc2004f9fdc718ef46d9a0c9777d48c27dc5504f534455cfe0e05397dbd35da7c8015349acb85ca3488cf9c471accdb0168b07f14b2bfc23e267057baea66b162dd59e9c1ddd01f61e63f9a05b610c1249e763a1a63130fbd537dadb4c79da001c8c73e0e6da4fda8934a229035336c918378659c28e5f9f2f74e35f8382b11a7e405f999b193f3d73c68d834ca49fbe10064119cccb06354900d8305642f285a72d10742f28106430faa7c984268f4cd40c20a12c08d9829088168d2f425e553a5da41cf274a67032f9636a4bbad0342eacd0302f757479c718a4c8123df7908a69d96be441814711eee33ff4dc0ea10c46f9d4902286abfa1a694881808599b01a2ddfb1eb3a52f95c697ae6b5b9002ff242de8aec610564a4c10059a326d715685552307b104cce98cc8dc59f8d28c169afa2ead0e8a8f1a069c812669a5a08384c57f39f0bee18b446abd7e4f271a8ab70b80738659eb281acca121075de5c3996f7dd5af5debafe3eb6cf68f6791105d1fa4d6e7367be1fe125922c831dbd33bbe6d0ac1b9f7968f7f0350f53362561071e415f3a71ebc2bb4bfa1d872e3ac0f925452f99b9679594386e5321c15106e78ce08d5a5bacca327dd0be8e2f45f0b4ef9783533bfe991abd434090dc14bac3ffb8c0f9211c95c849bd161fac0b079e90fb063576db13b410ab44fcffc41988ee048938ca5884e703c8071d00392d00d957c8eab21095252c4aa4f0d83176ca4923828cc23a5e4fdfaa8f72f57417318c26c3ecaa9436a4fb634f56bdeda130c97058f7378f36364bb995e5c9a6960df8bc6ff2a40143bf6d41bbb5e347aab06a6d64b976d62bd1539016e0da0e612b2b10a7c58dcec622486e4fd30e2a6237a641c22494a9ef44c20b9e225cd9316830585e7407d1b4e98c107b48e4b92bd57fa643cbb7e1b11445bb00610ded6d5d5fd3a18e9bd4e8ae8a5a00ef292e28b49d18ddab9b2fa6dc3469c8680e0d7549ed7181f8e37f339bbf659e0571b42a8328d468ece0e9eec731051953d3ed152b55110691b403708dbe8b85913539fca2d80f16ba5257ab7ae8f47ea07bcffcb5a0129a6e3e5f068375dd73a8a41098c3a63ade9f1f441bce877069945c54e2a6783f874fe518deaf6ed9ffb5b599f3e64368d1c4fde3260a6e8ed5a23b58cf1701df5bf0a2451846d016c341723785606b22113c2ea70f81e9a03758dc08e8c2b76000290f50ca8a1977c5d38465da079707957f4f07c0d8a56e91f13c1df3a5edd0694a136c517e3cb8da31bc0637a37474da8bf9cb7e96a3a23d163f14761b6ffb5a86b91a69fd7894c96cf6da2bd3ac3dc6772da3e75212a422e78e470caa04103b08e90ad7c7643024b6090b02d5084fedd4e4de9d71b2a4d368e33b2a5827c68c536e0800c99d2f4fd519ba29278e43ee518a1d5c037642ed17a8087dc2c794c77d7ea16db27d973dbaecfaedfa075901c069574b18214d5b5e33ba6fc1102ea8018899ef26636c2c13b241989e2c66b6c764bfb4912fdee0695b5ae929b6c4ba7fcfc443c18b5790bab3bd39258da7bdb30fb0b5b717ef30420a0c25ecd380377833709c8b670f3fa373f6425a64add7f5e89f45280b437da3498485e70cf3463443be5ce5f1149b8bc78d2b25c1ac5e91c4fd66e903b4bd91923a6307e4c030f1c5b0d555dd48ac9b2255fb4b978749ba27106c7c6c047a844ea5926a6aaf363be7a87f3c5db679a859f8dc18e71a4ee65ca3fb9904452bf3453da78be81a4a76389fe74e32fa0dfc75b8cd257982be99b5ae1b5c6a1101d1cea61ce67197a97c1233103ff1b6698b581002978579cf17bb2757e9083bb698469fd15475920006cae615bc6151ebfce85feb7b1ffb63801013b1ea4806f40518c02db8003f6c96f66a18977758b6e501daa73d26f316750e3887ad68482143c3ed8e603eaef9d9baf5d0960bc2fb2171b96ee67ff82d278ffb942d49766e74be24f88e73b2e8f3d7c48cab728c00907ea3d596bdd5442e02bb2b9bf2997b9bf0f183d24d28d4bec77e8202dc3d07d2168bc39da334bdd52aafba0116ba6db3149b437ee1d745bbf6b4cef762b5ef4527c235f882c877f9813ea0246dbb7839861d423dcb89bb505db961ed34dc37310ee25748bbc54d8d10c890d1d87a4282fad470f74b1ce9f929d0e61e1551731835b8e73f55a29e33d1ddb76a61f3a8d1f63191c36ae7791505b84464e6420feac2134e39486afef9ec0f6af47759a6bfe2d6caf9b5cce01b5e684aae20e4b814758f778aa461339139b97e60267e45f626b7f1b3ee937b48ff83df53c74422995f778bc96975d491a116332711008aec36e1e61b99ca3ee7b3f9732ec357e2007c2cb6abc92c60b3340ebc0a93febc7cb7cc5ef43ffd4d1774de16c9f24eda537cb9311b49484e867d606d2e4e2799c8c8ab43f8fa93ad3148bfa22c10032118a4ea87452033dcdc18aa065689d5d841d7d9acda75d766906f8e4b1a44770f899bcc27c36f8a7309152914b9eaa2f722d2dc0433d7ffb6845f38726aaf2e17dbacc3f62aac311b82749417d76344cce2b676e6a5b842c413a119b95b68e5c0a76ee80c195d8cb55e1fec179eae43bb3dba864273724ecd014bf86fcee0bedc72491eb75eea2e5f98d763d0b13882d87bba25d01593dc64aac9a92d6f808f3d4d29c5c2c8f56d1b771849afa6a088724ac666edaaaa4b2b66ac046093d4d5961b18c85f5763d1055e835a4f64c7eec96daf3d27f7470d508c515f4a00c216b23199f2513cb179e2530b467312a87717565c62b5055186061e08c271f396afba14bd9c6fcb78a239da4ac45d64bdb28839c3704b08ee454270213353cb30448f46b5306bcb7cbbd5f1c3cfa25c91b55e1150a4a9de4cd9b0198dc6a4dccbed2e60d2413ae62a912f4e16f622ab463789ee946a62cfcaf9ead10cda0279086cf9a3cd2a272b605712555d05bc2ea8803639dd8f955e8f8f456017e25b65f6baeb0a6049ca5381c7ab67b2927c8b148fc51820430de9f9268bc240d7a3e6acab3caaec0358124a18bf9c8817b53237caacfa8e52a72fb4bda77b65ea0e4b6a8ffe99ededb1e009a5f9e5b2b6c8c6ca16b2b3cc73dd3692e39504493ae597bc548c977e0f334ac54073619ba7d69ad7b82b4c01954c4c495d089f9620b99cc7b527d15915ff462afb4a7bb3efe14abc982d6afabd81808196c9982b5cc7c49dd7efc05ca49a05a0a4094366698a443c91ee38812439e720b0484031a1682c916877e851b8ee0979d647ee684ab2b96ffeb4f44ecdac5c4a97b33b9984ec922ac6082292aafd6492c2caeb164f84d1dc8aa16916511cac7a4578aa54ec3c6802354bc36c55bdddf154601656721161a56e28f3c623445f640d7802b595dbb1a245d47829adb542146a6c08a880aff1b73fced2338bbc3a1781fb35c6ad0a6d3f801afbafdf5cf65c8c41444c27c66c8e061ca828b479c333b5cbefe4f33a62ee28017a17f7d8939355a88cdd8ee313d46b78481d36ccdff6c79e6484ad37e8a5a4e02ee5feccf3578c517effbd74e51f17101c23ade85480ed229c72015f4cd420b780f6d8d4896f3e711a2d3f9076a791dabb73a9b1dd5e3dbdc0cc7e4099babae6c359c2f8dcc39a98d1a7fe785692f574543bdea49426692f3906e607704cb271bdd179cb9677abdfa743041651e6df2192ed7641559de9cddb0436e3190f71b65522dbbd3ea84ee1006a4e0471bd029f134ce3702513baf9328176c2fd469530bfdeb3d048858d6791f5b3ff235e162289d8a39bbc9cbdd17734f9f90e98911fdf9b024aeab58da7ee68593c73cbf984e049ec89daa3a0c227713135a75d2b4de5937b7dbce9aaf86e59e23a0c9ff7a9dba3404dd7a0ca0c68aec37b3b222557d2a35a216ce43b488ac0e1071b6cb6cf90a6c01134cb06ecbba5e35bff44c34d0cd459d63d580fa2aca3023567fd3e7756129d958224ec58f7870314a5b57a6eadd8d71779723ac87eea9ebd893272eb3cc6ca5f3d4f1aa91a309eebf46eb2ab1fb50c8b26ef6d74d4cf7af85fc57a03354adf51e942243a503c46abf44e0f8a854dfbf3d64020867a2d5c6bbd12502d22d9d0712feeeac5eac97bfbe25f420eaf13d056158027089cf3eebc3d0a3572288f491d0aa9369a0ba71916167630e0aba929e158b681ca49e1e725f8ec9019be6c36032777b4857f44d2861b7264f0279eea94c64fc20e10f0fdf15a8842f86b11581474a12635b3876af87aa48ea7fd9abea9d6b974f51eee9614098f72eeaa7dd7cacad5740e5119ce5d1986d6043ea470c0ff5ccffa27d5118dec2bd114d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h23434841ecea36282b76747a8b451184bd8f9a622938335195df8e3d1d4e22a494530a9d2c221b317ca3d5635b0591f16f7f6c35771bab24efc025005520c9cb7b1951b35b3d10067790222fd5743459dc4d5caaaac91e51ead5ec5bc5d84548252557df06090ec1fa90eaa9cad6b07c25eddd1106fc2186505148a530ae511380510bd5d606e29143ef49fa0e9c36b19d4f23d502cc45e5e53c84cc41f774f7b7a418e8b19687f2c4c66c704558d4b9ab5e6f7d27ee17c1a329a158db61bdb57f6cda8e309b506daa7e0cfbb37b9cd68a869ab077e6ada79fb5e85d43a583b5e1fb1b397866bcb6fae8bf6a9c8526994806ab3e9f5356397da5051187e231f6c3d35ca9f18a90aec8d340c6556119dec6c199aae0e22b4765d5025799154bb366e2adcb9b169916124d01a6180b6147fc45293cc8f0496b13aa6d6fa5752cc6e7d57a0593b6129ff0f0dc44cf2736ff3fea2dd1998b55768333158336048d9996437fb4961c3630220c2be168c8ba5218d1aa6e128a7bce516e0370f55bdd7f9e02184a4d6ef1a0e056d5a7e9dffff9f155ba2c26020816700c9d66864ef58d94d92f3e3ce828b35071f003be3acad65c2063af3cf0951cbb08d751a5d8b034a839f17f7fe30c8dbc8ed5ecd234651b9598be0b6d9b8e561444b56dec9cd7d4c8cb34db3a9367ac23a124c4ffc44271bb3bead57590d03133aeeac8b6b1a31df1dec0c8c721921d6b4586f897be620c3cacd26f5268f7a96053bc8c577a3488fdd24a7c1d4f4ce65f0be7d1444e3ccb948554d8bcee22ee8c954769550041ee2c403af1a8aa3dfaad35903380c0a28d8e9d4bc7f30af28e4a2258997ee69381da0fb3bb90c86c826a317015346afd96e538b6f4c8555e4271df632e88f497b8400c7f78c0482ba2ae44dd21907734d52ee323bd124cbd6fb56fedaa0a89db1c48ecc8aaab3198578e6e778f604fba40688dc9fa9c697299ee9a2bf26823311b42636ce7d7474c65b1fc092259a518309213df4b10cf324b43fb7dc33d5e54eaade0bfe607c06d0be73e78e430b984852d7fa25b5679084f950ae4fa85fe646a47ff11433b3c04fda4dcc96d3b501b058e5efb271e3ac85677f7b84b3448cc1d783b1f68ecdf2c621773acada41f6ccc551f2eb786fbd358481fcdd20965f5a3824ec28fedf60cdb21094fcbf6a63eb4847d93a0f6bc33d642f95ca90fd554f116ea2709631729b84fdf40399db1bee64178abb71fe80c24130f20c985b7598f2522e5628d7c7ec99dad5f986fb488cd7361100b9cea7db5fa910fbb7c0c29936dae456ba236c3e6f917d50535ef160d729dfc32aa3bce159017c3adbdb67d18ecf9ad97c7437acfcd570f796447e2961492f127594a46f1cdc9c7bf5935c0d155a118a3d9e6ad0fc0103409adfdc7040fe97a68b092a930ddb134d082685be06e4f40f408b421a125672c77970aa125e30ea1a233c9e8eadbb3e6fbe17aa791c2e12be02b3e372419baed04d64df9547c38773aab7eb193ecb1f5c6ad41f73972af5469fbb8c9ab3cea295d9b320f4c2394dfb886ddbc826cca377ab03465ea2a2da5203d3988ec3fe5c9a9df76084dbb47e10923937a57c207179d0e376b5f7d11aaf5172eb416c95e4298a8eefe4b0180655fc6bd8c11f7c1cc58d675504a01c771de672e73a9a710387a2673e0213a431fddb9c3534fa952a17e944eb5f767a69cc0e33567e1f9cfb00f3bb69c46574374aea6ecd575b58aa780e84430cdd6a8a9b0168092809e5cbf2bc15e67f8e3aac8b45c53559d02ed0d60496af72fe9e6ba0b024d5fc1621522d51cbf3c6160206eb1b72ce850c11820422735ffb85e6fbd0a5e3ce2ba831d422ae4199ea633079495f7a9f1b5cc76b2f2b6f757cbd9527e2744b0a3b29ca567e9605b02846555941854c2a5cec342c46d1179e6c836b3edea0682ceb0225632d2947765b1020a2c21dd0f8be1d838c02eba21d2a75c3947d7965d939e4f3e181521afcb61203eca190c05e40bd32b1badcfd495c529a2c06f8973cba122d0f8bf173afe8a2f733c44b3fbb0a3faf74e4ed0eeceb1cda697cad5f73bdb48a8b336d288bc416c92ee883f22b2be9cf97769eb1ec72093e7573db8ba65862fb6a6a5c7beb66d9328db421e5490e597740cacd6f6919f55941444875ddebbe50b383a5ae87a096c110e6b9e1cbc9302eb2eea68da31cd86d521de9bad3caa437d04bcef6f39ce99978758a845abeac9e29494cf117009971bf707bfbbca3e507ee5b15f547536578f2e862e34e8d0352606b358adcd7677f7bd8200eff3a41b751077a60d7ee1d7466e03e6a19df8f36360b48121506fbbe7245ac820a19be1377367329658fe0a0baa42b6e83ab9f21263fc72a9b01e3d8d93a38f01b6f8702ace6053dffa6feaf86874c66d6640734d40d73bbb99f268982dab1f9da7d23367c527f353962ac8e6064c203b92fd308ee19ad5238afff42973d378394efd808a8982cf9086a618e8a8e15a62ed4107b374702b6a5f5794c615aac89b9b05c45168598a65f5297978959a85befa9be893af336e8ecb9a2a444c6f030f1d867f9b5b83bd61f6f519e8eb6004074cb8f4754e292c6ef9977e0eb09323cb2f9d60d8807a5394eb5da098258a56bd23ac9b0e93208d59cbbc683f952dd6121ca6b3967ee2b88bc592f5639d561745e314b2525f374392e1a86b41ed9d5497fd67b426abf74c221362f15553aa5768ad65946f87647ce36634de910e2ed08e5a8a0fea9d60bb5825c02113fd6307f5e3e72e6f9f201ac88a17af258899853d0e37b57ecc58d81c620ebf534548a7233d228f2264f1e8becb4c46192d68ad888fa2f7e16fe35ca72aa6341edd6baacb2c06f8e962625cfda790ffca90fb853dc52901a89b61079519e8816aa0dabc54097d832617a2f728b3af01897fa007fd3f104b15a9ade5720eb3ffd1be5b62154280d771a6e502eceb57913c31822ee5396550b3a972de9ef47d1b8cbb5a7acc162aeb2649e632665f5a66184fd0d2346d7b0addfee023c016474ecf64ab983f97c8e04d532d2a3b7addf0be87d279dcfb5538edac42e1c66ae4f97ab20b8514058ee27512435c7a4da53e4dd39ab1bff122ddef33299935ef3eae04b325de508e85752f55ec84a42801f8ee751b4d947b0fe25b2d42ef81cbcc957a24dd85133c5acc1ecc37c6edcd5f9508e82b77d4a7f087541281392d92841ee226fa18bbbd332ab17c42cf59330e89317b52071a72c4755cf37a13be7059626b7ee5505b123e90438bcc8736da4b7e9ca0ff0f50ae29c0b5bb10fa2fc506d893c73fc3e7c99c83ceff5acd2afc35f3096b07302a9601deeec403b84ba393e4189762cb109be5bee505048a49ba406123e94aa423d44b4884db7a30e0e39ba92d09179baad5392fa3707e56468c8a07679fa806a2dbd6f2124f28ede34261edb61019707062b457024405e4177b36c3002e4e1f130fef7e2c72b290c362d9c5549a122e14ef2161a4fe238488d4531cd645b7cb005290ceb67db88a2057b9e6210fa506122047e66597f776656cf5e2e412f2c904bfe176ff271d058f324ef68dd5a7cb7b91929c41cdcf419b8b82e13117d87bcca8a22664c81876e2a5606afc40ef8b89424078852e5481ba4f260324bcea4c7f4bbfc35fc33d666f573acd189f7b60953ccdb707ac7f88663dc78e944ec69002a4216dfb507c09b7fd7e1a10b098360965d3718fe3a33f565dcb9c8f8365b70e4b4b9ea5d3b036fd7d39597d20bc8523ecf5612d485f6aaef112acba4c118c40e7a1289011b7845730780ca52e51eebdda19483fd3854f9c79c8e0a411c742f276e87fd791aeb7bfe7b4467aa2b4f0a74a6391c8a4f0a77093146fc7fb96be729a17722bccd6895693dcaf6a3efb9ed68535c7c5e2f37f686e4682368423c6c5a8b6ac5918c8f1781bdf6560fc36569651f7be4038cce8ae208e16a2a3b05dc9ff0d9cb88b148efe01d0388ab92d6389b7bdaea0ba61a6a039beef36f68dd2109c525e1614614ff82aa0c5b3d550eb3d302e54115877c0d9daace59b5363c848cbc1079520f19efccf26109eb23a4414a924981138632da9f8bb24c04c1843c00070e9c9a30f7e2a53a998c7511611ec1b6182a9112fbb47ce170735053c98080360c517d0139d3caf38a526b1241743f09a45d10c9df7ac7061530fd707a2f4e03387b996ae3cb32c5706acd1a051f89eabb5c5cc26b75663bf68dc9a303b225b8e6a0a4b8a78d098dc5113153f9e233f51b12e34e2d96e0151bc271dc1d6daa72a81a831bdecf2bdc96de33b94d71d6900e8c00047ca04219608badd4423260cd9e02d77df53c13c7f3a149e86ef4b6232a06779eaf1dbe09097b9731f7bc4ef3056a1df522f57a7f615b4ad818f22f130665709eedb339ace76785b200c731bc6fd00daf1648b874c9d362470838525813171cee698b0743732a9eaf5fe7a9c5375902f9bd38e67d81f14285273d014ef49d0fd1d6191de4f8950f6779d72c84fdbd01e337a1ecda39f40eb4cf76fa29f2a6760a4d0974bdd7d13bb84c77263399e33cd02032f118de43a656b436d7c9eadbfef8352a3bdf42c5dbcf3526640b9b45891444cdafbbfd0628aa906758913f2f39865b6446bff8223d3a5d1176311932a5cd51dd6d5be94ea277efb8742b342d70f2f0a78715a6bf24e5a357fcdabc8c22c6ba8a43839c29d72f42933b097e7cb643ba02176ea2d4ef58dc33e90f2b3d485caf2b6e3764c5bc78fd7b1863f84d52a788657afb2f51fc3e37895dbaacac88d5deb720a9a1f88ce817af17f1bb869d9622eb04ee5b928d3a8786e49fa26f1f8aaeccde593a253d7106accbbaf58513b663d8d2fd3ed70853af0ede0f7fb21a1130c4e53c1f1d8e1e6237dd8807d2a6eeeb1ef1b0c40261e78eb8737f0cc57d4a5f61e95a96ebd458f7184528e9ce95cb3b5e171713db30799f7db1755e1158e6650373dd78ff70a58e401fe7c97e0f6d3eb9b336957174c5d1fde6517ceaf98c1ed55e3f6bf7d2475348c3f140ae371f6494b0356964f47a00ed90c3eae2fac6b9d89328c8e8058846e7ee19c5cb6d8d57fb278b74ce31536e65d58de80022f11b03542f0eca93a5eaf9cb481a8939496bd96af8fd2348f3753c29abe3e7f5228682f963ea035d474a90814dfad1bad38e69996b4baa4d3a122d4a4c31c83113b4808a55333dc2f9255eaf785e180d91459018b345a93c28eaf8347ab4b1151cc5df64b07e1d5f5c4d32d82e3df3eb24bc84d1e49bfe3d788c23899f9f765366970ef9521405cf1ec738fb490c4a1d4a223c3ce3e8aad07245a883094878492405d752ecb4427d33ea2c77ba20417464bc5d614b1c6639828c9877d18e16c0646fcbc06c458e280542725dbc362d906e11baece46f9cea25ae0c13a1e34ed64feffccf5201672edb2a1936e0770597d130594f1f63f00e2f6f322076fe81d77117c4cbc64;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hef35792f266fd6d0f0ce22affb68b81bd4be73dc0db7fc3ea0686bb8c67574666e8dff1298f3a971ed44a824ff80d32f653eee499535fc053dd88daaa8881707bce8f5a545b553f34fcc450c1c182524e9966132ee5570168f1d9882cb55e8e0d2f4459ee4d9c53d05f1cfca6da49d370ed18ce393ae6728965557e657fdbd5f1218d94176ec65dc4df4f342e279dd6d2fdeb37abf8256a5b1f0a0c78fab759d72a8540c4ee2bd6fab6f71487b37cca8ddaaadfef60a0bfbe7c728a2b61e96011d09208908e4a885961e17c3229d1951c6746ed68c1d83f59e9d90e4979b6c757aa320a96a0145e7857758add8c0148649edf5acf7249caba58afcee126c3b29b25fcfc0ab8015bf943d50233fbfc640af053aa124764bd6f88d665bd362479d6dd12aa40f7e8d2b465873844fa3d717c89c6ef6a6079c690234badc6b3245282f7cb249a96c0245d1b80d1855a563841caaeff4391cac772e8ecffd1a1c9d5e5e4a3c09ee51b5d9793dbad5f0864bde1d818078b21984d1e17044e46b514ad668294149e67a1e176819223ff84009f05b4a6e42635bc559c725039bf755c2a56b58e40e393d8b983f1e3820a2a55558b321529b322353ea3332c321723a0c8bf0435e1ef25049850b0e630610ae4f5b74ccfd2808cc8a1dc4d06660eabded3251afad8386e1ed2734f4883d123a4f477d4ce4edad2488b5ab4788429efcf824fe57c49df306128fb4b9d9eb30bdc1cc460191599914aaa481bab745de984ee7beec77a6e39b27a6612c4bdec1b1c57b7c59503ac2959f135a09dc2f512aec835b383a6c076e5ff07697e661be4e9e37dece53c33d0aee3fed04e9071d549fa12472238c4b3a2789f5e0534c5f3c031a42fef59b698b2b7089b71c50b8e6c03b3f3193c2d8b1771b4cd30f650deb90cb0cb65b9a3dcb32af663cfb79ae83e780f8c122973ae4e13ce3747f4b4b787002e3063ed0cb0f1383a74d1910fc49f6d45851252c6876169c9f725a374abac4d90e7a248e2731ad7dee79be59fe5bb0f9bc01ff5c414025c317f82c673e6edbf589d034734324ecc556f226607442ea8c998a530878c2a13a111de728402087415d82e79e6a19372acdfc45a04a6ba03a279207a7d6933ae38ba7decba5cfae0c822c2f7124e64fa0a05ca152c296539f1c1e7b4b3ba07b4e96158e7b0b9bfb4fe13db6bbe0669a7cdd3e0e7c5b46f124c52a58e6492fb43b9c04b1b066d46d2084afb30de1eaf62aef45226b760bcd957202a707ecc68bea381ddec60d2af5b3c0d5eb9dd8ec3d02e282924216bac17cb91d788b057625ed2ecaa3a87882a57ee529a820540de9c7ad3e97362e39f3bd0be47bbe1de17f4cffc5800253ce4f667138bfdde7428bdf8ea8693347e33ffdf5d8d6ee3da85b71aa0e2a3ec76b48b5587ee594913e120c4836cb0e8a8a05c6b49b8a88003783f157447e8fb631704a4c953708d32e6ab8abcdb72af1e0930b9d0eee20cf21f59e96bb9e281426b9bc8723762486d378b135af7d9e26155635ef384d22a9bc6ab7bc08bf482f8e4cb1423d2c0997fe20d3bee539407010b6927c0e1b21abddbfb87f48953bef35cd1106e685546b390f876624a404ed570b3f35cb22e6c32e97de54941c1bd777452c8e8595047f9c3ca9dc330600e414c88c5250b9b9ad37808b8eec70181538cef576366e5858a344a06fafebeb38171e78ed46a8cdd150cbbfe2879504ec494e1fedd1e24f2e2c397913df67a2dad68519677017ab83e72db5fa6ae04684552e44c032fb2eb926bc814be985b44809be407bfdd3572018514d83683bd730fa667efca227640f92371fd689e8385675870c47fe65c665b0901667d49388070146621fd0eb5b802fd389d01eb911295f62fb9cbd7ed2545038984da5e1a9a36e3bae52a6835644ca30849f80d60215f68d1957b0a7133072187dc6b2298475dbecaefcf39e1d0ad6c872bfbba4ed309c4c2ad68788756c7251ff723bcd454b50244abca5f92949db6bf4e3d86c68449e41f8958d68d0546c2d16b70c6981c3f86e31bf25075beffac67b627179616df27929a1d80bb7daea6e11a4277f9dd700fd17c52db4b9bd3a3a8e124cd5cc770ccb32077930966babe5ec3811d63c21ccadb82274bf117454e6b64c8842acf9a078f69c4e4dc02648db2a7bfa0ab55662ce74e05c19f304dca9b1b21a8acaa2bf8b221f81933e207d26f7c400e84e755b813938e03ed56fae1892fe43223094ed40191eb87d16d8de105704bfa54309bd43d9d7086a45cf953005715a12575c4389236405e190f11badde7aeb32352c4ee8c178bf315dac48bc4706d06ef22027e68b76112058e2b99112964f71a256575c7bc892af2c16a75153b9eac8e8fc3e86d5ba91418aa37f7d3c39f727a7fa3abd43156a2493480e90c0ef13d2a462eea6c4c2a55c207adaf0f2f6ac9bb726723ce7a8930cbeb8f440d5903f7422a1cddadac89ab2cd2ac064f0187e6c2577ee528ff08d8744beb4e18dce135ab03b795027cc1b4eac4b826b1426c5d947c0d27cc2001124051633e14d465a74616bc0194b32e84d0f85878bb3113aa87d70dabc3e53f91fe16583ecb54e3e4c321bc720cc569404997164da8412ac6d214ea0556eafb5a44cc64db6b3509aa1ee0a0952a2895a595166e9ae5a797c3c2ea33c1e26b6ae42166a5a470cf400d916899e56aeabfddd061fbf84c24cc41aed2d8f7e23675e0f9dbb1cbce9b9f6bf95613f00b76dc01ec5efc35fb80350dc8ec02c7ebfb14f6ef27a62f60d83200da661db1c2316fd054a5cc36f0b973b617589b4810bbcb5450324c48a4f3e04e8d792af186728c7380b97026ab8e208558f4482a09aff423883317fed486bad41639eaa741f691b05f304c39d77f1e96b9a276d5306f31cb5d6b405cd22e94dec473176f9d694269b2c2dcdfa4bdbae48b4be415cf9d53642d91ce64c6dc66abe23369cc24fdb6990aa3c020f5add3951fe260dc1e306cbd081891afffd6adb5acbc155d9bdd781681db03bbd2f9b2ef6d7834e1c53ad0bcb3d3071a5645b82042452fd7299c5a0e48e4883eb39c1a3dcea00aa39cc707e05e10ef12fff2e8489afe5bff5a1f143bc9586ad258deed561d5059e9f94cca7318f09297482351bf53d9f4847fa356641ba6ed118a71a7d85f4d3a32c5b4d22ef49049a8baf61c751ed9ad790fab23a810e021780232f5e00a42b82de13391690cf2f384820c7678e81428d4c4de201ff250631fbce372f0fcf9bcfadb41cc5a138fbd380b6b19b63b705a0524d1a0ee573c553b24e6b8cbb29333e949918c2b1a5765b9aa194324d7b3964c0fabca76964e4f2823b1e44f6e012e5bd14ffc6f391f13793457a9b8189680e4d066814ed1340b94bba1f5a2646138faba4bcdf545c1a00f944f8a6a7be9d6a32cee70275b66d8a8f4c231761d363ac6bb1ca4bbf21f6ac8a2304ce78bdd017dea978c72472384f07d67a247846e9f7250a851fe1d1254f9a48b36ab3289822b6acc6b25b6a68d0107ed462cedfe0999de5665c32ba4d4acf76583ccf5fbcd4fb6a8662bed67776f3bfd02e27e6f56df12275fab573351f109768c9cd1ff3f457fa86e76a229f291eab8a79ab7ac09c880273e5c7cf6f419f6c1dfb3aef8a327a953a4a9113186f8670bfec484144a291dca3646a9117cc8e7fc19a2e8909938366424f811421dd3cefa8f193fa4176c5a1788c3f7cf089a3eb1422ccf9304c14a765da33921e8df39cdfa6815b78dcd7edb013df3d86788909f6a7c122eae2e28a0db9151a33e80aab718dfa6e7a61ac2289a4d8dac25b1f1cdbb9ca1a2bb1c256a976745a5e34f77e24038c7651bd82156f2e97b5735383747f88fafa1bb4e0b20a05eb756704d784deabe56db79f8535878c7f3cf25b61ea5cc9d76c8d2d3c9d8cc21be0c7c8ca47d54544bcac1e1a5f9db61b044b922311e6db1cb58c06c224de9b746d153892c7dc0bc76135fac99afd98c77ad436d63aaedf43ae58e3f63e9efb25f212103aa1592fe629a63e25ba16c5d65c2b26322f36fc10a1e314d942ab1414ce0bb7ba7af1ad929f599f43e42339e9a2fef0027e501d140ece2a58ecce11fae6b5a744a37772fc0129765c22d0b6221326c24fe0d878d1065ab40f5ba49306f8f8ed2ece652ffe6f253d41a2864805b18194178ef1cb9218c8a8924a910e453fdb2589d5b9aa066c2e134fe2c81e26d685fce28cfa9a728728fe608183299ad71f03decf5d07dc3ab38aed7c9bc695c7887c3dc18079ba0bb72ef26fe60a84a73d7e20ed96cbe6e76e49db7306ba8953b33269528354c6fdfa95074f930bca70bec8902873baa61869257e4b8790531c2c9d72b4a73103c66250be31f7b410e93e5854ab6845283531d3f100fa5ac89574eca6a3d4226b08b8a0436dffdfce42061e58bb444a0369c2da9fd10980b0f42a99881be7eb1a35538ebe601ef6b2ff9ac9a7fef75ebb2f2d347eaa7a9532466de015bfb2965d70fe51339be909fd5d719308e0c8c3f0dc5236a6d894cbdee045f981d3c1419790f647b39ee07e6c5c2949bfca6351468468a88933a76b7afb5fd74335ebf75426c4dec83fc99274609fd159de429dcb02438fc1b8e8023d04f47a43e7562759fc76acefa4633facc012b698ee7e1258baf3923dfd6bb65ecd595f3ac7e96392959dad6597bf6ab123dfd5af58df9e87fcf5ef7f533ec6c02c382a53ec89eb726589e0b7492ed2a21bd9b0964ec8fd4bef7e77dda2893adc2865b093f005eb02ab3d05102205529172c0df3b24af4864dd0c1e43321cf379b6c31a00a6a957f90546bb3ca705b475338affb1b3e88f9064283bb7214aec5258cc94666dee5042743a7c701c70ea8103ec457aa44ee675104c26a47c787d840f0d6b00a85e9d1cddf50d76a14d99a5b8db7e2f1013e8a41ba020079fb7c91407195c980b4c1395e645275e141672ff62ee66daeb3785bf3ce50772f82cce7e3e981aa7b63ddc4025bb93724af10b46ac838776d41b241dedd57cabac724c5ff23986d57c39d2b3e3980307144460b675a52f5c308192037f022a4a9fe6e32687caa9e3bb05ab95dd2d21f8f9bc7313a5fc0012fc07150becacc1dd016abf94c50bb08bf9f6067814d9437650eef704a6247821b65e265850f7e891272a48b8576fadab839a23eba54727ed4166a2901f936105258745c8c6f5adfc11df5a4535b33596f8dc43f0996b9a559fcae9d498c3f3a9d39f103da5c4fa0398b3171a49d9e9a292cb804501f5de2b18146f6c7defe517232ccd428b04fb5bb756a1d266e32237665be334eac2d592a8240cb9690bef4574b583b77d666d321e452e2024d0f25c57df76b42ce30844451333cb74ee4ff37872dd3a0586f73b329f37b80f16ecfba2e3e7ac7791858fee28cec3bb6b35404cba2991ca7992ed04cae718d584e9e020b683b88e52bbb3a513177a132cf11da30d6c1e5befe0e875;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h65e2f8a12c7a466e57a80d73f82f5294a0d4a7405ad45087c2103f3365b07b92e6c3719fb2406d5c8deb5cfe04b335ee6a6629f919582d8d634d51ae95a938c6af66b3a3c9cb29f4b541043cc51e48cf9f681f72a752491656c2670f0b993f372fa78e0a874352ab0d0b007dda26e4e8ab66771f47144bcbd9aae3fd4a5db550fc00ec33f4ad46a431d75e1b3a26f350a57519b5a6d89b9aca59fae37201a4a0d263214e4f056019c117d93113b245c6b1c62ee7dd57faa0f04518291a25eb196ba117a197a1a19b816cdced143c184217e7928968f6704caaeb7be6cdadbcc4472aeb3c02e47a0dfa22ff1e991c7ae8b8104d9bc0b3114deb902b6b5199b0f866c231146da1cab62ba88317c54e3dba7a60dbc3fefae473457861dc7ebb56e3b9825a280d772987fe1870736cf152442dd7a9fa1f00ce0536b9964255a0c3464025c54a83d118c6dc625fd7ff6ef9e9f5e356c7cba7fe31d15c7e16124753c4f1e314a60830fbb00206bc46bbabde99584d0b9933151dd6e7d4730d4add2f8f6939048e7861d64708d8c95bcb5cbf5909087b5f29ce560405683e1bdc9be6b59319d2ea98898ee71c21c1f9b87de82e06de21ccfc179dc0ebe16006bfd03295d8ac9dfc4c32f5957de50b5e17b456ce5df5b8e84608823587224e0ba5eaf90ec06daf233e7b8244cd2698f5373c5a955aea84c90b8369d6e1e74ad8df183f247099a445878f9e1707320d709eb1951975a479f99d09b1cbcde08422b3b13adaf5d97a666082cc5ba9e39528da0e208ab6294149df73509fe275808d88b57f8335f250baaf19b131c11fab33426ad6c40d14cbfb3ca1e3fac6020fc869e85e784c52a0cc75364449722f5195a81496100486bb276854863efa1b877d7a4c232964eb3dc26237b0e6b7ef87f2697c3522e2f3b32259597270c5c39c4c2b450da0d4b35f7059252f42f23e4ffaf15ff57dd1d5570dc6f4e683230c60cc6584f79dc1a41185e3c105a3a4171097a45e6675b074399d7f015323f4200a1e18f4fc20916999c4f6036688e2509db9e7bdf8e053b3bda956d2e46e1cea275e73e4821fc93aa00fa10a37a29e7cfe905759bedbe42141280596e9ef7c9b5a4ea83262d633255b72617d283958b9c4be60e6957507a4f81bbb8c1e0449c1a5cf8fe45079b1cb48d29512a8e0f801185d2023351094dc717eac850716af797a5e662c8643513e908302bbed8dd2c5eb9451c09e98891bf2b625274ea8f912007392b0036d7b7cc55f0d5afc1ee6a9a2efc263f79a21d70ef99e584946cdab6ecb04428f12ba1248c8072eb6b0bda2f834c02eb973c67c219574f4cbe2dd425bb4c2e1a206722617ad27fddce75b3e3bb30e808a0c4f37f1abc04c98a9aad4257c8d36c8523a96adadb0c207fa087cb814f8e292986c4106d8e671ea3c15a9802ba4b518ee35fbbf007cc45d8d6806e9e5ddd01b004bf9b95077a3a852c8cc769f63eca12ac99a665fbdcd93e60f4c65b891ec20a9f078af16e544aa41513442874e3b4f38dcf161b37c1ddea3d9bbb841ae396c19327856c43d9935ab2e897f400feb2ffcea888ec98c6ee2c5f270b91bbce2c4a66634701c64d1a5bdf5ffbc0ca0c03c31f72012279dede637f3224a94410d1468dc06ff15e7a0eb42279ef04e0d8028463fd674d2940c081e6113f945ab4de1aedac82ead75ca621832c75298156286ad1eef5cdff6b41ffa387dd18b6d82c01c057f2f20fccb628cc37aa325ab85d5f07bfec2dd43158b176144c0d29a2fdad1d75efb3556f5219c9355f4d5a46e7ace6234914c4991ee8af13be5e56c44d7b4f52c8f7e91a8c1b93d39c65611a62353bdf654102485b9adebfffcc5640fe4345b40adc745e41cf748450b882e943873739a59e1260e1ab44af249e7c9e074ca0e2d2f362f5b4a398b37b79143f44d6230146439289a05a6efd43350e585b4f1dabf68ab5bd5465099a0116fd7a128dfbaa8ed40aecc8e02f37b2aaffca9715d802a407c49ac3c092d3b7e6b7c458d519a650ea1f0c5707d1d73ff96428d58045396cf779261af1bad27595d5cef67415f7b61639c31e1d44fbcff0c5e75620bd6774ec6f52c4a1774879304a8d04577b9a4ff9b640a272526ac6b11472c54b915dd990b171c053d0929cb476c22c3702ee37cbc9d9047b213d6a3fa20c4007202f0d8223976e148234ef24bc502b2bf52dd9f83e5f53e59e189e8524637027030cf0a0c8ec9e55766ae321d34af0538ef381b93604ad0679e02d6acb0d3485fee3f9934df4dba169733b3a7c79b56351372c07b5b9c42aa47d1ba16ab4020732e059b212a4c02ef66927270c663c6213da0b0c804b36fc18443d98dd4e99ae58894c370057c8d8a2c3c8788dcb0508ab8d51942bddd238b891353e1fa3dc7a373465265b964731a0ee82c73063069802ec434f85972c3a3f5d3be3e27002cbbfc68399a52e55700d54b2ef160ae0afc40caca242c26e65b4f84e21eafc36e3a27265981bd6c391999efaa5e32a845eea981aa64b4cd6dc8498ff441e85868a512af2eb3b05b3dc523844282282132e18f34b58e6883e1d675536b998dcc6d7c83b558c07acb4ab17087738a9d86501a25ef07bc4914841148ecb6f7bc84aafd75cee1596f3f596461194bbb9852c20df93306d24b82afd71f17cc36a13e148a71aec0e13178717664ef7017989964c25cff9764d837039fa9e997dfb9ad621fe6df7304ca6c378d5b10f600394f7f373270dda1ab83d4dae252c64fc508a6e04100fe5d87316287cd7a2a4e14c839a04d1a8c6d1e015015ff6c324facc9cdf2f3b1fed8539abee31d1a7cf59aed95d1f06887bcda23bb40a5624ed71f63555b30447f991538710f97193510785a531e63c8c47e2d67ee57eb730bc8d584077a51223681179ea5a999a7f70a17db220c557c23a72fbc839e2cdf9673d6b6870c3cfec2c920c76f26e938b260ebd96f5d8a950abd1e77437eabdc584ce319e9276260e00991f79057a27725a8c0526b7528b7fdfa9e6f684abbf29644aa7527e17d20aac07569fee361ef10c20caa24f6ec371960e38f1a2b6a939bbecb4173118f06246ba2efb418f309d8224d1c7aeb50ec951c4b92621025d456ff5ae29162dbfb6f96a79e6cbbc9070647a3ac150b78735fa0480948f96f23c91b38244bf82220b390942331926b78d20ae57cb199570df07c606231bc64d9a13726984232c1a90efa6e4c056bfd9a8ebd7eac1023cbce7964a99d31f4831977a4abc94b09c7770cd7af7368ec49aa0b14ac0d98902f523cd1c5f9170a3f1d7c69aeb4783dcafb4d3ca7b7779577e5a5f40a5223dcd19e263c7f9c38f905d3a40dddd86609331316c3e78aab971a03271c935e207edc69fa7a989013e4b8f4cfee1f94b1ce185547e9a7f0e3ed32f5b0e4de9583131295971d6fd937c85b3aad5916e7b282fc6f4b40a6e115ece25c11db044a9a59e57fa70b7722ce06bf30c81674beef1d20d62034fb50a0500a3179cac7e8274c50067bf961ff5e7fdc766fe08e49b1ee4e154aeb5211ad9d6343d1948b4973fdb5dd2f699081ad96adb0b9203d2196f471b545807d02a51860f9ca0cb6cedc1f7f7e6f8d26febb810f874df11388f31ed4301b0a32c04f5ae1768efac4dfc323d9f2d81a477bab61aafdc7ec7252451f6eefbb5b150780179e602c5f16b05bb02a290bc8ea9d250f33c2ec09e0ef9349b661703339ab643888e636bc1a1e248f996c5469f5d6a93c5b18d9066efe877e92b40b4af2996f9e00759f70643e56329e3b32dc3fc61b95dfc4cf2e236b0c369510e06333aecc7dfc4160d24f8c59b2bb20a903e90c5bfc0e6803b04a9a679a019bf4e852de95221f7560d867244bd71110fd5165651fe4f732f45f8bce649bc7279a9c3b95cdc8993d3ed77c7bd0741ace22b8264a732dcaa8cd895fb34c0b3c0f0bc0b0e564ce3bf4a7899133e021f9c4dbeb9201dcf0ecf0d92fe987b93d38bcd5db1411b5a328a6a49601cd29fa0141577e4f52830b14f9d5cbb66b09b65641f634eaed441652dcad035d7b5215a2a4b67d5d9af01a806b5825c27d4cc2a11a7cf3c843640b521012578df2ae4adfc0c2d55105793e143912df4aef7f73d32d39ceb812f417e11e8e33e02d03402d3fbf86f1c33c725b6a02372c7de50b7f6080ddbed22cb3245a8aa79bdcab263c201126fa4b51a01b841fda378353e9a58cc3498d539df5ece7760c20f29786f5ea636dfaa5c2062d5114f5600046b3167d49fdc039d42291fd01876d6e37b4c6f0476eecb2010ba71d1b6f4f0413b3530ecd3fae577d16f5bf96f55ec974013446055ac70fc193a7a3210dcd6105a2b9c917a0078eea3d5aa0e359cb20160e62dfea4787225a00fda5ae4ad6268bf445c16c2e9adb3d6d4fb517870ab4605af6d9cece349dfc8d24a1c363aa72db5e967fe9bb4a415ea0691d7544bf1f9e1747e05f900ecbf813e66807b12d0a3694063f0cc801a33a1d2508e6e266689115e3428c138da4fbd41f573cc7116c337cdf4004cab82150ad0223bbe4050cb52a70f640fff22ad43b2a1667205df85286fb59bb319d2ab3d9035354b0ef8cda5e43c9dc98474a60661007a20605d3df6b6f5fddac4a8c118b9e0bcdeebdd761dad0b7789aeb3d76e8720a3b9bd437ecf1459aa4bb28f1edaf82110b10adaf90ce76a52b6033bc2727e18d2d8781ae37d6276b4419f49996829e412bed710eff5cb3c1bda79b663485977102d4a090c85f3d99e12dc071669798fdc6f9678bb88402bffa8e6200fcbfa01bd345c308ad89198c875601b79f42d63aec038c5eb0100796ae5a66baa782eb12c7f057b7491c9fccecd0502a32790a9b7fd0f9eab899a2044864c403debda8542ca4c2f7a45047bf1126bd24d3a6ed89f128a9d95c6d140ac8103fcf223475a47d62550fe0896835a5e88e78722bb1bf56228120b5ced8e8ad243d1473b24b62582abe23501c8350eada9c0aa3bc04368519bafbb288a671671e1dde6d37e89da0b02c1bce323b26ad3e7203a6ac5cbc97ea3938c642d9afc258143867dbf9d5052ed00bd6e3f99ab422de7bef4bfa69c39b825866d4c97704701f44454ec89b8c3730933f84e7251bd0f3d80d0cfec2e41b3daba7101688a03a546fabbe834dc2435f764112ca38cb39e89f6284dc89396737247f575a0bbcd50e487e2cc0786539afd1630e621fa770ae99b7a06aa4d1a7598a61fad85c22883ccd01dd4a73778fbc30df306015a5568a21b05d2d81ce2131be97c054401325b074606946279b4f16608e76c5dc55ef338921f32b25e4d6510ce750bef8faa48107c1c3d56aa45164edb788460b4bf8ba9cd6edbc330dfe5f78bea31ecd34fa906623471e9124c67ca802d75bcfdf840f7d8489c68f722878c98ecd69e3e1a73291b1356890077abcfeff5b743e663d2574eb3f8296120b6bc396b3c10642e051f8e14542c4a3a6997a0dc7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hb84da91aac25bfd0927dc0b30ef008f0617eaa6d5ce8a9ec919770c7e73235eed8a4d22390ebd112d25855d376138630418b8879b39fcc772a52aaf3b51f9f13b28ef8f93d7e468a92c5ecc56012695d537555a9051d94b3fe09ba17a0151d94e7daf93a7b24a9f12aa72924cc6fbcda183d9d4ebea2c37306ed495e6a364c58a2441b7ebf65702a6ca677f71a4515a5f783813ae5cbfb0986cfff2a69f87b59aac0641a22e2b0c0cf45772330b591eb918a1e637bb2278d54b834c2f9770b7b85e308f65afde71a08be81ea9edaf7c3263dd53ac2bc8b9e057e9ef2dd9e8f5b5768f96a8d099cdf359e4766375188f9b0dc03792130b088d2715d14eb32009571d6d2c75d51108f5e083829414684e20c80a093ec1499dc746c4fd0007898dcf8e41ec1018da2fd1cf2ff7c8a2e5d1bef82bf679ae5a38ce292d20e5833ee84a86c0142d0d340358a3f7ddcd71e58d25c16deb4eaf3c81fbbb77713b34bd27e83101eae0a76e4d5eda57edeaa1682007a22aeb7253e33a1e4e240b58b9dfd36db5f652e65969eb48f211ab00e40680db715c36d61fba673a31f4feef531fe818e168295e393f818a8987d782e24304306e51c25a87084e2add30327bf04b53494cbbb01733ae875cd984fcf793f7ac37d25c286657dca54f8d812e23e27e473115297efbe217177dd7d4a2e65eec4eba97c96c86c7aa6ab4a505f1456c55f4d867c00745537b6168372b393267aeaa01e9d6d93d03e3d1e80d9e6dee4b0a448d09d36f15b03fc95e5ac3a51a63d3f4ad70cad50b93e56bc01f2c170d32e09e22e443d2738bf34f07e35ec71076c8ad2cb77a3fcb8e04f0b502bb2477d69111dbe4305d75514767870e4fa441364d89f0f4e8b35b3f7175ead1763236c3b47e4403637b65a19575a3eb97c957f913d3522dfd0822465f3b1921d3af53dfbc7e1716420b6411502d3a6d94aeddce77d24903d91432b50c2c61809c0c19961e3f58a446ac39ff1f20a59bf987619fa78bc86dd89e57249d934b5e6ade23f6a0881b17fa35ce790a514356aa101007b47b0b2d933fd06ba9e6e4f9af5609dcfbf5f604213d95549067e9d9b537f9ffb34eaa67b3fc6858f6c049204c3c4038a45af1563a6252c8cb159ba778dcf4d10d14de8d5df30f92ff2b10b5139e6bdf64bb9516bb2ab36981da44ad090c46249b60f15d0ef5f66c5aecf53254b162935397f1c23fd7a1323abe7c7e927924080f22df24e9fb3d28b043ea78412ee0b23f5b3f2c45c959f4dc84f6a89e515a83eda12eba752f6572c9f84114ae16b057a64eb0c10bb3bff79988cc7b40ce1db7cc0b2283c8793162152af34c3340e8631ce4cf4878aa28991982aec0e76cb9f03f2ae523e11396b05bdf4b06454520b13bf7de9c074e4c0c8bb4f91e679130325ef1b52e076a49fee3eb87a886997e880b279d1ab6a57c319ebbde8e63030ed83d4d16c290c60d04640627f8a3e8f3b10c87506812ef6fcf7d3a0d9776ffe76253c3763938fbbdea071f42a5dd987d41422da1af755731a47d7f4558be91e308fc38d446a2e17f59446bde98c2f09e19773dc03f75ce1e97662bb303ee5eed9489a5a1417c9eeb13aa32e04c10330f07eb62ca453dd4dec2b3551997a2c3cba54309f5740a8fd8b2631022cadd95a633654f75f2f0c5bb8cc8eee67606d58d2d70cf93a3e0947ee4bf320bdebe7057a5b9105b59d71062b49f8337c84d90037fd949e48bbb7bcefcd3eb4c7185926e809a69923a839d2d1f91bbd1dd4fd6b30f0f036b730f7be2425169c8584bd6ab9dcf81717a8fb673579bbee1b8d2ed3fa2ee253172d2f64962c067b33f1dae0107b0b5f6bb8f0714248c73b982d29ed411073245c49410eb0fc9f8f70bb95fbe8d7d861007364f9b06aec4bedd5c38d2ecb7f1f4e8b91f0329369f2546912c9c22b9ac700edbbc46e2ae113a758ced1fe450bbb4fdbbe86522e5383056b14e473328b4d3d7aacee2bbecafbba99b562a8821cfd86b13a887504cf7a701b4e96f0f742aaa0d342e16421caa642ccad03625a68007985a8a34d2d0a4ce8ce93ee3b688d1ee8ee4557cebfc4b23a6a7d5cb25e625ece2576cb6b27bdc5a5dc7923d239a2861102076dbf973fd698230b2c87a1a76145453ebcdea3952f36b07333bc280a6f51dcb88bf1d12fce729641125d5a455abebde625d93f569749b61b82aab634133adcf1f8e62544516f24d513c7bd5c9fb48061964a169b0e9d0b9e07cb533bbad64f5b0eecd7fe99c9f5d18aecf954786ff0891f438dafd9c5755d132dda833606984be4b0840463ffd093d7ccd3e3087ff21c865902bdad91ce965e8e3871aaf061c24e71535bb20e6437ee7ff322b25cefc97490d358b4de9e63e3a157745b0c06cc377c418517a424178930305cf5ee96869bad5695f000912e4eb1b61a05dbabde4cfcc96fbba9f235bb767df8fc98f0e7cd4768b7d774345ab1a4ee5b81f15d1ad914a588bfb9a0bbc10080c83bd7b0be5760e9095f1cc36ad2e145deacc2dc37bd92cf5caf0ad23ac1260901bc37c800c9fdc64a900b05657fcb50f8a116fe7128e0a97f0ff2cfc69a32fed5979b366bd8254c98632c53045584ed86b997205c4c7e4a2ba5ba37fbc748812668eacf73f5bc03a25bcfb7857366492ddd6709fd50f25d45e112f4e24662513bc6b872ef354d50b43f0ec4cbd777ff40dad5a36e4ac3d2a56a6b0ccf5677e120313d2f538fd24a858740806fe17603643def6c3516470356730f3c14df4f60af3dff2d434086dbc5d35029c5ae803d1c244ed419b0004d80b8bd663ceb3b5a6bc6f053ff3dfcc0c2b8aa5840c87c3d154da97f901158ed8a60fa2f877d8b665ed9a14d5f2994cef89d8ac739e544155e24c4cfd5fcaf741a3c7edcf0634d722f6dde35e353d0406ece7388e4b39f96b8b94fc3eefbf7dbd83ac395aa4a81907f32a6a5d1fd04abdc03f1e02a9f702c52f4ba1df8bb091e268e8aa5876a6fab1fdd6865adac1477c40a02b986617be3cdf8a293dc3c24ae5b4b478f4d2298550ae6f0e375ff28731db1664a3c5537b29d5b2763791ea923508974dcc1d29ec693873241ba0693d5aaaed842d5ac0a3cb8443697db5fde2a75aaaa461d567106f6ccbcb71023fd38f509025e985ab35b9b512c9b3656fa5c9a620698be44ec5895c1932be1a05d59d8fbe84f48bbfc682332ba9412997fec85619be6b45694cdd6a9da85f24dabca4f598fda19cdfc5bff10d438e635ff052c3134b3645801888bc0b506e2e322224ff7a7bda33976d634dba2a1331d95515bf772a798b1009ba7f65be24f804618da83458d63bab1e08995d99ea38ecc937449916b7ae0cab8a7b94c2f4ffdde27a59498e814dbd61b0efff825058e4f767e39aec312e7fd8a8dc3b631ae508b309c7daa1bb8268df7b5c5f04f3f986bd48226df5bd5b09dbfacf7809f4c26e22185aa11a11fafd42cffc60fe5eec014ef8bb2a3bd92546ed8a1b74280d8f4771aaa61cd05d64511c2fad9d0846c3f46042ec6d381190af7cf91fd23cf0fb32bed1d9a746255c55ec5b3ed888e634bba33435b4668bd9d1cdeb38157e6285eb2edd2fa4d1b747edebd66d4b9b136383d9373740bae024e2865ba83424ca5c1b8dadb6767afd08fc333176265cd933b1e0bdb0d1cff065656d1489724618e55d4f78880fbf85f4607d5e3c8064489a3475c098dbc3292be4f880cb5aa3d59d56e107f0d383eff861afec8166454e4da6dc4b4acfa967109e0f1da12c074ce43a253c0077210b7a2c45abec474804b632ef96284a990584935ba48e4632f7f9139db4be0e33ba1e676fb47dd05e9f6044f3a1b1f8f0ee70b41eda3818db9c047d712a962356ed62d4fee691968e6fe47128f7f70199049e0ff228ac9399bb57520949d1a61a0e1ff8391c29fd7112d683d509cb079611a8626156cbe68f1f8944528eadcd82101c80e5f5f6623b4dbd857b4b1c504887b495483f6e6b2ced396aa931ccdb1cff404c576b68e430131a724a5fcff8cb9a3a068f16e10080c0a5766bf3ed5189588e70dc0dfa0cbea7194c9f1ec7fe6c743b34296d9e5c6c00a15959fc4e611145400905dd07625a1c4a8dd44771fe9d1c54aa0ea7c3896d92a019f11f5c0ccf91db691d808d8e86dddda403f3b631f121afb896a4fdf8d4002b8fd7d5a4439c10d18fb7c036f58fc99b3ebbdd40e6355a28995ae61475e63c981897ecae5ee42c2f3ea4d45ec5ea39c56425b816dd6fdfc62674213960c4d6709daa65e258ac8b31ad2fe90befcda9518aecea6c9082807a821fd8ec2229d7f8ac36ecdf9d152c20b673d71a3799cf8dcd8306f6d191a0aefd6a3f168705da1b960530e69a1768d1a3c58ff994f0139f2b8633eff4f150ff66fdc20e23e6a9937c3373ce7da86ed9a857ef9b0424b52bf70de58f16c60776412bee1aab7b445232be904bd603ad58455cbce5fd27ea8df9aef231b9fa599d8a5fb733ade9571bb2432e4d2a6f55c1a48e92f012bc6155ac521931d4ee5ddb2f03c6e2b240095dbac3923bcadae6688823546616d28cd4d13c6b91c9d6aacceb7485c8d0d84524df6547c46e9fdb9c925c4677fd88b4fe414fb6e9e2d29b67827fdac4052c3c1936cbca3ab5d07ca49b9302a5724304705b22307755fb52caae9bc16a641d763dee069b77fdb1d20d20b9974d1e7f48a0859d8a78cefac2b3bd21a77367771cebdf78d50f08f2616ece80dd443c852eb3c24988ebd1c5d73c9afdef9ccfcd8c21aa0143d238db9b77221f4c249d7b9d32106dd471b7e4670c46d26568e5f7a517d6aeb46823e84cb8a303e5da0887d35914b89721bd5c48cbbf7cc734e26f4777af23dcc0fa362d7ccdd24184d5266999a062ef03fcfff678d5f120d36bf8a8b2dc7fe8a0489ccd6f751040d4c5fd3b04f693a0cde70f6e3d49196e396795a7b94714bf20477e70d7284e416d151b72092e77557e5614748b13b15e3f9237a47a231cf78dc74899f60a9a65d9d9c00763f643fa002d977cc69edca7e08e2d71a956759e6b3b0dbaeff1570b2e0e093372e9961b622583ccefc86f3e3b05b226476adb4eb1c4e385f03b8e91590f50efa7b124aa70c30d0599f630bd5564144ec8eeada3cf59605eedd7da88428560ac21a60cf62585cf463987dfbc90e6a08641128a33fc05264cb21793855c22be9d17a6adc0377449467f2d1a615075301c04e296a0225c16b576807c9804d281cd02ef9f002109b25d0071fc67854adb4f0c0bd0cda435ab4af0a65c70a754250dc9c435e9b2311b9fe7585c4f57a479d7fd3bdc24b769c80332a91528aa32d222985f95b99017eac01630bc4212af9babd694018636d8cbfb330108975945d0de50d6fffb1bd1671dbc6df7c8cfad39be9e7145d1c448cc82adf5e15b1e1ae189a71951bf9ff696bf443fbcd788680a79bee8ec3d0a343f883bbe6c048fb3a0de0fbfbdef0bc08fa8f1c4a91d95b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hed6c793cba7100341f2cd3fb7394d5672caf3e96fa403bc38427b0c658e6a28310fac3ac2bea05f8d1721549ab253e363da1f534fbcf46236e2045a110ca8f842d33a2db936cc975bcf3576da5abd24540b79df12dabb9778c0df1bc58349b77f729d6b562f245ad3db8c0f80953e9093a259c9869e922b7fed4cafc662895f914ba5abb01423cf7960b3efa11c9603564c63e0f9a80835b77ff62ed510e6cb3d649562991ef325ef819e45130a4c15e05fd21ddcbbf74e8d949153b26f9c578023fe5688d5cb3ba140c7f64edbd9146995a55cf511bfee31750a8d669d0a90a26260110c08f42e4d679c066557856319d58e925ba5586a018a796800a75a0711fe0765b60557a2d7258566587cfc7d0301dee8436e55da67314b9c541ce642e805f3da919a269d357c5b131faa312d649ca0f02ea7559ca2733a63a31a8160e16d6fb088257243e24767bccb548bba9aeab20262ce106a9701ee6613b40b4bb119e7c1b4c388473b3508c168617340973be5c54569ac5a1a71146c0b837ea273fe3eac177f9eaae8e4b1a569503537cc8bbb24822ba4241287434eaffa89962eff02ba89e23cb34a3a246ebd05aaf928018e7585000663ae1a3ffcb87f17a011025b4eae91c58cfa8a13b286487fc08a06148ee2a7dca97c7c826f5474463cabcd81d1d9f19c97ffa0f67502ac2e386843092e2397cc3814db2729d2ccf1c6b47bc3eb65e823e7d524c3fc0c8da251eeb148d27be141c92f3f0ea5091edc9fe7ffb567d6eb65ee183ce91476a9d5a4e15f5f67861ed9bb318ddffa8ad261cd87731cfaf46b2a0d112c590ef2df221205e455a9f49b62fcacb3eb726515387121c551552814cc7adb6c49b2f9ca35d1b48bdb9695adc42dc81b8da5d0626b6d1637b39cba7d100d81dcb8643eaed4c35340916ac5950df35d15ee252d49da1dfd8d81786ce96e6525af31f772ac8988003404f2c5070d9ce4559b46026c4fffeae6948cc10d9037cab63b7a18d41f2be7a3af29cc002122533b1061e3cd2e1ceca84fe68d8c9a89c22f326c2892e719c2151553404611290d9ccbe44124a92b2a0043336317f7ade978233615e42f294b58fb391d60c83952afddf22b5c9bbc544d35af833536c8b20c91d42f12978280693a76734158fb0e52ba5c4a397f278ccffc86f9ad67b463ba3dca28ac2512a2294a7e4c7e04952a12fe8f142058be311439daf278dca58c118fc79a6c611a6158777614bfc16e9b1f5adf57bb2d75f39c0e762f5fa0025e2d4e6700c420c0f2cf10ee764630c172903770207b5e532f3cb514309e6a97f032daee646010f2211058c05b87f813f06d756210850a0f6e4ac4edd8979fd3c6084d47a3d1720817eba6b4b268a03232e68a7a83063e0f548e200e6f3258b732ec7effc736799397341b32da0dce099dbfe5a6f127693e9c19b932fa35d808bffb8a2deca838d8509b5ffd86a9bb28e786ebd2ebbe8f4559bd24f1ca5d85634190e97c4ae77ed309fae5df8ce36a025fb1e6b9cd2a9709948d4e0ca906c6be31c1af48cf45fe3fc465ec2d19d964188cfea2bcc8e0b13aec3de264e22047d1084a49c48c515cf12f931475b034e2cebfd33683a498955c034d72429cf62b8a4cabbfcf67b8e23cde48a233ef1194002ffb5cef89d1f4e5f13544396a66ff33145ebb02db7d4b8b2f4d489711e2401cbd9ade7d1182e8c6ab5ba662c5b86037f72cbf4c1c117ac4de6c5b22a542a983abdd8582bcb8504589af796d2cfe5877be9a355f1f48e78f02b34aa0cf9cf42aee5e50d840814beb4e029b221df5ca47d2a7de2221d6da9fa1a79fc7b092fd71ddeafec63d98e797f9adf605b8b326401a523767de5aa740474fefd89ce0fe0a9033a18a832adef30e05666e0dfcc8b28b26a5c438abd21204ae90089090a8c707598ad0030bc3baf692d77b94e80c81f462dc010ca6ba33c89d99f3e610006da8b74f9269a1b2d9ceb449a330d9a7f23862ecfa67f0bffb09a076011360683fb99fe8f3523f24aa7337a9422366d7e45fbddf52555b33cadb58fba55d379de521d42173b4994054c0d35aa041442c4ded65f2a67d06e3df3d45bf75b59a1bbb08f6c3b2a575ad30f73cf808a541347ca2f4f0ad72ab5743c77f21dd3a51176677bb3b3765298b689f9e062a63f010efaf248ea88fac3b5bca7a9cc300599dd1f2a6006982edfb6c3d3515bf240a79e3971baebd7341add5f22c0e25b753aa092a612596d0f3373f98a496c7d6e38fa275eca195bfc69c6d3980a361de3832dab9a50a10975da89090174bc4a689a59b5794101f50559a16504de16388433a7ee8493c2fc7332d156fe0d57a239354d7d405f1ebba7bd316e7f35d640a304728d814c931356d7a8d88cff3ef73f643e0f079ab2c3bd19644684b6a12d28badb87dd2d2458159908dca76a3c0c3a3f0f02be10e57167c26e3637c6eaea14df9b59853edcf0a20b6b6e5fcbc37a8d31eb1acdd66eea558686109554cf2ce2db63d71d73bd5c1aeed9c378a0330709c4f529b5af59c9c1ede583748263dc6c8bf84960fd230edfff75ba256a0f783df497e5f3e3990c0a9433ba7045fd52e69c10596001d75e5d227b48c00d9fc1853716191590e8c04125e0e50d6014ebe252616d9fa20c60a7d234d78c5715080f6e4855d9e6187cb2cbeee856e016765c7a9b38521697e59aa4cb77c63d3ae139239cfe377b19ff45980ba74895c2994b6a5273201bace02851b2710fd88af7a63c1c701e9212e746000071cb9840e998b79b9104d6202671db4107d4a82682c75fcec2b905ee77e015e9f5df7b594067dd2363d8ede794df15dea911f7090b646ff7cf092829664b4f10157c4c9207ef5fa3beef5b6b53ca46edf36ea23fe993530edd5fdf70c3e4134a977a62d39ca5cf2c98d34173c64a384c5920238e52d93092d64df006be6a25010a4a8e70fbe512bc6c6a7a09ea0bb79d8e068b37ef4b6961d904fa11c39b866ef22632d291113a001336421131b954b2b983286f83b2576008686ccd15dddb243dc9a3d6347a7f5d9116eb6dcb727fc73062cba71432c093a6333c580a32fb048c704c566fd4417226b4c7e03ee451768c8672143eba5caf235367fbde762e8048ff5b04468385de9aa670388ffe7a2f9566fe5478de9f4e9f3eb2c268b44cb22a480708aaab5624a3aa8d1705ad0f0a6f9920ca83079146c5d6cd198a90064c437164ae8182bc61d6f43262b89a1de7739567367c693da4c9b7d7b0a23d1bad95cd5249db4fecc01e1e8cdd5d450a3e1910806b2b9e270c4a2ccc9428fbf429fe9dfa7c7d0f9e8c228b2c64177a210ff47626631b68b2c9499f45b77fd8d56752060341c786241452ce8a0d96cf08600e66b81ecf70d3902648cfc8c8469bab5cae1e94567648776c44f2190a8f6b69211413168b1a79d48f321bb05ce5d2d302c430265a4769fcaea0b173d3ed5bcd7a528355fda35c4defec960311c8209ccefae9fd6bb4a9f5f3ba6d0d216ae39b5bc8e2975f3a41376f421bb9064d67d31cd7c365278e3e1f9c29a34f553aa78cc9f98972ee31dfa11d183a6bd81f5b6fb910675b46848a8ba766e39cf0c7388dfa8a94b820c77567ef4e1e24bd050872204261121eb4e466332ba308148926e4f6d0ac5ae0943770efa2d36eaf1b858e380ca5b4216e715324eae2dbbff5034ca197bdb5cb69412cf0fd19c3238e5eaa27c5733afb21f93b4c5d5455a87d5b477a12f4eed14e3798e1237910862a5cd2b55dff868fbbeee658c8ee0422785b031d35daa120e689e9249041db2e0d22b5a3bc14acafd98cf7d79122a3763e4d288e93cb8041797f6d5ea1b9face846363baf7c996a01eed0202e35f322dc814a21f108ed4eab6d310484b556daad5cb39c5d86a40237e3b294816a6c6ae4a3c19ef6184b70df9169a52948e7d39774da270fe2efe20c0172cd55482019c26959e5d4f613d39daaacb7b70b41e72b84f86eb1ff0e59232b27164753627ba7f2d2c869a87924b4f0253ed0544b2b3c83fc01b72dde37d82b173f083c5094d0f500c655dc43d9a47ef5adf553dbe2688d6a5d2b85cb590d7559cb2224ca1fa2109eba4dda0257c22a3dbfacd64b58e48397997ebf14b716d05f623c4b1247725ba6424f9e3879c7ff6708a5ef476233fbcd303e16cfa3dd69914d66904be5264db572cbff79a8d5b6132597d2750c063d0fa0f0a08e0fad4e3ddc2a0d4484d99027084cae22522088a82e2932f3a0faf25f9bb3133309a85aa7a1c17969acafde2bd7d8e3dfdfab8c5c3d3b31b6cd113abe4b27fb728fc6adebb943b52bf1676d6c2b01e15b2f6edaaca6679c052abb85a09abbe9db69a426a7ec7cbcc376408116abb692ee77b2ef082d57c0efac35f218f88e61f7a7f2a68169b6ffe9b7b556abbfac51039bba45bb814fb744140dac7a18476a59227543234a727596dc6eb29b018e8845c190fd29bc938acf38eadf97e7e7fefa000d6bfc482813f7303bbdf0048c285ac183c932dc1dc130b70e92c2391b9eb201e73610c885b892fdd556755be39185f170bfdcbc7677291505699ced3cc64edca2f211e47d7778cc54520a424a21a3d8de9c4ea6aa8afa5b06d5e47e87199915b63c91b64ac67912ebb88e77a81253bf73b6fde69a62b15faca0efe625a8eb8f7c7ef88fd06b52aef946daeb6a4bad7edd4fc8df6dfcae92a8087d0fabcd636629030ddd41e6ff3e0e173c45389c0b3757d7a08f1331ef8fab3eb0e8bace3a35983a17e5b45cffa51286099cc0932a602cc94e2f84fb33222a1a15e4771de932d47c500c42f72220b28037a4fbc7119044bb54e4bb4aa15409f8cccf99151a4836ff01afdb6319213eb496e6605f3c15f72eb95fec0c5133b575567cb8c25a1a326257ef1be0742d00db441f75cbf0f468f337b090141eec2bf08080504d3463557ddcbbb0dcbd45955cc8d7003f0113c573db77ce0e24cbe0d2b3bf90bdd8ab6ed58bf508c4a3758cfef395b90ff9437ed2fbb2e97295037f22b735d398a6d71f41a400899cdaff8136cc9c5924c045f57d19dc8d797087e8e4f1e553edba0120b3d0d8abbb17b7e415fa03b20969bbdd639140c3fbb804aa1acf613b9b3a40ca9dd481be99ee9ca10f1d93160ff8f5d573bb1a8caf2feccfeeefd2d15fc88d17b90be7b59435676a7b6506d8df1a09801ffd09274cba2d59224d1c7c747b95d01657caac3f59dc5b25f98267aef803ceb2eab8461c053b06db4c6834c896e516c6eac1ae531c9220a8e07797192675906e92806acecd2fe8c0fdccc51200a2c86a51d7ff0719cf44dceed52a3d42a4af58369f798dd287826f99a44d9db079e74aad153fd7de4e8277d14819f7a04e568231294f1cb1e9b8be5fa83c66b65c1b524b574f8c4b90e48395917a60476f30335b580be3f99ceb0d5b299280fd563bc12611873c971933942b5b1946a14555961d51dd8e5b81d55b05414;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h28d8b11406579c81b4e857cd762a3d24833c3a58d3b3af38a1ed56778814fd83805a67bb97ef5001c396d5f00698ab20b478fa8cb0a99a605bae6dce6958a00a05378734451937f3a9fd46818f74c0a8eacf56796fba307a965f0510bf11d4940d14118aa2c9ccc7199acee88a4e132aeaa0379684896333ca247ff0311c66b859a049b63c117e0b82edbbb5b54c9e31774fdb39f1b372cb9758b8357b5d677df1fc795ffe5b2b59112ccb1d0b1eae74ccd6a66a50f392fd8a210564b7cfc803204404927589825c2f81539abdea552470c618e8f8cc4caad89c6bdef8afe751bc3f1ec2737500bc0f6e53f8c9cb4c3b5d4a70f16bdb2c541f960b6331024a7155d4b13c7df409f00d4ddcee39f1baa6c2ec82229f00f28097633760c6311c982e4c4b6969e202170290ef99eff58f057b555d4e82a62b34cd2ba24696adf9ed48cf0ee4e2b528f6f607280d54134831a0f1aaf4dcd6851d4627bb10a2b78e84048efac5972defea1a56732a5e17ccd14d07e2c449bbce5396a8f6c7f2fa7de6131319c750288c1157bc0164da52f47128357ff70c00586c853bd1f6d6bc678e7e023734c2e3eb0bb5ec58bb7591e244d7a5f43741d489123c430c050670d12f5f9687dec2b39c95308104742a5f684193b59f36b1a7e5452416330e6e5b57101952a4dc28035a9d8da2e4b6fe1818d68acfacc72611dc61c811cc5bc7747293580b4567f37466b73fe9299eceb71e602d0b9a8a43b10baaa7c4cd8cba94f38bfa29e4827b97ba21277c3c4dd2f3750db4da86cffe1d5071431d70ecea30bf41f6bea43e455b331df4f1dfbc2428228e5c49330c026f7bf60e9dfff9d3aa14957fbba86607ddebe32fc9b14c1b471555a63b0bf418b1fd3b17294dad93a7c2effff5cfd1fb8374f803be343acfb68a291925db3054c36d183e3faec61786c34ef9fe43935697594c0681286666f95a5e8fc8ac61dbb7eaac09485cb130a4b7800854003f5593a710542d1765593b3a081909b05fd2b95a0450c48d748950525a34ee9e3e0c5060b00af9b5c4de21ec3870e9c640abe513d1a9c02a43c02fe29cc90cc7783cc65ea364b89e6945374bf7f4c185496ccda81070b708c6a8f8cabccfc1922cbbdded55b4a14c8ab050614a790b4c384fcb25a0987947e72a595ea5b0e5f3120f138c0f3c80ee02d8d8ef5323d62f34bf9a54d8054656663dff30059d2f9f21b9e9b4ae7a3e79a74ef1bff5a55df45884f31b9999fdbb72cee1f8c5fc95149f72d93b0b16b526d2998de922b9c2ec15f1d0033d97e2e7c59d4f871073d155b5d2cc43159c6afa0b3b4c6d26741dfaa49d3c5ca33b92c06fa6b37ca2584a059989b9951a4f2d31ced6f85dae3c7c520aed327f8dc9d94ff142f99df3ce17fef4079d5259537b421f922d6f5e1fb5901dc74bd024a718304227cd116b86012bf26e85e4a938901231897df031e414f45dedade5c3c5287c74203525daa968e5a68398c52917e4af1b78566e60920b715209353f886c44b9af41054be62d7b16f69f17aeda74db70b4cf9be5f8ea35e1487be5f9d34f5cc54bcf72dde848f68ae815b51b0362953cb91dd07f15c63265f26de1df45ab10444b56a69f7460695fa6aca32c52697b42f4d93c392624f6cc45f626c407603547820adabfd29c023f7ff71f295c191f7d69299f5dc42cac8b8ba4ba282fe3e57d706b07f6d51b60d1aeb7815173104b1a6866af9a5af7935ba878f507a357b38cc77617c21d28bfaffdb2bc4ff347d1c294e06bae43f4b5b05566cd1e5603923156c2e7a405a316bc6fd0c266a17933de9d25f08a97402f33f55cf47796611e74a707e21922ca1ffaf758b69569245407a82d17eda1280bb6d1762c0462332cb2878f2a22b7452ccb18941472b57920db6897e0a0dd259cdae1b54e2af8510a26016469eb92ed735044a7f2aacae17077dfccc5b14d569b5ade944d65ee012e0a1334555214ee551659ab3674289f5da696fa2f5ec62053b9f1ed162336a64aafbbf3d07337e06a34a3ca326b3349665c64b2d265dc3c0408dc266c0d4d7850915cbdd068418ebedcf922a4b4922b8fc38d6fb3987de92236f4b4d9829181586f3f3f482aafe62e4def0257280f3a7f9a1a0ffe56a657f48c159adf3dd9c5f3c397245c612a81b786efa88d46b0d164a0eed1f030cfa4f935b2bf16cad359e3594ee0c73c9a76da382eaafd95f0cb36cbfca3054d003282748dc570619eea03354674b885e2d3c17ee412cdf16b93a3aa36954250db1eb56d23b5ba5c117851c41dc2022238a5587b153e01177260b44518c2344ae8cae77a0c48c7f7f25e849f9de1fb0bec1f61c770ce08461359d34fc35b3d77ede6f34fa37a29e238227bbdb357c60d6abc8c9d672a6fe9d4d92d0a3337b67d8b82f757b784fb0a5f2d05180421e4a90719be327c4b6313cac9c32ee0c759cb1a2326f5060600be7a1e6d25e741a15ca31166d6f003332ca0c22cd3ab9de5a657c8c47ac91704a91f3008b040d4238e617a935dfbf06819283a31a63089758b88f1debef67412f5999fb550e7c4fbf7d163bbf86061ba0278d19d4b19a341548b602c23f4b272a76911671fca139e3047c81601a776333d5806f26cae414fd4427901285c0868694a0387958cc8733187ee7424e824e9f6c8300022c0f5da7dac36c6e6ddc77acc48d7d35b9d9b51bf67f9a4943e77cab8a4e4a84c287358bb32cadc93ee4eef898f3c1004ab5e0502a2021101e0bce2420db219955d10ce3a6476df0ec2e95214972ee61ce7ec16e2ab1e4313e4517027bd666b9f5c3bfd8f55b6da5f93895f85411119876f36c9a9b533ce5d1fff117fd55e0dfb029a8fe5c21667f67ad1ffac06a58909f18aa3e4a32cb49c3d9684a302868267643dc191333686a9d15b31ea49734eba5c0259bb69eef44407f07778fa5e1f61c34ce829101fa9606aef314726967db133f6e87748d6cbb08a6455156f160438ed04e362f02633c3bfeddd11260ce5e7b9a93f59fec0e004b4918504421dd94e3607e60de74e49c3d9cd7d69d9959ffc9c436e285aa319da5d874079641b4c2e055b90db9e1e9627d633adf9203088d77c654f1637a1075a4c759525167ea032648a6150571db801b99a048c13244a348298c2529e1754efd3f7ddba0a84c5b7724ab3db4f52fa22d1288081d3a3d1009a324a488e39a70c9e67e213e1fb7178ca3146bdb3f82209fb91fa174fed915753936db4c2c1fd6fcf7abfb1328f17fd7b1c902e53df52433cb49d7bc802111e6dba46277df80a7936041b87af7ae9f0cdaf6e09d3ad4e1d416a4f868bfb5383d12a59cc32cc90a8a9245eba4810080846a305a84cb5431bb3dad56efaa7d211e16b321dcc942f79b5fb69d3cf2b2bce6389d825be9b9f550c83ba66d38f12d40db4a028a1e0095fb360b034646e0901e7dda6a100d696ec77dcdddc5f47751f21d5fd940e9a33fcc8f86be34491d0da67bd7fbbd1c27d3ee768fb0b5350cde46fbcbb477a06ae4ec8e93a0bb34894a791e9c79fd95815a22f225cb1420799745af2f34f1f3d39f27d23dd4c84900b060b44cb8c0af08455b0451c3b77379087c466c04f71210d3c91cbd7ba98fd0df026f7289ed74e18dcded1786bad56715fbe28dbc190cc08d508388e245210f78e54c4ccb8fe68d269f29244d2604e62144cc8ef995b400ad8bf95c60cbc72e1b800624977e8fb39e778355bb61de82fd41a4ba0a9c311c97ede2881fc87aa3cbf147e481971278dd631033c4d3a276b6b3e6663b5a292e2d64e9a0a6b31260b92877585a13a6419851f9a27d1b42ba4f1b720655052a8f74291d3b265c3174385ce1ce3a7c42cfd909107818d8a043827b91da171a9a2d5fede9ec7bb45fbce5a4a90e44242412852270fd9cf22a116be31dc6ec02831b41561e83dde77c0c123d20fb834e32af0bbf850afd41509c1be89ebc726bdffea40d4b2e2269c041b933a9798cfc79a6f907c64e7cb323ed34fb46987990caff87c4cc9bfefc8f1690b965738663d5d3ff672ec99c05f14f86cbe1078b2ddb1ef3ab10453aa47bc6df2115e7d8ecc9bd47b5fe69145ce1b88275bad8884d15db4b92c6338699caa26c0d09f9d852003a0b680656a911065d142c0a7017a6e76b4d9d3ab544e2bcb9de15f867a60389f89538a7fc2b718578692eb44f9c344cbb46ca67549b095f6b30c2e8f421329e2c2027022c69057586a7a17d0647a4906e1dd275fef9b47906cf0c06b2d2ddd7f7c4b21889b9b23bc379a2b08402742c4cbee009050069c72cff841dcca45b9ba17afc55e67bf3889f898b9ab1a1ec67604336f656143054affd1768ec0c2f7a7bddd6fe98153692d66fb3fcd6ba77959996a8d0efaf38c52873d7fcefb07a28ad8889c3b8bd4981c81b0d042b1e213c6e00c90c274b308fa3a42f8ae7029aa13c16c02bcd211b9c4bdb700eacdc07bbf1e864fb092de2c9e45fe4f856ad4e4e68ea79bf542b335b80fd4feacc8e570cd0378b4be393bbf336f2bc495442e89d27a24cd5b0926ac3222edfe43d5a2b46e9edc859af0ba4ffe461089e6be61ed938e34f0344127c6991e73957dbbae5c33824a7b0065e561cfc89ccfa86d895ee8e7b8654fc55c381be1450c84565b72882de35bef66edde62303fba84afc723417ad5dc0f3dca0aea11eb50c88e1aed6dbd9c7403ef06585e601bb96467a69f561b55297c0432b761fdfa4a15e437f1f557b18c176760b42fcbc376e78a97af8b1948210b62aab5415096570ab88ee2a9903b0f85fa3728d19f8f70ba38ad9a1ab699b1bbd856324f9a778f9abd3588abef08db2e3446c4cac3c36f9d9502638dbd9a61fdf93841f54936f8ecb66d0ae38a312167ed394251f07414baa37aa7569c12cfb0f1d9d66ce83633ff110f929672e5aac6e1b4976d338b27601ec700f4b9e87f5e93bc004c0731a7acc5e21dbf9121d421dcc6a7d9eca7ea08ad495c05717645b86ae50c12012419ce549851960211e73bf9a73dee3d3d4b5e717560a41c4be40da7fa569c197cc434ec54adc1429f37b9192b6ee6654365c88e0fa74831bd01ff131bde873e1524d3a2330189ba93e6323195c784e062dcc854846ddd763886f955c60dca265029849fe958b2c203b7252fea941b60d40775f8e3f1bb56712f942f1849889b94e7e164adf304651f3c0818cd0f94fc4b3235dbcb53278cdb8222f2e85aebbc830c6f3dc832d141f991a63189481e2038eb29673b31505c5cb21e517d848372b6febb38d6450f09f6ecfe5bce5a8afe1ffb745f0fe5b664def786319212057d130a034c6373c9ca35b620b11b0bbc20af62ad1d8b60a3b4afa11bd0bcd2495509eb9bf40b9005db19d1b70bce1d89fbe41704b80b4653b8fba21c1245e7a1225fa6e82eadea8295db890e86cd86267efb1ada00e026107d3535d0ae1e9f67ac8945e28214472d15234e1cd52fc30343174651394b8c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hcddaaf244b4547bf0151c17d4b5661c097bce0b1a3fd5d150e11c60051716b90e7be8eeeb1f0e5c35f605a133edbdce7f79427cba1f03a90bf2b353d57a2352050aa77726100167f4ea85a8df343becae25f0994d6e0e1f7c5ace6d78590758fc26c520e634e1af489eab999eed3dfb6a86ae0daf20836c104d8b34dc7887f456d497587e19b99dcc2f06f3dfe990345c9b46941069a2718203b748d294f8b17991b6879809adf3698c8cb3b559761719139d9a6735d1d05caaba4b0e291b44bf72c5e056134600f6ad91d39be8a8ad48a7b039f9b2b4f3f9b15632773f62134757aca1ffa7965a3cff41ce50654e55f3d9c4c74fd4fe946121cb6500f58db66dcdc91380912f605efbd6f591b23a8e0ee843f4e11c6e391a031e26ef3293c7ba68be8d480666489859bf02fe54b9c9a12917ccb5153cbc9d0778248443fd5a9e823f4d05bbed467a1e47d4e1ef6c071e7e2870c354548b8e260c7c4e9de4227dbe8ec4dc6117b86cceca4ae9e0a8a9940d40a4872fe5f69e9632c3fbce9178fb6c8ef3e812ba47f7f70f9b67edd4f5b917c113f44ed7be6cff19f91a07f113d736e7d8021b54aaaf9b872f213653a94615bd372ff1649a60f2cdae5c85f095bea4d8468ae03bafc0a5c1c3aa1191177b2f4d25c9c7ae73e0e54da3df61e5ef176271d5a9a28e1fc62aa15a3cabf840badf236896f3d81be3ffe4ff292cbfa6f3fb3bcef756b1e816e02cc90884956f6ed691613a96cd56a49948dc99c18f800ec40dd75a07aa53d481890733493a4a353934d6f5bd76e5fddba1b240c3d73af24b3443b82d7c0c6319c315606c3e00c0982159837b09b96d54c6894ad052a4d89c99baacfae859f46436cf8c9fc280fd7ef2e4e53a570d6606250122f53867f1213f820cb0d729490976670fcaf410b9c9687c860b56434b7d883038d45aa7726075097f333ddad3ee87aa5ea2283c9579a4d90fa8fa06a0c33ff979506b61420295c82cd07e89a4dbf707130983ba6255b7c1932786b513caf8427f60d334af8c708a0ae6e5e2d36db35673f52f242908248674303546a69e28de53348dc58365a2f2a3e4f98ff207806fb20c735dc284ddbea2e171fc7cd374910a7ec6623e9d162d454e222995dbec7015b55822d568ce42d686b63b469f4d80a034cb721a42f2dd88cb51bb706fab77f0bea511460d5d1809654ead2352009e32cfb64c5e0b983308f0c6208d487166942fbcde79f8ccd3ac15ffb84c1b11299d81cbc9259d076d13b8b4c3f47ba414b06064c0ed14ba5c9ddee713b3c4f0e827dfcb81b38f8e5894025e92e3ca48f3c86525d4293b837997a7ed9efcbbc190c65905f8c42d8ce2323751fc982803d5997931e3aa0a9e3303063768438380ed92fd38ced2b9e7f89c26aca48634b36abacc7dc54b7f2817b554a356073bd4fdf2042181a17a559315303cbd2a401f47bb5230c9cc1826476fdc4c5452793ca89b32178b197e029d23c40d8b9a9b389198e2c5e908b339e403a862ead5de5b65c17b2de797efc80daadf322371bc9339624e88d887fa319e689f8d46a99b9f91837eae5ef48d5e1c68b5d2f675ac2213c6417495fdaeef1e82a050b270dbe34d5aff70864c9971c28afbf10be91835f0618fcf33c21778958960efe24827bb1a039a7c4756c1afad918885a7b5ec6372a64a4a63f297f17d9d4fe9c9780e26f4fe6ae397970d9f52f563fb2da5db6e7ef09402044c729ca327b750637bc58d3697e5f1266b719fc9b90be126ad12373fb72bc9fc7ce488edd1d34512d91697be2cc76370e6deaa4d8ec6c75d1a917914ad7dd69c7052c7d0e1ce04d0617d6a7d95966bc2bf8a930c170f366984857b005e4c41127d138d6024632daec9711b3a7183dd29cc52580bdd69d2fa0204068321b130b1ed0b11b097e9ab92cf89842810609325d01d4e494ceb92d2724778999dbb6bbeaad708ba39fde6f6be70e1014ad34a902e6afc090307947becca135fb6440b9c6a5d0f41e7c07c0f47e170f1d3d5421faecc4abc5b7a04e84f33cb8304954aee0ac6427853c5b5bf4c3afa3546cb8bf0b8fc0ab4ee40b975679d3991b24632b81577270611bebca2ba2a65a5ce3e5481ec53a1bd198e2aa65cdec00b0a70cb9e93b27e1f218c4dab67c458c6186af260ce7c75a9539d736f5bcf06ca2034c0a44579ac9096e0f3d9dda4a13dc18ff84c2c55efb5765a625f35c2f1b657becd17b0f2ca5ddd6452090c6b7d0feb5261f17aef7b03dbb4e8054459688467c3132695d03170809147933a5e2ad3aa382083c13617f0450312f5273e8cae5e95a2177a7183d88da45c7ca3f0d5243d96fa58edf2580704b1e7c7bd1acefe1ca2c6f0f220676bc7bc5e5f348bb28f0ff56830fbc604a52666649d357b8756b1c746d6253c3e167dea95e181a55e75442116f2f4f2481ffd1bd518ea506c762694c6b6cb3bb0d711922376da67a5575bf629af92b087efc04fe62b2d72f63ebf33d8706471b620026201c741a197363177c9912e385b0cd1d2fffae253bd85ffedb28d0dd30c07c391beb900d91be51f1c5289b8b89400560f0d2550ab2b095bd6c395ffc5f1657245512cc2f4335e764298ffb27f6c0ead24764966105b040c00f2288c2f39138be69ddbdfe4bde14f8497de30e49084f4078babe49ff8956f5d8a51e593faeaa5d85d3fc5056b086ecf9297f7346c7b39692ae23b85c2b1ab11839ead046f0c2d34a8205bc7f862a72f8ecd37c9c37336f47aae80b29932cbf253b543262c4fdbdd1dfa0365bd87e341a8963e3aca61dded1b91a6d33bd99fd282a10413e7533156ab77b0d38f9a940069a57aa6e036316fb71d34a36b062f7a01a6ceed2618473f74bccf173cbcc2a230473ff6cf39e0a5f44e49d4cf9fe20adea491f07b9c46b1ab6c203086bc5b77ce8d608bc62b9334e59b7b6cf73725eb27351730f3e4a2d2c4775ab2786dfee072cd1a437547616c2aa42739c6d73cba2634e1c19e91e2c95df14778f8b0f4cf2648d60b21b85f1114d356177f7dc9a8756ab22367148aa8b07b509aac23f9c2fe7427429cc8c966bdf1f768a11a338d9fa7b17ec553897176f08ffebd158a43ad1cdbfce6b5db396e96f0e15dd2cc16d47d19dc6416359f87245b1e21ee17cffe21dab3d256c8b58744c57f74c4bf3e7b8ad4c1089e17d3ec20e862189dacee3df2d28db8d73c5a5c1d6ba13ab20470f802e0771829a6853f3041d2ea6c691118a1728ec8b2b8c081fc49eb82e6b6dacc2eb6802bd3e21cfd362f006243dbc3d4c635e46c627351ca200c24fd8410835507aafb73c421f4c8c65946052087b3046829ed03b787317a54f10193e3932c6dab98294820b65c1cdb3aa0178d369233b3f4fc2a3c07e4d75c174aca2b6cf3c5c974ffe1e77e66494044bdbd2dd6333ad0b39a22f197cfad6219d792cf7d3dadb95ee86d7595b978e8e02f171f17374d603525c3395b933b4dbd4acf9380f202eaa4478a25482b113ade18af18b0392994d3a2e957256f7f26f1512604cddfec90be764bff18dce7935e0f4fd1d62ecbf06322a1288cb547f3138bd4dca571e6eca8ac943c19b2a5e8d5647bd61f8200d8568d7317fc5df0e931f2b4b50ac943e0296baa5ff844172dfbb9449c12e03d0e1494def9285f1075f2deb571e450f6ed75780a3d662f9487f141ffabf54f7692cb31b6f9ef0dd465d4588076dbc0983bb4c33b537bc6e305c6518ec2431b929b47c5e002f86fe592760d66044e649effa2dd5051b9a35c92f474f694489f194058c56970cf44aa6b67916ea45dc33b5a51408509c2dd2c951ba5f980eecb6cd087bd22f3baf2fafa4a7629c2b645f31105d9dbfd7b5b2df73df62c1e690ebe9b04faeb9e2bce3a09b8dc64fdc0a268ffd1685d14d230efca655f07f281f2a9b8b6430b9a13b7a9e1cedfdd58059c2de8b1b70ebd41637449e0ac1296a2d58795ca8f94bcdb84d8f3b5c1930f2462c95927afd87d7add643d5411c0c8143819b4dc1ec74f2abc6bb89a435ef4b045e574a8c1dabefb3c2b4aa6644c777313389b531c8ef00c115386c816705d985d46ec377fee793e4cddd20e5033da56b98417c45f55bea35ea99100bd778a94b4a1ebcfce1a3975aef39e94297af6abc0de8c023ddad45382fddc4fbe34446e916f92a9f1f4c566ef857efc65667e39c37eca56608df1176cbe40aad1285307a879b54b81aa292946578d1a9cb90efacd13e0cb6e3a15b07da713cc263e3f24668f4560703fcd88eba793dee94f5d630df0a841df33f835841a83ef4f3125faa3d7b523d0fffea517d0a637677b903668a4cbecd41f2cc2bdf09b637a081e8929312087316679de443002471c7596d375fcfa19d2b3d46bb1665894c9462b7356144ee81e996dfef4450c5cad31fde5c5948f14890f0c6b66d4d1e7d23a0068b051573b288ba835923d917aa6a0b98e976e6e3160f1bfff5c384dee39ff951ed54c7844878d18c7341c37a0cd506ca842bd8c3999b82c11e1a5f56f9c79bf5bd74977b3ee4a49fccf8628959c9755fe25ed3f7fc9004d49a733f092e3a3ab1c94a3c65e5182ff215195685e5882fe3c833976f7fc47f40a33ac3921fc9d90648c06bf79175addf92b7801108e7e611df036a6d0411b76875a4d5c2f01f0c664058ce4fa5f366cdbaf5f3915a54f4b669497a188c2bf3927f02931b95d4fa7f64fd130408a2eec9eedad7fa660631b600da5298c775bfd492dd9a4dd5e9dc83216397e2c69dae4a899ae5d4830e174afe07f014fcdf3d6c2f12f1b0ebe6021f853eb9be22cf01eef08430c230e39c1012cfccd5a3c008accc08af08dbe2d2bb8d65aa557e2183554471654620c3bc63ada5a9d49569d87a155e6379c7bddd5f341f77d1045341049f7380b37c4c17733f4cb4ccf28f68debf4a790983607534c086ecbef6cef881d03ad5734f5dd9caecddbaccb75a5b54094d1e99b8de3de6a7f8f91bb806c9d32fd8bfdfdb9ba659431812a862eb8c31ba04a8c358fa574a49196987ed7fbcab0d3534c9c291e937ec779463b9db268a7c83d02b8fb36dd47e535fa537655a01d16bf96c12a66bdc202d53e59c4a08937f718434ed44ddd628d731e484b2ba781e3ead9c5af4bf473fbf3c30e3256261e7929633875a7ecd850ea1da4122b439c4d680928efe3097444739550c3a2e2fc9d7a9ad06a144bbe1f2ffd07ba2875d86b1e1a63346ac5d68fe335254804eba624701e48ae7b3c8586fc708ed4cce54962e5684be719b7cbc68dd26a94435d033871a3b3af031479e4fbc0d9c3dcac3c41aa1eede1d56310c1f9c4b892ff4cbad730ad82f1ffce3276b82d68448acb32141068eb6fbfc1b21cf78a2087c89f2c58516b69bd218eae3d46c29dc99fda033a8970bf9e6e620b55785067959fd13e10ba105daaa96a9f6b50acd2e2c03945333147d8968d63e16398404a6ec3a36508f3499c2ad802d3d3dd904;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h8a58a4f67feec5bbcb87958684614fd85c4d1fc73a824cd727ee6fca648563e629a05586c5bfc9e27fa182f033705335530d2751dc0863cbd36b6a8377ba643ee647a15e80e796a0d59f1e4ae06336659da7a3fe01a10ba681f0fa4eb9cf11943fadfeb8ff17d81f16e2c6b7e17c3d648f4abd5b5f916b67b3f14fae97d2ddb45505591cb585d3b93784c8dd468e9546c5b0b167c4215b4cfb2ace27470f0e3e21a851b64a119ee5217e4ce301861515ac8da544ef2d26ad22bd3098f4ee3ec9d51cbe35b8ed913befc642872aab4a5ac23bb7fe6f80bf6881497420b438ca147c57e62f354f52d98190535c0e3c983ad7b9a8e67d174eb8fee684835e268aa95009507929e5cabc1a5c2600f5229f01938a18a5bd9f0879a2093eb148926ce735b18b702a5461f59de7199372f0dca400da23e4bfce98ec28306f1e4dfb2d0ca02baf5f4aa73e99a2501d9200b2aada20912b073aacaa6adea0a8f584248041c3ad5b0e74efc81048c75e28db374dfdef6901f846b94425a478e05bf6b543ba1a6ee2ab3e5fed22461cddf85ef2de4aadf6dd91722ec8f6e5127a0577938aacb0069460eeb31a2ec0be058ef689cbceae1ae690b7c69894554dfa1246330d86d3482c1bb5716533265a470b70aa8e04a8c7fbcacb3bbd47c7b3c86a683b61ae5aa5992e99733f1d2c781f5e127a54de4eaf59b060d9756f30564c6b2f2ffaf6fd06fe69319788b87cad09bca6ac053fe47f324d3753d975a0930facb1824e25339eb8ea5aeb1e2315164affd0405866c6f262feb44b9fb48ea468fe393594cec0230e4bcc1106e5e031b4dee655713f205a1ff9cf4ce938eeefa91bb9e838d310228a14a545230e8c29b6853ad0b5f98efcb83599b96afeb87ac5cc482a50a66e0a2ebd72605b5a4281ff237e63ef45be73f880fce222f6ffa1af588eaebf691683d77a607ba25fbdeb6a691cfb5294089e67947b528b16714cbd6e7348e5eed882ab23b2c7350ae2f5cbe2ae4bbcdfc8c22644953dc8f2dae98f4d7426afa21fa2175e62d27a873fea64d8e6ba65bca8aa3a5eaa01d1e489e36938bae90e51b34cec3e22b25ae749d5ab3e29e33c8995709dfa8a4c1c5bba17fdc75d03f551ea80c475c3176b01ed62dab1a4ed2c865156f9b1bc9d6f64aa04d19cb0a29b829fe61f5e34b012d1457cb3f162a195fe3b9d7060e5ac26694ffb476111f70bd23b751c8847fd6cb770d62427406f2d2efe312d43471a0808410fd5f231049a12f9815a3dd680014ab9d5a3a1509ed5e30a9d46185d3d617e8bffcde25b02847d7b1c2c43c0946d109f05f3d4ed16a81226302af95c44e4ed87a8675551bbe6dda89204023b09f3e653a073281df0e84f21b3605f4ae2f8d0c51d0822b03e17ce1f785a37ef629c5ff2b9d82fd38b340dda388a393c66b21704139d1c099642b1a0426a030fd1cf68f1c5c73d9dbea77a9fe1e934e7fd6e877666a1e061de686dd121bdd341fb9caacd08993704a1c85f4823c83947be7bc90d6f41f9389959e9048c6e3a45d45665085c095c671fa9b218c2599e6250265f65edb37608ff8471e3759a63d8ffd773b87316c6d6784b92327439fb0a6e78ae890c483df6d3cdd30307228a2833028167238493623c9a6a5e0d6a2a223345d287695d9fe5362706c05832ce0b7f4f722be11b3f98921966eb7f30f768dfdaf00612375a6e5d55089fc9ef4aa59fab11dc7d800ecb385d19bab27853aeb9a35ec8c06c0c5c45aa851ceb0a5478c7b2f0e8bcac8f7f4e95784fa95928f39e93a8bc3284be0427d331851166c3e80bc54b9a371edbf9f39e225e4ffcf0957105a6cefe894e16252fde8168f230aa44d0bc8dd4c2159bd73f211bd7a0cb5c8f68cb75422ef4bc75794138972fd1a4cc8ee46745988ee6ef5587fedaa668e36eaa146b08d5ac6dfce742a800387699984ecc77bb9031169fc822c2974678f9dd1ed6476f65feb45c04128059a50bb4b83e0de48dc3357acde326959e8410b1e2aa3995fd2670868ad09fdad17a8de1ce53c05be8373b2c7cd85709ae2ceed03cd2946680d469f7a6ee4b95848df4d249467911079d04a3f680bf188897b6e17d515909c2b73686de204b177252f8bc9479d68401e07f8856435767787b34e7a881ade3db517961cdb281ae9dea03bfafc6a6ff64bf6ecccb618a2812dda614a4712e79c7ba7dc898dd76b1eeb96b75d44aee91aa351adea747745361f49ce15e17c5b5a02bf92551c9943589c7fe45768c01ef96debf4c3dc34b9bc089bae8fd58f9b2ab0a82b546586a79e60d25c54f8e7b41343f36ab62c8335c1d4cd5b529cc1cc96403953e95852ec1394ef1d07f529ea4fbf8e3d094eb197f2b0f59fa9d8e76c2fb93150b8a95ecf03c770bfb5812012cd7784dd15c90408d5e7ebedd4e3a73897c953a84933f83e98a0c9a7ce2f273ceebc5fb9f9d88988bd2028d0459d51f7ea6db940dee6d0c052ea24a00e04e981d96bf1cd36a48c31e7b23f11f2afd8c7d768af38a8eb44ad491b3255ea3b8b22199ac711a65baa539a26b288350aa0e4e0bcc748a2c3a3f9d3a764cef24158a4a0fea7f6a4037de82fca44f444dcfec871670ea292b2b6d2541435ee63240d8a4350012157f059c2031923e8de8c5501076c56f61656afd4d86052cd8a1cd7d6b6de72851c0775c6fdc2aa60d7e47efcc03d665460932f3a1d20913fcdba788c96c9d5cadf009af2870a4d7cf1afd4d6267a5d5c951ea4847e211ec604974407c3242d9f51631dad3e005497274fbbaacf130fc599adc82b5eddd54bf114e27cdcce88c3b029dace07956441e0a717c2f7448f9cabd3705bf85d6d2b13066c4a658ea207b86dc4f8e599f78b74b52b6f3b5019ac74c8b70e5e6824408bf2009df2e17b60b10ec6507d5cdcbc3de994e8d5274c7b287bbc1e74ed932bdd2939d19859d294298a71c44c11d9d15890d1423d9c7c5317d471ea3b0a02ef50559ebb154c4446046a8f6105b5a539b093097a152f244e0bd178bb085265ba9fd639a936ce8c1af3fd2cc9723301e00d49209d435127a13f133c8e9c99b660e88f7187c9c2574755efa5a02686f5bb17a2982293fc8477ea49de7518f1c37e3ebe4eeb4ecff8a5d0a08eb72e38c4d4ca01703ba576c27660f3a7e276fcc39e313a30f72e3f3e64036195038fca0b7562fcbbcb43eb44b2729070bfd452400f0a897b20c784d2b9a74aeeadd4de2e7832da9eb8483f7c875a6499e1dc22f7d3a64201587302eb7e7d1343d7c9650cc1726c8f0195339b48c00d4fc15e69897b505c0c76a25c2ab8d131958900fd2589bf6d6e2b1b5cf53354b662514c21686bb4186b58371d9a1c793d422069b63895df8767a03e7f35ce0cc7a302acd5100cb5666d022a82185f84d7c06fd924e5ff1297d1c7e084b2174601a0fbf886c7f8440eab5504bd7f4bcd78111291eb0f2d43204642ae4b3978f629fb2853511a1e78517324dfc12eeed3f6dd2c28ad8337b3489490e7d872bf1d813bff4ca185e16c0960fb90617695d13ca963cde9d50d03321961880ea9703b5a09f36a421cba4be14e756e27514611a5896d62dc84690299b7156603939025617ec99145202f97b7d55d623202acd151f68edd357a849d0d81eafffff338ed61bde112538802f4b1542181d9741f5c63bd8aa65a4aa35dcfbf849621cc134d8beb5c00f23b9b3e348f1155b8ffc9e3d562c0b18fd6b001a4174c190b0e65add1c60b620d1a9020da42541230ef7fac24672a71b552b18745b5357f83d8cb213ba188c7148403513d8acb631817612c63c4c3fec319724b03ac2ed24275b72fe43c069ad44a057708e47178fadf4a5c97b3e8f1276a81b1952a83e94f4530886768f51e90623f376ae4fd18f80fae34474c99fa8ae66a955647a6165a5c36c8e508c013a8a5f348958f99204681e9e41571958f8ca70963b8bc7ea68a8ceb2a21cbf5a84a83f47b598806bcf39e6626f1674eed62079b355b07fabffcebd79a996774ef2267d5666e2a7120927865744bcf6bd5c034f899e46fe3b8043e34160f20585d5834b0d6fdbd05d1d115a413d92b801fdfc420c267a436bb6de3cf6a42cd0ac819c58f7190347eccf78a33c36108a8dc078c02d00086c308e841b7eba87c50620f0f9b33fc6ea0110fa454cb7e933d2ed74c487ec48b0e64c4d7e9b36a0c97717396f94194ed74729db13577faa71ef71abd555006afa58caabe5b0990f4f8828c3df4c7a832040bf370abdb253a1afeee1d8423033fa34940aacd7303a4601b254546e028bd1ce6f4b64ac4ea941310c8ba44ae6d940b3c18a6fb8c8e023c830e8f544ad0a028ce053f3b0de9311bb401ddcee31602aa99557c93174ebf2253d8a36b26abf8bc2e2342f65a96089c45d1b7f09741ce2a94335e7cf74ffd32c522846f5ace970392b957a5a0d4d085907ddfdf2967a615de8dd0df50c995e32a439a3909af0248adf5c53378ed71681ecc4463c37f55d020d39dd69b843e0c5bb2d0d8ccd1980e1d6d8acbca62636e603a542b2c67a8e3c21e4a8398a504ae66e2b59ba702967147167b3361620685d5c2473b13b555ea507f9acfb2450ead889080003ce89c76f6b6b6ed13ba00d047f411519cc8b4a3d92a7a586ea563efdadf9a360f188ae28a8d4897769385c3c94d9d2309a728af6bbb66b715888f58857be8f3cfcc1f052806df717e6d41916f3febae05fd47a4802cc3e7be1e9f268396853735eab6cdecd7d044fce5aac9bdd526916f6fb6a3cfd48a4174954912fed61bc71a77b66a56c27bef5b80ef9c6e8ccdcc31e8b68e94d4cc2f3e2c9edb8f6bfa4f129a08ddebaa84d34745bb90a6983ffd679425bb9f652b752994b7f17e1ba46f738b709731fe2561a99439b5c6d4e51b72999aa9e56fae2a394146ffc2bc027b82fdfe85c9c3520ce35ce80cbe1e32a12c6affd8cb4cc19f9443f50a5e03e57e3bf73f380ede01bdf83a9d2d7d190bed2c13fe690623407efcc52e8d193afae5faedfce6984ef9dba453da9937b99cc28ebeeab694851a0a51e433f699361e3b448e778e1d06c44b709fad95ee36048a4ac8ab398e1365a1031b73fdced4d6cf78d6b0dadb335086cb545a7ff5db5c7ac2ae33b47f5ab4872756f49d05b8ef1158c8e26639bc08bf50ec2c2000160ff96cc6ff8b946c4c516006ed6993ca44f480010e3a56738bb56987ef57da96df2fb6eeab2fe9e9b292507416db24f2774a0d92a3f652331c6e6b0109bf3c0d076d55520754c6c7a073bf66c34a69cab9a1288959a1168e4f1ed2151367cc3bb14f99beb6517893e342c46a3160d6cc9d986a0d03d0c5df62906cd19fa6a658257f58e91a99156548a9713fdc3d232393cef533ac3def580e350803f3462ff66ab48bacae3260f7987765906d75fbeded05e6ba259167cf4fdeb3d8ff1f2fed611de916f5b7775714c369edbb63b816edc46510079f41381cd6e5c75c3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'he81b0ce666a1074a978b9c7b943c6e46eef4da958c6da4317339c2eca230551a7b6442e59d0716813501a078de45ba822f6ec19613a0c122980181762e15cb0778a6866475bc0b21c39f337ce6578db2796aa26c7856cfa4a3b108fba8696c16d361ec16bd1544002750860865a0f0811be1126239424aaaecb5bb3e7d0e6e8636dafdd4ff3978aec406075427c9d1c8f432a2b5af57aab87e716a8860aa40548996734ed0f9f53d0ae0ea25a32cf68c6f5e98a7da20faa3f54be5862fd8ae8a89813e82a5aaed9c8a31badbb476323909664137be661922888bf91e0a1395cb6660e3d1608a44676f0b4f619e78a6f3084b45be0d089350898c24597d9e6ec657a4e3dcd2401dc54306b2c70d944b85b24686160a34d849f25f3e5b069f23f1b6724e5b493c302ab775a5300af8e0c3d459f974eb09f349dbab2409453202d3421efb356627239769581cf9403b88d5328733d3245e8f07aaa3824d2260f8327e03a3036b68ec5162967004939f68a0ed2b3b233b37a65d05dba9737efe3ef87905a9d7877ee1a536a6ea0c347a8c862d129c8100e51553549122b4d9f264c03c99f8abaa17f149c4ffd830cff6f28e773187b857c32b5c74de12d6b4c291e1d28a7f4c5ce174b904e35dbc2893ccd3a59de5c1da95485ca9ca505f1cf2e6cc92c35bf815b9ef14a254aa0f05cfd327ac76b8246a103b51237c49749a613c2c5f9844bd3abf1869a95a6377f2a7de99d620dad965130df091910f688972ad8af14fb721dd025ae0a95fcf75293fd2783e7c7d59d37658673c41b938c1a129c12c0c38377a769fd93447261b8afd16b180625a995a60a5a8b0fc87ee6486ad709fdc4fcae32dd2ff0178f57334963d8a19fc1426d35b84f225b0415f0fb3d9d4833cfdcc8b00dcb29d985f0507c3f763092df7fc39a2fd0ba31c1e030b5af98bb3a4e4de6139c934a7d27d2e0b16b2b797900eb6a5141fc488cf82ce22c25700d9c47918ec898132f064436f70f0168cfd0395d716a6812ba43b07cf6415984ec2a90b0689242b218a0153632f0edecd8644e06a8f4ae810d939d5852b433b6cd16501e4538a3c2de945a4e09b604a5f84a0626f774a6e332d64b76bd64f7e8b4478d3080a495c530f9fdcba143d4fe23015ee7b8955b34fc10f181898982906030ab3b530773a101e0610172d974ecb4b70a422dc2b68124f3313a40b49846604b96b1f3dca73d2503aefbeb53b08c230ddd345932fcbcb9073f00765545f16908cddbf3de5dbbce64c8ca6dca2b40e3faabc04f72268357c6635aeaceadbe79097a21886bde5be25c56fcb1da105514abb63dbb261b050372df97ab405b77a0c4ddfe6f02eebdc0959e53e5466f7f68707531e1eb9f3ac6f7c23e703ef40068dce9be1015fb33224bbb8098ed543afdb695bb4f9d3c11ff3d63881b09ab419d70b10fc350fd99afb0d5253a2390c622cb0bef5102c8eb6b762d6669ff1ef6bfc794876ad9e099f2c4662d533b151ee1d1cc6d3490dbaa4c6e224b386993ffa4977e7e5e7fb2e093cea40706d50a09a4962678eeb65fcb144e1763c739f764a4c30ab2f685ce49f0651f894736f087b1f26309f706026ce02e2020660b59e8d8713ff6e046dd7ddbbf92519ff5c003127791b31a9707fe03df8e32c77ede802a71288b8ac2e799be47dd693933cc50ecb9647cb8a9a7496af037ad1bd0cf730b8d9514de9f26c9629c77d073f7482cfa20ad94adbec3055bc0449d1e0deda192ec35390a3f2a997738c795576b72486213fdffb8ef1f381f5707016bfcdf36bec8824bdc9a36adbf78ecdd154ef59ff0e7aae9b20318b206038af609e883118b812dc52cc6941194b82fbc876deadbfbcd5c8c064149f6130655157dd346e4cfa56e6b2687778d20ada3174c3629f0f168e7d3534d231dcd02f157945acc039c97ac51ebb9581c02906ff7f1e3f116b7fd96e20ca56bfdf95988ef7ef6b538ad85cfe35b19d4fd5fcec65427a76e023d4555394780a4f91ced338682bb015433c3fccf464addbfd93201e2db57be78bd9dc8845f05327e9235eccfae01cfad1728841bdb01d9937e2eca0f2b9b03f12c6b07cc296fc33e42a66a1b31629433b0de15668c05bd1594c2ce07b66e7061079941442fcad984ace2fd3598d00793daa08cd88db1f2de210d23fda0c9b8fd88adc0043e900ad2b840d0540a2398222bae8ef05b3c7ced611ab73c01bb9d0a6220c10554aac3dcafc584b2ffb79fb30a9c019a15d40cf4f9b9c5dabae0ef1c52a9637cd087fe66b8f2500345e785c5717ef8118666526a6decfac3c37c45d1a66883ce87953763dc5728cda2f4ecf95b98a3fa4432cd5a0d8762e8852b2e4e64686c29952a12a0538511af5fd82f3f948423bf5d19ee5b90e4066ff7890cbc1ffc96a6681d47fbefc42cd63ddcbdc38f4d554b16b771f2cfa4155d1aea0b07df256d43adf2225c394f6e6b31f165b08954a031c35864996eea6f06d4d331f252503afb3c41b8a9ee391f7d88294ba24e386100aa423039882b099b284ecd781f5690da066d3c7b7893408c4a56e3be64216c88cf35bfb9094fa8a847c19e96bc4d7c0290910947da8a600ebeb9b89bdf4c6dbc377c412165b8e8fae6b57092d4f9d88a8cfdee023e76eed3873273bb89bdd50bc68af6aa2991cc58b7408c966d83ed0aa9bec2341a724e34c2cc3ab89d86739b8af0694eb589a7d00a8272fe90e4f864e64385648c20a7734a32e404f36cbed9fb2f2e21974ade2aede3af725b345bb0d6f1241e1c94d5d2101253e06c5e53a6e88f7eeca3b8a722864cae8bc05a56e33d4c8418f134da6c3ff7ab8904096ecc80e453ca98b8b2ab2941d2a6972fada7e97275df84b49189d5832e8f5cf04f9f3d6cf44b553bccdb93ef7460f489f586ed940d7686a02dd8402568ab7a31192cd7aee7c81e172f8e555ffe78467057dc6b34a5d50941988a26aaf827d37b7f9ecc1e08c92436cdb1c32fad81cc93e7029b47c49aee8ff0f81db826a9f182168ab4d08ae49882c2980d17fa6e565da81513004e328e70d5d8ca2da99c0b8527cca4c02ce22fc2c90ad415bc539c5a9f763b3237f6ea8c11ad8a338cec5941668b08acfdfaa0f040e45a1c71fe74c08b2a487e9fc6b6ca6bb38ef3dc99827fa370cd0bface6540bb40ed33ec4694c77aea404d09768aded5be68d1ced667cb9014d139b7854d11dbf244daadf7457b359b84c06cf51b3774afed0b1580acc44ae9c360b286adc26227920f9bf269818179da062164245652655082e7bd236a425d0b6607033ba6b197a9d5ebb69052fb429ff4d2d36524fe462c070c00be820691ddbbe2f655674dd0e71d4bdbce22ce28c3bf2513e051be45fc5361dba6cf0cb547c43ed1a75f909eba3797d8946b19ebecb0b8eb6fcc24b5138af346cb4fee67ebba25d5456cc84a205ffc9ebe5d97961cdedbd190107fdd474d85ef44dbf83f37af66310880376dc7cf2d1dd1889b3bf4b9e9bbe3cfbdb0c3b05a7cc9f2f75d34627a9c01b2d5ca538fc5cd5f826af27102de0ff3e4172db1cf959a6ab1ff9be5ef0845c8fa2722d2c33fa73efe3d1146faedba923f2ada926153dd24c75a8ad8ca5d51b5c3af7234756c0d1069270e2d068036ce0b81e6be9499bfa8b85e6a425a4db860eb2a285f9d4652c954545caead93ab05982fdca518d37feb6eff1c9fe7dae4fca8196bbe52bde847af973b47ac659e8e4f6e0c83531df0dbd183de92b84f0944381ce78483063479c1c472142504ec10b17e4a9628b7efa630639929b85428cf8b98dfc5be765ed8c02c5a204cafa5a5fc9637f81f7942eb6ba680951855a98105033a15de19de15b2e33bb489f4bdf164bd00df6c49e04165cc862092034ae85ffda9ab75ce92b08704d6c0faefbd202df4182c78f37ef5469131ec0e0b7917a9b107eaf7e92fdd795a805af8d49e25ef5d47c325702c6ca4977bf2b1fe8d6aa855d36b15cad7d246f857bd66b8f959d8115d9dd219418d2e7aed429e3e3c18af5ca351daeac1bdb85d3ffc3936309cac602c9ce50f423db557438aa86ea32d305c83e2eabf254d620a0e33ad1f500d836b236314a8258f18b9e82276c3c8c8818c0ee33cb7b18df81f1779738d59219e78b5f619e0a874c0cb62deb0e929a5d6abac23d81a71a86f468dc93a7867814e2e6a45bc46da902cd9f6a9610ea24194eb458dd204b08477bb1b1cec98d12c286f83be19e61bea6d169a8dfa2b40d10225cc322a870c4ef743dd103170971ede4810c850de21e56af208f8b44e7fda22f692d2e061833571c570c94f43b8c0bdbe1b78cb14eab5287a6741825ce3956d4686f11552fa7a4c0a66381502f68bbd001b6a35257fcfd916cc3e601b60b2c1831efaba89aa2400bf7cc6bbbcdd15e5665ab2025b16158ff2db2efbe8e6d71dd69d78d156560f41fe3ac3b21c40ebb35442382e0e7c7efc063bbe942f6a78bf002799c1c21ed35ac574af16c2f9f96d494cc14a8e7e623677e2966252d8d14169e9f442eea25cb52d3975b15ac2a29f4ff740adf74ab5e6e6ddf9b4dfcd41e633d9b529c26dd5381a06973f992ad0571999c818ebb9e1b4ce1af735227ffd850a4d81f4fc26fc2b7e7379f6b7790521fd87a62b127592dd0cc5f74958e8820d1e3895bbc34878c6f48a63b3d9c8806a14bf8be81bff77af262eb2e277a2153d738b56b2f7d2c0e57c02a7ba08cd6e08ad243b3cbdbd0cd4154f6a14e808263257d28ec04c3e7c1c9d4a47fbc8a6b3d6128638fd61fb97ea36cd683bba71000641bd55acce4870a8a8ad81d38ce3e0fb65ea2ef7c8bfe742cfe1147ae907fe8a0105fc94f9c8ebdd782939d46e0ee5f1423a982ad37b1902e25bad836e7f4dc385316931a251be4b2972ca291eb54d607c2e33aba25c3e92132dbc9a02141dd4d796d4a83da8fb4b065ab2e8f279e28fd758c392695744c80b1a97affe80048afed0d67e57a43840907b0d82da4af696905ec5c865835866408431248025049d80617a4c98d8451e1a398ef3770b4120453ad7fdb4689d6f78ef46de61f162624e035144d78a24a06660a0de3e8925423cae1eff39c660d8758e2ee9aebd763612d942df7b3230a4e60c9ffc103931004496c4d3646efa42f1b94c12add667b786e095b836e7a31c08188aed23c77b0bd653d7b18bac88ee05d969c9272aac7292b13adec6b1917abf0885b6db62d2427fd72bbab2058b527efc32be46ef6f0cc8678dce75fd6ec666282792091edf515cf0f9cc04b17921c5e1f0a786f321730df85e3ac376fed723e08ea1e1144bdecf3863e400963671f9e32e49c8d1cca9381effd6dc054eb97bed797cb218eb04620ecdebf7cae9303a28a09893182e47c80acf471d7ca7c089f3d6ac4f1ac41640a50549726b55f17db29d53fe4f2cde2a47e8c641ee518cf2b36d73c4e4fd60553719c296824bc4a7b62c52e09166bc5dbeda294e3c4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h3cd329948b9bca609b51f9fdf0df2b0dac4e5912d1d7ed2b88fac6d8e2bd7f2f595fb4756d30e4dc96cecd4067a59f9da31f03d5a9e6ab2e178ddefedab0d90ed5de82a1f84b69c352e7854e11eecda44b767c5c17508a65ad8f1bbd8616a5ffbd4511c6a75bcef8640831d61909e493cbab22c3455eb07cf8ff3c9075fad4dbfc13c94f99813d872967036d4d38eedb62b293a8a52ab36098adce9ec82f755ce37bacc0e3cca78c13adf5d2bad7749a8497d06413e19fd4d5d6eaa9044c81d401ff6356c04f412936b5fad1b82cf5a7299a1cf9032ab37b0de3708d263c49fbbad7779bf528ff3cbb72e0c515064e64f91eb32444c638c812847d5174aecd6bd6a6d91bd8fa52eaa77c0f81bef5ab1764160b3a5d68bf5c9747c3346d65cf45171a0d6097abb71fb34288b913ff9ca857966cb3bf832d4e9e4688c339eb92d17941677801dffa573fed7588451456193a5ee78941a54e91121c441ef72a84cf2960c90c91c8b62bfa3ccf179121a4d5400d14b5f82966ff14bb8e2b83d36ed27d8914b022e6cd82d8b4dcbae13b36984269ce964d630702cc8e769c498e42c0ac561d44f5e9abdfc9e7a0154c22844c720db1577de93ac15f5120709cd85a827094f7c9e7adbee6d97066a2ffea9be0e381ba55bcabf6bb514b56dc834e217d3d0f7576b58b7bdf15ed446a6c9d91b4fa7e38763bfa733e47faa39454d707497c5891eae76ce423803c805e93b34183d751e55a7270630b57a5600ffe1be00cf7b5b5b41b26dc8f9bea9e2645f20d3bf270ea058f34065d19d200ebec24d54c38e4c74e232c027676b4b33f12d36e859cb47ddf0be0276a8ae5756199efb9e41f112fe22eef94a6e6cd327e443e8c4765f762b28e58f52c6d59d2875f0491ae4c470ad6c1d4a394a8f5556489d654842be3eeb311518156c284670391ea76bb90e5daeda425c4eb416ead2b623ea323066fb58cf975ccead3bd678365a2b0b292744c4d33adf74e2567de8f89cfed03ceaba534fd63d9336b4b9bb255e5f55234b8bc35bdf6f0048ca61a8e7c1523b50c5a62d06d5f6ee9aec269eade250f5b4105e82b5d875e7cb42dc7f026492fcac295c8d1859e966264beec951c04fce12430be8a49b7690de909a628aff59a84b9380afcf68224c65b1e8632b336d4250245539fdaffc2d499dbd7b7edf13c2a058e988330ecb02c15734b98a06a39b6e04781bfc2b4a125b1b536534f32e312cd0f42f3e67a8e8762302f777dc7b1226822712f1e006ce7cda388029a3163511c49626dd80ffa11aaac17c280b9c0675babadef6f5d959dac66fee5f4b1d30ca01c0ed9679bc0788bb100a492c08b1d19edffeeab7b79221581dd5204bed0ab3fafd0df6577209d47346040e384f3d6e22d0995c1751b87a194ecc0995b6a178eb0c037c307d6d06cc96cf2762366fe8431e3f3d74eb78dbb35d00d712955532ec0052cc8d5c21b5aa19013df3bc1a221b555a20fce36eb991390401ab45c15117ff539a615e11ebce50b34cb86e56378dc75dfda1b4346245d722a115eadcab83831b55f528cab77a0c891fffb8e22c50650517ab0a9c320af4afae1554ca925861af7f9b68264ed6f1d078a43cad1514cb0f5f2ac10c4cfa1d57a83894861264459e38da65ec66e5a69a9e3268441b125f4e1b035fc887de12b04194d984ec83661c6aeb382baedaa9049818ccbfd9e0e91b36e99d3cafc3767bd00279a67be92acf4847fa436e05a9689a4a8030a2f58e0bf98a44247df7db345624b804655f3710b8553255f1e1c44b366bb0ebf9f2f8baf26ac35d2e613cdc1e48c7c31a74e6ea72100f0d0b8d26f86e192a07d649b9ecd8ccdcc012c3a7a1ecbd9c76771bff8443eff975236a80121a6e7024d7e6ad0a62c0f4e242389b7a6fcf6395c09984faec10a36ca132a351e17bd0f19271cad1e0d26cd9acc34d2d7273554d56454f0cbdd49e87393f82ee0f7f73b5f6fc72d08cbeb92d4d365917eb5e195bcb381385d219cbf5a01cdfbaca18830c143e934651c62e114527dd3918c7176bb998562ba6a94a0e2ca6157a7baf894f172eaede847b8c9fb1087c29b43e2f5bef028dc3f9c82c00b084e97d5cc0ebed5d3e5cef4b874d1a024a0e883803ebcbd821520d6155bf4a916d38b8500878bc2335cc776c1be2d9344f5ba5d35500ab053c9c0616a6b8fcc7290b27e645a8b3ba0b82d23834370f3bd00b236b2c939c73b6b7ca008d1c817f143e26084d8bcee2645d7e0b58feb4b82e522c90d4668ef00fa7432508eb11153fcdc3f032c47d1dc7d0b0145ab677c137aa3025439a48ab8ac348ce150b98a1844bb2160e1bec6fe56fc6d04c9172fd3e51056971cda60c4eee0f6592fce81671e398b82af5f42833f0179ed034a8d92afe1bb232665c58c740ecb886dbbafcbf85a8e87d762a9cba561e3f279244d5d70edd127982ba23e80ea1ee643f2c91f8411ba61cab7411dcd176537faee12f8cf83cd29eac64d37afab0ba24b9581681aec3793fc4a8694e44c41abc40f1f434711da2ff27333c7348d39d2a21e054a15f8cd54b1832e0b579855e391ff635a4a679625ae4fc14e706631d05bc38b7cb8e07f02601f55c08baad043741d5521d40b20b8689c4e731982cba692454ccc031388d2c16ddf906bd4f17e0c3e168a7ab7b9c51b6a0c20c739c669c2b8b318a3899015c360c36fab5348bb8c9063aa7b2972c9e206d03ec6695e12bcf758bc9fb05fe6f4f9d0117fc6be7f4083c6ada95a46aa7d0d37d4e1cc1bc247de9b0aaa6e42dbccaee328f158953300ad2ead5d7c631587b9e68bd556b38d89ff248a6223eeb05d6feda2daf12c74df02652e4a9fd44e5519823a8924e76eff59d51eedf29efeac1b252956ead8d00919bbfa410c6ab040b15ee9ca5ac749a3f2c483ef81519bad003bedb5e35bd0cb36d4759669030047ac220a04ee31ff0ef40d2d4d0388f8ace6779b518fe42c60384d6f129158f705acaf6cb7f8683e6bd3aa22a4dca5dbb719bae5eecb6795bc7f6af28d02d3060b632ccef5bde47aa9c6b751228e80525f3d0a0704e40cf3b726e727d1794826fae9039945227edd8f05df4448b80eea739335062da35de350f5efe981855bc47214bb2b3eea6cfe30e4a2e997de5d2872cf8c891a241afade5fe4ff3e5ee2ab9e11567e7b50e7094db21719667d283a8d65859f7fd487ec5a1a906f680ce270f4e4d68001377f401d56e369506118c0b001758a36f8e616cc0d50d67e552764ddab172779479c3170a078dd4372a9a2671701eafe83f95b4c5d1dc9874b10ad87687e14cb66e3cbb03770c7fbbebfca0cb6a3c113acb9a4b2eab9c8d59750187e912bb1145b4b23de18d65c082cac9c4bd8c981cb96f8f03fbbe06108f2248640f58ea4b586aa816888f8241d40dd20839b574cccfd66992841edf1389578280ffc3b8b5ce47575a466a217d64b004d5a1c4b9164d022b5fe071e15846f5e26f736425f4b0ce31be8a858e91fa791253836b403da0117f3c5c29470f3f88944041e82f10623f786625cc0acab7753526ded0da3b0b3e29d16ac9f7e016ff867352bb334c35da7736d6c986756e6742111f5720ffe10a72883e9cf30604daf3a749463fab60b61ef036e5ac42d88a69ff97341fa4206fac78bed6891f2fc4d34be0010e7ee2ed2d6f345df628df47aa50305e4b4ef9f5f76ec961d395cd20bc4cdc0710e0c8e5a31b8fd275d6c456f33c9333fa29e6d149602f4c43b42d0159c234a1ca3ec6ae13ce743809c0d2a7644a457d359fda9ef9bdf1ee2359c414c6e82f5b49899a2642e1a7ba18cb6076750329da87f4d5c921b1f91751d6a242962ccf0f7ec6899365b8aa6dc0a8fde146f7cc12f0afdaa61c364f6ba965cba2f89c74c1f244321de7e27705a0d69a31b8892574193c2ff9fdfcfb51eebda2c1efc8eb1a09f86b74f67338e22ce2320be77ef99774d4df221c04f942663c8ebe630f3b0c1c2e8298bbe86154f62a31b85e9160dc4baba8be1cadea90313f7aa2e7a09795ed0f9cc1c71570aadb673badb530e49c2608fd73c24baae209486db68266214b2e3212e2b2d7b57c5c43d22fb204f4f937dd270e9e8174d14c22c2f8781766f0e810295dc7bb99b7a17f3701c369abcaf77fbc97483059dbf8adbc3ab034cb0462456bb85d353f56e1c72d4e75e3b93c75baee83e294d0633d9473e4bdb9cfd71c9f61d0fa3624c50bccf1b040a1a5677624b4b995148520b7c5ef1e5a27f1144dcd9ea35c181fdb4822bf2918cc362ccba386926cd722d6aa81aa0f65c917f1a0e0c0b95cb8f0576dda81d94bcf8c65cc4c20fb2d6e09f4b852aceb7b3d6c12f0a91a61b0ac3b3fbebeaf69241cc8ac94cef6726f41ffbe25006cb7270ddd4ee83928153241708de53afa6e608f89d78aa8bb55564d346ab2ff473398504af0ca15da3c8844a2f91def4f8416e1e8ed6c4859690ed8806c461824bd9258011fefba1c6f6d4215f808646bfd6358d02ac6d272d1b18f203757f72a03dccb87335b2ed695146a78dc481a8dc844bcc084c694828fd8911ab37a314c8575898c345368240beac90402bc548f02987ea6760c574b3ee80a4f5ca055d7eed2a1a7f2e3dd51113fdadc4044a229fe95fd44b7353c00b1d2dc2dacc1b605e5819e42324d1a5ab23703a4dd0985cc35cf7949571dd7e4574234ce5e3b9c1e6f85f894ad63fe7d67aea9c2be41b8a6f55ac05ba20f3e959394305f79b4f6d1697a8d93f369fa97aa9c5288460fbde5b54dfacf83b2d58d4e28e762000284a272beb1d253dfd4163e6680505ddc43bda156ea1cb7758e982f4bdca8ab041c2c31337bd8fdacc3cddd7f209c0110e51a2e5cadae4b51e11ede7944d9626a4e0a0b2b557fae32be7332ee0dbe3944b4fdd61ce5cb73f154ffb9bb59a83aaa19ab5069f086000d0ef5a5d2d6cba49c769397c41b64c515be5ee9b3dc4a61f4da95ea8b8bdc24c000d4d8e745e014dc7217fc9c07227d2dc8514d60de6b965b61811a71144a4bda48b2fc791aa2fbf2702d93ea0ca0effc439d390b4e4fb5d17873f3743b90a7ff1d0d83f6461264e41bfa2487a144b8bbe8e5c651d6e3dac7fad4559a43c5fbe57d42cfd724c6ad8dfcbb984ba24b559f5d67e40051e373be0f6607c23e447bd6b8f48d1c49e8995622f63575b9987c381718aa4d7e9789e3b17e149e6005ebdc83173d23ed74d59520ed406d0cb439d6ef0e46f6a4af08149a78fbe225ab00a30d653debca75c9cb3b9375df6656d17c0b6345072c9c5af4dde0f4fc4f5237b48dd13bb4deff895222ceed1f8c59d11c1e0125573f1e88fc2a3e23519c382ca7c48e99e318d1c7138e701ef6aaf163362c57580896b4ca758e77ff917747d2ad64f39f172c41f80b48982831fb684e427b64751576b68485f44fdf18840854dcb286a796fe269dda3f0d9e1b861c7ee61f4603692295077391971fdda1b8488;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h2dcb510c5524b221c71037ea48068a9ba0af44b7da47a6b269a4f89419495b19280235412f352777df8dea1d28dc262055c1540ed94f6dbe6e7d8f3d7a1d39bd69b01c8d2f58b68b1745375d6adfb26388e241bc16a0ef419f7fd20eead0e02c41fdba3b30c962f2c1809167ba6c56cb9a39b5039211509694527388b7aa14e224e45e34b34c0caba29b9401b69777427b34136ebe2dc12270df9dafeff23feb249920ecc9946a7599f5828e0aea3ee2b22013a747bf6d735a37271f94733fb4bcb96280cfbf435c47df0101dbfaec567544cf45d912a358adfa8bddfcfdbc5132e7e91ca957ef70ab1b5375ef66fed7ef446a9812dff861e14518637b163b679474a4e578086d2221422750b416bd4fb1762f13c3274f4de39df58dab01dac6b2d49f4143ab0a066d74f7e692ee195928460d35b9f8ca85ffd877afe4d843df851cd167b7949f52477d52850119a8467519d3c3484b4e938439f1824b84472b5f5943ca1bb0bcd74f6081010e227cca9e004c5030966db8e2cf7be6929510b312d6ee7ac915824ab9ef616638399292c2dc48e234b780aed9d2f6d08a6231631aae12c2136c724ebfbd4539fbaa000d43fc9b6ab345d24e0e69d094abcaad4f46e59ebfa6c4c6bccb817476e0c9aa46331885be04b8bc8ddb6a29543845de44002d642fb16f36c66339c2b417dc484794c691372f9759c45fb51015f20497445da53a7ac4d91f537c4cc43f2cf57845fde539ed2b262124eb15ccb54618b0eef89f784ed5dd6d604410642fda94ab542d58ace0800992c27a644933942c3c12fd582de1b21f1ff3493cf4623d52b98f98c4990fb59c66ce6abcb26f1866c162584c83ca8a3b7b1763ea082246c402736da1914ebe5941c3717aa4aaf91f3dc8608883e1eea42d02ed6de397b112f1ca2a098076d2f2f1913ad1e0d50e048fd4778e436838bf60441a86f14d8fc4e2980684a5b1215fec2e53e6bcdf38d91f915759164d4fadb374d6bf906065958e60e796f07b963959eac2cde80d6071ab6c5d3a727498a7931cb00c74efb7df3d9a8c9e12119b82bc9b077d3419162ffdb061a707276b3f4830a5be81966f8bcd78f7873748e602bb767c14cd0498a0d27d7490a94f36b3eb88fa01675869b519b5d475bb8d86d8711dcc1e2b6576b36db1fae8cb613eb63e234c2a1e5a59cd040916228d168728a6f7878a005cd570af7fa306c87076152645c1797590857217a71ce07c0dc2e09c2ff5253ed6dea951ab0c78864a57c75bba78175d9c859b35c5400bc1e79450632e899122f439f889d896531ec6a851306d4a49fed6171f6f186df5be2ed4956cbdd48dbc77a507c163c8ffa13085967ec20656d376411bc82aa5939f10b722a0f3f93409a217079e469490973843400fcffc5b2750ddd37b5471c5cb03656baf330018b549355d10dca87aaced6ae032da161a08dbd65c9a8b5014f5838f55c32796a240e2f3baa3307808b72abe97988167a858b19a3f0d7c84e5d8a4c049a6f9fed0d5e2cb43e1cc894fba0f6686fc1327421481a6131be7650074f900e52678e82b61eab0b74c65e5287dac1a45d77652ff23aa09c56555d6a75d50b07c8164784b7b0fb73defbafac47daa01af687d388eb98771da09195d483c0ce5487823fbd58f8b5bdb7e35cee31d9590484fd36c4ba587e73adad42c9332f680a755d43fc16af4373708ce596d96d9a9cbcffe6cf1428d31e97e2b27d0ead1279f7e68234a7139fd32b540220e5c899a5366be4419d279ea06d600a1b8b0235adc6508a950dd17f981cfe9ef2e2cc1a589d379abaceef5b89d5507e7f3418d8a09e170521b7c13460af0b104992b76a43d58d5b6158756d4c3651a909288326549778643fa1f76cf616857575d28a956c5d94beb4426cb4a149fad93daa51a108971bb6a20d973fd4b98b5276a04cd64b0eec5f642b2101e6ab7dd8a75e3419b5149ad40c40bdbe9a45d0f6c31e8a2ec373e14ae02bdfb6765d9fdef53626ddbe3d11d3d56a908e16952cfb98a973b09013d4b8134f340d9ca13a2631eca8a15275d6a35b64eb1a69002ee45aa76ee82a681c5f31472ce239950c854e87c38571fe2c4051c570491f41c05583e291749be63a143cc1a9739511b1e772273fef5155d60d05eec4bbd59bbbf11ac47c85b79d76a6002e87d786ac9e8edab584925dea875cf363b8694d6f8fef76a0cb3bc6c52d572e0d0b1c508e2889c9918a06b656df969e80789685af60b321ea23070baddcd546713304e325328373bd49948c12e00fc69956575382234c693f7f8f51285df33c8d0ce0b50ab70ae32aa3dc2838301452597df04e20b66926f8880479e165506cd1657bf7a04e142f74efc33c54a9a1d1529291e5ecd76d231cccc575e8d3041cba45ee1f1d79de08b7f86adb0377a1effc8f1cea1ff412c1ff8bd2e875470d172f913cdcf102f643d684f8e503f05d5bce3b84c96334476b36f6ebcff90c6442e81cbff4daaf27ffd8a8c31fc01a593773b2724a1352b43bd8cbf7eb09ad8ad2f62ab6480c95128d27c029cf48633b9bd8c4e8f5c819672bfcf79cd2b60101e243683190261c55d6eaed507f404ad062ea0d348e57b6036e968aaffddc71dc33b06c64554ff9b2782387c4ecade5f24765341d6a85fe71e5f7ef370a2287c0784e61f0f27372725f4d7c3e3a455430be9a11d04be856f9b721193de350019998d3c2759082e6b339d92aaecebd562e45d7bd48e66846d0b0ab877eaf71838e8c9d90f36f2d2cb384ae25be994444dc3bca92819e8eebe77e5a5fd1f2e31357580df06acaed30c3c685778c9da06bf4e648f25a87d9dc02088078e42ef5369f61ae54b9a185c5e83c5ebbd02308b0d2296b25cbfbbf2188d21f6a95481c891fe1dff327c56e4e2dae01b278fa6047684a686eb93bdb8c01d42f362147de9150d783ecaa4627b57b53ebefda400a966e1a4b14032932206a77094a110f0f229950e446117e02375bba39b8045a5c1562a8942d0da286bdb3ebf7a25f92061e4d5680077f583d2a1ebec7162bddbbcddc3d3090d00036fbbfe3fe248b9c61914c699abd7e0a53c0a589c9185325e1c3da2c7b54a8472659ec0bde12527e592a586d745ed3302b8d37dc6ae74973e4f39d734616a89c7fa3f6c64b751203f69d45cdaabe84478096b61db0a103fbf04a843359b2fc38ee6d247047bcd110bf4e747ec6f7f7deeaa76066625f74892561f23d3c929b6097928989774e7d7749c1c62766fa38a047812c5e3dc3bb4f8aeaf0f938aafa7d62bc27c3344338aeeed3183e91df46359e7552390bcf9ef3494068a0fdcab60adfe47b9dd3f113044c9220aba5546d1ce33206d160147f4a52879788e41c4bb506eaa9ac8599f634c0b9fe53b764de18e8d2cd364b7364677eaf9c38cf949b50322739a0810edcfa256cbe1262ad92abe2c4366576d24709ae1af566695e15b22fb2054c9189f2e17b0d0b1ae78250a5ef3bdde452e231ea3d7ff98ac24da5ccfb01b9511a24d0490918d99611ccdba76a1fa727ed8ef509b65af75fff4612a97588aa11d5214bd3745009015ad83631671efe4d429633a07190a436fa2e84c9fa73dfa5a81c4dace19cef3aada8f658e09f7b2f0ec5652a668264d094c7f3c29a343599cb491d36b1394173304737dcf017fedc0dca1004e076e9b33fcf4b3362e7da71833a829bf0057593523854581cc9a8379cd4e4c0fa5e9925b859c3967d0b993f80df7a75455e5713fba5336c605c4f732575feac0d16267ea6f89ab5bff5fed9368e21fc2599e46af5bbaba8b121aa19c128078e9dfa1afffb888de32501c39d98dce63701adec80e823609587f3dcf7866574723c293168440be76cb279c558edf9fc4077f71b6b65fc5f6f6e3262de3e239c9a6372c29428476f42515c6dff92891ed5228cb80eb10647c30b84284c210c2232461f13389714186dcb746ff3d6df8f12004e2d629fd5c1139e74fd6e34c3c6d97982980ff3cd4d9f43dd57dc54a8ea45b89da8292d2b510388aaf8cd6dd9a1d145c4bcb5fda46e4197159f493d7596ce00a74841a23863a483d4dcfbb2f484fa10b1463d342a4d81c7d81942f930d9a594f810b1e8b192d75b169c0f1d67f430cdfaa923853d3314b411dc23fef5eedfed66105ebcaf6b2ab09871532b7b6ba471d5f8f2dae724a0959c50a52160503c08a643f7af9eb4a62b74b08542918c5d455b7e936fbb090c02ecc877c1667fce60f2adad33dfe51ec4df8f9bec8142f1001a070e81971cdf1ae1d4b995cd3abb11b6ea82a5cc2db6eb4b1b8b4a73720b32721df768b789af9c99fff5b9a298eef48f41c563db71b90297beb57812579ecc574d83854a2ceb921884a3f35c23802967be86b37a7bcdd3a3b9d8c8e0ee3768adc66490c76ddf77d0c7b911ee76d0822de483a9b16ab835c8d7115b4cd3bf502a3dd338c662789d260fe2796c1028bc9bb3fb44f4b95603cc3c89c6d3ae458ab1d8e81e5afd8ef6856a1b7706f2f84200c82c220c559291b82b76961aa8a0e43c9284a9c8a498f11deba5ec79fa4b33637f4c80856a09436f52c0964d1b0f63854a6d8ce1b401e89e5349aaedbeac17594b44f2effd8089d8134044aec33c67b3d711a65b456cc28a7c6a691baefcf19fda17440e353830a80923ff32c6753c6a1d9027d76f06ef187dfaf1fe51664679a918ce72a1c304ee1516ae7368c2ddc04897e5499cbf2495d9e6749ffc0bdd395ef0d8b535063cb671448279c3be1682e6f0f469329c362290f31e9256382addd876bce5f6b8e5dab30c7cfe9523a791a1326a2038824c8a746cd25dc3aacaf902cb19f22e59cc8e13e379d8e25de508a5784e0a60ca2b92b2d926c120a323690e52c6eb913086622a4511a2b94e219cffeee3e49db9eaa9141a9b2284ad611ec2993966bf8a4aa4d7c865c7e3a22332df0dd1bbabddf88c3c411f65ab6036a0b42f990811d059a377acb0a2f7cc7b83d22a7f1fd66e94d96f62662d2c59ebc008090175f6d3183edcce20567bb025c02cd3f0829a33c1339651ed17593fb8cddfae25b94224ebd4ce3260213463d70f81eab7721e3ad1d05a46954def25cb6ac436ff2e08d93c2fb02c46b0405e9d822f240f91073bee624111686d637df96007445514b4ab8eede03a3a96ee3b391967f270574eb93c333314f0f348e302deb6e9e7cc10eb33ede8e0851910d04d7708dd64a37d10690cdfc671d4339f79761cb32e58a45951d8dfa37d8947d2290478651fed637b531fa41bc34880bd4735d4ee3c1c93b111328e6ff1dce843f83c23a1c21f66cda94646125b9a9cbe12b901f5f91e05ba41c8ee3938686ffa6f2e9c561d00f31b1f3ea199ebf4bab970b2e2a360a160fd2b3c5f5472069859b4d52c6244d384ab0d3babe350ab55ad9821f70efb8bcb660dba3b4ce0398c49f6e88ad7a190a84674bac7a88d93ed86f9a6dab5c53e3e51802b9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hd059a96984e2a64921bf052b30e01bac1a4c66200d68113d130b6112afc4fe375759f96164b62a80b31c87bbdafc892999366575b8e9be2f67e9347cbc19fd410aab42dbae2e94b6b6aa03efe7e1f746cf5cbeba26516298635cede55dde04da9b178bc7ada634b4428b4160b13efed70338e21060cd38f68b54012ce188d8a36d72814e92489ddf24671ab3b1778b04ba6e88d329ddadb386566bfbc865f19e5c7bd2178d5f11d9baf9160b5be378c3d513fd6f1a921636c20d5863f5b3ba947b3133afac57f22670e3420a485c5ca516586a96e3d634733c0f958298e23475a864fc21aa80af5266b4faceb90c373469d4720a606e7d2b73392e171a092c532f768946c0381fc0cf1b082f9b9ade37755ddecd865daa32a3752e617e104cbf71acf1a5cbe53858125d55239de8de879ab9cad1fecf2786352e562d658c0c68f25dd5a988f8368ea1e43b2f8bfe92807eea11e711551b1f07ee62e424c8a6f33cffa8747027b2958ba5c1ddd3ab7b41e098667a326d53974e2b7f14754d81ff1f7a9ac8afad1e84aa10d47495eec057e59b59f94dd2b1020875dbfa68c292ead41cc94db41ac2fbcbaa39a515fec9f3b6a88fc9de300fc2fc72439d52236863d17c4252e1fc1eda001df30b409723566fe4c8a7658ac1e7b153d4afe7a45b80d086b00a3ba5e2f4c3723b2ddd3a2f94525e8667937416775d155035f4580952c3911eb57a4b46b2a40ff42d224ab7e41df3bcbf6a6b54cb18762fb595f6fd15cf191a82613b912127ea2d9cf6896b0473254fbff7498c587565b528b9899685abaff6f394b938677b57fc9fe486510c4b224f6bce3024653046a2ec02e3b3ae902d7c35f0ae2c0f5a15d2ed9b7f096daa92e0f7eddbbe96283c714b65240ceef532088545acc7c58fd9f4fa948ae2755822737c325acde13346d5dac1d5f7f1a5371a95836af5c6955a932e362b17c63d495f94ba96a3d5b3fd48906315e93936d17bcbd7c4b853836a4d0cc8f19f247e9a107b1f72a4251b0e73cfe59afb991787f25dcc14b8e751f773fc7b17b4675639b33fec570e247f00fdc9c9762b6e4eb2fb067bd1ff9cc778bc554077076bb066afcbdc11e04739ec13ed7b9b6c9fd890ffd7ccea9173b42413cfdfb6595c651cdce6329ef96ea21dccfd0d846fe80396c1d824828efb849d001323706bb77b9296d284dbdf40688713e617b787f1afc20a730e0f9f292337b917082655aa13fb84a2f9bcfd80cd69c13738f6a2bd849749106c8ec5d6fb294a53cf247e1b1cee626fcd32033db3e0cb462778e2bc5a2ffa6fcd7dca6dded62fcf21c06ae3ce1ea12de36af4737569d538079c9da1952983c8b518b4d3fcb18a73344dbcd6a890a0ddb129c4dd2c0d75d05bc222c3ff749a38c1f1b723fbb1ec1fc8664b8a0db03f5f73eb644b57fe6507b49801764fd6c38662a11fa50f9e4c9c53e814ec97af6ceaea827a5ad60a2dfebbe779e6e7577ec0ae9857911764ceedb463f6a2dab596ac765793cc8c8e32e562c66a1b07450cde113751334d3b418c26bc2983ae966d37fa003cacbaed1bd995ad8eebad0517d2d1027a88c79a915535486fb8143529a7e03149a76b55c817c3071cceb41415fa3b34d274d80468756310817d6d8d28e6135872d68ec01aefa46ee3a8e586e62654126d1a0848f29130048ae7487ebcff3048ce4ae98d14e59125907ee44e715afdd1b83fa342c445c6ef9f8e6b513dc4dd222dbeb07ffaf57aeff32fd5101942d034eab79772c876c17ce65bda92f3b6aa702e8e4e5211772c0110dd652e558a645aa3e072035afef23623186825c082edb148ebf87aa82c7464bdc560249fc0b4447eb959aa760216ca2b7de694535fe3c359823aec8046f206ebbf1dfcb23dacb0884c3063d7b5fd721785dd00e8314d1bfd2b453f9df7ad8b180908a3b3a8e81431f9e0c1b68417f80c6095a38fce3ae04d4f0e7d641bb9de301f5263fcb092203cbfe54af8789d1a599e29e96b8746070d4e458d20c9c29fa9fcf56446651f4ccb8a004457d125e53620caf67845af7b75611c89e8f820d9092f7b066e4c06b89c6b9dcfbd94b99dc64313e2a7a9953bc80a43f964ec143ecf76585ab58a6439b80a3db2d008dc2062eff21a9403872182fc3ed3a1cd6265545e9e620738a1750f54cfe34d441abe160b58d75989cf79c763ffbd408d2877426581df982c7aa60a1bf2ab8b2df1a6382181a0e2a0a80a5c46767e7ab17d4c619e1cf3f4e4b58943798ea341ae6dae548e807af21cc623bdf87ec28c53f5abcac20eabe2060b04e93384ff827c4ea8b82bb6dc378ee9f43e6c0b3f6116018e9bbb1f871b4fcf209fbf685392a067b11f138144f38eaee37fe75bb2f0e3f297ac13aff746fd3307ec9545a337da60872533a2ffba81bae5a39437dbe855f5c0b6206a3368550ad493df286c8c6381a8cf1fb07c3ef7276ea8e95b53e94bb473b9288e38dfe9e07aa04c7f30bf18b452ab7ceb855c079040a5589d34e1d68a914a186bbf677b80aa59dc7092c286fb2691ef915fd620c045bad56ff07242af2f66634bb409f58b6062af78c6a27b11a455bff35c555c25a0423aaee83cf96592b06578c0f661e9d913537b6aef7821e35743d8a573f63194588d449f06fea349f5ab5eeea8cc2d514c3d0b229dd986807f17e7d716d7cdb425c6d5a717f2fd169854bca2852cd54f2bbf6a8ee622f805c828cba99fde197053f45395b6940a63ef99153908503876c4e41d1afdcd11f33ce294ee037be42d6e8e6b7441737a734509635dd4cff543b458e5b0f46c6077a0361e69c771e00cae70a964efd5237723e903bd0fb80b2c0aa1b825e911231b53e86d02a1490b0882ffbb113d6e1dd930f4501d6dc3e157078a4e89edc50d14eb3a4ea423fa3414ab8bda945ee417612e10604c4e1df3487031027d480a0ffb2eccbddadaf7519d499432399d9af7e34e5d89c51ff4663d864cd8958d090fadc6c00f29c1754b2db586bf789e6257547d3fa1bc11d45963a6201de3ea18a1831d9ddac38d2a21d9df8890a258c8adf97fac1cad6f6b3808eefe3f2f52f6cfcf30a5e4c084987763d73875e73c7d0b77b059cf62158e366e27be33f14b6751e3ac13a9152bf552511f25f7b0d37838a2634c7a96cb5c764b873e8c6883b46b3882de7ee1488ede7a1bbdc0faf45e730b0af59b7d222fe4c7dd075910f7be4a149c7bc6907f0d9c041d5bae80eb1c0a7246473b64ea3e5047c32a35641885b2a2ce1723fd780578ba4c4aa5c9b77b9d2e2a885c7600fe721642cf887b019873edf4b8adea01a13d6e70ed32f9c751be90878dfc39beacb671d9767bdde1497e95d76e09d7ab93e51ff362ce4863cb1156dce5cec242f1b12c9c7b65ef812b6e745c0bff19b6ea41af47898d74c8332d9eadac4ee139410ea0e717135891646a7b38e4c85a74e57a8cfb47b22d1672802ccb7bae5df8e19b83bde7a6349cb4f6fe9e14ad5d35c943e8d12a99d6b9732bd0e13cdc1e315e0849aa6b176fcf8ff2e97a993469f31ccfabe8afa48a6949e0d067eebea3eea6a6bfd49702a97cd0884fe6efe2d125085d55ecf2ab9f9fc421ad5b82d1189f4f6d1144614392faac32a447871bc3f222b2b621776881c21d3767b57aa512849825c5cb844df137bc001b179b26155ae91c9ebe4e15b0838aeb826dfb9eb38fb52a6d9f28b54ff2985b46446cbfe5bfdaaf649eeab0376d78cdf63d9a965b0b884d75968537d5e81cde1b4384aa2608b3d31ed5fbc2acc34d7367aed510471ad2018ca25f9af5628f68587005cea1a110ad6429d86f28e7a4ef3f80ea54071fb152a09a2b8333862754058ef21fc9947f393fb28f91598f0f2b8e1e26a957bad03df99e3e614c72dd65faa2adbf070797365f31c0266a95f92f7cf50ee493b0a61990aaafbc517a630d9398e7ae0ef37b603709d67e54153b0aae073c3e22c8c8112bd49874f6c11725b787ff1fb629f413415e1ba4aa46fca91f604b9f547ac9cdcddf3f1c5db69430e6863b95ad286365ebddaaff783b69ddbc527ac9250d006b2290b4c6f1ae93e57d7a5854b106c096bdfab0a51429b3b92d8ac0c0dbb93895d92b1fbe4339617df42c46873650c6b701f30247a71de4aabf2495016e40614888c9e03eeb3bad413f61a41f15375d449a173b07c4e258ae7901f4f921ebacde36a5001ef4a380b319ad775a8a42b54e1b0d1b19f8e5300ecaaba0110f4dea466690c98c708536d0538ab6c951d21c0c91b9476d3dac1f8197f64cf3aecb57ae39e42f4a2d18f272913069dc1d36093269b4e1e6bc7daf3c0c5ffa33280be9f5254ac71493e5496363eded7696e7dda9d12f14da849c4533752d7c958975a134409ba84e975b335e4ce929c6173b05654a68c83f60426fbb47ee990e12403203071531279fc88dcb9260fcfc76e54515aec40a310e6fc47846e1315f278b72d8ed8e43ba3bd559c0a0e7bf1f05310306f865d7a423f47d4e67993f57cf69a06a0618de52cc12c4e1d3391f406245b27ff8bb90874139bbcb96331e441f69309b2671e92d8f6295fe61cf5942f93b124dfd96907c893fad95144b7d4b88448c26776a35e23723fe1c55224f36d8d923ebb10368c5fad3e8452cfa9aa2c8bbdd0d2d0f1c7a3e7939a92cc6a99c5f393748e6e8194f71b73e24f37e3efe6ba67d6d127ada8fa489932973534bdca1c1192c8c5a9bbc95c1a636db29607d8ec0e8189cf503b2ce5551de5265c65aed91cc1d590be1a70d8c9495425b653d63b74f86d6679d4fc0332888be8bd7e507e580734e79522383eda3abd6010347686abb60e096e96e34202dec4104d477dbcf15d2d335bb99981dae7779d7ace371ca4834b9fd40c33a07e5cc517f86aa2d06d9d9719c3b2e041c57eadb9e128ca18a53ebf489df0c79de1d58b861f82fa4fc11aa46e638a2fdd89c6f7b6e791c4a89733e5e69b044eed5e69ffd6f7e309514fec88ef53a2478a1a4dcb2c33a2fc92f8e71e0778839987d5db1ad4b434a73340dab32b2437597c8315ce63e6280ce798b55fbad9d7fc57430d5e44c359947a4b4541d04043d8f2d409084d2da4a12d915d2fd9cb025d2ab7523d416a50386fbbefa0a1eab8d11ef94221129842cfc5bf80fb86b88a73532bc8db3b964c1467acc81387336c68274ff234b1db956ac7686ba9f04c6f83ce36a84bf5a24c254f5bdc766f140deaab29c59816ea427b472051b924954e0b60e3f184063e49f37cb4435e931cc8048d17bd7a87d9dbacac4735ad1518e43cda5ba9770a54fc59cbbc30fec3f57eabf347c5b449a7e287e5ea3cd9bb05a3a466232a1ed10f7d622cf2ac7dfdad9c98d3f6c31e8d13e8949fd71181a8835038c3846f936ab718ca6222c669ae08522e8779ae4ae310e9c32feb32e096e9ef50ebea3d855e6180c71cfa70e693b9552a7a00a35540928312b34720fe180a57fb3afa87aec5852;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h54169242ed9cd3e830f49f5bc2adfc0270bdf91190d26203cfc8cd14be77157a25b0ce9c2f17b7175d18e6de5ebebe5f57d49c799404e71219b69af695e5c4a7b89d62bd7ce41ef9539b79e05c6143c2c8c942024f1471a89330e7a0563bba47fa19fe5e33e9aa31293967b52dcc8edf03b3e1ce80bd5d8ebcc71843a015d44e9cb17a1e798045a633146b7f9cfaa1ca9cc2fc7c76e9c2b1822ac9c3f0ce2e2a6aa1614b7318872a2e42da41af1d57a42b5d9721b2a25b476745d3d5b596fced694d5704d2e7b0605f7c0b668adc58a1afb9cd25bd833734d7210cad43095e9eb1f502bd82f3b7621d53b5bac3655374cb11758ad3860933620434ca82f4f617beb7d27583c41c304fd92f7743c898b3be4754075f24d6c12b275954b88be9c6b9029164418bc77614fcda2792ea725994dc9040913f5606b30a223040b1a341c2e212a0a2ffc2b649d16d7452fcd60ae2dcd6211726031df9b03c9a8e3f17bdd00d1cf20892771c1af3354c8fc1bacf6bc869f23cccffeab8aa39b8453b930a95338e0083433c8462d64c2068388235e077ae4f5b85629f444849e9410f03ff39fe5708580d0ccc47ba105be85ffb9b0ff36227751eb2256817032a7560aace3889fce517929c0dd83e09a0091963c2e16b096b53ffe67348e59ccbed452608216bb12831950dbe37837d1d10086e80db4d505273649ef78895fe4662bdb8a02e2529fadc969beb837989094d37c6375aafd7cf1e180aa02149fd6562753c33806bf8eb37f3f212a3e9c53980bc21e21f4c89f9bac5368342801eeb96a8a21a4ce7a77fac7b45058c53a4332be52bb70709e891f580f7f45d049bce2cae96929ff5c2564b42acede4ff263c433b183a20902b34e0a2667920e75efabe04bc47097fccb6156df1e4c253544cf706aa360fc1ad5d255775222456a891317e500c78ab6ac181bd6cda5ed95d7351f8eea0ac85ed78d3557d4d86d1848a63b626d90cf9dd950a3ae9c56f6dc8ec01be150b156211d0ce5cbaab1b61bdd3bafc3f46b7d4c54e34cbb60aa827491aaa8bb639aa424e65704765048c9f6d0b16ac0348a6adc5f79170f87bd20f4149481de84bb1a27d545072ba68156fdeb7fad0d9272ed0e7fc57d04c62d6f57f9b9bceed5b20c87a2037f85292b74cdd77e2db24e93d812d0b2f7f6b3b91a3767073bde4372c9e6133d0fb8f81f3f5b67b3367ef1e3982625cb2ec7da86271de18144b02f8ef83a3153c484a56cd87308213f027cf50a93b46efc4005fb2dbd3dbe5abfe6a54ed2056f2b01e29c1b88f7b873c9d242e989f209c1e0c17b3c19407fe37a12e69ce7e1a39b137d5c8b1f4a43eff03a08c2c2c5abcffd68beb64581772b9fec5f33382f30373a4c34e56780ce04a1f0f10d40244276e9e77c8d0e7330302d3be5bc7783de1838c5a9e573734accee1d06bac0782726a28804ac4b9351fbe99efa19f391e92b1ed0cca3e325ff13779a03ea783026a00023c900c342205da0c85cba73abf048a1aeb0301abf4b77f66cf40878afb00996239b097bf2c6ca195941c14f73c537ec79456ae2a730e58b219e32b0e9cdfcbb90aa8f5c4d493895388691412f325278dc8f856cec609ed9c681a08d037fa90ff966542ece41f0b2aaed81d10d7507440a74b7a750bfa388661c40dba7bb90e8b67d6ba1571a37e73e618ff9c974127b5a38a461229db9a590868b680c58051bc1b882c7c26354d5fb7a6b5fedd6757d4e4330e4401ca2c0f8ac5d4f0f8e84bea425c253b4d08aac81c7305748ed273028ad09e85d0e4376311bec29fb56a92b158874fddc7ce731de0c3cdf1ec52edd35903a617d0fb73d80e43a772130d62e2e612873b591ca2979f691e5343cddde3d71c12a4b96265c13aa04bd39774f5655023fe7b46d3d34e793c108079d10f4af9ac6aafe00c5a82fe343878cd92538020b6f412e232fa8ab81580ce9661972b34c51487822fbe1b083e520e5a266fb7dfa917886907c47a192c9140f100b540a15decbf39ca20d677d7cbcb5ab2d13d4c73a07ce5d26431ba748f9cbeeea96236e108386eb512190a541996d948e713061506ebc151d90d2ca295316453be70dee94944d7e6530c1a10de0c92307941a68b85ede34ad6bfb17c38a960eecf399c40f58d07195a498be8d6773052ef4f5ea01b9c2296dcb2be62508fa659997ae5ec126e34d00c85fd597442140fdb8b2674d0888e314586d4acb49c6df916e020731cfe8fbdb290f13452847a614ca4574e016f508995bf9adcd773f1095feb5d875c15ba62132ff45d8fa2838e072b6940b3909552b2e46d455f2ebdaf4930d4226ad1ba35999843cd8ee02785a00aa4131942b86863037be49c260f5d26e989484268ee42a4a1f36b5ac9786e68bef626f5ac56171188cfc94d5fedfcc5536aaec1e7f0ace463855eda2a7fdb45b5634a2e57f8427cfd44edb514094f8acbb35eea60a00c4d112f357e9221f50b43e5446f9e239666636e0ca04ed4ce2755ccd6154cfa7f0e79eebb19ec5b2a1baec307a1655e251df208e7d560c91f4a93794ff9116786cdd1427fcc58d3292c8770e337f07559cd98456497948c908470dabc961b7de65c9d88ad252cc38aa1bd813e86178c1e648d5b986eb429bc1b1df2fedca4f24e0b42e1d562289048415f7b7a104e0dd6bbc3bbc75e0129977139896fa93032c05242321a983a0e4db85628779f34571ad08f37e3d00882d47b6dd843c5b2fc1f5d61a21390911f7bd66ea9af1ce03bf3f05f86e7a463a446555c4633a38ce124801d6e845aa1a6bfd9c301d9a757cf90daab28977642f06c4057a53f5d1d746c9d0a3bcecdbeb4ce285ac32fa543ad6fbb6dfc260167bba9f1d41515417867394c1d0ea13dc5d29954803044559adcaf02b566341ddf23a8ee9f1a61fe66cbfcca6da1588f09caa75ca26744f2325fd5c5cdc03952f8b187b8523e470f24729172c14a7eed1ed8970f9da56e5ae615888ee73c52d9cd9d84c3d6c3aec9af97a22b5faa0c41a99de20fec44081a5ae64de5715723a472030b3dee387cda2a84e384c428946f6667c0e0d5c99c36500c072c18ab73f54f10ed04ef8ee6db0a39fa71131f9ede8ebeed6e0f64890054f3cd6ed8d74a0ecc2b081b71aa657b084787db4cdb9849708ac3666471ec2eaab85e7110c3be0e46ad5d8d3ea497386b446a5e97e38939067ec2a8d0117130984b61f414736797135023d4a03d13b2a44e3b8c74822a3d48cb09249e165eb6c728671e66540dfae9ef277a3cfcaf4a7d5e9fd90f03681cf87768ba2e3bdf4d8e0865a75ace384aa7b3681e80d19e8dff61187aa8ec49aa4828e57d904fa0c92f66800b4c4b9e390fdfb940b30ea3def9ec840faf464e9829e57081afee325b26f035740b2c8bec29fa8ea799a7c200194df1623c22a9e022279b31fb774e099d5dff8172645d65fe685490efe064fcaf56d07c1310d13f28f392695b43d46d58563fa1963f5b6bf97abc209576fd9c559e9b0a9f66df3d95265d186da34b808d92efb12974cd0a9f00e23792582424953b317ddfc76b65e2963a7cb6cc553f7bab7fddccccf65b2f0099f3c424364f93abe3db2c32b34c6b2665e22279d854b9aeaa131def5fffbee89c3c06993e1db21b75d5522e9c600e36c1fb8bef58004d3ae200d625a0a421b32009dff6616537d0b047235abede0ad2073ff4cc539b81847f46029b6a4de4f364cb3be1769fd8f7a2bd1c915d93c81159915a51c905f5c145956d95db2894bbfacb8faa23f2bcc09e3a804a5f40d60b65a6f685af61605ec38716759f593bd49269ea8090246c48c820186d40a1cee21bf87b03f84de8fd77ccc67b247537c0d84edcfe7362c2eb6f92429f068054b6690ecb1045946f7d8593df97454444809ff87a995e3918d34df68344b53b3f0144549cefb8173ab2910f816c8aca6ad1a36a4c0a2631d30b34b71cc7b3f32e004462c57a63b38d3a055b0749d79b5a78af6397b30910cab072cd51269e0dad6f4b9140008c75f297a7b923d344a371ba2218585bd9ac12dfa8e95844c827b1a7032fef0e02751e9b37c824ea96c088bf5359ae4bc0592089bb317d44bf91b149f8c3440f9d832a2c5a796f59494adb963e854536832b31a549ce73c7f0bb7826ae2839a6edb9f8a2c7aa404a42be2702e161e4cfef500ee76677ae5da734e4aa80fbb6475d30efccc1f4c59e1f88202039d062212732ed893d05e4726e01c5a7c7aa0a6be8d5384bc3a012e8a8547c273fc7bf514a3ccaf40e9828004ede5f571efc863f00cdebe6f190e0b9b911719fa699f672110dd71ea84851083966c0c4b8a7412429e684c17d3176e38392d488b7939794f3f9299e1cad366f75b45dcf997e45300a2e902f935d3d510fa4fd5672782ec81ad9e16d87d8cb1bf3898add19964ed0c4efbcae969f8b0be912ab14bb196c691cb5fcf0eac4df5226f246471d39ce06c23ea09a77a2667c36e0bc5fac2d5048df88922d6aa27d31cf5324c1c8320f4b6e8719af893ca49bd8621fbb955e13a43bec1d4755ac558874d035a521de285b2e6af8e0c47fcaa538e53ba5509bbfe0ded39fbfa885017967e8eecd502f7337252041003a595f673a972507f48188360b17871339f5bdc45228e5ebb17d2991dcb950f9c0831451e4a49476d21ecab53480d771f86ae8582b28ace8922c01332d21d4cac28fe8f342be281080efd15714b2a4de9847fb814875cbd26d6b5ad85f3a7aec27e95d72de5f9902a6eef7c1f865f902243bb86061d9747b01deaed9a45d430e61ff3a70d529672d397a333b8f6ba2532308cda7acbe9e51058211725be7fb01b00c5ce5cf7806916bfc788ee99f220cab59b9e5dde8a079afe3caafe8e2a874cc024c9e15e066d9cdf537b2010e464ef5cb4490f15fd3c435048feb438eb88f11c35db5c0c74839de0d4d772799266f265dc84a201028d6854a7efee2c97185fe8319b12276d917ec66233e165181ae626e573c82e3155a471192306114b3a9de3c6e932dc245828b712541911009387b0b847090b29e421b3a389218b926113472a7496c696f8514f54925537327502c6283837a63ae20838809f14ea4e63b831eff123a45fd8034d92971e9c8f0e2ce200a8c945293369ce50f3848121c8894dc7496a4c116bc0c647bd47c59a007811587cf9d0b71ffcf316ce9fb29a3c9a4cb1f7bd563857d7b636e4af2d1894acb933519b6334fd4fd6acdc0d2cd912ed840d78118c0b954604aa012828b4373f78612b7c00da45e67da2087582d2900e3c399efc22b036355fef563d035070e4dc75896df8957c31624351a6485a3f0a2cfd0a05b89eb2cf6a5ca9863c7102b26f66b5366ddb7930e3acb27b312cf800faa6bac4f761e8c2e954ca2fea40ebf4d8583e9698141c89bb61b2daed003b36dd85760c1e3057d7f801f728707bb37642413a887f44cc5428fef8f5432b8437ea51db;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h66636fc127778c817fae94ea44ef4a18fba170a4e51f6fdafd9e5547d594d4b373650c372c4d580d0553e1ba0d6c17a0f432c5a2e5344aa6f4a5c248a40cc73c7b8a667af73283cc12b6b40b8214a08a57cd18a15269251afb3e4abfa8f6aae42378c8a6e4eb88a88eca5c24b2176e453d59a9665df99f3bc3b22a96e2c5f1541dbf709d8060b5323e139ca9e83503a4fe3f81c4dfbd9dfde9bb89b44b48839505c425c2bfa71dfeb7a03c4f965401f2141651490c2b6e5e7cc0eeb74f473202ced7a57ce021553dcd5e08e05c5839083bf4908a8856a215199c558ad85e9653c55773fe22eee5fffa293c15a0b8a468916f9add11cb72c79de67d71a7f99c04042f45d06b6bdbe2e67cacf37e808dd980b9f219a6a7605e0dc00af53a221ec9f8f15cb10e0cdc7104ba00d51a516415a3a13adf0db9cb56a4e673d12d76b4ef7031ac638f0c817b9e69c6b6a4ca89ade3b11c59cb8463bf66407dc07fbe84846a86f84d9b03f55039ce6cf53e35f50ba0846ebed1cbc9d3fb819def0314bc3257c2b8792081015cdf8c8ae34cf0a72b0e018593512c47a63cd3488a53e33182f683c1ffb76d7954dc55bf853b5494a64340d5b3fcd6f7d6f348827a07cf4732ad83ae78369ccb4d4f1adf193e9fb8fc4d28606feec2dd0664507ba7fd28186dd7907a2d9d3fdd597693cfa287087848d6630cb7ead9d8f07407cce533bab00ff401710aeb823e6bf0a669b94d87eabdee2ceecedaab96c7b1645ee42bee08737d87468243eb8bf3de92747a9360d8ad5212ef85868996e1d6218a16a899c81bc4a3be98a05e7f1d16c0bf685087b770f9f2f5f4acf2cf7381480852277fec568d8d500562982b15a592468dc3bcb8e50006b0f8511aa237a8ccc06c230032cbab1a849f5cf9583cb0df6f1a115d690ae4ee611ce345ba012ecaa9389e2c01e1b58673fd0aa5c2e1f371ef97ec47352e276b14cc950b74576ec9abe538e716eb45546fb1c2f8fffe3572473e5a232bad6b67780bacc80ca0cf161b528ab5efd6696b903c068b7637aabf3bd766bde224f8f2a21057b9367523bbffb871926a725281e182da3533335bbc1a3efde15797a6e9614029825b72a831091e30ffb08e1c90bde87570ee2581176cfcd5144f808ee41ed7e8f5258b53f623c1ef6bf772ed03ebbd1e2bedaf1d4cb4edc01520eeec68963e14085fbad36c727c009a682f6d35bf2343aaa1cbc977b6f5d13c8e6ad239e828e630936a99b926806e1f74cce0b5f4d76b2076ca019dd92539d63737b987128f0522843b610ef448fe66f1a4dba99c50d11941a6731f941acea65f0f892b149b54fe4b44510f32dcdb288d2b9302afc821d60af1c4f8fa391a308f0bc6c76be36ebab291f19a7239d6589a5ec41bc0c863e4b2a676807c8718167e02c868ed67dd192d6953dc4ee2fc9cde403ed78101618fb05f6c6f430f39a44d7816ce65502db50145b23dab9f5be0530900199ce3fa9a14d5f839715561acc8fe3cc5cfdb7a7cd9b5cdde0cccef70d35a499f66cf3336bda858f7e59e6dec80bf3eaa1791b24648a4ee41fde34100b26cd85a56d8124e6201393c04dfd4124597272e4259421cc2d041811cf03f877750bacce28c8350802dce75dfd2b1c299a4231abaf7ef8f4dba8c8d369dd1616f024643b6b5533f0440d43e81d11eeacaf81fa86d03b72d320a0207b29c4ca04cb60ab5d867c2cae3b06d90268c068358cdf051f89091f757009934bbca4f82568a9a00513bc22e4a9c6cebe052497cc3256a4d4d118085d2614237a619b10064e1e90027115f1ecf7124f6dd9432a7c36ff9c2545845dd9ca803068370661a81293d1d373360fc618ff51de3aa6655bbb186ff462277a59471834eb5ff6e41b8868c5410b57bde2d94bef78013a2c5a66127c8d18d0e7eb4851436fc6dd7f4e1c00cde48d5cc795ac5d6c5042edaa491dc1bfbc1d09fd6e6c2dced7279c2725ecd57100a36f87a2de3b41a91ce0f88439d3f4a3314491ea9311be4d0cb1e60a408c7d500ccf54cc17a0f8abda5627846f657124a46dac509f0d36c2dc78500e0cb3d42c1dc7af2ca495e0fe8da94bd31737e765b64425c0569b54d1ad81834b38ae1b34323ea876e6ecdc139ab26c93f831326ac11ed666b09e84afaa81b558413d200ef2f665075d05c32e756dbd36c6cef748cb2da9964b8dae5d1cf0b1e9260716c9db172ca45357105adc260d00d5a3c47661cd6db8b6d0b9ebe9c9e6313f06b1fdef37b58bb1609e77f0643e92dbeb27ad203a3e0864f3917d1b650c377c09c320760a39389ddbb27b0b51a3afcb6f952c527ab31e23b85b068dd765f2a5478721d2f73c67f680ba4c2d80eaced6c42db942ca0e00e54315708f2075c859773c17fe7cbe6412a47e768e2c91147381866230d6784aceaaea86f2d53123f761fb5661655e7f9b5b17b47a1e5989bca673b65a0ecb2cc80387f8c7d2e402446555aecec4c14330601548d321dc714bd9f22b0d3ffd0b825e28df8e829d3f2510705e9bbc507ee48f55ed5c5b8fdac848f66a2696ed6b535eff020bf80cb8ef78783670abba6aeb3582925b0bdbd08604fac1f6e6569ba3c7f82875e19ddb7e49f4a191ca6deab0d9c607e33e271dfd87ffa4bf13e10d1d5c971e3fc215453ef2d8fcb71c27c8d5896450ff7ae575ed6c3863e4425b10e42a4aaef8bce831765bcdfaf0eb8baa7342863f46ff850408c6d18ac7387f3e4cdc2f365887fe4ff880e6d103f145faef0b72299ef2e177dfc6a90e0e689afb15656169bdf32a3a86f947d87fa5f4dd3b6ae1e9b2c99795963d8b9ce077dfa1614575a72b7d757e24c48190537f27c2622d391959456b1483968e52e04fc895f8c78b4667176a15b74a26101eddcfcbd56701c4611ef6571a48d51f62d3be7d9c2a824c69d013466884e5a9af2d8bbbcd8ac20605fd6bbf69a7f742033f5fe2101367a76c39c76d9ff8e0c33816ad63886717dedd8e289ddbfde9690edf3669692f90caa629f6aef310773aa139a4c197297ee0d464847a571ff07752d44e68083fd517e7e6fe266f25a863645c4484df2ade84281deecb10673cce86afb9bf79dd99b209d7dd8c37a837c9f0d53177cc620a794abacf52ab75289fe9d1dd25c1e0c457fb87209dcbb277fade4d0205f98d11de04eaa1dbcd9b1199b9eb7693f4d41996e53b9ed756778119cce9740cbe1d56f8c4bfd2cf5973783ec85770b69b2f2789cea2c97ce73abc6e594ae8d6e3d5436840cab48b0c6e3f4375b4a44e4666c541c56c2246e91236fa0957f27771fffc7e193443a82367ed4cccffd32000e487f42dabea85f7f253f0926484f4220f3b1b2763809a337f7a09404963c89aca5dd2b07e7eb1ea3e26f25828e717a7d022a499178f8f29c0ab33425e203bf501eb8c3fda4db67391addefe3fc5f62c6bb21ac0f1e9cd191ee3592cec74d6aec75afc9f2b81f3f57f9d51c6a8c00c20a60c4e603ff192c2ba37e5b9567d82412748cf4125d1771e1ca3490fad6b938d8d01c11c54ee881caaccb707c08bd9ebca14f12d7ccfe832ecf66b34738ef621101f6043437aa40f57578ec8bb5b4d43545806391986c3c36679d83c260c432826fbeb45c4755cee1871c88c9e43f2e5153344e222d94e30975ecab24aeb9ba4ef4f13e8567bb27d2423f0f7e72493a9f07d55396d2803ee7b3f58e6ffd2aef538a1e05e63376223b00ae1ec593cf3ea1f30cfbe8f950978a1c8ef84ba5318dd76318f77ea750f9537934d53458fe757a9761f1388119d04f253ce9d22b66375ca93870062c52a8a2e590516ae4f9cb520452e7af95511ab6e200c43f253760dd2061dbb4b4e071458ec6bfb6a7cdad11e998b88d3d656647415e7f45d0a020d0ca8d7eace52dc29128af058f07f039e87b834cdec26a47175c148520ff835a87e4e10081f12ded8bdb4ae1b72d07f2140e835d1440b0a33b7992ea9d4b5a84e6e99458d4d088ac1d271b469eb11ad349420853843e86fa8d676c606d206288065df5fe4aaab56fc232f73d5ddac2f8c2481dfb29243406931be690d02cbb520262dad57bad3eaeb675ced3c0a8245c94740ff92dd8c112d5d2a1239f77ec17ebbdfeea4011b63906b6f7183bbaf77e2b1f385d03de278b0ab2cb630a12dfd12e31982b9191817250c60d3baa5fb90a2d0025f66ad8455f6937072ca2a71abe2546d2e024b0cf9b5d8ce768d0ffc041d147ccb820b096c5cf5f2cae5194071acd68fcafe3549bca9f2c5a1a2c4e459e3879d44f79912420deab9ecbe212b3850044e132ea714ae346418fcbee1f183a91df8f0eb97296a06eadc27f17025f7c5a9a78b6b8309118290d705eceef7489c2dcbcd81933b936d21a04b8c58ba7070935ac2c8ae4ff8552cb5e336b70b38b9b3a5228a4da90fd353ca71672a1b9da9a5048c8d63ba11f6906fb5ed94efd6c244fdb55a5c9ee579f296599d38d606878d674720677995688825ac8c7bb43756ce0b8daf5682a3dcb71a826510f36f874abec5ec5d8ad75fd8259b679bb55978932b629a3de3bee21b1b5d7a13064d7147265426cb7b511339e4dadd0b6614f870b7cae03297d3f079f3a6614dc445bea1b44964121864887e536dcc6dac9b5a22d8c4924e6571674aee56e6339b22c1bce1e0d03cd43a5fbb8781b84f1637bb8df97aa4b407146ada3fbcfe96e5de221c0ee7f3aed43ccb4ab300ddb7cc472792440ca5e1ad3cb71983a507a00359c6df10ca21e76d534a027d177df8a1c9ddb175b53645ea329b8abeb431f84b00c29401bb61707578e838678dc3ed3035e71dc69cf14445a58eec47d4147a75245a2d621c5b8ac1c0490b32fbfb2a447c05bcfbf3cfa6fde8b6f2335cdc8ee86430df0002f4e8c3ac8decf612b91b34630f2ee319a5158a6752083ef930f6d3d3dcf00e8bce4d84c1a70d28f128fa9e464741afa289e9073ec44e001ec802f4af38b0b7a8f941107976531ecb763eb85731c0a40502f36d6231f7a950fc7708ca5fcdaeec025583477d67c4ffc1ff3ae72c578e76470890c24e85ca5aea2f110e3c5c5c9e9b93bfd33bb63299d506a616985863e7fb6c9dbf0d3edc8b5adabe3a716da250f040b44524d723eabd8bf735bafb533281129b227fb67c11162f5e3588389ccd0f390097deab2b408c4b2655a888bf9e8f7ebf300cd3595d1b48516b3978a9bd5197a90de20f423029d43ed1a26b0b48a8de13977f385d2836108cc6d66fcf08e3632fcff617ebc7fd8af746e833b3e86e0a8a6938c42bc0a59187801bafd5b4f776062c5896fb07db727488e2998ae3e9f1f32bb86140ef6dc442b9b3c2e5263fdb04160d97efef224c4015464c2b291f67e19f5e8d0d27b395d491fdde2b98c358dd9ccbf84e53aed76a558508102557e2ef9bac319b25709c185f392f2fedfe7da7eb04a33aab7cb7028e329ea392ac7cafb0ac23aeba5474646f1cebfcbc3e362846451;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h9dfbe26e90612b75dd21386aeec51fe86fe77329e858fc0ef98ba5f58f0c3b44c56ede0a7a7fb2801479ce029ebca39289b6316f17000ff2235f649d9ebf8340ddcb0dc7c367c89c8ed9d53b9ddbd8ce580de439de51e8fdb12818e549ae42f8a96ef63b5928ca31c67940ff599c9b1e2f8ab81b09614c7294d3c6cf7a0c2c09fc89f2b9f6ef41c87c819613ecb88079f9369ca843038729c8602d4464704881d07c188467ff6e35ace89a787bd44bb7239988898f1a1e37525a7824bb7a554e7843d8013706553f0042f9bae9e59cf2d8fb61fb967a8aaf650556256cbf2dc0a7a32fe4509d0eea7465634425b6eb319bb3a5f4cd7bbf1172c8d58aa242fc3cc32f64d0506db7af546979de39b422950926b13efd83a209df1b8d369413a9e70df9a767359990cc83bb25c30a1a4cac0f272d4e5d665a3c648e51868ec90425ea2c3169dae51fe0fb7131493fe16a5f248eb322b917a362f4b0bdef8f31bf48f8f3ce99b947c80ac470ce0af6bcb3fd98d63b3ce3d6e3c0c4cce55d435da8bff14e9397ff4d73e86a2999ee04b34013ed1ffaffc120c30aa55b2ab4e0bb27251b930ed80a618911d21c2fb5cd9917ba8075a03abd0f0c69b5886f9ce141cfcf8c37ea9e8f161587170d9a48ef7edd6d0a0ae99a03557bd51401d73a27d8eccdb9661a759fe1134af691453e704f7b0242b384e0920293b47d90e80ee5623a17bc1ab816956a22e8ef90f9d94747137f86ba097b763408d14c81ee30a638fdbc7cc6d9dc978c47d97d9af8d59c85c5114672a110128641e8a2e8ea7a35c53e2242b4ad3b5941b543b1813ce9c92547900e2d20b7d2a61633fc7908baf5909d10e8b9c12a0c129ce773eea3af4f2402bc56d53d7c783a311f9233cf33d159c16cc9ba7e0070adac2552ef593b28b0d83d5fa7cbee377987df5d310a9648a0774a8dd5d4410d95a6488317dc9d70c44af896c9c9a0ae17fdb23a35bd44fe1c63323d70c05b7cc4187e9be734af3c94a1789f0be3b339cfc11aaa7f7884e780c99e56ba423e54ce153096a3184abea3d8eb35faa4fa214313c7bbe427bbc58608dd8337bc834ded3d0f99d8e8d1ace654457e8a2c467b9268e8a5ae879b2226ae35df7f902d80984cb0388b4b4a57ff78ea67899aab7e6e55cb38c4f8d02ebe3434f9d6c60e3d8be33668590ab7da3165750dc53341aa2facf8d78b13ab09b3aaa8709ea781a38746d40ed5ce35986fac588788d3b8917883da50cc120a6796ffd8803aca43e533b218cdb36c2f374a5fd3b52bf99f6addc5790496fd89fbce5f3ed11438dfb7c1d7adf8c2c305b61011d2108065e84d757219a89c4c89b9a686380da9eff984d7386f47af3b8e40449a84cca7a5de93e479ee54d89e5b7dbf7e097b445d2d1511253a38c903b5758e769a0e1ab8fd8d1ffde4ce7b4662320b3dad94b3bd9f0df9b3906dde1f8806cfbeef891d599572a16943a1d4072ac723bac1bb4c20261c4f7b55f5030c389fdd3ae3103400765bbda8d58db0586424bd62c99ca3fcea228ee1a3cabdc6a4d985c08c7907cc36cd1c5036a2c8327cd44fa4e42556f9f092a331ec3306507059310c0b567353f5c93ea8a3a71c219c43d1c83e89f0285940d0e3673bccaedc2ae82c05388ef1ddf7427bc566b7f0df4593a66c24a54b3786bdb996a6ace40af966b2b04c6ba6e632cb75ce4f297348269c79b91e31fe978fc9d241b10aa5986ace9c9d387e87ce3453de16ff2dfcdec8a452145745b8a6b83108d1f925e1aff291e2ad4b0d614248c7f2297dede0227a4980e5eb164bdb6437098e1857b8068edd33de471ecfde6e662c8e5f0b2d9aa661e2a37a83cfc7cf361a967e33e5a5025db04d4a2c7dd6c13cb95e00060050a568024a30a4482555c5a8753c67a3297699aee3ad4cdddcdbc86f2005a8f925ba1fcb25703286cd0c4571595ae2d047cf20cc6ea38bc645b5198f2ed4885cd83de7a00d6e4e255953bb702bad4ead376e59deb163bc719f7aae56ac17195f51ff60528fbd3e099577336c9dcbfe2f48d0eae2685de7d9817ecb10fda1a56144a213edf1d7255eb2d72254b25d8ee1bce1c2e94d8ddfdbdd656b7c8afe730116fd0f670045a0f254b2ea318a40aeb5a2cb1c7891dadfff6b478f58138058f2f22b2c96912feb807530b2fbeb43c85173c4bbd9574c6257a427fb9b1b47248cf76dd3ddb7b3c108d764d9e94735eaa1fd5422461bbcee1fc1a0be55ad64763dbb4c6808ab6321a07bc9e037f3ac1fe6b327efe557f1d0694df69f02f0b4f15dd174c88fa57b155c7e714f727aa587f8cb735b8b03cd465e15084ecb8bde192f8d899b800a64b9a1691b148e5bf31855f6f2f9ba65cae20189e3f9784508d2996df7d8bd9648f0992ceeb2eb5665393c643d75afe278287838953d8e0e27871c6e8b2bc95d438cc7e488f48842279d4a48386eb0ed04f8f952a41bca904aafe9645a78580aede3f5287023dcbe12d09b5ffa728c3a1186f897f09db646224870214dc8c59d2bab1cd52e515b770af7a47db3b3d267857a1c16536a16e692fd1732f5e7143877ca2ec510a9a55d90e1c28ccaecc71f639fffb2411c84ba5a3cf7335f23fb736e2d4e932a085e5b7505f75ba4c8b76dd4221faa7c23d12c6f619097cff9eb6cad0667f0392350f1cd77107c5542d6b24267e4a9743c2475d31eeda4ecc6c6d023391fb619989f28412eebcf7da6a4004e0b649e6888ca538b2d543dc33b42c75da58921a2d822c0b6c4d0abeedad1fa1b6789dfdf43388365f62943c40df9130a60cb292fc69e1a6392a41b2548c1e217eee1a5101f7ae34e0c74f63d0979524a6d4d89ab5357d544c933e9bbc3630d63f8aa75dfe3c2a7e3d76d386c52b8ef367901ae3ceef80d7bc0fc8ec0e242d8bb6e428b49f45f70292747e3323e8a7d5804c195a2fcbed540b3d7795f0cae169bbabf78ca27233fcd7dce103e8152e065992d5289135308f7fe611547b2973d2425d7b564327b6726669f4033aa5ec82cb94d60ef5c5eec4a96cbd40998b76088891d4c754bceb8c654b0b7e03124afd66a9c1603948c1e638390fd8ee93dc88935c76127e1cc9e2d03497d0d0af38fd8ef3348b91867834a73155bb9034b2433b33706de51776c6716d0a308a38837381bcfd1f08ab1c8938ba83576c88db6dbb641eb224107695be6047b2bd783a16d795ede3a4244d955d2fca277dcd287f2455febc5a7206185e74314352d80f0a1ab0e4f223dee19ee66d60a332b17c029997ebbb212c98f9e634cb17b769ff44dbe8b4a22dae3d6f18c6872ac56c4384376a278bd2c672b860896e5d39f7def77aa487a96ce74d2ecb77411bd30e0ad28cedfc74a26367f60ce31ce21d4d6e7410bf4f7de6ca06421aeec6187bd4dd158de4f2e3eb9a076c44c5b6e4f5f1eff0cf6f77f51f4d4a964e3523e2bc4f4e18715d7dfbd2d812f9994cadc71fc20e77e26b40f32355a630142af119878432af8aae5a8e178afff1d3f62bf8640fd201e6e6b793302260b4177d0366d69f3f2bb8b39e6d50d5f4508fb7bdb132f2144778eb6dfba3522bc4704a4f41764c3ed94e7c9fadf74cdfd5d9ce3e1042f414b7ae6715cd0f29a9a2105d3f853396a7651ff3cd4d9b64ecff3ca965b29297cf90ee7ae2b570cebd59c98b43ff141eb7d813d94fcc82366b0d700a82a496eb45457c758a06079392fac26688b9f169c1d69c330c98e60ff2d21f1cba58f5b28dbf436ebee47f2770ccde2256daee5f52a6572052904efb85fe9053e77bfa0b61099cf3ae0a123467f4f18c9de96d8f840145c2a3ff51ca907311c827a2afef9a875c8043af953c636c0b767a2e5613f6e29ea0fbd9b29da0f2e5d8282aebe6ee767dceb636b517de4f6ba5fa9ffe0cc06692c34b617076a40cb6cf25f00e9c248d471542296040c23650eec1344beb51d9ac5344de40a3a3d98c8d03aef7a8b5504fcab3c83d38a5b4cefec5fc459bdef5ed40715318e394c6bdd9da1721b8acd3fcffec6a3837f6e6ceb11be6396078bd6d8a9f3e06fd8c1777989bac8280743eab53ce9763986684a6564c53f897a761ea6e2e35576792fb6d0a6e34848e24c47af08c2ff93b8a2b4210e018089c5cdb370c011924642762965f5950c6e24364439d99476e42b18e5747da70a97c643ebd8db67b5eb1f9e3a54891da7d3346106a24710f2437b74eb544c03ced47d44bb97c71964c9156cdd939632fea34bd5a43d551901632e2c70c776d1b0f225b9cd91b5fa91a1fd6bf9aacff267d6038b5806ee174b3858a41e5aab3e516a86a88fc72e86a24cb6f49b2846c1efa1aaad9157c934d36c07e887c90747190d68aeeb1f1b8b5006d1a86ef469c6f3690cff73100bbab150020f109ef116634562f7ef3e8b61f84a7ee215995710da528ea987f97a1b1a0a3ada9e1571c89ee8d2328ce03e67dc9ca4627ce28e60ddeebfa7f886259c2f1dd2f2da2d5a460f52ac00d8ef0820fb8d10e65797b66699772999056ad7373cf3b7ace37856ad278046adc81498b2235642b1e3d9c8cc02f422a57611679829e1988c4f4d8543172999884b62e66ba3bdf3d6317025c5f31c18eddd2dafd251bc73c586cd48f948229692500a95298702d755609aee988ccce428bd87f93a999553b6bdce4447be9d47088ca4a915972a06772f62c33189a8a6704b09612061274d278aa823d57c5e425fc4bd617ac4eb87c4c48b976fbf2f5e59567610087c04f1c30b6f17babe745776c5fe0a9b016077ec7ba98582b7a3a577711c0b6cc9cf109e84f50936715a14ec1370c7bc1af4e60b39c7f98380cfe8ce3aa43cb9333774cf83e412bf7b2694bd5cc8278a707de863d3987b702319464d74968254390a64523a14d7b0662864c12c868a6d82a35b0008e526a4d9532ce99950a7dbae523bef945fda2308b21518f783f5d7e9e1511c6c62c6dcb614b031ce142d725d10574bf66c67dc95350ee8dfbbc329c007b0c1b568527cad85db921671a31c038db427708b0fe464f96a69b5a7aaedcdacee3ff99709d6e3630faee5ca794f309b72f854e8cd1965bbb2a0d0b3cc78b96bc9569d71698524532ba4ea4d3e0d1102de0e9c31518abec215872bc7ffc841ea64322da5ad93a473fa042cfbb6b94147e894e4891d1ba9ebb3f0caba73bf17aee35af8ac0791691ac542bed0076b8f766b6112a326f729e96302a0fcfa2ef79db7e9eeb092c5e57c0ccbbc22fa168c36a67c007531610e6bc7fd21cd6a6aa82e2fc53aae5720eecd99c3d4a235cfb2235f0239001b167df980a8dcad5791a4806ce582790559c861e7d3c3bff03007cc0698515b836c761c902f76621950577d88f6b6da2f5d56f7febb662d6efaf4c27a0037fa46072b29824eb0eb1c24ea2479ecc5313dc21091a43492b5b2a99aa1283afe5d3f98bbdc8ac0f13456e966b77f20748e754a9948bcb167a56a9e2abab5532f457b470160dee1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h3a52b4651276f65c9b9288cb978ca7227e00895a9118de9071e127376bf915b4aa1f0372db78bc56598d551f6d8f714d5c1728e0de1586ae4e365a871e1b537f221763794fb4fcf0c314b17cf2f85229ef5c5da62521f3e0167375ba37d0295a31edbb960327e94b444790bbfafa082382ff37a4cb7aa7681cbf6273b546d31bfb9d000ab57c17bdc14d7e822bff0188881fa7e855dd193af77d2fd3abe74ef06ad9f62dda804cce5d838f580391df8e1e1a766b98aaefbd84f93309c4c986657d73abcec3276cc80e7dc2105cca0697f9bcb3cc843b305bea8fc41589e84ba3f99ca61f419ce0814e0c8d69648fbb4987707c589ebcebe37495e614967a316c262dafce2f207d0dc7669dcbea3f108857076c6f2685c42d2d306c0d50da1fa9cab6df815f1daf51ebb696238acc6ec1fc26c11538e2bce04b85280c8120aff0239adcb32caf65bafaadca31d178f66a32a9913f36e337f795978b83e57e0a9bf305ae1de5b0376142cefd4607c177677f215f04b19372fb8bb78a7aab8b9e842d8e34d3be73c7a5166aa2e563bc102eb6d3ead00861b150eaa4415f2cca298caf32e297032c6ecb1a89fd6610c3547321e6fe573393723babbc6be894adf48117ec9c13d01d186a423fdcd0b27c5f5bd1c29b8eaf90a6a9e57ac537f1ac5b704de0813f6953c36b5e714c998bf3d9a5e6119a764a728cfb4e6c9d6829528ac3e46383f417d43f3334987096ed3c7e98d798d689efe8922ee7df5dd32c740c532b029e07852ef72b44ee0002eaa9a502f92d77375b2e708be06d325fc5c8857969cf3734a500030a5371b70f562f0f505f797b16129ccfce8002257bf4d3004b8debed0d33cbb958b4362649f2781ca1d3225194761146a55181e10a30219eb1d6325b32a0fafafba93c672aaedb726eb75dc3f912f404cf628c6343d01841b90b5fc6d0a14966f399bd410e851adb4331de310080eda1b1add17b4517b59c57563d284e49b26992ca8dfeb617a5c6be1a01a34f958e8c8587caf63f6171c79c16b8d4398861a009279d27e2bcd705ee85f33837900d1e05d8638f730a8ebd00ff9206073b8dff78ec880fdf5596edbea12ce3710689adea0a0bb2ba37fb4ca21d0cce3f72cf6039d4711c6aaeadca68ca2d68fb26c0f4ca12f63828eb6519e5f56e8bcaba1722bc4afde0e6ef0fe0cebdb024189d01f4879b4ed138f4c378a91abb0fe297829c46fd365c93709f722b7d127f9432e8febbe984c3b3b81f62e3aa9f07414f09f4fedd8b723df1255b32ed15f8fe012f26c508e15540e48faf67e6ef5de74107a27efd84a2feb65e48ccfdf2985e75dbd9713488fa41d86e9f0f59cd43212b9d671a11f48a1e6d38d6f473e266d3b978a686f798096bc04db4d92623336adf45e712ce49d4fd056ef931f39295c92e54b973c5d2b5a7e6a5752720320bb335772b61fc9cf33a802f90202f3c42d25fab000f6ec74c6f37e89ad9cca8f107e5193f6a0d7e92da3483a672d19d352cad48a21a8e1b520920a337a39f6f922638114c158e0b5ca1e875940388928196155197fae9e0732f622955d99844105b1de5dd72fb4cb2d1240f4973464a846a25dcd1ecd49810ad54d138fbafd8d3086d155e90f2ba152649f043454b470e8f63b6a9ef56d7fcae0a28168a4bf724ed0d548b3bd41b4899f89eeaa12f95aed625af88213e47d5ee51cb6f727e664e3a90d33dfc2a3e31f51af3be533e22b95c5d3599862ac1a4f148f3474d7ab6dab944f62afac8065bd177198c13ce7a308c892264aaf37f01d52ef302403f58f012c0da129030f4dd60f651d98d73a756c522568abe47e83cf08051c64d87b12e236d0fbf99b0f8b01174715ca315ee5af5ddb4eed3b988f4f4cee01e614ae335fc017e1179c1536f5ad76f0af25c715363695ae1b1f1f07e445ad7ad427cd349545982fc5bd97fd6350112fccab25f38eb14a710168245126c51bf1fe50c047e78fe96d1cd5c986ca0c75c64d5ad71dcd6ff7e728aac5869dacb5df19756c39679651a784d91d2fea97de4c709c91e9c679159c8280d600d90c59cc3f963036a3a0199897968c33488ffc115dd574b1abeb4b5c166c0e8b83f800a7f6bff40cd13f8a2acd505b074cdd0186e514e7e9f892a48775903ab7a9d9219269cac6174389c84744114f74f01b4544b3cfc35afb57af157134222e529f082f2ee855ca2ae4c16a4df5ee849852779b1f08adb2622c269eaca60554fa74209128747b46997c0523d072a1dd8238d4280661471810df7e09a88cdde4b87e435a62f132d29cd1e037e4e19fe9cb894c9c119431f12c7b73462dde13fb963d74354b8b1a95079da3d6dd712b298fb1bf635e260775dbf53e33d169409f2b78c5640a56e543967253f65f241281491be131624b5af0f29d603e1d2220eff892806d9c36b72b24dfdc2bb58b1d46137ece8bb8ebf80d74e497e1d4e8604f08f5b336e1e93b36059e3c571421e6cbeeb6bfd1241a866473f203ee93b0a722cd16598972bf37e234a93edf381f9c086e45e238e60e4ec4987ca79322c12390354297f0530144cec04957b6219842d48ea51a40243d0b3917c9c43fffd0a49699d96d0ec1b6ffd9ce39d581b8ecfd2096fc5811d100b2ddfd7ce8b5d2ed135700a4de0f42069f0cacdea77278cf0aac198db481e5a4f78bcf209db5537f9d2650cb55827f921a7a8a3024a79580c45babb10de63b399fedc039bc0c8d17af4cf030c3adca7ddedb8eb896b563163289ef050fcd853c077384de6ab6e9d540f11105582c3ae0c4f920e023ed46924ffea6d2ea07e0467494efdce7b287d2a700ce4bdcee73e4321b4a074222bc936ed45153407e8c4a73ba4fba5593319f17583e48be693d94e8916ee9a6c2cac4fa16d59a6561e1c4284787179c464a691b0259a691beaa94479a2c5c6bf50b1adea2e21935aa2ec34c6a827edc6c8d093740cc4613a988aaeef81033306921a041d7c43cfdebd99069eff38203eb92c1a3ebe707a2e85a972d668cfcda5e947a1974c037d6bdf4f2ac5f09fe4891be7cc64bd1041b9988d7a5c9dda4299bb1c1ef12096e27bdbf1fdac5e9221c83a6ab47451135afc7d98b90afcc2c117da73dd81a03292473d8e4ca301f6b5b0f9d135f3084891a92ca434dd855f696fca07d064c0f1f0f180890f760d3e0ecb54a2dc3cacb132fdb3b4244aa3af2deff96c3d4b930c89bede692162094eb1dd81d01eda4edaff3b8a5358072ab8a90fb7157a2c9b8f9860b5995975d255492ce38d2bb53dadd716389816d43dd2dcf68a1c4d744b190cebdec06d829765a8d5cad2d11218056afbecddecd9927712ec8818a2d0ce6a6448473b5f3b2f24b615c9d2ac4cc510fde0e7cfc6db75695c59e99c35a843d4071db91e6e3984ff0873cab39c73ee1fa0b72777556e2d5b5b7e90f9c280192d1f27bdf5208c26b22c28c7a1821fcc7e9f7c33245fcf9ea3ddc7d2410ca21762d92ff7690aef365e8095d4adea05aa4764b528b8ccb82bda94ab15e929a4fb0851408f6c3db5b879697a1b2c336b78f1f6880efe8099b2e01f67f2aeebc7c9ea13903b15c749002063a02206e5c11644b89e43b86dfb03931448f6d09fce8946547a887b050bcbd63ecd2ff8f2f3fabf4dc08f7e6553d098451a3f5fc7987c69fe93fa1ca4aeefab53c0f2b1e2568fba9a33f9810599fe8baf3bcab59c1fd44602a2edb19bafdaaa98dc2e773cac0f203e7cc98c6d8a4c28d87107ef15165a1dd983ab3ebfe0bdadea92b8e819d5e61cd0e7ea32257aa6aac2983765bfe10f8ed8dc24c45c04c23f6e3c6b7460f3888a0c7bbb0e883191a2b72450aac7bb5faddd0b7fc71d49bfa4c782cf3bd4ea35ce68c38c49e0c7959557535c66717ae1f47a246f548ec94c8a0b2377179a51a987917efd8af5734484d1e18c631238c20674930f9dc2106ee070bb98f6abbce278b6b84e5b5edb663c916762e890960dcf18f577f5c05117a2f9f0d6acce17f4beecf4b42fb0a9ce86fc3bfa2069e094c38db4818cfd8ec5c6ddacf11af8044ff60ec4fef05509c0e94cab6a91cd4233c625f8f204aaf033201a1f90dfac662428f170ae067cfaf6222a1434717f575b7f4568b6266dd9d0d20f1402876be9a73302a30cabbb0d8ff42115bc26712487b16115dac5734b0309e0a6468d18949ad41f4c9341df8f6ee4b6a68b5cf98a6eb84f9658062364b777ca5ae8211f9203d5a4e27f76dcf486b6236c08904f0286f67764f6871ffaca45e9a7f8a5627cd32b245aa3f98c509394d93e6cd274643ccaa551bc902eb7fbca2490b700463274f989e125bfccf05bf10d37676e7b268266a7b10c3c8ad6fbe12a47a71cac2f03a40a4469c282e188528116c65b761d820488a7cd377ed3f52436314b98712dacc0ed0e39ec5402687be9679a5f9c5b86e46a69d8c884684e1f7898dfc0f190eb64801312c49bb4038765fab10fe8de31cb75981103517474aeefe7c0ae76f9f210ae39656005daf63a996a1111aaa21d74cc234cc164a4937bf775e2db3f6f6547fd2d8f20528ae693e00508b91ed440c9f8926de3af6b55e3e31f4fa17658aa7ea033a666c50de031a04081b70b5436093ddbd4e3b1b18b99c4ed89b047d7fae891b47e47506f0219b0c1f6f902ce64a080b2e25b20fec8e9c6621af139ffcb906ff8d6b41fc9fddcbac8ffb0b494baa237932bbb06235d6c6cc85c91cc40c0d1a5ced816016a4a49f9a8b2ad32fd2eaf370aaa6a6359537f19baf33e3e3cf47c7e037d1d8acf8d320ddb82bf4a98f265c6361b362d1f8d754aea89c47f56a20d56f483d054e2d0e6cf3fa838538d3bd97abccab553d209c27cd8d05392506b99ab1d991179d11e37b8a6e765d1203d202934a0b8df2b0d8adae2fd017aa294d9ea3f17483ac09a6e3e4b454ff41b69a3ceb7f628245d665cf3895fd0e7e5f330ac2258ff4417e9856a730576fc16edae3a4993fad6fa97c6c1a84681d15c8f65f03ce18d42c474c81bfd391a2b0af653bf4ce2ca1979846655e3b6aa1061e42b8c5f72b525ba1912e08431a184de70e84bb1dd017786b2ec44551fab85f7309462eed7b6c0a6a4d461449e593c4db981df60a6684e9a981b7f80f8988f099cacf29b51c91a61be8141950ec82b0ee05d4c4dfb7168024633ee01aa8a16bd9f0a257543097d5c3da771b13a1068889b0fb30f773ef955f823d3617e0287b86de755e9e3e0e23d25a0d23a9a2f8e3d50bc6189d29de027fc6b33d56cb9a78dbbde626e91997fbbf5bd109e030d0755857e32f0094deb379a9335d990970f85ef5e049c13f03f325272c67e55875689b68c1aefacbe03768a8b0200d5eb40e91abed71fabf5d7ca3ae94535717aa89ea8b0178aeb6280d051194380cff565891a00405235e5229476ae12d96d183e41553f6f699db301999bc164c1d26e63907eb6ca4e67cdb77d52857ddccdedc400dbd73cde4e67;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h694c5e27bf3b34de0c2d0441b4de6a419e67be6d4cb072c0ef8604daf44dc7afe300e889a215699289d0ef82ef5fdbe293753ca516e8c4f3fb7e4863a193e5c97d1734713e554dc5b3f00c7febf7d5226c30f112a18aa4c2db4b0f9f497cb28c0bab7a953be6976253fb960d405e85c4d7c2aabe0fb4c45075b48d7de3d8542b8ea41de06d96b1689f3db99bd2bb68503a8866d52096161d7ad1feb270d8128f709fc8d055d8a97ff831f752cd7b6172cee33e1f32aebf54d9b425824909dc35789af3065f936b10e53ebdb8be1f3e783ecb3b9303e080591a0a5ad3be00dc986b664cf05b2d7746e48cb1ad51901ae4fd01e4b72460e3bffbde457a71843ded79f03ecb8b0388cc062df06ea278a0f76db3874824d2010eee2f90ee24f7cf8cd15a3a2dda38d91b096d68a9a2bfff217a9ff98118e0d06e187bb00ae9d95d9d39813932fef73caaf830f075f43f3cac47d4fdcc3f18e5ff90dff84f1dedd37e40a3ed42bfb56a35d5bc1889dc171f602a9cd79556f3a31c78fec0845ca69afca32d8a4c03ca4d6cf49baeb2789b0e656c1a251f51612713a0221e6185fd8987e580a294ccd9560ebca6396a1c1c32164661d25f8862864f27047936f74492064dd4f67bd00ce6bb585e2aff9d2209c6482aed964422987773bd4cba6b88f12d0067884cb02758054a44211c15796abae5068eed45ac2bbfaf64345138d07164639ede90c93c49cb01f5d8a6404561fa38a43b6d787634abfe360854f07c08db70fd39a634be3f1b98bb9e603c7be37622521f02cc31c5a6fa1099cd304f55146f26be0288581b176edfa347c920b6fce8495a6de8bf018431ddd5c4fa6e14ca38e1fdd5aea4efc3aea6f16602e3ab5baa4de06c38136a0b7aba4d6608765eb0bc10d89651cae71f8c80cdae4a456bb71a181507ece24e2773b8ab39130d362a7af5f7cf93d1c3bb1eaeee65db9ebbbc4b4a75348c454c56831d5c58719a175517a14d551e2f65311e1970b6bc32c228398414bd93f99d30bfd207edeb41c62d60cd99c44d0ce1fea12401343e53f33f4927809442577f2d82be5ead231e1f0271bf22dffc1d4a2d74823018a0c17714c498da204ce0f86534e272bb8bc8286cc988d7117bcb819679fbb7460cfac8a0b1f6aa8d281e513ce0637044694e6cc51fa44d267a4d391ddbd50cb1c51079505fe5977ff06358999deab24ec5d47dab0fbb9c9cc58e7a4001d06532b4bcf28248ef50a9e128119a02709837a6b1bad888497ffb22c4e6065ea50a30a40a5da05aff2d6b6eb8f152f59cdc141d97a2fab04cc4c4fcfae10cb52bc7c215b7dce33f5aace1bd9ef6f0ff7fc213325773629e0a6bf77f3a2245b3a92a1079c682f52802107bbb2f2b931e1a0a574191cb81505f01c268ec4ae98ed3d1c1229a53e3bd234bef484b49225917059c2e2e1c4faa7707049b280d81f14386c56fe9ab1d5d26ee1e4fbc72fa07fc8d673255d4c518bc1def354539643664d6b93fd5ed69089c5e3cae30e68b80ca09fb375c71621aeb08112af0f00297eddd6af8c822e1f1a9d45ae4c7087ea1efbe297cc25f660edbaca618a4122bd9045fd7797b75951f2f6de41ca9f5f68f3f8ea9d3dd258d51dbed8a529894ec3fcd523c54a049bf4e367230d8f95444ae9cc741f8fd05fd0db52eb3b0186c605ffcc167984a5c8328500026d34d7f1e4ce10eb871fbe759c342788f92d7d0b986b2a19d8b63dc6771224b2aca8d6ee4cfb91134caabbe33ed99b442cfa8df06163e70f20be0e4c41014ad683dc8b40a2324a9f8318a2995f8eff36105f44ccb0de700983a8a0a937183638992c9243b22f03b50d2519e092a636fb549cdbf34a3b03e0ded9141624ec39be12414d440a5ec6b190aff4dcb116543a99871ec0a8d8591d0fbb64fa3fbcedec0f2ee54758c699b23a3dd8e2ee1a4ed7c47e86b2453a9ed74fb489857259643ef34ae0937dbacdb151bacbb4949db0e6f052d8373217bbf45da24c84e96ec2f955559ced75f93827e56929776928564443f11eea68798fd299d60106599f31d35a8acde28845a4a8d04bb75fb16e75eb32e534ee864bc8152d85abf14c3f81f4666c63694ac180f9ebeb00c97c24d674acd20dfdb348ab53be010e7630af0dccf70652dca93ccdec5857333c6105ecbb6f0e97383120ef53e8e3b4408619799530616ed6c31b65006bebe9f449a092d4a775ac6b421a7f74176a28e450d5da9cff3abf4134a18e2d6ba0fb1c4e1aa4ff2fef9e615939f3ff08def1a4ad927f8d9b9f3c3c9409a508ef8a6e5138cbd6c3941ce668cfa81f04421c8bc0977c35416b5a27594bfb3b4385e764ac3bf9a3776e2819dc7662f30be37ffe0df6e7fb8752f1e97d77768b344345e5ca38aa45efde726c267b1dfe6aceab64c58dd80c12a3064a0ad0308d3da68ed068f5e7c3d842b9a025173763c4be579dc0561b05e838317fa06e3f185beab001ad0227ab691ca28817ff677bd710ccfd925f5a205d07ca27a5d2e17a114b4f821d7bd88f87fa9de934bcc9b6fd57e4ee1d3436d32d108d40953f57a6442ec9ebb9d92933fa5ad4c5ffe4d0fe163dea59f80fccce9be5371139b0a56ef42972ea62841ed358b2b53442b0af53bf4ba0c27f6c517fcf6231e7dd2c4022f909c8f34ab4d44ef2c2ebdf63f2e0345b27345d15f4e26f3e3ea4427df420abd00913b98502688fbadf08c28292857ae4c0405a61353443d5d69989a91878b975ecff18ca426c27ba403ffb196ce357b8b91e305c03c7ed8a66a0acae07e66b3a6e1140a70f317c0b4c76b614f647f431ba59bfd3bd0a0f761f91ad9dd26c0638c2a927ba421c2c630279873334536ed0f8cd3c0c3c27c9f1e47a7cacb4d92e814570a097c8607823f97d9c66ae7cd3e4c09410cb9ed98983dce2366f4c418b8e99cc65ad27b43a6909b6e59df7440ce617909beee2e40967932816c3c3c7c8557c1a7d5583651f7d26df8add77066195a468db1a87eb2955492d87aaebe9e0f26f99650e17f408ebaddca6fad1d4e0bce89ebe0ea57630298313fca463d32c51c592e1578ece1ddd72dc469adf602b4c3b4f11e202ac95a513a41b8f8b304aadedb1fcf33001d035e900a969dc6c78cbc3458c822a5b65180a9ad19945d8f2c82942a310a50c9da0542d1f10320fdb7aef68a70ead9549da491d49c77329eefe98e22bd0fec75c540146afa29eb87e7b97b6bc9216be15d6233417ee9dc3e4091e9b742331e582c5a729e1452688506cbcda9034ea8415b17c5ef716231b81cf53094b28b99e85f90b902ae3fee7c82694381b7bc8e2f1dc94f5ef076dd3ea68065e0024deaa12ee194902232cde30689f17e656843cec7a68d049501925c3c3385dcc5edd3ba364222c1ad45d6b1e1224c091c3ce8c2bf6a6241e50b5bfafad8cbbefb2adef7038c4a7c2ba8f422838aed506140e5a616e1071bf19306f85bf1dfc6150b8761db22da799178868e485e65b5870684fb2564c9a83a81b8a5bb2a6feea8d6a75fcbcd274d603ec261fd92d24aa7443ad0c450e0f2103d343b7ef4edec6b74b718aa143cbfa5febcc86d416919bd4b3f3a4e24c1bd7612eb501ce850c7cb51f670264b1f541763c7429c5e63ac001db86bed71c5579af9f30c3b0ed8fb29591404a4eb8844b184b82e4b0cbac7b52446a7e5602c97a693b4c8aa30a226fc47d289ab847e004390347aac404f09d00d98ebb6d9c8584ae291a1965aefd9dfb2b50c9cf5e76d8bfb8cc2b5facd0cc367cbbf18c6a6792a3c6809f65cbb47beb6a696a3bf7a9bcdd6978e602bdeb42cc21dd269164469312e37e0d1f75eabed7de7068c0462cfdd04fbcaf82d776581c391a8d95d69c8cd6e429348b04c63a84b03bba68c28c0559c3495ac28cd0cfd9c1faaaca3f43a0b9a877dcb9e49fd72b8cf77db12d7eecc0475e38364ccebe9aa619dad759954bae434fd180a43be89a7683e4364d9d24b1b1b17da245d8e76a2cc0d032ac39ec1cf962c7ce9a0632fa7f0f7d4d68d14f76af9d01f4e047ad2060d060e340ac9ada8add7079c5769ea3714c7f14d36ded19ebc7843400dc3aa78e702f70c6bc106ac9d33c2ff52e6464ec2cd03613427990508a17cdd985c6fe33eadeb644f4b0791c38468ac7e917724e6dd3433c666bb5438f673c10cc9132adae187fe48444c8609d2f7d6bf9dc1d5dff3ab626f7065fe13427976d04a2a0eb556294e21c783117f2e274e8fb3819fcc6919dc2ea1340ff119052523fc9641b3542bf29e22d2eda4d011312e9ded7d1916edbf8b51105dfa322179a5602c5ff7d9c6b64b80049983b9d89b4e500387a7983d152110157c405d784f8c55868ed835ff7b64ce537381854cf1dd98e472b864832b3a5ca3bc157994e70c5a314e1852985b4985b89030c54611d7b06656b4141232d0fed3703e5e8c0de48476e67120b2672d60e3b34136a95d8840cc2e369ec5099ca8d6c552110681799cadb7cb10587a7ded6513d1ad5730c247381bab2b589ef9a269f01729d6d243577198eae10f0805893d3c736ce1e95795956f8596efc03d1b8ed6687a2f6188c2dd25eeb2fd7d99ef7130d5a1db1a563641be7436139e81f209be7dca2515b01888f07811b997cba6f0211348264b932f81c740f8e8627e269c10c811e21b876755515c03b653bd9ba62226c3c622bedfe09f524a37d13027ce86dfa58fc4151e9578f26d03062f8764f163e6d10f28ace06257518a703926bd2f842ef3731ae4614fa7e99d605abe4600db64c9454bf37c2fc63cf2e6b4cf185f4d9af21adaad2a77e9aba011604c8a3d12aa9055178c7e1fa1e20206e3e8cbf6e67a882c1ec8961a8c0138ce55bbc00812a9504464fff02cc167e8a83727e2857d990b4ec9d8529039375d861eef26b8e4142239b1bb47591d4ebd30a1322e297297b22becedb34993deae9af30703f595e83853f1dc41721ded22672fc41d35b9e99adfe3835ced068bc5b31fb20d8fe3d34ad983254fabd1fc18743bde5af205f0bfbb542ae3d7066c11f61a89cf88adf2571e21e34f156b421a3e65034ec6054de41f812722a8f2062a8ca459f399e9dd525f8b96d82b80035406c68087db5bea6f9fadfed7dc8a4ee257fad659c05ab47aa643760c653c17bbb54aa9535e93ce95103afa6c83d87bb8eb92508243b189ce04683f72eb033bb05145df7d7fde818f9393ee1aee7fc777668568bd1bb01fb0cf2848e928a3ae25035e1d0254f1b1ba10ca5aa35aa0131b5ef9064bca088b02abace00050ce4c0f59d56323b061cc28abbf1b217ab4d4859a3f1de19c43c29a8b23bcd5702f1983fef1a55efa1cf44af33106fae9e1f8ef5f8677d07bdf6888fadfcbee41281a68c0ba107eb86f59988a4807fb225de8439e637c6de7ecf5bb768e75ed7f8e4fe04ebc20096e28b64dbf335b22ad2d5656e11a1c82128e14d506f327b006cf2609c0e6030d4f3963376ec3728574;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'he2bf6deab1b12dba9d0d0a47b3cf41663264b2650feb179d14ab3d68598fd35a42a686603e7f0da76f47db51e09fd909e1b393a75ecd2cb578ead9f51e80eab5bb7e5093dd2b8e1868dc7464c92f0c7d5993d83c80fe34cfd75d5baf4f68ecf001b7c5dc7da8b3e536e452b8e2eaf140e58d5ecbbb1b36890d2a64822c03d8acccda019cf10b17c3e8368086c895d592034fefb8876810d43bf553dccbb1f6f1abd18fc8336f520fdd4927357eb2ac099fcb391555a033d0940de02c6d942f947c3aa7952fa0452e4e425941df7bdb9084f5455cfbccbec2e7945fe5e83063ef841571726da6f405ff67c0207f19055327c2d3e881092414858080e3b9f4f923832cdf19c02e29d846357fdc36083be80739a63626b32b74df5f2c9a1767d671e0069c28fb43d822e19dd35e7e2e3619fda3842983c88f9923c825695868d6612bc21f15f01910b9ce0cf96fd1af0c556648678cd514504d4ab8a7e5323e06a329050a4b72c9535a3820dca1c6a5e75863b28e6b543878424e7da06162f21b453264c0bcf520ce60b90c1081f30d88173d73cbc46c5f933295f852f919af94163486c7fbf08f8d02a19e875dc364b9f4d2b64ffa8a105f69e5d9db462968d5ad3e00aa8b7d53257ff7147ba4fa9b6f824362ba24b2be35db8aa85a1a36d674158c3cbf5be0eba12324fa0e9e71455cc2f4a1092c39909b70314e6b23c29b69364a280cfa357db5db7fb51107b7fbc3d3368d4ca4f97b6e4773079bc1ac8b10f0b9f8db7d82ab2974f36f1d4758aeb04ef26166109afc30be9b2a6caba3c005eb752cc4994bf2599f1871b057adf6f314a1d3a3623b36bca1178fbbd72ee50cbeff6f91b0daeabfac7b361470932197186d12c22f4ed0d0803368b242f9c6bb6a1d97d16553fa6c9a01e662b0b50381deeb513874c7b3a59eed6eefbadc73ff635afe40614a723c21bce124c9eaf2562f715fbd0e5006aea8882673c7bcb128d2547d3d7ddadb54084618c8f4a0689640385e1d48185bdcfcba31508d6be00326130db729cc4fa74f193111f31bb4f8f2cada870cff1045e964a7271d720bb0ef1f17e77ab13d10a9e3d28c468885fd7e465c32bcb4a010844ad39ad0e3bf8fdf18097bc1ffee937085cb7c95807cc3d4b0bab62f1bffe0961886da2ad2d6a0f0ff7d290092a52acbbdfab901c2fbd6ffd868101c308fa6557ca230e3c6c6c270683b66cf516b14b890c1e4f9638fe6911d5a7ee351768cc8ffe9a68c3078186ba545d8185042e21f893e7fb7268ba040b321800913d98e88b82c96b75c86e71d741080c02564f9a597c37e56f62f23cca7934f8069b80170d75f28f39771d5c8222d40a8796bc16e1361bda240609a770c1854178ecdf671d9c402a21d4694b53584004af4bf0b32c768cba90ef16eb555c79259e703f4330df8defcd3b5e0ecff80e1d701744d4467c30c62a7098abd207b8e823c8e59c980d9328522cda11cb9f7ddaa45288023389bccf165508e0be6d3f57de319578b7083a6e5a05ab4af522a19512406851ae4de89db734e54c2ad076639f0262bf4b54b746e2d0bd568d74151136640ae3d96a1ffd63509635fd3a65134f9ce125d368fc8bcad3824ee56bf712a1c8dd492f121a421a8a030d3088299181676df629ff224b22430964a688cbb13eb54919e44e33f3bf14724d3086a0eb52e2675079a8cb1bbcaec37cda32908407ef46b38d4acc4a508c6e049f1891903434f91b2534322122e321ae264f2f7f80bbc53a5e7ec13bbe2ade6d5169163cb3337ba0db1e8c24f5aafcd3d84cd16925cba4435a889505fc27698c67ec0f285da92bb3e4f619a26ed645fb24a70afd6669ff58a6fbe9409c13c8029eca57c662270323d890558c2e6bf6dee0b3a272746e4495c829c8bf2f804d21fcbf44b50f54fd643ce93ade5f9c096e107ead2ec23585a5274ef0020c430208f6510925fe05b2f659ff0eb17b84fb8650ed7aed96e786524addc5256627b38524e8e9c9f9743adec48fec09be9a78768efce7b5f21253d391bb8e621e7308d19356ae163fa5f4bead2a6c2cb12a1be373f916d912fa062b805870d98e3ed69ad04d17a956a3713271b3b23eb608fa4d8ef7bb301a64ddfe3177b8e46a9d995686e956f2d85c1c237be111aebaec5f555949d9eb6fc790db06a37452f24ddd38bf928fd88697509fed8bd28d8a2d278245dbc882b678a631151857203d2071df42b748025778b6d24ebbbe5c386dec20db6da2f8d30688af1a624b024bcc3f7441f71e5bb5d63d97f0cc22d5833ab6ceadbb8dc8456d2753f1cd428308a9c7e788b30769e305ad40cb526e0aa97fb50fa7ab5bc67801c829f5016340694d09d894f4d5651e54c77cd5b9e4ca4dc5fe3379a2557788bc9ea9e52eaaa0b4cbe6d23c6704875bdb5b1387bbe8b1744fc7c6f473607b87feb684aaa0f1694c8e4acf1e28e2ecbb62a5b738d09e7f8d8ac24dc479020aa02d17b9256a1401111e46692e8c951a865bc0162e45f7bcce292b646ba54e801159030bac749e3d7efa0af2552fb974447fe08a830a1ab6fb17f518d08b1ff75b5f4774943dea3784b1f3bd0ade90e80057a6da38a1e6407d54def0e07c95aa027feb37ad0102fd5feeab50142750ae8221097438d5d7c0976023281c54210e2811f453e11eb4b587f91256450013b257d40bd446ff70e55e9c2e0598b34740163fb91889b1147f62ddbcebd2aba896b10ba1c513db44e698c97e52581cf333e84b913417b14b3d650496107e5461e92c3738dec90e57b3ea4acb3648d04c6049c517fca4917617c473d52b6955fab2530f61dd3e54e1f08496046a26adc9ce774b720147115a3c2358100aa24f286bb9a2367002bc06b12c5c14ecd178bbe7e642d794ea8ac07427193d24ef2a919bdacbdef8d00c4da2f30eaee2cde7b049c7f2446c6d46e867de3773886f5f09643db8588c845cbb20876714609346b000f8d9fd9571f982be9c8d36520a38dff59ae8a605245bff24dad197c569ba61c39d2455a6d95056d9f4259dc55ab3e329d6eed818e9a588b8dd81a1519f800b70f2bf4c91a0c7c325c82d8943cf06790f24b8186dbbd01be97715adf0801779cdfe1a85eb40d0a56d793b6e943668d6a6763d5d3f35b3e7ff598693a1d9ff73f3eb1a39f543a5ca170e3a4f98927706c4aef0c17fc5d3d77c34ef88393f5fe6d5295f65614ddd2bd76ec17b44bebd2ef5ef653928fbf83456ca33240b245ef33001edc212f3ecb8505e28146e92555dc9df6e7202b1995ba16d693c9c58efdae9458c149b9357fa05c68f694a39927ce63c90c42b0036ca4ea5478ef79b29223067a3de53e3808d4fc5096b3986984d11e137fade0a6ba16a867785ad0b55ab51cca2196525cbaa3d832dd8c98133139dc467984214a168305156b3dda201ac86fba59349dd5bd9fcdabbb9e1cddcb962364344f54cd873f8836a6eaa1973f3d706d27f205ae93d039614ce371f83131a0551fbc367b9533afbbcff43c4860b82510d330c0eeb85b6e1b805b60d382673423d1230985a464448dfadb71bf57dc7efdf11240700c8d857aad9106ab206d03379c479043ff30b30b6c2a0f4e366f18fb243bf8a4465d5a5ab215d4f78d364619f33424527fa4bfdce1de48583c62c0d77a8129e6cb0a51766a30db00c89750125c0035b62cf865ee774937c6be9186c7326b1d8c5aaa0da30065c9f01483a47e54ac970d4ec4c7e757dd81fdf582c6633daf0913c515a35d3d49726a41ccc4cd0691a8f20dad38c160385f4bf7cc13ee80a9f86d0703a50813bd131f9a5f90bfd2c6bdf44840baf9e54bbef8811a42bd76b8e0c29066a3e7ad2a1aaa79db2ba628ff6fd9db788ab9162e049c9749f37a1abe4843d05abc92cb8cddf194b0275a8217bfb4049ec59e3975d88b184c6f2d46702cb488b92534dea14a44176fc72166a0e48f783134da16a32dc43ef8b3bf4ab1c865779fb696908bc589369e47e44a1382a38800bba105e4286db528705371561d9f4df5c933ee07589a36fad60ac8c1ea418663e843e9c1944108b57853b649cf63052b07446ac16e1243e65dbe76d15b721f5fa2bdef0110a3c8cd3db2b07f08444a3f5d4cc33c8e1604b5897f6c58e30ade49f3ce98308c0bab64746313b3268e855cea1d88ea39695c8f0155807189ae2fbaee393825723313495299c05457dc63576936ef3bdeff1554a7c522c85d7b890d93859ee49e049ed657b4bbf203cd1520440373fa5192aa34419e6533f81beb29c05c6525a64d35bb832003a350478232ee2a2359a655be8d06a913beb4204bca44c824c09346c3d127fe3921cd5c44c61b145003ce1a8f23d66fd4cbfcf8105f29d1ece791b0854d9c95366faa731c492b832424d72d8db8bb18652cf4327f806c1c2bc5e08897f7e8e308b0160f36ed8da016bce4beab68d514ff4b1b79b2b84527bfbeaa2c1ee19e49913498d8fdeb436fd0fdb3162c853d2c4904d9edbdd4c96ea88a958b2e196a45958d5d6a070864e10405fffca6de290f9cb4f3d3d202c3d660396002e18a25d5e4e8a1ad18b4be5aea4ed531d9deb8942fb453ee7149402d8cb9e6e2d0aa7c17e6bab22d987a4d4ead76bd3ed24e0ea2dfc3b4e18d497225b045f2643bd1ca9faf120e0c625cff349e511722eff083ccd23c51f7665c6e8316c079d6480f86f4837e2cbead724e153c1d2c757313adcfc9903b0ff7378c61b40e39f528933bb9eb5f7333195c942c37362228c03732399bff36c737cdac5afe5db79686bfcab60a8f5d0a675dc0d9886457e7d117a973cd51621f32b32b620e41b7adfae0617f6fc97e46e0e3363db2ad8c77bed5f6e25035c5096394d276c3000118a94d29e10a4cb9ed484323e8a3b99a2a9cf1546be8132fcb0d494f20804c76fb6034a823d25bbb58bcc6ec21ce33f000e18dc7a7a5139364ffc0d87b1db22cbfd56a4de3dd29bf533248293fc416c9d8549e5bc81bc82c5a0dc469bc2be00f3510a903e036a4424080bb0278f83132556709c8b8fc129b33ff537e687825db232ee519a3840b77096a944f183bd4198fce4abacfeb19e33cc0e56a2bdb327698fd1f78cef095c211ef0396b5791a0caa7ad4e904d872108f842ff24f400e9d89c80e2d28459b157659fd5cc5598a98b110e5ad31db1ae7c2c848735509bc15b1ff3f050b646b9e11358bbdcc8bc4c42074f42b23a99928ea0491f28e8e561e52ea8a5647947c0a9aac7e1feb774c2cae940e553b4284ac8d2e20aaadb4ec636f4891e2e1f3a9170cfd67671cb59ede26d43daadfb9dd590047843a60e5b56f8a284ef8692784c587c2da69fa69eade88717b3fd250a9c7f705462e67ec1833b6ed7b69d3925d24aabea3047333814fffdb7a21f0c394cfef020d1e5795d576b829c4ff726b784e04d2e982ea39698ef47891f69fa3d5b863864ec76c4598b2181f225b191962c7296f1456e4e51e72;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'he37a72475c7f9813348a61eb7dd363ab7dcab2af9cf27785ac90a8fab35a6032130b5053fae95ff8961778aaef9a11d3a25880f311d0c423abcce242235d60cc43bfa9ab2d8b1a1975c7428f7e4b9df610d224dcde0e81bb3d9057edd421dd4dd769bc8249344e21b8fd918596a994893159d8c41df7bbff312bb3832d34f7f6855bc11ea65ff5f69715babdfc772077963200f92e5b96ba15a1f08c0f147bbc88b4ed88ff110b267335fda9be714f70a32aea36fa62687870bc1c331381aee7455f58a9215c54d012c0bead15a744cd0eba67c3e11c685a428a920a3eed7e100b242eda45f19cfada92d23ebb381b001c852a4ec2075f469d651aa7ff440acbe2597c9d1526bdbbeec74423d97b39a2c3356050b9bc1d2ce67f50ba03a1c9bfb23ce4bdfbfb7e29dc9693a9e3dc379970e33597630858fcf187e89786d34b1d16e108cdf97df7368dab81555f8cda3a3b0ba2c9580d8b3ddff23319f4ab1b6fc67dedc040b63556d95557f3f33c9a114dde0e010b100331e4e1eff1bf1dde42bf8ac68e5ddc7b8a8fb295766c984e721ed0be7d7446b36c57fc28f181e568f7c698595d88c7042e52314f2bd25ead68abdc91b778bc683c9341dcd068401b0d8e66e490f558af08ee195f83d2ed25d21c54aad311954034bdb2b73ab5ffb0cd914742c30e2e9afd45672d013c0ca4bc5f07070af425cb70cc55350162e2ae9921f34945364d3c54abea5d8337bb882ceb34c8d02e005cfd04d467ad85dcb796f6bd86cf9a239f436d5c5897e026d67b652eb08f7215a18bcba07d4f9f95562ddf708aefb191fdfc6d0ecef75e53936676e31a08d8ddd326f68743c825a1ee191a52949200d4b719172ed79c35ac2591d8f8903ad89cef4a140009b5e16830beb2e8b271b88bf326a444595cc3b980640d2ea8142d6f8d287494816a7d06e9f9506609dc66e70703225ec98367f7f31d40898a3929a3aba07bafc04b04d841ae0924c0ae2a799a4ce6f60f6302f31e255c593e8dcda05897920cb9d57b771163cde9500f73f522bb158c3ed16e4bdb0567ec43461931420d89a0248c82d89c4389f1ad6f6f345962d00f2df8a3a6ae90adb168d57f06f3ae83a28408429aad0170a80889a7893517c937a9b2cc03431af278a270a37996066846e625328a6a36ad7be3cd92f765b30f835152a1dc0cbdccb8e75bbefd22560cf2123b90780766f9c4823efd18380402524d6d49852f8a8583af16c24539496742df21a00701defaad11b918de976e0a98c814b4cf6a1ff2c0cbc37ebd2e4aa2c379b4fcc1d0e108690489c2cd94448b7df3c2b27698a91b687f43ede32c5b229d52e1f87711ed0af9f8f963f41f9a1d9760489a3bef80ff4efe0ea8cc38fc655bc7420ee67a5bb7ae1ee3b19e86f1b0910c3069b98acef568a4f5b7f04469e5a3964e78d6f06a77494966cca50058d672f47f97d72c6923364a3741e95bcf63966720e120b9e3e6a5baebf7bfcd68991e68850cc3d366e1a6a4e16c0ffdbb26e6b177cc3162c5cd072aaa4c3e7c664643cf063e25c403dd095098e0ebcd389b59edd45708068dfe1e940cedc503c67ba5c443bfbfb2b3dc5b7a6f4eeceb54871b461ff2777a4b4ead30405c1c78959ebfea683139501e092b7423ddf1e0523e632caeb8fff5c5b211df94b687facfb3c8963e8b35b02b4b7d21ecac1372d7b5f15697a9a1d971766a3628c669f785a00177c35244fbf575b07d976ee678ded4f5bbc1ad7da70140199e5637a7335f47ad7568389ebcc3ea9229fc5aa1840e51cd8cc1d46db816a8f446b8e5a8e3de72ca21f5fc5854935ffb1f8b539c25085145fbcbe8f64af86068ed8c4fc184b4a96196dc950df3120ba8a5fb036530de414e6ad414afa5c6ec425ef8a3b68b32667ba1eee2633b6c577c3ebf322ad06726e25ec1cd3bfa7f57a00613866bfa0d12a8400e207699fae79d5aabd41716e1015dad452699812083fca99e42950b5f347cb364cfab3183db662613bec8deeb200641e49f5da0920b7ba66e0be88b47751679a6f6da3f43b8243a0cd87d560f963458cc0f16fc8bf2a8b6c851179b7e23f3c5545294b58c8675eacd21430a2f4ed782112236d46ef1fa2aa180435a1d05e67180dbda9f460a0d23c7543515cf3744b62dfe3d46eecedc137c18e5a4a7e7da5b27eae2ec348b0bde6667955c158082982564f642b47f56e230876d7c74f4c7642b4b25a1c4245d3ed265307e17ed7ddc5255b37b513f445b8f55c4a83e2ba33ce483a860b50149be7d2b02dc24c2627ef86e8402464f8e4f169c9fc9752747e53fd597de8606e4ed315e24c1695aa5a4ca162e325e5f4f90124eefc4899944bae5c0eb8a14f8c3b4c4b73df1ddd9f3137cad6fcc7e2c8525612c6ba387f013a1dad029872207660f38552051210a73c9a294a3bf0b56c9e0682d72342bdff2b0cef50f2a90993ba8c8c6c6a5585dd3af5ee445005c23343270065b10d35980a42c713b383c85d6891054e02bede3ee99bac3f98bddd2b9b69a1fce515071ec8b396cadaa87238341a1041ad289f5aafd090e36843cc8ac37163870d64c6f6534578584c872c474718b744ce1ebdbb30ad28463baff88949fc51a0a4750158616ce214461edf080f9f6e1ca70ae5804ee82bf1f7a4d1b26b1c21fe72e7e82381d872ff755ebf70db93d0a7ca7d255bceeaa4623d9c9d7279d0b8ea9d4309f7fa6d67b090d9f4ab0b56fec6c0d183fd96018b6fbb2fce722a4804d74c9c0784f4e30f0b619381867fd68fbeb996e9ee50537c960cdf204a6683c05b610ea86d3fb816a1249bf82a525e70ea8fe8ef5834325c1dd9794641e4518e2adfb09b6ada027c87cbc0ba9bb8d358a9825ec4d28cd0498a7f66a9151f04fcdbd5da9d67ca1c2fb481801eee4d7e0c1c4a3f07a024562be6a0d91703e8e02e17be7f92c1ee7a7ae7f7de1b0666141fb8bb344c02cda5a3ef388e6d6a50bf5cec9a33c08fa46e7451a6de4e623148cf17bab8e45a80bd64492ecd1bdd5fa80ed5baaddeba3a32fcd420c32865f7c370f9b6a5482636e66b8d39aa6957456620e1448356bf7f608c6e537f8f88a599069f9d9fd5dd8b7431c5bec603e08bb9f87867adf8107adba4d58f76944808b377638a71c7f22d19c5cac7808f14d75b0b57749a5aa5d101bf6793ea61897fb1cee0ff058ae85b4fb45509fd96740e1d6acf8d8bb33fd3eafc8ab3628bf309fd1b6cec62dc56b94313058d71cb04154f623a1fd170d70224cfff13592a75bf8b5220998f1398290f25955149091ca0095aea2a9cae20187e9cab95282814d462c169f3837a4d9bb16d20b8938f98e8dcb0e25878c4e6573667200cef913ae35bc445bbb113a67c08d4ddfae09adfa7197abfbb3248a4ae118e4b7e22d58ec5985a8bab4b0a3d2c3b6bce9592b96fd70a0a7dbf57f948909bf10e5d0e1f07331bdcfede16621c9eec92a5123f92a059f697766e25550c04e31e36653ca1ecff8a4ea877966be54ac76865968ef2d80009e0781f0ab33ca0c44ab4aa6ca9b3ca01a9112c397ebc77882650bf908f52b346eff53c05ec4ec22dd91cb3a58a1952fd7d5801bdffa7571638e26891d712e7c14fdd214972883a1d3ad7693c871e2450bedf344c38df1625fab1b8225ff9894734891157a92c099ba88157d0df41fdf6b9bb2e40e6e535a37e5ce59c836092b359371c4469d7ccd800df8f35088e6746403aae92c151930239228686c17013f145e6cc023818ad1b42510fdbc04b777a9bf0763b9b960d67a76f569d48b068d7b822b4626dcaf80670af5ad6bc33755e10661eea6c621e60b91998df89a8bdcdd529fbedf0094378af1ffb19f9fabf4a1b319838cd61b9dbd530efff41091829384e6abd3ab5ab9c33a57fbda53c947d576ecc93e52db8b120d4266f8356c0a93bbf10f4213feec74ed205f37eee864a273a73328d47956d944ab4489d9a9f7cf4930abef7f955b3deafbc80787266d94aaffee8b01e924e5db2cd0bda9fee5b8313e895c7ada0aef41b9cb19c7ac9b8ac7fdb39779a9456faf8e24a3432651585489ea490195bff96ee6e2339b92fab398053895c433d39975a6a9afa0764312429867e604aadcc9437a0e84bc8510c45930fa73cb3cca875fc3e78b57775da1edacc1294f4a8ff2249fd05b78201bdd74d5b825f41afeb8133078356feeb61dfca8b852793a3a14a916b0ccf02db9a9c2dae1eb0495280354f0c31db14d84db82e66fea475a498bfb5def7451bcd967567a09c7700099969b98275e2ed2f9ba2b729d7c17a7900ea78d6d65be4229c950730d244aa90a6a2a8228159f94daf40c41e70794a93e14d17951f8a49667aac12b3b103d20cbcadc32f2e1a4fb6deebd00f8f8be930b29b4b811765114261af931c91ac33336345dc644ff259789b7341a5f7ca2f832a080d3139878a71897a4442943dfe5cabd51ef816ac88a9b5d43679747bb7b3f1719f4afa3fb4e24ec5438b9518d753d667155a1257a7f59f736d7f74090befcdd728604d8199101e20c16e58cbaf6db0ef1afbf47102d6b161080ef161f4b71a84deca12ae2ad3f2af87a2ca1596ff44b483ba2e6e52172fee4eddbe91917b9b74585c0d8657e5593904ac5698cae9ad9630e3fc6fe296830e2de7609182633d36ed9383f6495ee32c7fb74f9933426138a0abf90df8120f076514a2221acb2b87a249fea220155ba1fe726ef2306793b406399e3b2ccb2ee9fef8a31882ad24d5400ae2b43a5efb0c45b43b23e2f6b3051acf0854fe7bbc9e9d8b10c6441dc8e86ce02b69d4a9663b0776e34623020215aff49bf6630535d59962cafdbd52c609e399972605d0e10083ea5a68d4880ecc1020fa5a08eff52fbb9739e11c26e6a5225ef27afa1a0e1ca68ad2e9e66c5ce342faea508f955fd1853d5a6b95d7a8e1c2f2d4527da3b4b88ff48d54b83fdde9affa3fff87da57ba21927c77d8dc29470347c6e5ee8a0d2fd5a4e74c5c31a6044818e8e90e2c15547d9915a58964886deaed36e7c3c4ac7a0aad0abfb3eb2a5276a4c7a7b230a9571138a332ae72aa67d6526aae8f09294b90ffc10db8d4865e52e69f4f242885bb98816b1433c846a38a30eddfc1e966edcc2be8ff07ef11a443540efec2f779d00179d1b5c60aafd7c23b6df1d482e95a2c5c0939b4f71f515f7252039366bb3885b45d10227a17595e5a42ad2219385126650c1b324e05a76e4a318276b446d452712ee514644735da844e4def6ab0b0a9acfc991837541a0957841c082e40c585fdee7cd81d154ccf9b62b18f0bf1d0516c6d3bfbf778d99e550e225c4126ec9a46cf285a6651a4eb3562b1c889dd57ce3d670673ebaa0605b7157da04ff27b653502a858e906985bce0999a6035d196f8e24001d2b6a55db569deaab31673a546e5864887817d80466159896e000cf6faefd4adca5fa30f69363b94d878a3c11037a29d02c6d9b5e91ff6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'haf88d1e307b9807322fce4aa0a69727276009ebbff7e6306e6cd519229047106f6fcc1fcb7e372e2fb55838a656c6d835d741475df2eac51fd69f7af7a26eb8cc9ada4977240a26d5519140085e861f28d052c9ffc4d87bfd92e486b6384fc373e8b5eaa059040090414b00fb6e8f1754a97c6e0d65d8708aaa19094fdcf79d4708aafe447510fa33fb423b1bcbacb0d57060fa275c34d46fb56f70db60438f731d932a3b8876c29ff0a4c29a018b64ea79c33b2aa054273ce3592f4603996430c81650cfa9283873563b5e001af715cc1553cbc86416bd5b697665a6b4716a2aae22743968ab8aab7d46bb9ddb781bd18add919f3de57e26dd2ca8f3aae9db39e00edf92201c77a80b18f3adc0f9beda2dd1e4d6b23fea034aa908107448ed2a0837d5d6fa70e8b9ba1c58ae24108508c015e1620df9213afd7b101e8db6fb3508a180c9f9f6557dbcf1eff881ffcb1c8bc34c06b232614756c02b086ecb27eaa375459fefc2a5b20e323d09a4b6b117c1accc2e240eeecaa1b5c04a8a214a8c926285087fbf07b6b72ff781d0f69343bd9144c028eb1f7f80d4afbf5504d90244d8b8d318214b2d5bfe4e89ffc6df39fe7275d6890f42046635ce800ac965bdf144272d417d791cdb32bdee1478ef95711f212f163dfab736212e7238ffa55d6b9b091e541280949515c428668f51b273021b8032b7b2a78a66da269213eaacfc0e5bd15f512cc295334c7721ed3df0ca79a7e5304872c037f87eb155cdd2d1107ae12d61e307297bd5bf525e2d4b4cf64f949827e49c72db17b8e23eb08c4cdb687e3e1cfc5fb80a53027c1db71abbc5e091067c9a67fca7ed7165d0db5b0298cabdca5b3379d8eb228ede19f60a9e663420d6a36800ab01b58be7cfd3f44e77db9a82a6ee2a4f051a35f7a5286c35d3fd0bdfd8c327f75e882747cee0da0a7d5f4620eb95a1579640e03d529405efc71672aec9d4c90f7f706fb948035456edc02c9627816557f46f9b9ec276875d4dfc6c9f97e123f7fe8d9289c4a0e4a8e1444bf499d35d78699eb5ee4413834c29a8f72b21ab5beeb25052835ea3e728223950e02af518b5feea682d93f4c751d50fe78cffcc248364c189a5320afb69f98d4ce06c970b483a08c6fcfe0934692262d8fe40b9e7367f424b843d3fbefba0c6f5002cf28e945672243e905a9e12136627a43d2e3d71a273800b62f23a8ad9c28baed536279eeb1462a2c5df680bd67a84e3eb98b3972f407c50a8de56c098f0e5259fd41dd4bee047ecf3fbbdace698e247e5eae8ba63d7b7616436dc191e9ffa6f1e6152c8d66383aa72f6a53647c6dd2cdbf8fb6020c75a8c104487e1fef4b6e2139f9db1f835d5f4102ea439ade0ba9ce59a1f4fa2d7ca99f5b61c5c7d03c8da153444cc01a553f4329699314e59b49a83fda10153f887657388506bc6aa4cb78eb1eba0236d83a0de1560cecef56e07ce389bbafc18d84a7caf67acce2f9f494c34b10b61184beb97ff7bb3eb0954d491b1a71f3e474ba834fe1b5b9cfab24c50016d7a9ab2427ab5a24955e2ac78e144091afcd248887b2becbdc1e37a05e0c0effa9873d1584db7f6a5838b8b08c63c484b36418fdfb21a9fc079ae6a3a35cf9c57e26b2ccb884beb60463cbb3fb62616ecb6b9d466b8e163b056c097a1cb35bc778348ad5fa2cb2f2ad6aa5cea5fa7ce5d5449fd1b3f3ae92793c132a04cc6f550c4eb2d771124de088bb1fe856a8ac8d84a82bce70937e3becdb136514e08d07f86dff6cee8709c7afe861865e18b2dbec2f475fccf459b4a0751b75314a55abab43862c54f0bf50d8a69a269b5eea756384b9ef5f34e9f5522c4c0ad057c5ce0d7aa61d3922c470a328d3d2bc426f8c9d7328369f0fa5cdcd1c00f6a978e9a3db1add38bbe39bdf1006ee48544627e74e1ba958c1924dfbb167dcc0ce54dfaaffa349f35b69fb3d022b4d77b80e655c24a35a5f278f3f98664a46b7b634788d95ee2f857d9a75a05b1830bc189d934f56447e040020b8de050b84508a691af995c0c79f8928b603ac13f51c860184ce8a7ecb3a53de07e630301c017c2819784a9e5634eb410bdef8abd084b1630ca224f238c2ef7adee0662b3a55bab294d5dd2d0ef60d099aa156be349aaf23f55cebe10443339559d7242782711452a3118d89c5c6cf29f04fcd89c830979a55eb3fe06ced7fb8dba082eeb370086352ce720402588efdd0f5e2c04dc13506fd2e3ae6f4650b9cc5dd1103c672312b0e99522f0d2714ba1775d93317946e78553fe7eb4a8917fcc15e4ef9afbb538563ba6803769e791af1b3b10ebe9767953189dd5efd93320d2eaff51d3ad3d456b56322e8518b6aa5bafd1950cf9d0ae3848e310879ac65eac468acf2db1aa3ae122e3c227b18f1203e09b0bd785288d434a452585e75884fc06e719d438d823e5a270663833a472cb56de34e89c1a8f34ff0b86dc03aefac3bb7adc6418eb6ba8a045dee518f736e272520124072b17851ded873093fb22f5acc1a8d63c4e8f33d695ae7ed8af593dbd3b1e434dfe1d6f3ebf40e6d2360186cbd8ee1ede78cdbc413422d0c3a9517a56bf0060776b76707c6e998fa5670c5b659ddc2d1335816caeeb90a1ffeb4dfa8e3efbc55611cc51acd992591c67c6a150dcdff9df151983bb591655378a54b3e7a4ae5206872c804e8133934fed796cc84c01d4ec804df3de5ecfb25a43c672e61c730a71317d4c7219e026894b216a596ea47428655e0d01240849123be3c7ef03b1174b8db2a5171db010773397154075d1edec20143c29c27a23899dfc439727d52098d7c62c698b4e6233e40d57788a2c69bc696b2001227a1d83c8dccfa0e3085c87931acb20d7344bb63e0cd4e9b9e265ce28b750b8fdb54164616479e6473e44ec1f3d5493e3077c9291564f83ad82939e7a5b3fbcac8a9b725210b7c3049c4a15cefe58824f69a97d254682391ee2ef8c328f96bd74918667c5b0f8ff083a80812d7b3e0c1e1d122e8d108e9b6d087b6c7f67e1544016030f4dc44653031466c3ac80dd1aed4a7ae633969e39684d53d539771eb0e3c5a53d0f935e6c4752a93d81155ecd387843c4eb1783ea7040893540ec906b9ab3a2c578e67278cf48f3e7acbdf54db628d14649c40c70d1955dff67853a003fc0531db3c6154c14a7576db1c1afad671f8d6a0257b54bc31f79c11f63bb8876f04072f4f55409882d63e393be4f86198a7b23a98d5bcf170e427d5518251766916ab3885a8267c439e660cbd744da04bb92759da4fb248de2302aac98b4799c60103e3033144996dd540eed93a471912aa3b76e49005546227f3829305207c429b81d6650f8709ac7102637751872f6ba2a0b10e09bd5567d837498825a267a5f9c822dc20853141a92fb62ba3ee1b7cb724a5716cb4f4e240aee3e99a8e68bcb24bddd9bdb9116f5552c74418d65838087ec0385986523f4ad1df627cb231936dbce263e010da126b4345002485d9981c41def67c1eeb2f4646cad7452b41ca9c18f2a5ec0ee4c4b8eba1308746d339e203bbdbbd5d0be127cc0d5da486a82d45f50209e5b53fd1d31911d82e677a4aa196ae0299e484876c483cc72c910d6c9163e81f2c20d1926a2843b2cdf62f0d62a370f735e48cdbd93311f739861dcab15b1ea9be96afbf66b7422270e9d14242e73c99b0e1535c89e70e3214a64805e4c30d0c6ef498f9861deef2b0f4f85f9b431648d54e2922b51496053b0e21fa5223331f15826315a9d6b32c7071fbc0138267f301bf58230ec67aff26e0d237168be950a9f9674afb6c14e40e87bc0bc6d879c67681a44bbdfda1b915c8d87d86d22cee1311ea691f2c3347c8c80e440e20a711849daa11a03292ea3b617d52dee0d6eed54b70b585a43a96def139a5f2f1ab9855fcd79401ac8ba472d644647b7acde488a866b083ed7e325030ed585d9f6dd76e9819df21c5a133c8410e561214b99ce93fb2e4c4af8420280519f375b4e6d6e8e1324ae7beab39618bdcb393e1eed70ec4c5d47aaa8a2e8095075d1088b14829480d8e3d2c69a9ab5ebebfb60f6f0e77430af5e4374b2379f540f4017bd5e5f8c820b83aadd41f8374badf17a37fc8ec76458fffa829b06d1288f41b9f2e1f24788f0eebaaf48e558d3808de2fe58df27fdee57710a2d1737e6fa34ad598d89577a25a1fd98e81b15147116ae24fca673404e5281df4088f8dc56214aa42113ff4a56ab2c8356a51549817b3435bdf5976f02478b47c325a2cbcc473b752fbb1f6daca553bc74115d31517e358029ff506aa032772629a42f9dc706e6a7d9ba21aecee89b2ccf6eabf067d1808a269fa435d3c121bbcf56db7309c5d8e919847457c5db5fd29d92a0867ad484aed6ae950290876db2ad177dce74cca12999c71aa3674342322bc4a7fb5cf57fa3c98ea6d8904c13605bcc1df68341308036941debf759f556fef69d83ec8af98da234e0b452f14879fdc35b62cd125cba105839486203d8b43a24c3d063b2367f02a262dac0a863848ac09a7383fe051afecd709222dbd3b31bec7e814a95306550100912fe333463595f689a66d33657ab466c2abd3d85d1f2550bb51ee5eae1dbb2d2e8fbb04590c52a62c39e92d17cce6c018a53b98818c12d5f7f55f49ad35a80e7ae911fdf164a8253f10f6044a49f8ce8ae498a2fd8c9e18a509cbd765eaa7efd8254ccc45498955ab2c956a7acc05b8b547d65b0e40db924c7795af88963f08b4d81a8cb125710efd94f76204f082057ce62169ad327639b7d6f76f8ba03eca37f649bb7bfb1be96ffddc4e1ca308123d2e843b0451071c59440101d8b55b9f5ce6ac6e69d471bbc932339598466d7128def848b1f51436a042fa1b8cf754f753786b118c6d4a78e184429d368a8977434dba96d07df0c397e532565e26027a538000dfda01e729b9cdc8bbf683870835bcb7e382bd1da8bbaa1e16b8bc05880a2421dfb754739b673e58fa46f5a61fe7e7bbff2d3806c8f604c4946a8bb099b22fad8e4fb9910eee7980961c76687ff9b337d3eba1a91fc353e1b66c358dbce7ec5da7ff86f2187686dcf2563096961749be97d26635c8a9651155d7e3751cc1a3fd3afdd99111a5ebb24df24412637810d1921ed1c74ba1fc85238387f982a95a74e2edb7cb4154bcb33c5ae88e395142570fca8533224dca8ae51e53a776464845f5b3a1c77aad2d372f8572c07b2dd20b102f189c1ec494b8f4acce2f10121bf21c93575f755798a9517f901840800dd09c9a8636ba9d2b44cb123328dacd8ed42ad40717727528b9d179937a47b2cb884a72ce8a5a292b18203da48e20c8354d96b35c591f03f4e57a37b55766cdca4f5aabebdb0cf41d6048fd45ba147d2ede7b98697535a4b6eb218b1358398aed8fe00e6f43000efd17e65f4b48366c339e37756af09029215e160eec4878e2dc6fb6bf335745edbca425ba697ec0645163;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hdb96898152a5fc74029f68c67d2cf9f984c574ac266c2e6365ac5fc5554e82ecb985327976137f49aea01cad5b46ab861ccb69b0490467b7b88bbfe2606a52ff6b23b2c63146513e6e32e10c108ba2c2855493caaa7550e079ad9a6331e7a761d4f7494606c29e60c447f835855fe8c4187ae0bb8c9ebe33f3f933a2919a692ffe0313c9e0df8ae5b276d7d88fab1fc340f16465f16ed38c512cc2e7da614f2ba9b285904f54a569659a4189a770b544eb3fcec61c9507dc70d9762dbe00a57af65acb18a914c9021c303dc86ea816771ba9390e4acb0addfc7e535e4cfeadc206acc88602f90e22cac60bf9eef7822a719fbdf24cd552d1881ad066be67e1a738bc0941bfa04a642c0fa1a888f2b46a78ed47c9493678a730d3b6aefa509eaf3b203d419330e9349929fb6f714b998f12b8cdf93579cbe28579599b3c518876c959b86ed5bb9eda9a7172a468e5278abb9c7db2c9dae0d7f79a163394029d8c2748fb684d0ced443bb61cb02330e93508080f6bd554e4b42105488a101d0f8d7dbb2d98d5227c94d413f1311e02c610365a3302244f22d91f5bf5de99e0bc0eeaa97ea8d942851a3d2c713e0ab8a8d2a572b1f6e2ccb6d54c854810726a8dbc8bbd21dcbc0725848f2f1965d55fe521a525045de1e1037fece9e1496fa038deb04de0bbb8d5fd8a2adf48d8681e1711ad9428e81a8339ee0362be60d421d540e1ad935c757a866eb828296f69f424ee1d70d2b022dabaa3dc6b4090a3bb41446fead87d9209f67cc02b9772e8ab19d34ce08dfac6fab86c4d96c4f05fdbcab1adcc38c2a1d612b8a17665286a0c086daad42b5be6c897eae71b2cf9bd7e0606aac58d50a95933e67a9b7f4863d6c1225074aa089b576078b32d23f76f8cf5388bfe6c4b0aee90f88d5631b4e8589a7e712b0257ff49d24bd31b6a7d1ea2094284507df001fc5268871b2f17fdfd775541cd0171fa2211be9051c017375ce28f8556f84eb9a466cd1ca91445ebe5f239bc3f1dc29fdaaabc8e19ce823ce7afadf8cfd1a383884c1cfd971968e0f88903d94fc602454f0a4594616240e224701fd00eb82382faa5e22811949f5e1d7beaef1d905005d14eef499fd05b869adc1e60aa01eeb63158863431adfe4c8013fc06a5e2b10a7f2017c02151532855f0d71af8adb02134bdb739d477425bead6091e89ec4dacc32a55009b1652c58818e3ac7aad0da5f6b1cc2f166799ca86bdc1b41566479cb145de8ee218f0d5c79b524176a6cc144a19c06a06b1bc9c8f52321de1f5decc53b1349a116927df470839f592d6000f29423e8973074ca0a4a49d32c129fb411157ce848d6b9b1912a5337d924f7ba59c2dee637aae8a49c34ac0b7b628bacd12d7f519367352f9dbaf902a6ec25cefda98ec06d6c0f74b03d4671ffd2fe41af85ae24db73fa88bed60264e86810b20966b9e263294a9d2642124dcf70ac093b130e08e7c0aa78058dd8e8ffa807abadc1ed602c8fe69522c51dbb1e625e4c7fb527d82785c620d85f289ba2eadefb8e53c94ec781723de83d2ba864fe1f3306e8d60616727ee4268020cd5abb3c0b6ad7ecddd2ed63ddba0a1802a95fceb1b4d1b659bf94d0ed78655ef3f1502dfb36c17a93b139fbe36333f019b8a574ebf909d7f8b6a65ad184a5f87cbecd54d9937a76b14a45533f70eff07703968154077a5a3fd3ee271d359cfc3bf1c3b41718cdd43ec18947a73d158fe78624b9f90cbd70357994cc79fd5baad90fc46646216edf364a54bd4c2c12116a0ed1b823254bb27690753232b89f6357b66f87024edbc302d979654d25622c04815ff8ed1eff10a0f824f71b302a60f94fd8b8be81d06b6832670773bfee492745089281c97baf6982af590c8710cd1cef2af5d85f6bc427e86a782ffe89f8a8e620feae3aa64068d0d04548d836b20ba332fd6148cc54bf24e55ee92ba78e77e632f1beb7ca127e5d79ac73cab42e848df31fa44f9c433a065ecf5c617465a53d6d52db8987f5a7ba5c63c51c5b5a51108ab0d9578884af4abff5a012f9b04de167445beee3f62f8f7d56c76c4e7e4b6964fb3e29d875921c1ded357ab2f8ec3e3089ebc7ac859ccc1b2d0a70784894c64c257c344cdee2000b19efa305d68f019f0938233a8beec115868811f847367c1dd50865f6b3a3b19e7bc1ae0ff57c811f822f3b9ee2a1a05cc08a2b12a223c5cd218053ea875bea2f6e163e15f9e104a184d753924de88388d9a79978805dd5437aa002001a39ad0ec34d6793aeb2bc3cd4c51bf1541d44b85b0521d4b152fe4656fe8ab41caadefdd2bfb8d101163f2c1e7acb8cd400355b759d8e3713a89b5b9cee58d09e03fcaf42b4a9215b6bb8d50864982c47ff58b0eb744ac5b37dbefaf3a568d7b2da95fdd4911666b01a4a2ece00dd088e1167ec8d38821a22832bfcbaa1c768ee1e16ea6765fd2b9d84c2a5af59596545ea212bc363436deb687fc7380509b8f0e630196864b8dbf1ac76fabe91f50be4802f9061e4c5b61887c942c92b05dda66e245914bb677f7b302292eb4c16a1a1d17a03149d2f04b9b23eb39cf403f57f531e5250fe34865908117d2ba3d95330e7cc96849ce0f52d11a4c2697db79e421d2aea870b54c77f371efab64badb5cf1c94be161efc415db9817a28b6bc9585d30eca110ea64d6c74eecc4dabb2a1e959f54baa12638236850fbf9be5f156a55b6dc6989d76c000e8245c669b6497cd2bead8d0e06731410d5d5615ffa1eb12a3629d1184a89076b75ec41964c89b3c8c77ddd58b6909e38f15806e6410f23cac9f3a44c847ee2886f7d4b4d24679bdecf016801810914ec5ecdae8ede35eff61823789ee8c013e3e77fffcdaca1da2899f75502ca56b14065ede97e99412748d927b0ddd154fd0454e05b7c6b453cecb297449383fd8bf0348d93d829ffcf72f55619367f78639e584d9b41a37df227392609d67f7ce5e5a9392750d868a2105a6cde4a6f32984809814f8bb87d155db7311c128d903024d40355c03c4704c30a7a1323f9ff7ff0a6493940b9168cde96742df32d02c74d8092ff946717f2af2514ec52cf53b189a1414b9ed12deaf62bc130dc76641c3759ad62f0ff5ccf12b32f26228ec077c2a2b12730a5e63c36aad21c459744722c96bd645f671d9ef35304818a34d69022b716d28c5c060f53def4af03e11c5da4838893e48292eeaf84cde4a9347159a6de9ec3d4a0888cb4441a3d4ebbf87f6bad8096072b39f43c0e72cbd06f19be08d6e560c080861cd96616547616258d485e510a8bfe267cf4aeea61636742c8b931eaaf0212865a0c1d6eb5593fb5b51702cbdee07aabd6cc8de39b137253afa1b741926a1c3423c15c090d790f79d9e1f06249fda21441e1e45918e16406d04a046b8382a4759ea865c4735355f1dcbed3bac3061e1299c28377e35b058313a73e75caa81840da9bdc4bbe2f34a302ab47fe940041c650d26e62b8122421b53263873bb6a77bc8fdb28de33c69f37f964f16dc33d56920d8ad2c8b7af3e41913c7a53050715048e026c547ef63e8f23042557e0b6ddcf1e8076d8584068088596d735a9def50bbd490728f6d14583d79934bcf309073caeca5a5f5161c15dbe45a59c9e22ad85692e8bbd7086d85b65884c50526a0d019569ab7be80204738e1e19dfe892c9fd27b57aabea08349c029379bb8b80067178b7eddc78684d373379cbe6c08dd59b3cc3afc0bfd9df639b70176bc8df3ae2233e0719855cfa0592aee4c46bacb1a712b0f070d4fa015fcbf14b383f0e3f4171101a00e3d37a4258c2815768fc140ed1e149dd2a3409c6d2c29eb295fc1dbe01817cf423d6ced830d08da61cafdafbf4f30acf2220bb80aa9f0e7576abc3e2f6f55167514af6bab07a34a0979a1f4e78483be023fe616710cd84645c4bbf587d8a078fad8bbe008fd8272dd7ad8ec47638c5b0ab8d8479875a7556632779ddaf5317934690dbc7566653382399878db4b82ef05d84ac8af99b5990c9b30d84f7a16d14f823fca351cecfb7e3c790256d36a286fefd9cb3f27742ee53785e863734562e949734bafe5e2c82bdc4c05b7f25f914af54a45a5ce59a5491721824ebe72e16e673006c0dce7197c5a92ada2b7f18f8c7a0c498615c08b6ddff53cb3cbea1135c75d288d63c3089d7822e3c41c700243965a7f56dc2941f4a91522c675de40a9cbeae46da63d7e35d8083187f4244b8349997d770e9fb3192f730f4a630422ec97aeb598ced0ee548f44ce5d9d430f9d772e31118e06d67a5bc86f7cd8e8f503ec5949afee02f917b718a83d7d3ac39aea5d6e1570e0f4166b132b62ae5bc53a6cdfd1ccb86cc9948cc38fe0622f6f69d4ce7f3a95604513da9f3d2c77a7c604157fa1e9b995f1a866e060a2bb24ee27f8ddc78246547e44541aa84472c7ede6abb2556521d818c5ab1b588b4679d792339b3093c883c397733417c1150da176145bb37aa9eee34eb8698b79b3bf60bce918e2a3f707970754464b9782646e8bdf33496efe8c113cbc3f86a1bb500479080dc7e33472b675746e7a1bcae2de04d55eafaa8c33825f187672a92aec84f52db43b096aa9436522062610818534263d756ab6de81c0b5d7f943d5343588baaf1f0711ead75596d0bd609a96554e7d601174fa2d718ebdeb300dfecc906be5d729422214a86e3083d67f4e15ab34434feee97880c8608ead84fe0094c7a53de60727df8f45b0176a1c2e0f197158acc50a07ca2a9d6d274316a7265a477b043f68a8f8d5f5bab03753976c11711e2fa691505dc4a581de4a5680dc93041eb63b16642847617496d99a12eff32a25b696bf043ef350905138c46bc2946d00cc18186228e7523282b3d1724c698c833726f6aff1c34e430b7c106db8e929615950aabc7a9d3f617fbc27e211d1327ce8b85406697ae78ce1487dd46c5ef00331d578c8c8df8d9689f06523608268bb6c1e5f5fd5a7012dc114e2c60788eccc7327db5f934ddaaf0421c1463db2a44129bef6aaabbb9b942702c72a5e20ec734f3efd62cd3fecfe04c062459fe4be586a33d14074dfe3c369ee347a6995b3f2f4fcb56f8aa999061f3bd74c673feaee0207d99ba5c258e7fede6bbb442d5d3940fb34594e80d2d98fc957bcdb7290c6aac6208afd7715a95e38eb9227828ba94894b8dc88498ea04b40abe1ddbd577c27fb7df8c12f821a9254680bdbf84fedd7609dfc68685a66271c9681375d7ba42541c0959d39b3f6190c4ad9a7c2203c13d6b1d1d84ee5db52bfa1f2c9a3da91aea642fb5fd66ebec92a3eea20384ecd83a18da97991359de16c9978294618d6a7463b57779fe3abb13e7b2e55f1ae19094bccfe6721e3f4f726cd04c9a35aa65403404eb503cbe369be009360ea5e3ea1901b5af73a66e2af5425e1b81bb91695d9dc2cb529af6f1e8e9e43eda8d9d7f740669052e5478ee254a4f0ba787f171d5509a3b1d6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h472db9eed5dbfb6cae059c77b808e34832197075c46a5466a43bf83ef3cc21772c4684a08b58a88062240436c5dfe21c6c6acf17451e40166326f3f4268b53d4df92a76891170a70e283f58f8753d4d7ce061fb92129549ba10538b87c9a785acf8b7293e61c32c605ba40c22ecfdd39239a8e8383120139551b8f46016d819f1182c2f6a815187c974b4d03d34812ed9267e58e393c2646de0542933819876b47f2754ee74e69b76a831c3e2748ade2989e727cfe132d558d597ea4dda3dfcd257da0c8adae2f49fce611fa5983ae80a2681471da2025b696c75247ec070d7c484dc1cf9fc8f09ba3b2ebf81ab2170578a4a0b835378ba9ce6909a09731c9729372abf00416177b2bd2f860a3ca55828508f9d3da81c75e97b7cc7ea9b30411e406dcaf65fdea3a4dd469482e380e9c58245b314cf566aae3d2c02a647f4650f7be7a1156fe1d06cf5028ff3b3e51f60a1c0c41ad199ec644581084a470880a015145ffa235358eea4542fef67156fd67be1c3f42a7bdb03933334b2425ed8d86519df4881650777e2aba52b1b42a18793cb2af675143f7b927cdac86b2d07017605d21973c2ff1176c5881d44b018425218abfc198167c7f9ec5ef62370a51c045dda3918b045a87b203133a2ccc305bb3461893a131e65ce04248684665eea20ea4c6179e63e1d919c6bd7a09ff40ab9e80ec097695bf71f6c3934b28274d85e7b861c4b10f33a79d02e313353ccec760551b1b67e554dfb9095adfe09e8da1ef7c4885df9d46d4ce0dd8908575d5efb76115f123c06b9971e4580dbd95a63394ed9bdf3ba957d027ff2cb237d32c3ffdc5e1f7669aa9b7a13126340d70889ffd41c2aa0fb7fd6d3b1f0953e90af7a65456de68dd86ae4a9430fd19ba6595ba4bc9ee1d86a79e1b738375f05356d396e3a3723e570ebb0299fd29a5c770b195e4a3edb7ec2ad77511d27447a078133ce7b49018a1accd7a79d2e9a2e67f544fa396014a80bc3feccbfe219fc8b764ed94694e734dc1bea1057822c705b6973f3d8c64d554c0de5f599eb68914372ae895f7c969051403c863c8ba9d72cecd1506180d3e584a9bb4da0b9ddd8c29071f9f984bd5cfa65cb65b49811b0dc1da016e1c54a8c723105bef2a80ad63b5c81236e51ba20b650a317e3cc4c68c32efb2d2ab81f94782154ce135801c2301a5abfa112d8f6b72d22df60c3dbaf4f7ae6fae68b873f8468835a0c993db523b23183e3c74a84b3d91e322db6d2056416f82c3c2853f91c97ccb480f50c2e278fecd8e4518119f9709022d5b9ecf0234451a269395d02eff6147b68c26734487457e5de4c30369284b014e1295930e92f9b7eafdae47466347907143c3dddce46b575ae03ceea8ebbdefaf1855a240bac9d10e5327381ad218f74e9079056f4b62b2a346e8c510339074a32025700b1e8f8c4fa9af3e24a33aced409032f6adef03acc83b66ef0fbd9abae8b250aa7dc6f0a5212b44eb24b4d695814636c1157463f63d88b2971746c6edff3dc38ed035dae9f443a5bb204e0cd17ad06f9df2d2e62090ecb8b86ffbbf396ba20877c98030e1c4b92608e15e599a5f9b0949b0546124fb1d7d3ec4be082fd1da31c38ab828ac474ce6890f802c760471ccc9f132d783f7e814b5f7fc8201decbf6df2e5459f9563dc0b77b19f7dc97f2f02aa4dc2591652183da78d93ec06909432994f3b0c5b22b08777500599b782bab2d2a8e7130e37d52631c6fa9c4aaef39e0bce223b09cf36fcfc167e2abb90c4dd11c3c3294d06a9654b495323dc050febfae7b6d26c5dfdfe98c8ec85791cd48a1578042ef0efc4cfa125cba67e13ba71abf7edf39ef51e20baf007dd46b3b80702dd921f01654c55f933f7ff9a1d216b274bc70c495be284c0de90989ebc694b0c514fcc877c3105f3f8f2f04043816fae35f91d3e2447109a67ca380edb70e0ea25aa191939421850840d31d6743e2d3fc9287c8ddac8b68d7a072b307cceba2453323d54af2674d6802705b7938242cb20469df5054183fbdf02dd7c89e44c170798a11eba9fc65ffceddda488479e62fcb18e121f32acfb5e22757a9efc1222a65ceed99f2aad86d2c6b2289a89ef66ca453ade6ab19ab5c0d76e9d194ffd45eba0d197e8a965a0a243d26e0752470b6a0eb929fa5d00ed25940c6215ed6df2b1534fb24510b40e58789299a2fdf60a712fda2db59bf08883246ca245f1d2b4362df978cac88c0a010da4bd0fce67f8a4b215fe337b305cc57bec3091f492788f7df182aa4613e576f43eb81e0f5356e1f0bf95da32ed6a998c531dfa0b77c9f193e878668ae4496f8dc694cd85395c5eb4d41e60671127d6a0684d3a1217906079ed4abe6793d59c51102fb7e0ac6d6a3608e28fcb183a84b6e91d2c3097052e49721d814d86cb8e4060af618278ceacd2c728c20d2d528870e3d1f30eddb9623eec7155d951e9da9241875c8c95b509388a2775e70b455fe49e2e9033875fad73e02dcd7594d05ad80d1791a7a1fb31d6a4b97aca4fa25fd945751b8dd32c7e0294137704ceebfe372a05f467ab85570b00a3b6e5c3a6a8c43642705e1abfbd75ed47cfb07318dce7560a3a96af56c21675836af055b02b4e5fba6f7ea6e189da0ad4c76efdcd0ca5139031b0a829a9b4934ee70d937b3bce8923ed58f8b85118e9018364f5b340c2f6a25ba052d24a85c41861ad2b368a302917d79994f5a43d5b56c43af6c37b60087cb66c3096ee63a37fb732d06a55b7a83ae401e2ef9da5f00babbab74053dc6dcc49c482e5819845efb18f08cb7436f49a99674091dfb02c7a4f63cc89ec395bfe00f0c9f3c2b10fd4be5f30cd3984519771057a0c6bfa78a2e53fdeddf90affe93114b12c9456b00b4e36323d1a4a0f80d24bedbae6b42cb03e0f26b89cc6b1a56b548bbd441661a8e62f8c1693bd43f1cac96ed305cb6c0412074301a4d965eba600eee9a77551958fe69a0ec5caac029bb93c07931765de950761fab628f78a087708ca066307fc9fff1805424eea9e719abdf18203a90e7197316bfda7754c97e0bb6d106924a328abebb032d3eeba07ec5ffa2ce66503877fc453f7d937357ef7627adbd35ab5014309c5ec4bb30ed13ad94ac81ca716b67dd808b30f2331b57345da900a1b8bdefde8f167bab5e8453b6e1d9bc6307a51a112b40a3e60e5411b9720b98741c98df1fce4854004e1e79441230bf76412914127bda958767d7405501d1d9b55f5478c0d9c194c627e2c8ff863056f521e912cd8be38a04ae20919f908d7c49085f72a34813f14184fc0d95e031b486db684f4eeeb2b93d495866553f778b3b283de63cbeed58f5d89c96a24b78080141c4765ce0a6aa53a9477bf4c022b61904ec2a36b9c4ce9ef2855685aec969a088a0e3840d29156e43ced21646506fc83b38db6596c9224e9e6eb0b498692d21e806ea3a58cce6caf496eedc7cc9fdbfbe074ba003e78e12d547df57e88fc7b94b30c050c182379ed5a1c73457d3299cbfcc0afb7bb9f4c82c1d70e465495f88a5ec1c55824783c838c88ef4477fb44f48fbeb57e073ecea858e35f392a79a52b3989c4755f0501f30c6e10ca9c25871605e93fa71e2b364f3187b6aa29b7487b093b3ab81eb7dafceb789695847bf1ee9e782421bf950d9f2bf3c4667bf8cffdfccb6fc8d86c502b410eb527dc960eb2cb2a4a3c80cd5bff1941240d146d661470dccf812f6bbe817c15fc1241c6637ecda25c506d2c54f3531c71357a062491c7f57b6b7b1cb05e1e184b6c3ba4136b27b68dde6dc92807cedcb92defb21559f60b2b7b05b933ad923bbec5c16e89fef25267b107dfde196a6eb1bff492c7e57983e95858ddbc14bd4b5abded533709261fa959912272dca3ccb8b93ba80d958f0d6ca550cd77ac47f4c3866bb21660080da0f6f2ec2185db7f787449424bf56f472a6319084b0d5a0ff486f2ec749ee918f7014b71691056123706aece749e14bf6d525d75a38a0d4fe90aed48628e3c797d1f223d958ea2f79aca62783ac94d41adc28b6d38f340e7dfb68ae2737020598ef30e43a739b0264d75b87021ff91c2506281842b615c433d89a863aed01857e335c8a9558c91bd958281fc52c7d82622ba33ae4eb101af643a0e0bec3a20f85973f4380c07143203b0ab507423ff0561e22baea16eedc6a311ee15432f1cbb425ae0117c86c478310089db68907a090c00a95abeeaa0bc2377c694a462642fd39ee15915cb9eec2cf1774420afa5990a382ea7885262f1853a4946dd446a25c83e7096adf4ce5915ce6b61387f14ecfc538a01c1a744e88626d547f29734d0c7099786724a3c23cb7f14ea403873faf022ae2ed06a3164d89f1d8adebc857d56045f17cf608de0b8c4df58abca514a9b94933ad9b09accbbe11312f1f37830cb206e582da1ad69538df63721e1eb0606c749ded35f0280f20cf51b946af0245a943a2763e620bd3d191d091fa38c13b3d237c6a86d4970f91f3b32c94a4f3973e9902dca8b94f0985caf5337de79bff92d2fdf214fe9395cf2654a9f91f7edc2e9ebfe0550bf0d30d50984dd4683e6765b368d5b892f21ea356bce6a06cedad03c22db849d0a14ce7961a2db4bf594567e39f9d0ff3ff71316f74aa0067f434984626c197d960b04066254f79c5af39b2fe757878a1e62f88df005243e1ac8979cc6c4031b48d25200d8ad3aa739249090e66152ce0ec554cf05bfae8e9375b4bd13ca6adf4f98f97f680b7cd8325dc215c2a94b28582742e2b391d5afbaf94cdbf95de0aefbe67f4131757da569220f22fcd5dca5997562e5b3c5f3649f0ea3b0e11e7e94f9cc3eba84188f9b4019d26988a32bf0230bdd3a34dc60ebdd9dec2d0749c130e188296f82a7c967a71468a03598c383f930fed86e743ea01cd8f292ab84a2a4d9a3479906bf227b3922a2c60fba634aad7d88f7dff11d5eccb30b42afe97480803b13d31229c3ea812ea310fc04eaf0a6543a45a62287325c28b74e6b297a302e4060c42aafeea39e36fd9fe3f0a7781def499af1efae9f047aa28520fbf844b32a9395760b46cac403519662526f509f15de7cef6ef0a61af6b61cf04575b38efbff215ecbe51f14969be53c377c70d6457b6e2d2d407ad531bfa1cd47aabbd2539aa425b5f4c1062fe669e5d16af7991eedf179a940f9706946ed22b0d3d416a0b31dbd24caac1f836708ab2800a6a08c72b8dde557182b55dbf3bd4bfef1d39d79ca89fc3fd76f86a54095217944602eb022adb9ae9b04d2eb3aa5a9154bdede9f143c299fd0053697171e4d490158ab5184859ccef0717ce577e728f6f7fe5589d347a8a88e030a88a50a79ee1b4050ade25e6478a94b97e2447b9144432dd983747049ef4b641ee6d92209ca4530a8d274399ded08cbdd8d867a32b609cc9dae612606e4408c51b85d51740516d12e490a8840ccef4aa6934e12380c31a38dee4620e439;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h9b367f6dbcd2b26d994f0789f7e907e0441ab367e711e349116639dc5a8df7a3347f6a99955637a63a9cb7a602c76a885d4e94ca9165a56f404334f605c145c4041d643302e2005051cb6edb27e1fe03ccdc87a05b5ccd3d0ef038ed0d725818c950e748630880a68050b2886e2cf03f75745fd2bacdefff96b7d00e768a8af508297ba0acb136ce66ac721a82b85013b465599b1aaede3fec88fb7824584ac1c3a6781780379bd1d6905ae397ee8136b590fe060cc3ce8deecc580397341c90fb51ba06b52eb0c2637aabf2b6999100f907c4bed01b3006edf6f7389a1a3e0a47a2a246eb12dc514393296e0c87015c4908796b60bfe5becae14d578face198801bc550d1f6e13b5c6c49597d5c408c20b82f98f71dcac0886bf24bfa553dade895333ba5e39b4d02828b79ad909aeca0535f97c9bb0e21a236679be2fcf395938776ffa0bdd46cd010aea4457df32b830f0a8a561e6c7cfd59495f3cf01b2febe493b64dec87d156472359b34e5263a064b484345505313b736df10366338a757a07736c076fcaf26d627e7d5317373cc299d961fd1582b50b6e338bb85dc2ba9a986e549156813378d16a3c07dfc5aac5de6102fe19615b95cbbda798b3098114ad3daccb5d11eaeb62d554f4c826db024f9332a146ab2780e0fb3037906a0acde895af03d822773d1c6cb357e3b480e6b6169a4bcb8a7fc10f924a1db23de2f381ba7fa7f337c995cdff2c8da67e21b42435c4f6776dceb49048c61a28950d34675775d2fdc6f31124196af9992fc818d55dc0af54120cd71ac0df8a8480784d312696dcd474c63ddf3aa4493e45ba71e310859843cc071187d701b9bb48c2a6802b4fb92132d3b88dbcb95b74a745960e7de75473264fad907fd376f86646180d79b53b7c918a7413e7ab86c6921317581e745bb22255b165c44974cd793be755a1ef13004f996ce10415f93150e78b8e602b76bb0e7f90e149e6fd6ef4e402280f0255cd16f18a849efd96bfdd8cb2f471c9637a42710dc3d2c6e85f0a7588dc6d14699243870cf2e5d78ffcbf5aa1b61499d0573a064f8621baa16740a5412051a946e34f4d0271c8563fbef99ab0cdda46f01f9f6a7c91778f259e18aed0e0945c59fed1dde4d828add50e50a355d8603b6d799a324ce5e67c32c9455f7801c47e9223eea9e5eb064db5c52d4e72a3e4e0e75013c88b2ba9123e4e9ff3ca6320c3a678c4bba60f57616cad423e2bf1dea1aadfa714563e2bf5c0a3aa5c4ae5976a24b9a919e32e90d0dbdf5fe914e99cc46de9b96548706b32187da9aa7d06eef467161ac7b3ed741700878bf846ee43f50b18bbe97c6769913b7b6bd272377b66a0949f99fd223d75bff57522e65670559a0a7b2a3d310558e93f1343c8f8205a7ae6f2a4dd3fe18761c790f18ba4757c86fd5f228531146a5effc725207cfc51fe2f4f5c1dcb6b5924975012513ce7a69a7f9af5d7c08a0ccaea755bbfb025b2d3e76b2da8899bb70119297cabf73fe95c044f62644656bb59015b455888e679e6b4c16a3d1f01c1dee7cf9dab172d56b65381c608672216d3717daedb49792ff6040b5d1b77de0f709041a079c34da0a25724ba24e7e2b050c6d0d12b05d879204b3756f0ea6a1c25e01fc51ec8800c33ab999875fce85fb6b24148ac56c9f4bc9d4e1093b60a90b356a8486ea07dddda33adda1e3e8602794c5f831a1c4a054e2109b5cc0378423924c2b5d52ed41810953ff55ba941f5c457c5fd4c7a1f8953ea4ad14f56d85d1179947253625c64c2cbf3b13cf6c5c6b5472824153460eeb8db692407491cb8d41aad327d2205244817b04170d768b9e4b2da0719a938507eba6553850defe045807f91db09135c7e6c04a8b3545d1d4c72bbaace6ee0a1d9008c25e7c15b1d121ad3bd7303f3e5f6e9c6445b71e777a6c604f08a8f00213e4c81c2c958b3cd4dfb60eb67c4970b567bd3b1fce1698895c4c0d792a256baa7e6bdacf1be5abf39df648305d47056e1ef38024883de8169810af98aaaac42d58a05813bcd4e9a7734da57d5172a09b94bd4d492457b2f97cfce354243d228320744b26410bf65c8ecbcae49064d21f65231f5e140f344069da0f4a96ec53762d1657513a8052eb68fdba6cf5e7f7fd5c1ee054e7b1b428099dc32c8768e42d4db821a8b26ca2f9a4c39f775ec5830b602bc8df60a46be02ea371fd386f02e3fac0af76c7d80663fd07665dd51c6b4b27be516c81ec88c204f4d8935aa63d71da7ddedadf1c188f6e60177c959133ca8d8deda446b0e4f58e53c026846fad1162073f0bcb04d84e77d6fb3daeea519a4a3669ccc524c794c029cb1fa925bbf9070bed473c4b589ca7b60ba671ee3793d2445c08bfdf8774cb0b24c95c20d5f1ca32d4dd6228634d76993e50867039eb015b3b99eb4d902e73332c5f6fbeb1049e1f3e243187904b8ceebb9174231bb660009815966354b670a1ded97f984640320a356124fa7a6fed24796f575391efd90a9e75076f7b671bdbb20e9d572792a73664d07c9d61557b564efa303ae6ed31a1ebf5d73f45df42d9476626efdca2796c5886f7b81eb7b148be839a551ba4d1fb6bef2de02eb488613add05a6dd12e3c8e7b658e0b0089d81a9999e8a35eb3c5a726ec014f89ff6a6f5001a7ab32b478911af5e5e0c9010960dfa56af2424a5655642cfa233b02d8dae5f7a35f2092fe0ab60356554d1c602ad1c212141d1d4d305e25b15525ee3f8c215ac0d389c489401f4b1869fdcf45bf635122e638b2b02b09c00f53f70d6e28dbaae4aca3798380de3fe584e6636ebfd04334bb815b161bb65cd597270d40ccee2304c049d8db6301b7b0970cfd463be86216783cea3c0c93d3fd39297bd635686ed9283cca9b412b20f3876149ed52da308969d6f1ec5e4e66c68a70bc741e13b151a9544294a2882675713a34a44e79b3481411601bebc7ebbbfb91fe6e9bde22a3d1c2e1015c59c80257bee71620842b51080144bb214904da1b687bbbdddc5ffe54f528f502655b965bddc62b11e24695ec3f149ff4c3f8aae3b3b60180f468d89c213f0bade0ac81a152332887b5ec2358156aae6d9026ba8709b04306f48706dc1b8971ef8e7951da66053671cf6f0fcda47b409e810d795c8ef92e0c026be59fa2d4ce421d9649167de684d832cd8e1883ce42949e846d3f55bd2b7cfafed79fd9646719d89a9ea66ed83caef3771d29bd2144a239f00436368765783867d5fe9e5117d0e6863cc98d52c7d4a24603e94e14f11384066b5c25ac594235ab4d6130ed84efd9aac791e1687a428ad2297136afabedfdeba49cdbe92cfb39bc2227965de9c7eb83449172e0dd6dc173a755e67ecaec04f59b92a0ef91d8ac2e1ff9523760b79912df056d42d420f4cd2a4b96f83fc49a92ef6cf77f525a907a4be735d5e4bfea09c3cb68d3c020f42dc8e3b45588363c167c9ea12b07c6c089834532e33b5afca31ee4c3f8c27cd9281a9e1f708c23459a45b7208047a16b6f6449ac39a17fdf375119f7acb2646e466dfbbaf3e2a3c2a3b08b4b47904b72a1b86b4467d0682f9ceef9e1045aaba9ef7ed9ea7738beff7a4cb34ca840e49a7b584ee3d6431cf18a36127896fc4a0fe33e1a6f7e57373958077225f55c47ed73ab28a6de2a73e0931da71fef13c46844e8f22a4584b795476bb5bab9ec49ffd306c5123315046e3e2018e89b40acbc58892b3936184710b3a460bb4f26eeeda4d5fb88165b3a7c27e98c23699a8542ae31b122eef1396c13523061b7b7aabb71bfc1f55ab44565a6acf754ff3bd2d67ab381a5839d871922e6e1d0a1a4dc7290c5a92ed367abebb2ddd3528a1dea2aff113822b2cd0d02fb39663cdb2824ad74735f9c0999ac68093adf7be4635f4e6476c1668ec942ea1829b9a36245ec9d6f976f395071c2dde14deb79d14962176724cd40c886aae4623149a40ab727dfb72a2997794e7a150d699666ad8242e352723b3f5483e806a1170a63218cf6fd4d89970b1622c0852830acc8dffe07d0349f8f633e9608dcbc9b32114f0b2ae2645dba607f3803b481608e81127ed0a86fe39c80b612a996eba86c55e8aa36ccb02e2d73a77ab7a17a2727ecf862dc4ea8a1b08b480804bb95a1ed0f242a85d7cb6bf957dcb7cd73758d093cc093de51102494ad8921c8723cf5d1cdb0e6c7c027e0424781a2b965d4ee9b629833326d7b27983bdfcc1b1bf0b544757f4595863d99c31bb21659946ee839c8a320388f507ffbc5d5f1ccd6f54e9b777e286589a30f33a6d268fb061e4f084ad94745636476af7e120f7fdb99686ea12285adca339235dc6f27e94f9b7d4d19722d06bb65ee409cf838620e259fd5a204b169d65fcc25bfd54bf555d66d86b23960c7b6316480963097ca91aacd5ee7a3cc3aa934136be8d94df364f9dbaee92760107b6472382b850dbba15c8e3ba3212c8a80459f762408dbbc211606ed69728dc1d92a3c31515b9d2ba08211702c7f127940dc03e0b43cfb1f90d45ee98e26536632fb09596e12cc58ab7c5e689157c7e75d3cb75bedb87ebd4ad6aae0172d8eac97cf50a480b3797d29f2d86c838413c7b3c4dd2a923c170a61a71ea3bc6e3035e4110c9377e661fda9467306f6ce83ac2a6284879de3d765948a2207c0ccefdd6991324b2f4e82fb6f60358b200fe0bdb954b42921bdfcb04ebcf3fa43f09a973f0f1155fbcb35305d8a8404adb42aabbfcd5433932882083557c3a05da55b1d27265dc34ffead5a1c56468f553a20263b4d5a1fc1f5436bcad07533471690b66e4a6c0f1dbc0f96f50e5da80e0c27cb24c53989d1a2b501c1f3c5852dfac158caa27be9e98581945d2bfba4139e8bcbbe705af970557987e69912fb6fea6f484f51f8b87de351868e69c7f36f762d2ae9bef09298097433e939331c529a01bca58e815aac02cca4237f3454de5700b5123c6e27fb9b89518da62d6224cdf7a991ae430a887c4583fc6b2ae25bf7ac701bb98c34dda5df9609bcbbfb4c84fd4fecc7b98d1d689e6b914c3e4cc2e1be17bba9e9cc617e3c582b8b8e00ef2081d9c8fdc36589752cb6c9e86a0fe1415f54481ac7abb1ec21271e56c335a82c7c7b4a33d1731784a7d10dc94c7783d33bd0a1f804d8a36654307d26fac21247d57d6131336dc24b268efd410af88b723c0c67000fe10e0f41383011fc8f46136280d404f51602f971e662c52aeb36d9f50eb521b66a327cbefba6faa000947f035a1b82ca105edb179a2c209ae8fd48a50a9a8c0fe42ec95447accce8ba1ebde2f6f9b09167b5ac94a8000e760e69127298f63a63d4c042afd6563030323c094370456480664ef8a95e459dafa9479476ea0f882ca83ac265ac08c652c09d5156682c864e0e463ac191b65a4121f9a0109f4c6ef52b0bf39776d9a4117ba5c0b40881492bf6a59e7b84a89425ffafbf399b2ca8fbdffe0e53552600176100573e3b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h7cc5a43dec87a2699226bab38297841fe16fa133749923d4d86245fff13fa81eb9e6cb5abbda396a0a13b86ecb6e578c254ed3be59d20f40a69c9f4c3be89a2ac7960faf36ae8b6cb47cef974230ecc3150950c828d5ac28622cfa23112104698218074102984e120a23b9857205753d3af63aff229ffdfbf2b5d2df0f75298b6bdcb02bc6fff2a0d099c187da8d47e9abac411211852fe39ee81fe57023b482493586abab18c4cae2a6f94915f4d69ce56f27fcdd8e48dbc3d9390619f18789f83d3ba8a49869600016ca360016069ffffa8e462ca715b587cebb74ab8d610cbf6fc8559e006b02a621fa20f459a283af2d30c1bc07e5d24f8c7fa1b470c326e1217f76c3c95d16f4dbdc5c9fb3beedad20b0c2c40eaf0272a7f7dde9e0281ed89facb928f239112bcdadb4e6f32e6ff905d49214f46bf742f94271c3a410bef74f1959a3a87ce6884318dc49177bfafb7aad52a5c59f827bcbc1ea6f54a06026e12b760803a3039d1c427951e0802a41323f95bbf9a93d8610c05b3b18dd6919fe736923707f05cad4af9d6653f275e44ba94d39d0913557826e0613d92359012d396ff2e4576e38cae7352a9bb50d133b705d3000500ab83c678a0a056306508278bc251c4564da4e294ed968ded1b389e801930016ae4f4a8082bb926e20a90b6dd31c82ad508ff4e56f44e08f2b900bcbd2389e778b441423a7603038d4c2ecb97973ed13937ae666132f62f6e9823fd2c49b418eb86667a9d0a42de489f60ca72eb6823f9cb59dc78456fcc32056b7586c730cb1e8ceef85be1c4347b05d0371465c981c71f6d63a5cedded57180baeee78d5d9f861a9481b5c448da957f221034fe17a41388dac27d11f89727b530d6d7a2fe1c64a9fa8f0da24be3a4b18a28ba2b9364d6431e944c5fd2c399a01e58a9f2efeb5b02b52c78bb60e3a40d92aaede62f05923d4bcf1fa2173767d818fe7191dcfcb6c97948235f137cb54b422d8c7e88f211753282c4b6ee4fdfbb542e05dffd4626936063a8790452006d285095062d865fb1c62dad2530d3bf696137c9585334ca46cab8775a8fd6a3805b8e55e602e94b89e51332359af1603d594a084726e9e24f1d106cfc826de0a36704ea22a283e2a8384e568db55a831f7b775b6400356d170518bbdbf1ad872e091043f565d9d0aeac723a95ff54dc745cc5b0e89af30d0546236635e41154f6c7882d16c30f920dfb4fc97a7cbf2d68a0fc5a2db15704b16d4320fc2fbc131243907dce95fcbce292442f0181e90213ab62ebe33127c8a2f575da74254dfd3219cb863611c74ab1a4256d275d1804c67f7a5c9ac2874addb4da3320f5ab104e478e993d2d907803786995b7b2ccdef37f0ed2437c684d8810da18539a24c8c6d2c88b48b6f467c903faebc9f38028d44de004487ee9774b819af22baebd135aceb7121a2b5b65d6f63e9a047319b93a4a3a887f1240336be52b51142d244a17d4554e9872c68b7839e2d634950ca97edec840d553e2618e84c65b56d07ff49aea0d581a7db93b556e61adae8c45a696f3983292d46e7dae5648fc34bb1b444d629c0ad9c03b071adb24bdc98a8467e3a07e2047c2757a746a56a6ebb907e177c7de5398d2f3a529cef718a7b22551599b0e6e0cb5678a944aae438524db411b9e1041aff3626886b11e0f4830b75df48b849c4821577cb6e5263b096bf4716c391550bb3f5aae3cb385ba190b7e384ec4fcae0696eca32239473e5d3d2f1acc5f272dde3377b9685f1908e3403d7494d5a2356757d96b4393c0dce58338cba69dc20fc6c343ac08941cc590013084453ddf6292b7b33bc3dbb963b588f7ff5cc3f292f1ab341a643966e655a13b61a87e8408c9aae8523d9ca332faf06a12be2202693e42fb3ef89a3adf8cca7741f53f68cef2a8ff4757c6e93686ee75f99fcfbcff42614009dd923da7869bbcb03dc69b6a8e7751fd4c78e604db6c72e160c5c6c99a972e1e89d0a55f1debcde6249fcca30469b8f2cae82d209bc87360a4fcb7376011600cab9e268681b694119c3d857f44945d1f8bcf7f966ea2e17f4725fa2869bf4e3fa27ae27ebca941818f5bfcd25858d35e992e86f2e5547be7c149d66c626fed7bdecea8de34e67cf2d85f7a33d003b4c26900ac8c7084fa59ecceea9c3750013a95b9b4245904536e6ded901769c362fcf9e2fc1016c1197c0dcc2b4ceab244595a62a14f99df91d307aa5c5d11a3b9f29b5e3db6ded03a0be2366cfeb1ef62336948de93e0224e1f1b9fc06f9211d594ed034109a551437ff46b164c9335a289af3e8b920b93da0531a7eba209cf5a5f2a625f5f7be4919e36287e494dc9c8e6e18d64d48185166f39951b04feb839e885d437f85b2c91c2b8c2995bb0e396877909ac8866462602e3a8ad6ad5b9a0ee907fcb02079f4ead5ac31255392b7fe7a7e9badb10d340a925a186dd343284b615bf8683851e32caca8223bf6c197b74a8b43984f58bee4d4da4c9641ec6c552b6d276dbdcdb9d1e048d8b152c44f06234b3ce5df860ca4865b6ff705454264d026a603f82195dd120ba168697670caca481127411f3b8d04060614c0a40e3e1c55eab52fb57b80993ab14c689000017a893ad4d373c2d48f75322f341257c5a9bd94a5a5385598cf99bda9177a2a0183ef5c1886082da9272c87340d20f835fcd611aecb7df07c9766bf3dd8788f76001bb5298ba04a9eb08b2b9bb2b4f26845d8d5f191eb00d91db925b9cf4b611a4efb46fe076a55600bc4c123cc3e9d0077a3d0eaf2e05faa9e375e313a8c8d4e434e11a92661678efdfaedd050a49e929055c8b511b67e4bce5b343a22cdabce8ab520453a5866d8bc72b3027c6f7d5aa44cab3dbfbb3309496ae42ddb17f37ca7c3a2fcea3cba54abb9051e1f7e16e9e9ad30f4faae50c499bf71daeed670c1485a3dcbae04e88b54330f062b5676c4c83190fd549b7a31220ffa62061216a6f2ca590c67081e3f86084eaf72a89069ace948640c12aa9115b99c4a81744e662964ae28836fab99c9bdeb3bcedad6d329462db2aad915f08cacb60d0af42d9b85776b842c2a055ab4b54f4be300ddf52b3b8b8e0cd5ad12b3297f7367aa61fe6ae1f020d6600de2611b38815f86df617e721105c3fb62d8f5713bdd362464ed888b8a6fe41ca1db3b486b5c01bea360487f7c68d3ee52f452bee53402e6e6839a296869bfb36912e4c19b723365474f184183998aa55aff712c5adb613fe0a33feb7bdd55460f71946c99ae08f8f5ba253957ec6a66217a9fa53de61b91ae0279dbe64a1bc5ffc9666a217e265e413b6571ede04b2faa1cbb43cb1732f08092a08a562f373d3f8c0b572e837ed42dc845f6bf40042dc8bb0455cb52b4af569ece9bff78392c7a433ce5eb5f631349e3167e58313431b41eaa4cd44d31899f77db2860bf7b7fea7647e3da108730003ffcd4132736d06fb7dd3409cc981959ffa160e2f5c46a54c742a5d6f90b80b950e80baf8f66731b4030c4657116e7123615429bf31e6d9320f587317f8a1fc90bf56149d3cc4b44bdeab672af53e154ab6c9dec8767ee14faaa2947bce78a9f608e48bd9955ae6b35af16efc5d59c81bd4ff2187fc66e511636e4887d69485adf6d74b2ec627f652c8379e7ab26b7a7b1414776cc0cbef8f8feb6aeaa165d167cf50e6a75a88a3bf5baedf44bd5b651075abd249b1b25e0166f14e73a0f98e246109859bd660fc3b79b28547c5782e62a1c5ada54e792ff717b175bdfa852d1de3efc9527561006d8593ef17ea8e1b59f1f791e6117ea5820d1f228d476219c766a2dc1b7ffbf3f5787e0e4117d3461b8671087e824fccdef9db50d5b737e84e4f45ece6d9a903ddd4e66b5951fee21eb004551627b52a6c4eb2047ddc546ed3495ba16ff0134353dc1e8662150a2b756df81fb4b69ad4e7451eba5686bc01abceff68484ba62b03f8218c8e566b561c52b3b6ebf3c7233ffb533e7bcf9529b210d2ce8cf4ab780e8bfced932ebd44874206fce36b6fa3561fd1c5643539c209e58cc372aed58c64c637fb8e9774c8b2cf6970ae35cdd464f1fcc4a9761e307221b0425f1fdf90b03fd5961d77917ef9a0f0a782c618cd9c5a07ba89b97707cc97c944822caf3e3190fcb3cd7b417efbad8be321f25fa8743a1bed363fb9d7e8f78b8235ee6204cd1dbb72b98bfb86c616777b215e54b1a8793993104deaead788f89061d1ba10f23862a96572fb5dfed248ebfc6c94573326c8b95dfd4cca2122b742ae05cb275d786ab4512663eb0c48de8eb9c5ccfa2c80a0486f078c5136bef3c40be367c821a8d5014e67f92af99a663abff0a857c9e303b6de338061566ae0c158f76ec9374e1f60792ebae985bb71e325419aae7e6d14b2dc56335e25fe5bb8da97de69a4e689c7b2cd2f5d70581c53c98c453fc89862fdbc016f1e9f06d5eaeb2cd302a11b2d6462844481da1c72541612e5c97ae2a0d383d1a5d8f01c2974862e1b1e5f5188c0cf460b992444eee1c1709ca489dfe6f287a227abbb0382ba8385f57921220c4d3bbf8d5260b41ae1285141cec40dafdd73dec5e604dbe3d3321b59968cec71253d1db112cbdfe9c4877480ce140fdd2b8a586f9d794e0169ca4e5b029180d54ec2462a2f31ba82b41dd98a621687baeaf7aa55ba9f415d2e5d7e634b9df8a953a73fe2f3336bd9887a6ecdcb8f267896fddf3dc929eb54f48a350b6efcbdc2413bcea52f65e389b18e57cc4b92b56fc48e5e81bc63edff133584fdfac785d18105faecbd949a8b4572de3cd1080ae4edf1707842e43469286d8b9be879a210dde9829fde658f0ae2a4861d8b06dd62768a22cb064641be1f441c660d691c320a7f382b553b761e2ae5a55537e81f0c1bda4dbf7c4c86083565ba70eb01b2bc46e7f3ef1955bad775e29cb32a188b8aa0a377c7e17f4ad201f41dc8c957b78c4b9763d2060a618495b809bef593617049119ec962a91a4c5ab10ff4077ab738826ec283c3daa9cdfbdbb4295c1ce965711838ded4296c32ef7efd19f41b6d99fcc66a4d7087d53e5744120845b55572ac7e26badfb4d9002e18d1b9d50105f39cbfd33ca6f802c27f92d57f363eadc494ce5c55517f94096b31d7090284f50aa5c700df1081cd52137f1b34c488c1d027187363941b4fc5f3875add7218ce7d4e14b59eca685f925172917af84ebd920319d7bf8f9e3b091f7a5d68a418b797f11b926f88dfad8512c2e8011fcf5da1761ecd0a5dd910ee450e8e786746293f66bc363ab2e6a133376960c602dc4b8525dcf1da75412e6468126160b12efbc50e89bed650fce5877daa4a390d65f006e458b31812ae22c12a26775cb653252a0ee803cc2adfd16d2f6e62e3a2b21167cc56ad23c9e4ca7528a4a5f7b05d2d5e720402b7f1a560683e9c1acf5c202d897827e10f22bf90de8dbbda7b581c89cc6209634899b5fa660f9a12fcbae4dc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h785ca9c450458410e6f0826eaef3a7c0dcd0ccc8c7b813fd8c556c63ff8628ec2db53ab658e0c957e7c4918f954b75b22fcf7323eb86599babc50475aa5516bf5be234d54e2ce8b53550519cc29c7f3a5fadb9dbb49919d424dd8feb38c095f0008337ca12ff244eee3c2fdcdc4ecb0eebc3d7a39f3e8032f079b87b4999344875108893f822853e9f386431aefea4d774b0308d2f35241e490639117138cd6df9eb8fd946a20c424f1e514c15a1715677ab03fdcf348bceadf40ffe194c8ffb0cc8ada7062c0416ecd982a0fad90b983b26c1e57f194d999986a6da3f18aeed50ca425ef012d97dbd6cb94d55ce4a17b8e8557c7fb3f109e1de0ae26ec7b94e4a75ec07dd02024c97f040a3f56c21e9a039fac2aaa6a609e5caea67f3a49315861df81ab4f2bc7faf36c5f57646a40bc904f8d7d4b1b2ad627024d8d3c98a04b5ea665fe3daa6d044afac570a31b45280dd105449c7817e848dc87b154417a92da366806d20e0ab7c5a1032636a2987ed140cf87894051314994f81a92641cb2a45c34a8c89de47f1d326a0c5fa31ee08c497ea87ed554826b38660c0fe78a6c38dcaf69c2fa2257c96b64a634c5794063485adf8b7a28e7b008b84bcbc7afb09cee4c0628eb981bcf32296c663705e6747fd68bcd25e140d2d1e4d3e470be0b7795c56afa9799e6ff649bfc121b96a5660eb093c9774ac0e5a378373d820bcabbd029179e24bff82f3816337f076bb76ccf9b966fc75a587f0ec3e1d9f72adcb3f5e3fb5a2032f663945bacd938fbef5548f7459171118a3f124dd8e18f654dd6f258b2d1508fa50741ba0c08135c9c99ecd9d92644a251362c365fef66a116bc41a27c5149ea8c2a0469eb0b61e716846925de265edc4599daa0bb73b6903d6aae70e1b9555c707740cfcb1f47ee3692bd66ac63a953aa601f7942a8dbffa7c30b2b2961b7604fecc058d76e511dc19b071c7cb25878f89cbb269344ebbc988a8ac69de1d04875dcc98aeeed2b75c410f70ebb46d57ebf24d13dc2e9689781df5f6ad6024acaa1f0def3ac99e7367a9c2782ad029e02cfcd22a682ae4c27d398ab8a2956b0e9bd37ae16cf2224c8edab8869b6651e665c628ab429779e9685c30bbf856bcff994242d57a23ed820fe86332b69e50b77845970300f27830e0a32e53236d37062d3e9a1f08c6e14d722dc58359d1da9862e7ca54ed0f225d78ff9dde5a1addb0776f0676a8f8466a108936c78ee48891f37c1ea67bf8a7bf4f53bcbdc36f1f79b1d1513487cc911fd3680f8cda0b1d403fd7dd37e9b5322b95da881870a57a8cb1bd9b2262226ba584bcec4c0282c5165af44b1c125ff116624bdb6bbcc4c44fe334c83f51296ca8f6387b03f2c98aef9f2b7078d2072aa30b2d315c8b0d29791c7068859b97cc1a7ff69190e1333a617564e46f087b0e5b6b5534a0cd67c8612f3bed1d5804cbb37e2083d80e94a5f48d8dc745e3b53fe2784d58f3144e78269b4c24f435c6e81e21919b531bee241e532eea2e38583d426f2e65e9c2c44abb145cfac7b210d9b8cd7d2459375673c2606263d94efb3ec6864e1361edb11eb3cd1eb1dcf9bed7f5735960e541eb706c88a0498a9092aa0974c53a71dc688e132e23ccd6172faca122b3116ea587da23cb05c4b4cd3c02a0a230595b6f6d3220f1791cbbf583f74ce30559f9682038663d4f68dfe8700c014d79389cdfe12d50c3223976e27f0a5ff6e81d7958ed83d750be80c1433761ba544cf709678b90526d9a3b499929ba1df764fc9ad21747e4bb460b8e59c2890421d5d5f91c70c72d69e9529c2a8d943709b07297f534a10a487a3e45e5f3721f01ceac9039bcc71217fbe54756e626d7b5afff4755e3ea96bc92a348f5ef15613e51bf8215cec63e2ce982938290c650f6a4e2e436bf7d5640dd70d21764f7a438218107602f86523e463ecd0addc15e9f38724afbd14b55038d56f95808a65933b1a49d28991af98886e1849e0a8bcefe6e8785e1ad37f1bb491e59178b10d644561ad6921b0cd86d54be5c0666f8d545939c6d8fdca77989792615e4d18216a00a648b354d60bccad4447656b4f0a7a334f0583eea7651f3c4fd7c20461765b455140c1154caf157e2948b5285b4e39aef2ac8c88526cf599fe71f06a543dad70a47875f264355ef02b2b6204e56fc728ddba81ab1df5d70a37a27d3446c0a5378658c0b90801b0ef2ac07ab877385a282c61b48eca6a6eb2c357bd8f3a1109c993b57ce1c73ce09e78ac18d760a0adee6ba6e35d9153516f4a183c45ea571bb7d8df3e30236ed74ceb4badf901fb6e746a900d0ea601d335a5f28702c2e79963f901afbd9d3ed5fe4f604fedddafea73f1063e898502b14551f85caf8a172a64fba9bfae992edfebcff393ddd20e46c0f863a39cec96eb2f44513716ac818405b2838c9beb48d58ee0cfe6e840ca75f7244b36d5382a1477681a2e5f9bc409ec62d297a59ad713b3361c63710a0b31b6cd61354850fe513ad7454d8d9569dc1a86bc057093abe81ce93223a847145c8320bfb241eba4430f971fc823e9b15d3838dd5d946a5fc1b0b12306e92cedf5a739ed70b61b5eeb4cdd48c7e64bb4fe3aadce0c5f4d5a7830ee6e34bd8580b2e77edbd1c23fa843c0b4d0d5e1d54d8f5dc50647e1968c1681869e46a7d0351a294fd46857f4bce16d3105ce618adb3f63af5ab7ea2692ca14c836d2e53712b253459e090349a717b22cb0ff03831d59f79771a58e542943b82d3ecb01caa391583b352c08c27aec02ca03242c7326fc1c3b0b30e35e4172a5dcf3a4bc2a4aaed7c47fad814e66232bfa9915524839e4ce14c9e0083eb32361befe19fb8f05c26e240420118725e5f02b1d971a91f048d063b4873c53ddd6a0aa716856904c8d849bff4d1024866988fe3740018f1b12ecd84c102b275e56fbaf398e2a1db0e8e7dd0c395d64e28e5b25a39eb22bb14d002e584698a69e86fff8526424de1305b065260736fa10b44a9583a99bf01d10c478c47dcc27af88ca0b8edd3c5b9a92a834fdeefd2f540c7f2e294b6b58455ba8527953bc9defcff4a5aafc1291e49a5a7cfc5252b881415a742371f53ab81d323ac925128277d58f594020802e00a4cf8fae35e123df93405d9d352c840de680a28791a65e7907ecfafcd1f5fc3bd04a6a8c67012d5becef9bc554a116fc02b9bb661c89f41508412fdb088b111e353a313fc5c451f46fd1729f33bfde2d83d3b9d314c081f448c6bd0080381c607e4be12dbde49f423efe5b956cb88d8090c6483e8f73a055f80f548a71c03c126111f769e181d823a7f799e9306d2923e79cf4f031b63b8c9afd51c45244652d97cfa1bdef3853f7d04baa752787371c5c31e6911ed739013d8c07c4e74babe8b3d44ef2c80d2b058b3a64644c87891d3d694db4b8d158188b862d16f7ccc13045abf559b8f0ecd09ca3ae6141f6e676c53151c8085202e21bc354cb554982179a359fdcda806f8bc2dc012c7a6f28b2aeab2ccf9826142a3967bbc03380dd63b2cb4131695f1e3f0cbf5e6806b259e127f5b3f3ce2d5d719de10c764e27102a45d5b1d71b4c6f7a083fe55899589aac0f8382e523d1b92d61c427e78b91a9a6ec5f1b04b878034308bfb6798480c6b12c58a7eea656a8762e3d549090aa925003ecc98eedc78bc3ccdf8a73fa1c91c667116d9a81441128ce1aa0d0377e72d6ee74d5f9df47628f0a1af35bf61e91f3e370a27a7b420801782afda300fb6fe4a5157aef95bdbc96af8998bd739088b2f6cffd2dbb3f0c9e9f5434d01a2f823d2d14981031fa743c5a1dd3cb932bc219cdd40a05ce8a97be85b319e76390e9c369713b5ab03cc7bbf3de60b39a7332477ee0dce04a92b32a689e67f6183ac5cbbcb8633cfbf5f7a0d9d909919a990734c1a0c0d4bea7b74f6d82c2448d888ee369850f16d8e71e27de00aef198f51109366e6f0195de6a3b0a21c596d7fe0f35c63e4e1fa92a7eb4b588cf3d0f155d2109680c6da2df451ab09a4f5f6b0d9740aa0a2fe3e12fba5d1044856127ff975b63310ae01b2def0bc5504212f6ee8ec3724c9f05eace997b530460441ed1229e6cb8991716cf887fa60ef5704f266c9ff04f42b122ad3b63fcd91fc8d81804174f8aea0dbf0f95f04af9f9f67fdf17c3727a775968eeedeeb05aff36a952055b8c8b7c770458b3fb4fae4703442988005255f8c29600998edc3f52f679367fc90298c49f79ca774760e883ed1210ee6a8adea100d0a2d13268f2eb4116b9d61ec4e8b212404892c97e2bf9db28875da3ea7212364aa7f2608bcaa6d163003a1fb76ac02bf7a5fa28d4ec95d3229b38d70f4f47f595dc73caefe536f03ec342128cb65f6cba394b85471d0876174a2a4943fcb9680c3980f752532f3293e62a9c2be3f2496465160ce95947dee2a45d7d7242a7fa6c067da8291df6c917ab9d6fd74e3a3708cee4aef7949c45b904abcfe11492b5947b6d9f638854c8d39a27ce233dfa4e5dfed1ecbc9ad864fe87eb9cbc981321fbf0212547aedca072cb9b4d80d42546134ca8dfe869b93d93926cd68af3c585777ac85444e6f741141bc4440b2f7c9b83be91739a06872b398d22e956f4095fd7d7032d429071d04afdcb37b1e633b5512cdbe8ba847d2ab4e02ad2f00bd5b39098d37d26d393b8e6818d62e4ecd6cadf1183ea68fe1e8d7f6b3ecfb5a121b0c4c1ea7bba522fa989222974c2bd954098519efed09c614e68def06746f70ca010acd69682f1025dd78c46431faec8aa391560a5a18af395e1d4d96c1afe8079785e4894efb2701f1b4c5b04309e47e6619a8b184178abe97854d8a888ac73cb26fd2a892548f038918ad10d1a01b7068a5b27613cc4bc00ba3f5b4b267a673273354ae244017b1d61cfcb4ac676303a00b5bc647fa56a210f40ed3c91612348f6e93d3a9f3b528f887cd07deb377e9eccd7c635976fd9c3c681f5f4abe63d6f1a4d897d8d7220abde47f6d5aa0daa972eb2741cea8ec1467660ad543c7f71149b4ae0f66b31598af5725db01da5ae082a727cf657c5ce0533127aadadd5067bfd570f8c3193e3a98558de3b38dc10761778d953749b5e5d3ddd09ebf134fb966af43c9cd2e4068917f0d44cfd5646296ecb027b7d531cc24832e27126f2193b2d8f9588ccaf819966cbb03af502b4aff792ad5bbbc9be837bd45b1996de5498f152233259034da6dec23269a3fa497b3695f140ac4b72af73c15680eee06469d9c530028227e420a721d747af3986b0af14ba7ae2081574cfa1d93c308362fdca8e9cf28c6d4f7f614770d09d5f3bc6ee033497441d63e03c9a286a501f641dca5623f986bd56fdfa91beb36368e59a11ad3424f6ad496559423dab841aa93538943e380cd288fc93d6d258b463fc86bee6bd54755af059597c9145a381d0ba3a4544ac9be61a15b1feaa32986d11a8edbc8dd9fc8a82c6da540a496ff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h2168b0f5de3fba85bb33bcee1e8141c52f909ad8b1d3520e4ed98f32907237ef029601d88b261b7717c9c384f5f21f394a4c39fc5e2369e0cd508d00e2b6154af6c423c48a5ddb003135b7cfdb65a5a7541c3f5905de3b62f71abd37ee8c7001100f2a9bb4c13086c07a57f5603d842d6f842373dcf4868b3b547cffbd484ea099e366dd1b08ad8b8d9f45714032cd3c217874f6122a7b454f00d6fdaf1b948960734272f17cc01ffbf3b58ff1e1c4ce9794c6ee23419a6836c78ca897565100d1abaf83a9354b324fd6a1c8e1b19196ed5c71518b1006a572432333e73f0f13b705d01a1bf7ae3cb584ef3b7923c545102b5890d11df8d072b93ece1687282c5b80b1c529f04a63ab2153c2e52ae2832b87e3f539744b79a5790686269520a43d012bf8d56d5fe875ea6bc01995fde4c0729555b7b47a0b19c333baaa082bccaec85cf33a264cec7e0ffd676d79499857752f5e81019dd5c243795d0b91adbe19f970ddbbca70c4d611b0fbb058417eb4dd65560e93956a02795257be22477145285ac5a1a2e8706a57f4d1aa0c9192831724588f554240b934b81ee832baad94129ec4468b27db512f89f81ddb993a7d60e72a550110337be221704c28e815f5f965830397cf27b6237e5918987de0c140debdf967ed3c19525dc0fa5676329040dea120a861c3bd6f7f76f66eec4e2ec59cf38e89ed90436ef31165654bb125f0075f0abc4186023eceb3ab7ee045c0c186214ff3d58790b183539235f047f6b8db18f15e4861dd75cf52652d2ebdd7a0a67ae81328c91c955df47487d1fe971cd3ed11e260b23dc1b4601c49b8d60cbf4bb45aeb2eaf1401bda95432f2e62f2e8c4d433e09678858a74334b1413080210e8b5a5708200a62e2aed4678c0e751e5b6ffa50ccc007642358b45d12e00578a43f2552f92b66c834986710f515d7272a025a452c7115896f4737b2ac7d0e4a13c80a74e86bcb86314ee826a8cc18b1cebf0fc8bbc6abf341a9abfe705ca97458b1647c1ccc7e01d1c75aaa40d2de8ff632bdd667e39e7fefc63122ff29016db1961d8660596c164ef1c6af84dcf093d3eee2908c48806c14b030095b51aff50b4ebf6c31eab89e3d924fd05f77833a00752515edf36777a3426ad1bc9ab90c69a880133b475e34b1bf51576eb885f227461dee1bd6f5ab46fda2a0c9d25fe47e3c1a3059873c3c13fa727abea1f20cdeb4300de5da7e5fe0d1fdffcc1a50c528fab2f18b23cce69f53f76559f170e98b9403e92efaee5113c9932ad15152276a1c38677e7038d23d3f5cfcd158ce1a29e234f8035e85d9af5338021fcb8edcfa3943272e454bf3c1c74afd41068d436b680e06ebe3c6b9083e12ea6123812182de173e352d8f4503c2705c7dfb74550b3af3bc498691ab28641ae601ad3c7e58360aa4be15a64e0f6ff01a4c89e177afbec0600101f7de29457c644c5b13e607aa66af0414893ca2323cc36d6bbdb9f7373732781d66f3d4b044769796b674559459daaf1791b0baa3d0d08da9a13a23959e2f329d89f562f56c9f960fd04b219036ae9eccb7451b55f614939ac529c2eb36383f9a32fcb655fdbe3af793be14de79a4abac7859644d20d31882fd082c3d7fc2255d2557def3c14f41d16efa8fc21e53e654690365400d9b5a64c79e57ea3b60d7654678eafa59d83317ecf4bca8d951f6876edb6c4f80d15373cd62d803e34a6d6d6051bf883f10a9c1e0bbc05a9c391341970eb676ba0263465a5c196ca791ea99fbf2b0342e5dc6ae994fb781dd4227109eef619d8dc240d13805d985420ceba607fcf28c1b7da0bac4cc1a3ad2fcf3b085efc237e5859904cc99336d1a1ea130062320eef56da351782b8839263a05e572508181fb8ff16b0ef638add646a381900167aa4aff58bc9fc12e4fdcc78d8051819acfb67593ede3fe34553bbc67d25449f4c88e2bf11e6f1e27f5a139ee74b2dceadc9285fcd39cde5e79fe4dc1d760f50caf39174a67b9afe842c9d04510fb9bee97c07e0869e2398cb802332c07042e268927ae75932de873b6d416b08addf3aacb989e82cd383b4d3e1e7e2047589d5d63eee4932df4d720c1b42dcee69b8eeff41a55c176895101abe9c69efc8da069434cd52346b785d05fc8664c5b86fe2ab7086a6bc27113a01f7182741787d68dd26e84e17411ba9280e7cb6cfc1aee9b462c9c6033b355c797d7d66838bcd6629e69ae62b5676a17695243722082d31eba0d58a796d0f62d08c7b5861d515349500147a0da508aa84125f614010d7f8cc737b82db4840499ee5c6f3e1acc72a240d0eab7bc71fdcae4630136b56b03019733bdd832a39829fe0fdcf500fa08230f56683f00eea6ecfadb82f1b276e904d3faa7cae6c74a963cf0772fa0fbd028cbb3f766ee1dff4c9342680e0f699a3e3d04ca343b54cf0d22b18bcae83b27276132dfe0e4d66098b78ce0b444a2e4f3fba81fef8d94832f8dfee2e0838aacd72bc6cb7649d1ab42211482a3887f5dd45d4b94d16a975f7ad563765315307e8c0681630a76080f87e23002ed6dd6ec7adccb96caccb8b7d0114009c4f8c708034888596e199c4fd1ecfa67ff7dbab01c7a655401577ba834c98a077f227a3738931c9284a57ed33cde794d3b74284b57044714c50f93a16e1cb460343a4e6b3a6bf15ce82d6afea4ef438298f5b11e95f4c4559d2bff214024601eec63608b791c32238c3296520b0938100d72491409c26a1220fb89c2c322d28a75c82405c308f07aa2ad860b085c1955e9c55c04506d60f5bd98a0f7b0c19fc6e4785b6d966ebaf4823780c83962d3fd7dbd85b0ef37b39428a860e1bb57f5ceae1a5aed882c3c03b3167cc7b1a18841e4cc4aa23573fb41dc133c666f2865c982b184d0563ffa8c3f4a2329a5d0e10bb351c983d5028bebc89d7ae5a0462a21764b0d1ba25c44816c7687a8bbb77588780e642827483f128892e240d5718aebc78fb3fd868b2b8cf04281768ffc53a0a332b8a3bad33ca0aba9d8e47e2e89cb9889fd94a41265caeed7bf76c1d4c3a2783e1979131f92903cb176a47d8177faf9283f8bd42bf310e66ccfa233752735cdf2ec3756cbccd363dd60b557ee9266c5659db3ed6350477f07b4af2bf9316207010d26c1b07fcf521e6581e30758e8a1ff161e4bdc834628bdb743f47d2a20d1e45024c22f12d8a87add168a04fffbf2aa2739fb420afa49dcf4e7217fa617080bd56fdbc53dcbb2bf3c663a86932938c1ed9f0b55f06fb975f19b191c4605d0a46808bea097da19e42e1dc36c9d2d3b177af2e5f4c0bccda6923e9874bbf8545d62b909eb0aae196c9c7634076f9bbe0738684fa6062689942090983bc3fa75eb9a4bfdb6eeacd0313dc8043614a8fa01ee19a5140b8ccabcb6d1073ee130254735c733bcd780332ca1e3ccad8433352fe50395ca15f2c518df574016b83b09f0b5e7c1cc2920084713a884fc724cc436f33f21aed62aff4dc25bdac4c0dcd757c44e350c4267d9e28168bf77c9b05e68fe6bdcd4b35259e3ff0f8e6d85e487a2df11dee9888dd2dd2995fa0550147ce2c48acacd77403efd9c1378b7315df128163fbd72b02033d06e382c0de9e02fabf2bdb3f40f2545be4f8b1285dd8227c291a160a2faeee5221347e97dec6f5eb55a2edaa5f7f034471815f8bc191d50b329afc3f8ffcc7b3d10442d36e87b87de62c46b2b2da0458e9f51faf82819835f60c55c255b8fce29cc7e911fd6972013014a35a05f2d53f478c2ace5820b839ce659eb3fe40b3693ecf3c8d5d1294fed3ef34bc15c9e2506c5375ecd26c742cc257640a363c52bf6c5c3f011a90dbd6e21607b66e50fea0821735f8c873a59541a5f59400beeefa6758356271f1c9fc139fb0e6df9bc2f5015df89b76f9716ae14fc2367e2990186fff2a4a38adfa7654cd573c5111da25b4d05533b3c455de8fe32c33b33468dcb6e2c9d3b5910f301b0ca3e46a70a0648a23245c2af02ed320803b0371677e828aca83770ee2daa74f51021d8915eb356e09593a24397abbc88f39f287e764d5a8a8a0612bd0fd547821a493cadeaf91840a609141e648451d47656800673e31bdc2f3d9fbb27d5791c8ad890dbe4a30ded18a4013365c768a5140abda9b59682dc6542e35de9a5ba43db1324f351e77ca95ebd5b5b605a8a3d93a49e5b8184b928e6fa8fcfccefce5a99e0c95cc4b95131d71a8dacbbf921827ad6eb50b962be6d7311ddaf066262b9147093e1a9c725898f6c6be145df389f0b8952f194a0eada66d56dc75529c691fad26eaae35fda1a9cdcdcda3e451c5baf02dd860d456d7044d4ecabb381843b8fd356abdd4c86d03ae95be07d43c5b72654d974a460d04151caf9d3383272436dede0fa5c6b213310c00b11e6b6e816761ffd216a6bb3961935607f1398c9df4979c613aa0a13d765d9b057de97b8320457e716f65a16ae1ff3b301f76bc55eae50075d1fe4f28450e600427ac033d32feac811d0ccc5f5a585d46b053c809d993610e03d4c705e99555fc31cdfd98552ec0f70af68974738c7c7543292479a31c4e06dc4c151f0ffb36c0e80a5343b21a5bdec048233b775b2312386f581023dc5e8d04a06f949b33ad23279679d34eb63d080e65de8d6ef318ee6a218afc5f0a70424fe0efb0cea579e30623568067066970fa73e3bc288b2345edac6f2b2530376a1ead8f76d601214e0b37531443685f28650c19e104ba9b72fa452b4b20d554e0987bce9795695fdb4e023ee6dd362973fd697e637da58a61110c5b673a19110fa9ce8cc4592bfddd8a4ebd8a3e6cb3074fb39fbe9d1d0cb570fa8d3e5d8e6cd1fea6f706f237a85c116d6667072d452866f8fe948f78c2d4ed97acbe3fc42e11b42b26893aba1548faae0889f554dfc63742e64fc5910e564898a1448474c5f2e020d3ce64befb3d4fd088e38a21c4a78d78a15f2c7e02b413f9cd4c470e19669d4402d45638182501866bab8484fa579dc79a39cb814b19b70fb659177c493f8ac4e60f5e6674325aaf1678ce11a7b5b9eea56bf2f1654f90ee7d7967b33eaf32054d79be24e698648605ba8cec3a27d65d0a5464ccb0945ebb884816dc44f854a15247936263751ea2cd8c319a52e7aadca1581513c3a3a6c86f14f2abd19b6984a903a1168688f7104c89d7dcf6fde07b92419c061b05ba9227ba632bcca22e929ae52447c74308a82289d3c45bbb292f5d17757f3687f471ecfd708aabf2da2c382ba75edbfb7b435f0bb5ed1a6c4b4f8821a1d4f7cd3bba253dcb29c4e377d5d51c307db83bf5b9ab7f9af263a1532371441715f2c504d51984907a68649e966a92138b2c5c4a5e7db7b02a095f900317b1c74c7c4a86cc565ecb792d8de20392734a88a2113e7e24a79562de0210c16bbe1829e9b88e6b2a64ac4e8e87832c4f948118ef77d9d8003c277327634e729ba445c00e1ea5a89ac85153042032578b6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h14c7db6ec8964b04d3d44b0dbeb70c54bde87eba30db19a9c49d0c86d0cb0acd8f6ba889fceac503d96b66f088f15e2969fd3940082ab8467d3ea84b5049635b6b39f4a94333eb680bb759450951ed8e6f230ff6e9ee83da22bee4dbdb3229d36d30d6fc21c5b0995130c009f335d57d94b58849cf89eacbdee12fadbb9409d54b865365dee06ffa542b04f6d996e7aa618bbd92aceeba5f5880f684b9e5c6c2b0545d8a3553f5f301b2506f329cbd45049890edcbfcafc77bdf671e35d5802db58ce6cc06bcf4f952e29e5c71e79164170e8eea357456bdfcf036e80408d0af5ee30a31551262daeb03e00941acb7690af54993fbacdeabc1e3bf69b66c061cc662e6cbad959c151d6ccfb49c4a60ad152b9a9c70f5e78f99729faef2f237614eeb6c764ae2d2ade3f9d837b369523083445e23c6efa6a2ff0528ce53ee4b06f49314c99ffca0a30e065f155a074c0abaf525bc51bcacd0b921520d3b278a46e430efdda31546b5ace39d78821a52de98cc6c1de4201e821fd4fdbc23081f0d3328394eefae23ea58875cbe1315363f0cce0a08f6dc6150680f3661a3a88187176ff4f9d5221b36943d87cd1461a9e1088c92ed63237cb38d3a235703ce086c0ae38e0c007ad1ed961732672d46c087a159aff5064a083f43a76762b98492c1c68ec439ec0a7a29766c8c5e174135699a22cc85ba9af05090921ae09d437cbb1ff24ab778a8fbc8c526a46fb4ac15248fa504e078b436bcc17c21a55e5befd8751a95191b9560f9f1304cb5ff3c84c9df5d59d7046e8119766cb73e4524d275dd9b4c7a87f3a103c4fb55f13409d6c85b651276cb6c4aad4843acf4ab13b66b1e728ff6eb80b76973c810527fb72fd5771ff6581de9167f254522f3ff1cfc8ac105ae23b27de877f8c526bac8655b9d4ec7bf3fed39046e0f9ce55bcfde14e6f6dbf409254dbf5a95a992229f93698f1065c7feae1d6bc07e044d1b4f1be41f2990ddd0e580d52e602606b29cb45b5aa2319478b20dddc5cec5b4ef3356e420f07635dbe63c5292866206f326a24cbc6ffde1879ea83338bf3f148eb415219b0aed1ee2f26552178ab66a79b2d04f9319c398baf896f953362203a2ff451d7447135635bb72f26a89805d7bbb2ac61654084476f2eb358afb2f08f1c0ab38ccb2bba968a5a5eb056dc6fb525ca57719da6245968288c6e29d31f7cbef6361b9e304e50cf56d2d84a38767ed16cfa8e4a5a990cb22e74d8af5968658e3203284237c1ac7cd5e3d16bfc0a54b9a359d62df897f240fa2da65622fc38ab0c6109e69935855a56314e0018446d227fafffbda7402a7ae56f90d86f6b6befeff3e1863c2bcbd0709779177d668bf34bbff1d0ec0fe611216c6481a32328a3783fb0c44ed7e543dd737c6ed300f81132492b09f30c2affbf4537b2bd6c8ce9ac7f7e11bc054129a7e02a0cc7126020add9d2de8827ea51b732f7891c82903b33001b9ab011bc2b5d96cf4168e90afc0f4a7c637519f4b8b2951566c4a078ed7852efd20ddad6f378d961cf925fac61a41bc255ccbd78e602deebbf3d6463971b32adb8559db81e7fb97cd249bccc6626b6099ad5b0914029641f04d19f8def505c48c5372748a880332d91e02837c39f2ffa5e6e44300d9986b57b1ecdd11cbc92f74496a6f795d19243289f65631c10e6ac3dce19ca2c9fd0f3df3e9c20655e9c9e37e3b6757606ebca2841f1ae3f5002d98c7aa18271ddb1c376d9f6bf055d1a3fd2e94fff8f56b6368df1eca83bb90fe303eb31894a70ef5ee4202035f83f1fdc86d3d8acf2b3548ee66f111a37b77ad5fd21b042146c52c70f30ddb859584571ab3c51063b9a47e74f70a1fcd0711b9809b741bfa29aed57530cf290c9bcdabd7c59813eeaf6cf5ffc030060eeb719302172b93c6c9e724c8da57ef7b249846e796412b2fa636d5aeecc3e6f9f855dba97bbcf27ae2ae4a166195c93dc2157b9d035a013a69a85543c2873bc55d45d0afbc4bf0352cc4b8ecb6209f155cd7ff5e1632f2d3faabdc0e6ffa368c6c11107fc7a39c6149efd810e186f3bfa40f692c8d7f952ca66026b1e5cc74845aed5b963c302c2a9cf5d9d77befa50b459c1902ef98d14e4863c8a7c03147edf895ead6628957012f6835314b16d75a8cf0be2c885279333ec275557a1d134b4ac30cef55d75de6cfed06bddae60a3983d13518fb227f3d9996e6aa3a1dac1f0ceb87c814214fac203d216ea77cdf8cd2f64b2a792f4380c33c3ccfb12e0443555522b16c8b70259a6a59205b167ca4a794465b0bee5c69ca2b8829ffdd378b843f14621f6c7e83c06bf32b4bd366d53555d0f7d8a48ad95cdb649b2d50c15ac5291d9f9f110bacfd90bb4ef8a47b59e0e26f974ff3ea6442671b11cb896ebe07fa41a3d500a5779c2ae7eaeefa992f2c91f9be8a5881fd37aeae4da025fca96d413eae3e2a3f8aaf130bd94e7c992193625ec15caf8b0a8a0f07a59d0922b36c4ab88db0ff2003e755b11486a6307342174a868b287279a0e37f1becbd7737993ff1b5bbbc5088385014847104704dd6ff0c9b8ad9ac8fef87c33ab9f56660a2c534b4cafca7df2cf95f99fd880774576e25ce3d561852e57474547d486896fcc2959d46f1e96dcf14c630c5af50b6326e31bd7065bd8e3c7e8667a362624207ca3fab6f76975497ce26363579c1e9df46abe30c28a9db3418e34b1b8813523686c8ffd93a5c44938b6bd73def7eedea17df69902f48a402447f47698833c882436df9a273938c67e3778f56110fc4db4aed7e43bfff7f033508ea9da3e0456630d3371d42085219228d00dc7f343a63b562cf9b43bc3837af4ae4b9aaf09af2c4bf7f0e38167a5601f54b08f592499ddc749717cc3ee6b22685342689442194c06e5199b73e8738d34a9cb21d304cc66e8feb1829550de2f163b058e56fb03ed11d12d67880dbefbd2a5ce3a1fcf2a285d8ffc695ed2452e85c2ca648a20904bd476c599abaf56fef11687c6d5ec8bf848cfd75c1c6b5da5b542e26a24f4172c4ae4919fff3d5429c09f90572b63408c1398bec4c31eb17559201448baa7565a2c89344e19ff546cc15a338830c9bdb8e76baac77dbd9d9092d0aa0e9f6c9cef4f75051894baac39c17ffb1f625bf3fb495102a005019bf0eb0988798bf6abc882d117c90419f4bda10b3b1f68003f1825aecd940b3aa7e58c59e78eef6eb1e57ad174b957e5a44e682f1dbed9f0cfafb7e3cc228a6a38a24b13b09589f804c1ffbae73e94d167012b83a95c237dc433d9cdeaa3d93741414dffe7a78c09786c1694f000d92ba18708b35eaf30f8ee1b7da0d64dd1d5e4993b63fa5641656216d218c908e10feb131070db5b4c88ed72a3ea6780b69d386ab603d21063c58b021c9f6584d91242312a985e85e64f3af115274fd1d3b24e97ff54b70eb341fbce5576e572d4f0f8337f065a88c690ec3f85d04990fa73feef82237d700f814eda64c0f25743bb754cd9f321f5a0d29dfc04c90badc2e79f419806defaa518871514e18633d7e800d709aef1915ddce6db3d0d306eb1e3dc08e65d51c3dc3a2ec78e62e8b549f563a4a3caea9bcade801b70b57f885a059ce748344712c10e05ac46287a24d4f0f86b2a8b00b7687f86e138605e520895e46dc4222b76871cca8d0e2dd86aa1eaeb3047e9579e45025bc0aeaac791264ca802b6b2841a7131500b710a623fd2ab2f0915c6868c7b1cd6335b4840a78eeeeb76f1277b4d70dc9064e242ee1c54b23932091763e72cf3241438b77ead4bb61de0dfc389f30fafc3f11eef88c0eb17e3c1640599259a69e183a471a096d12f0aad0e69f7b977e43c4f45469de1846b96fc9ec6299c0e095b4bd89a9bb7bfc4cf6f3cc006fa9274035623a6a74eb0199ce32c793e6ecd799b0f22e25225fb79a6d83abf708a47316e312f480b99d3166c6b5e4c1ecbd098fd696f64e9a496a31283ed4a54beb3d502e31f89cb9a136bf7bd1ca885c8caf34f773d3442b97d3e7f42600d38b82e26f0096578326016f94571a6c017c1193361ce909b713af94b40f49d4fc1a3915f684e49738c3656220d54b553e26477dd481eed0b7ca20cd3a24f94995a04ff99ff06f8e5de7a0c78f1e8261c995b322c44ae9517d2c68ff65d4c58784f76e212a0566900f22401435ae7f94cf6f9553a5ef135a9bce07d2fd890effa04149b211d73885f74c3cd4a9629892fd0856a80ba4af0dc03ed158ac787e286866acfd1d89a3de2d26e01f374936cde2f2bccdc439b04b37b8bda805239def42c5af6bc83b0ef91ce396a5076631da154c4b4505f858e3f57e8c6283c23ac656b8e2d4cddb5f86503ea7f094e1fa2b49532b88d754b1d60d324da2c7e209f4865be5de364324f6d7af83feb743dc7179a7d7b5f7fb5187ae2268887fc8f820259ee5eea283f853291182a8cacd15efb0e80f3811baf87da55031c4561116f285eaf372cc18a46d5bf22c8f93058d45c5cf08bef2de5cc4a5d37890de9a8f06b2bce57206b5a2a26e3ea38081b9642c22904c8f12de9f06e2a070cd17a6ded89123a5b89076cdeb14057b339a07331b077fcf0252c343badb174d018da5f02912531e8be8bdc35c3bb657d95a0e7bc9c9d3d7d395c02df44050d7efa59e4840f6c79b0fee91aaeaa5b53ec16b68acca81500bee8ebf7e34bc0a238e502952d33bc17a0cd07d829ecfcfee26b898d9ecf51ac02990adba85cab4b2776b8bca87fa358c1eeb001f65c224caa2320a36a3a2903ef8a794362f5b5ca6d565feefb4edeeb5f7eae5ce3836f3f22394d889c804c2f708caac4fc46836b4e70e65aa2dc351d478407baebd348f2cd06772fcc1b87b3f721af0a3a2fb46f78e38fafc6753bd37e2915cdfe5d9c43fce295d4474be1d126ebb1a0c96ef3f8e3e056b947c743c03130e78fb5e0e082f5f243c1d4679ed9b5227a685be5846eb5f42c2cd4cf64a0dc69bea20f2495b2217deb0baeae1b6ea7f858d7e3089f2803816189268c18d0103b79c136571039253efe2934940ec6e516a053cbd0862e02b51ca3f8d12fe1ddca78fd3cc497643fe333c043787d47645801ed66c064f652757a429abce94df06d9172c448f9673f28e13be212432c44d3ee031be71e81dfa724ef3c3953df9c7db496ab15aa7c3648f2c593ddaeb051a4dc8758f855f57aa36eedbe8da15b2c14b2ed87cbf15c4e6e45269124ef75491502e36ec38d0516d538ee5d144e4e3733dfadd7a94903525059846a94f7f70fc0f1264a8d31955c965b2889d04bdac5892e1f501688e11df2e4692f1206512368277b0669b3cf37ce002b093b271f2a49c47b369823b5676cc459480eb0bb3d3fc862a4967d38e7a498cfaba1091adc56720eb9d0fa86c41060254774e45f69e2dd9792fba0ad07b99c6229a875a4abdd29433448d55369b498eeba5e45649ca315e32856400fcda95bb7950cf084d321748ceba0e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h6761a273b5b3d93988e35590674f1bd25d4fcc9461e7285f1f3fe03e624a78621ccc82b9eebdf2216bb80290295ab07d99070093f8f7c2ca3187e8293b71d3738dcef276bed31086b7aafa449a8d52cb37d11167cff37ee78052515e259b11ef18e207c2a1561095dc3b411f533676602685d88c0b65cfc46daccf4e0880775f3f91fc18e225dcedcaa9a74655703c5574674fb7ed5761a6fdc6f20e2bd2d59d4683331728c90b08dac555a7cc94b004ff7df7676eece71a9f986a923fd3e292e88bec338cd5b4c2a2a8b11920a426b0f2e871f1f2debb7d63ba4578abc3cabb88d505723e45d44866e39bbd4dad719a4954109097b9389d06d7bee8807f9adc2c07796aa560cd91911cdce8f9f32052e42f10ebafb36d3cf0463e3ec962a197925d41686bbcd40ab70c3d550a243f498ff42c0b597be0dd091e709762861eda8058466978c9100a9d541deadf7da1e950c57cfc1816f10de19828269ed2a89bbb013f9d5074480221863fc1f1176b04cff46ee14fa3298cc40f5cfd771f5c1b109fc48691079298c1f2b6c58ba2afbb54e1c8deabf08db04200395a7fdb2e120e16c2addfad6ed31fc0b09d87cb2c1ac4927a5e66777f61cd7d6cfa089abc0ad59e58464ef04cd1e924f6a334df88d1b5a6ae905bcbb796929808b2c1dfddd48b1d1808b998b33e11e0f00f01236e506ef3b6b78e3ad1ce05174ce4d677b5aa9ce6620953c4e7614f23e54bec90eae3c995180771ebab52cf48e84385b38166e9503a95d7c179ab5fb0d9b003ce18529fb99653b93968b91096a8c687b30d2d6f77b35d7da886d0a7d1e6dd9a5de353635d2abec9e0e90771fe2154a5c5e8c60abfb9f82370daa450572c8774b774ebe5441c6846256982a7ed9ba0bd477e04e3599be1dc7e61d758ff053c23e89131e5c58758ae8656d713ef4c8ad66b69c1f8bea4732a44ba9856987cd8ba23b48d55767632e78543d8b69f115d0b1e047839ed9e8994a3ef5d9c98a09a0915c3e54a98022869972548a97970a158624537847c82163e7ad91e406eb9dfac8e621a4ea68b900ee6e087abac768b92320c6e55a0e5cec15e0fb53941fa4f152607b6a902b1f0dc2efe3dd9ee92164cc30c233e196d5b7247d3191b7686a13ccf158d3f8d7ff8e96d715d9bdcf667f09f84c23c6489cd24630b09905b757a13467fa679a2578792a995035a55fbf09cf3c78f3b0cdcc9ba94271bbbe399610fdb974ea2b18b7b81ad5042be8e396721cab939154585ca61a36be648185acf935646dd3a1a395975c0f2146e4ab1a5acd6c44a42b7e1261c517e98e6bed0ff28d6df7d4dfefc4664ed8a09fa3f070ac2f643ee837f5bf3541f33108d64804b5721daac84bcabf0fe2d08c37afa4ed8c48d229f66a5a37d1a4d1b7cdf4bce02402964392a3d6dcca0892ccf54a9931c8f46a38cb1f0ddf3b9849bf99ab0a79b438f44b39efb6ee0754e2ca8a0366777cab9e88c37274759973707152ddcf3ed2cd96da05ec9a478814cfa0d8b8862efc81e09105a2afefb7f29b83d3427bb6b4598f31d27f41aad4bbf5f2b53117ed3d2aa6fc6c904ede7c36260d9a2ce65217c11618a949ffd0bc44413f0cd37ee883b3f9a8ce5b21d163e98eb4f6bd1dcf16de96ca4ef95bc10c5f419fa861c93d1224da656ad99f301575ff1d15914daed93aafa0c19b069c71008d0724ea09e52292f0706d4b0e1d268aedf2e11c54ba5527bc013c818dec22adcac29813a8892a343b6e1ca1fabbb475a61ee9ebaeb0bcfaa5d1889efd9714878b5cbaa7138f90bb21c38fbae7b91c1cfcdd0e6a1c78f485e6e5ef93210e311b9e84d8b5dff1c3b57484a63f853779c1c4fbb9737f2ebeff40a9d2c82502b14aac59ef10458f1cf2540bbc7bae2f9bc5f2cb8d8c497b117854a071f3cfdf9363727f45be462ea21e02bfb517569e663e1a47540fda63e8b9f298dcd8f905d96d5afb58fd845a82c36b8ae5cbe0c6e19649b8157dd8196d44726cac2c004567e3b730289f81831edcd064740a328245ab91bd37d5d0c421869abd8c0ece7fd60f58b1a3d4ac4562ef99c3d4b4799932cdfc935924e77b85fd5b9832bd84bf5edda58a86d4a04b08b42d4c7e450aa55d9081d9e36e0f1765eff313a3ff27a3d0073e1682fab8a6e7bd52db1121d2c5ba08d061d5323829f1ebd07276fedfbad0d4db7fb2c7b63dad5ac3a5b793f50b3eb91c0efe4be4f30e47c7ddfbe47387016819a1888b64179cabd1cfbecd020ed95a6f9b45468fd341b01562a3611a9b0cf6d6ca2f864ae845b89532aabeaa814997d61e8cc29e3319d64838223daa3343a9d3bec50b02889bd72ea7996c7edd96eaf67f148905005cb110ef45b8641c211398b74aae64ffde8feced1d8add127581daf9f67af35a02b25668619eebdbf4c7062c523bba8adec76c79d54eae47b9fb3fff5e60596d4c8ac8a9adb5cf365db9403101823433119d1b54e2288b907e7ae8e74620b8100faf04dab7e13857d50286463b73cbb3830ca40fce6cea028086ec9640558b4edb6fe18beb9f1ec05809b7b3ad2b7f03d2d989a79db00ade535c43c5f030eab05f4f05d041c61af64f061a07d4fbca52d9826841b443d98fce987923e25f03276debc27f73b681a6ce148250c5ca4d473852de6a22fc0f9ecc831cea3e6983059dac2dc15a98f93e5d4d4fd79c2792af022d823c8beb05a54b07bfdb1fef5a1c0b38a87a41d6ea778dd1505c893b8e7f8e7a8463edb933eda9352092378b15096739f8d583579a30e58c678c2a825487b425121522005d28f80fb25d1e63e871c994e086c802bd83355f6d3d69b18afd2f1ff650204b4e1376481eef999d9f124ee51458f88246f8c37ec3a702c01b4cd02e9482494ab93dace69d1af4def6ad4960f329f42f8d9e3ee6b521fff99fa045762bc9153660aac5605ba65a2cf1c3be0ca0634ec21255a2d06580113020b5e5ec9fa4c2ac4a048ba7f70bef45bf82668044e9debfac30cd0e37338a00fc9df8988f467714b015b83128eb6efe6660772d091723da07ef6b9100578b6e90be384ebf4791399e7f1e757cb7b748e6961f4ebe3e052db27ce11b93f47bed1e252ad0d4cc75e6c99ad4857c2c6ae148774df2c73d60124ebaa4aab58e4732b7d242f229a61eedbfbc7a80a7b8fb54bfdfb7f010b7b6ffbb4560fdbe49eb0ac8ada3038045923d31a4d16d550579167655c2651687d50b9bc416623a676e3e1732417dcfca42d3dc94db2cb454af0ffdb4cb8e5a3cd72934cc03501c1c1d5503cc9a43b1e31d2b1da9f492c4c24a5899043fffe8726ed51782af3f6d3b7e6480d3f57dad8b2a9d972b599b5239ae6e33ae96f36555b20a69c0fa612fd30c1a08a8e96a7dad9a09421b4fadc2b8d202dcf216c7606774c9ca023e4069f34cf199197ff02360270b5a2c1155e10589ff72818bf2227a3e29f2fbeabedc71d89fce60c7333708148e95e0f72bbdc2c92dede1415b19618bb1021f7dfb259d6b0ac6a77f01acf53f74d30c78dbcb9653a9e0fd8b0ad9ec9e47d93457e55da6fc30ee09019c106e76e70657335b753746272d6522e66a11a56cb4104aa0816ae7782d91bce0aeec14bc073b8df6d14174c9451b80522b4976de0dc74bddad73c37ba75ce0a7ea08c82e7ff2d03af7e000b22b36cc0d6e254ad5cc0738afcd844beeeec383ea28b625830156b91ce9ccfa53a16291746ffda4fd5b320f1f2a3a083aa1c8d94c76fe196c6d3c3a22f129aa2d2e5ffdcce98ffb53fb7fcef368ed88f0ff6d8484c10c7fcc5157fac0e137f0387606f33e5e0a4690fa1884e761b3213e3064a73a38569f5744bb7086fa3d33d5141bd3cd1a0b9bbfad5ec218e0f0bae3a100225ff5006306191f2b1cda4a2de5074f64c51bcdf3b7463a02f8b6eb0793a4380f043d3a36190736a2bb802b0bc7775e8c7680f2df22a817073224171ca488acc76758a79228f35da9bd5bfb74453e55239c2789b2376e4b56fa8a31a6b6974dd55acc13572c3c39aa5ca9b8b307fc5c5e437150f7a30fa31590deff918d70242464ce3d1ca6970f746e85e0f76f2248c2f16a7a5b6b5b527b37acc93bcaf20afdb0efdc1aa2bfeff8ecbf6134ea2991886f53abe55d676b0f51e8f5350b483f40e636605ccd4c1113e76b2a847d7831fafa3119dace7c987d9c86d53f506288431a44e237018024b762b717799f47470fc92aaf5c70e01d2eb3b633c12127e28a9d8eca0ad1fd7ab9f58fbdb86ed7eabf3a640c4e6626442725c3add0473fca38c62998c1dd7294f0e504262c399b62dc1aa4616e6def04f5d26ab8bd167421f02a59cd7b06da4e812164df9de2da146dc65c564d47e9fe2cc2a6de47555fdb47597f4c19bad509971ec2e251decf66de6eaecc19145b5ec7805c74ad1dfb8f2f4774163370dfa7eaa382d4ae7c9506d13d89c56df4cda46cd344eaa6c7d6c84e73a7fe5cb7f958ed0a278363e7c4f2ef91c1f31d3da17360626015596ee8a0b41c588c0a12756d89eccb42a917e3f25b293a73b340d3585d0504684a3305df77326c16da481f236cb8a636e26a319025707d46b167001b1286870efb851db8159d27e4b93f7d7ed8610764ffc8da8c78a75c532a59b2c0194950cdceaa40419637e977a46cdd238380aafda06a26e41812d22fc03edb7f4a34230c257708abc1d93f9bd7a4ed1471a91b504ace01d25dd5793ffc9f959752f0f2724a3b7081deff28354576a93c6363411ff1fb7abe1630f5f700212027272acffce8197ba96b51ddc732be07905aa713f25680cac20cf86dd728f9369f44776ddfcf7288d39f0aa4f5fd861657952fd2c470f5d2dd0ee2a0adcf7d72a645c888d042e3721ad1c41c26ac90e768062712c8517a74486a7c3e28f8c9ff90ee0d84bb79ce8d03dadf9190e87dae3b6c252cbacc0ff5696fa121f7fe7824a4bf19be9c654620958ba38d29d721e0c7079d2a092be8e203c288cedb64ced42a2cad39d3c1eaed50976ef00e5ae85ba30ba5a88d6efacd2a2336d00420975b06f5e071d569ce2cfa229d3cce809f914f1721eb4157009424e637d4617fa6dbfa6b06bdd0732ad2e56e3f02114ec6fe300fce8520841e351fefbbfad8bf65b8435762ff178216e58905948121f9c43afea6d51c4d5b47a12759a31a0e75cb5ebdad464bc7dd599c8fc510339036c6adca1b67dface3bbab78c6d63cef26f978c65f721c17e7a821449fedc3ee11fa96e96625cd93fb2abf49a17d031768d3a2473470ab69e3532a2402563b93e3cb6ae61ef0a8ee35eefcefef2f0a9afff94746115b38f7bb7bd0951653ced9da5548c714f9cf069d9f17ea3c2f009ea700a492882ab41890eb9bd72114be86959afcb5403615208ede010e56a032d457dd53c6de40389e8d323287e128840684648a90ecbc1343380b161830ae90778f95fecc4bbc21c93878b05fdf5b934d93511a5936422717735be3e824b9d2caf;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h21ec7245cfee037f1b5c60f8506c82d0ac748b7af25e03786d35296d946183e611a7803a1fe99b0878ba53cf54978a418e207544b26dfa872c8c21ca8e6308d68f6e3274a23b7590b693be6f8192aad30b41ef0dac567fb7d8af5dd12dcdaf1216e5b56c6940367b3c190648a54bef33455701477a9d7527a74516a49490771f0fd5776603d13ede759791c7cc5ea321508bcfb74fcd3d01cd0b1f780970995d2b183e2533cb420abf78dc599b145d4fe7013f2b853b530a411c64cd650fda947631d8f7604182fbe2f56bdd48f102b45ccfd434577ff71a1cc57f84345e0b791d519f684decfbce828be8596a0b923a2a80af3e45409a8db71ad46915005477707cf74082799adda0b06cd6fcb5f9f6f642ae41970ddc9b3566efe6a1d2cf28baaf5526203fd514176fa97cd4752473cea0c142a69d4fecce1e1f95416dee72bf06461d7447792ea4bd7107e1d3b137f5af94cb28939a793b798307e57bfe0c58c13df31158729ec5dd4946b504cf527addbf85b2a876833ef042481bb69e5f25a59189e7e17bbbd848eb428c92e119c346e80d55e2fe1e89785c2fc2a062ba7d574693940cea25fe6afa1bec0885f166a24f8f98652478820e339b299a7becbfcd768dfa11b7cb1d09a9d0eb6f2943960d01a951be709e866217a62b4eca1699f1d857124ea8702f0d1d812e5a7d64ee6bd15a3936943df5c050c841c5a27e1a88bd9ca91f15b163e5f56fa128ce03c7aa68539c76f67bb23ec0c07b74268f0566b597aff12eda9c5eb76ca243c246b176430e3b5349c80e28635f70f57cd1402892fe04fe5ddf4f8b3b43cfec9edb67d6b0cf8b3ea9422f04c24743f9633655995724dd7c38573c33042c0bef073303fa5f82c97d8d5165c4d11fce750627ba9ddf183ce69506dab5372065e416c2b171399fa354c638020c34bfafdb1b574ce0be5479d3354cc50802ab9dcbdd7abe2b275b5424c41d0013700342f32fbdcd8785e9776dcd2ea8a19b1cdbe176f00d580f624eed365b080b044c9686ef23f9f3b406766560e3b9bf5e8f5f8224b44967c2a2fd51758e26e65cdf5c5703b4021564982f0ca573066622f1fc5ac5aa71bbcdfdec7a2652d38aea3f548e1c729b79b06e5ce27ac3ca422e85b820a8261532327f1bdd7d3e23dbf30db2ee76645a6e9bb3c64f07baf74daf79135199fa6d3322a25f0f88783afbb5b95a162b1353c7b1462d51ab616ec1cf243c0fda1360b4463433d3dd2e32816084bcd34a8362e5680dd4b36c075ab3a48984c12f244dcdbc8f46bcfd26dd069d0fe2abb7c1e050333f7b49bcf2e8bad80247ca8f41b62f4f9d36a76178b3ea2993d731b52c681b76d418736086925ad771516aec6f8708351b68cb492b37725a8ff711ded5277c350afc585a08aa8c243265f7fd84c1c924c63f5f9f74ce56804621f68da80cc9e0deebe3fc840f8598754c6f2956279ed8a5962423569270225b562f5338381cd1eed99cab346a0a08b65af0204a6080e462860f76c31dfdfabeb7dfeb4eacaf410423b3ab7934162338c3efd91607d123d4969dd9b20eae2e666ab6fd4becf5cb70d16768e0fb929205bef8588f924ad0e3955b26b768b583c26879341956168a0aae1ea349a789699b8aa96c1d12ca4fb14598a361c2a170e53e2734a0ae1fe48dd1994dbc8e0ca7211d0aee7768f51cec395c5668481a45c627dc187b67e273e70d11dc1ce483c6f00984c67bd78e320602fe16d1cc591ec9a07b3e0026c413475c3b16e112fb67038f739b49af0004cce89a51a9a31574568f4a2ad5030347c11c3df5b2d91abfbc067c8775593a8bafb256ee91128e2fa628d948b4efa992e55f1db64e4fcd054309419cd3f5efd433d7d79f7d889f7ab89bc033efc478dd54a808bb0190677b74999d8c47018b5dbf07cf273719b64f9da8e5a25b5f3f14a2f04ef267f893d3d6fdbca1d2dd3662d74b145075dbe937a86d34da5b1cc919b78026e47de1004852a62e76a0c3695d942957dfc81fa00e9ba78e676322fa2a180d1841ee437f246d082bb45e6a43f421dbd36853f2cf4bfb03b77efd4838b2d096092e758538ec16ea760f6ec1bee06d581474f478575ea2d97d22b8400e4d735051cb5bb6f8fee82b874a5922b77f634295737d2d1aa21752bbaa5f461cbc779a5cfef600c3bea1549ad040523335d0248a8023bb5e10d282c4be671795c1099756bfa169d8dc9bb04747335863ea5eb5a0ba80e805a5682998ed3df6f2ecf3882841db9bb82c262a4318076562cd7aacfdafe227244fdbbd20c60146efdbb9cf4217e2a6bc970577348f5760b7adb7421b2959a103945086595165dcf91cb70333f23e0a4df2e204dbc933ef888b642cf0eb0bd207df92652492c05d4a4238288ef39e670c4ae2185b05a57822e05c2f0cd4516be168a98a76433885166d191fcb67046e0a16bbea4f087076970070d110cab6440ac1b624c7e4a210c91a475995a233bb6c1e3c6a687e7f144f44da778762a4c8ca0d54140b024a0d50a1dd3991e280a672b718506d558869690afb7583792f08d3da3ff0619207a9326d3a58226d266b1e69abf69dec5964ee1033fb017e7323a21cfaf38557d55b80d37c47464ed809b16c677dcf0c64a802154e9a40e324b579d07469946fd99f5d6db3f7869e207d4ef0066cac97f2e190009cda3cc431b0c704b38004a28339a212e93d11859e174c01b9d4baedfbcdf801dc02a48c39fc9d182fcaace5d47e1b33c24daa0b91d856b060269c20582d170f25f539965e34c3f6328a0fb6aec22bc9386cc9d7623874e6f3d359be11cd1c7a24e6d215178a6ed5a485918de0ffa944e3f310779078e362f199d288f8abca27b0312e2ed5094011eaf46be151f8f2a962379f38f2ee1e55df531fb6cf06899345cb30b1fb43fee5af5016a2ac60cbec4743c388ce4de43fee753a5dd53155e067cc40be97dfaf2cd644464bc9da7298b02176faaa1735ca1e582851b2d443f3781a6f83e38705f4a65c0c03bb113bb6942be10b0e096b2500c9cf14ace324b72dd6e6d602c5bc5876bcd554ac9fba6da5cf37bbda20a31930bb0a250b20f2658307d036e4b262c818effbbe9ad9c9d0a74043fe5451ed0bbff50fe898f9f70d4e0ef800fbbed072c0a253f8f7aa06d723554923082cc57a143b1d3e0694d02088ac77327ec1f476aa0c7ad177e015737f7c4375a7f463fbcd8569dab61025d25e056bc84873500296e9dbb34db9ea8c9305042238efb873f7f8f945cca65760d780a152fb510a1ec27955266655cf052f69a154949b108b852e60757f57d6a2139270323ff0587da7045948c042de7616080c110b2fe1f1e88142b6cf867a7637fbd421e0a96f8c0cb4b7cb0d07fba4abb4c3950a0cb933b206337533eac608664fd60e0daa3945a7ca1c5b4ebf5e4602353ce8385dfe3726c8d8682701d75743db65f87b5767d70c34cb239119ed767c7744a99b369f4383398d6421814d818274c9619ac5553ce8f4879c66135f42a67e34cbd20e607b9234865b39d8389f8690b904af13b05fc9dddae2b6091e7c1dbbbd3f9c9fc0f978812ba493e5938679a328432c2f58f01657c03f56eee4eb375f442766b395772d345fbb1df3f61f92a8bad767ebe39f995c9bf4eced4b32feb4a614612a5c537253857c6f44020a4a414608501ce5bf674a7e55a26150cd16a2abc5d1a29974443ce874651f4d7e64d693be760882c2592bb7fcd474e9c24ede193d0867eebd7e2c58ba200811bac1b9851bde66492846a2dae39ad0286d0e2625a6e27fadc7724fa1583985488c42933c6456b4677386021c340f4f18eacf02ef8c8ff0fecd91a87f242d19ba7c4b6c5f7bc6ddbb3c6090d3876530f0cdaf58e982c09b7fb9f351a7bd18e3a565df32c8b86b128239dd1a579b646e9b66b38f0f52725e23534655cbb1be891d09fc3286c326cfb72a0c0a84f83e87ac3cdec2378d12919a96ccf2249a671cd65af1c17479a3e64c785e3cc0180e8ae051302c77f572f147c15120388af6541e07d6bc73980f1bb30f6fd10f6144a3e1353de69f349d3ef286dfe73157f1170a6891ff741bbff47b7549861e0d9f615b5d181035308d6c57bf4cf8c880c350916372b3d3b3c2d3ab69377f8fa35f2ec4530714df479bfa098141d9f9266f748d2908fd27855c655cf039a6b87a82ea0d3171b29314d232f520ee66cc9c9e4e3b6b64a906d24b06571c2e3f5e35eeaae037c8e86da29f702bf8ff9637d1ec29692ddad50c689ebf12d604fc63c33f2c30ac3164535cac50b4d6833550ec5304b10ca81e8790f6a0efc353095bef584787ea25a47eed3e4176bbe140ef320024f9ddc4c9d535f4287dd1233b32f138a15378cb9d876d824eb4300d23c8a1fbee3b87e00e49cb9fdc54e9d1c15163f525599c11bd73b6c5c6fd8b512cab8c00ae859d31a4cd3da3bfd8e8fcd7f290737acca95c89e5ebfa2538220de3ba0e680232db3a62d38e0ba97e08cd0284b00d822f19b79c5025c6772768ee8a4911e9d73308890f195cac50bbb76d4479a34cc952208716614ff552174a8c12e62fbaa0455a258cdffc1fe4b6431fa5120a6790f949c0b21412a94264184619d7cb52ef85eabe709b5174fbe3998ad774ff495a4f1a4c6db8fcf27d690ca461de27da8ed53e0d06edbea1643937d15e4e40970d2bcfa1ef65d8fb621b7aa1c57160275034be822ebfa79fa697a1d5d7ea864d34b6554732da6907cbe994973afe6d9c25535fe154c6b72369a15f8f3415afd9b64d5715e77bff0a41bf2751f6da5df15c1458693659cf56c1dd4b793cfc88073c73714c256e3476eea66c79241639c093b3bff7d148e09290eb926d93abf97335450d6b6b82a546a8bcbb909bc80538b7a0e6125e780fa935ba556725dd61ee4c964a68bc3c1fc3e7fb5a891ddd199aaf4a72853572f64e44eb29444f4adc219efa7711214626599f87bff9901bf26fdad07882a90b4d29d446150fa677d7b19532c7b8a9a01bb213940c1e9db01c33c398fc907c3f0ebf5ba099c719912fb4bfda6b884861ee37c5a3bddfe862e4437e866a0bdd84e3535cd2e979d99aca654323abac7c449bfcce9af1b0c2db39d1633e6923f16f9faf40004bbe36531608a2e2b5ea718ab36c024d145df4936c7040b0eec85fe0378c153bf3a097df2bd51f66a79b64afc9f332d08336aebe1a3c99eb595c3d6ff6b4bdee2b5758c50ded2e036af32df4562d4429a9e3c52fade2ea58a0ed2b88fbb0c2f7712601aed1b89602d1048c9e42384a745a1712c9df8ba470aa9420412118814c8bec155a54c6696e45cd4858e650c5b5fcaa70a54f305a3d6dbfc2b818bec92eca46452838e2947cd9f997191c3fef46acad5461afdc411ff78191bfdbf6609789c364a6c82ce09c494ad33ab253be2585e6dce798d0a28e49df8d48a6dc9a6debe62e0dfb0094b3d5793b84a7a092075e7f72e8e76a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hf6726064e464b0acd683c6c6617bc07b6479d286618e4304ed7da762b7f7b809db448272f1a3f21a0ee0bda4b6f8431bd6c41f004833cd439031b0fa9eb6f3d70f115d795d54a2a4f966a5268c4c832f48d27271aff3e1ea25515685f51b297acc77eacb266766c5f0557f3a4b71d58cd12fc00ed131df2a09e1f08418819079101d99829b9f2c373b59a6db54131454780b0d52d3bd7a0a556a626d43027459cf075fb81d4dfc82324cf8dc7d68e82fbd7a274b837aff634265e57bc0af60dadd87245cd41b7895b883cbe4b8e76ba397c6b2fcf71136853c9be6b2b62352fe976aaa0685c9fad64c45ab8bf1eee0eef78ebe1d4aed8b2554f658c9d653de0f54f37a247f2408dff60a87f3fcf05a59b222b6710db534e3555b7e424c9bd9c299020d803f7f3e377695ed240a8f4d3b8767acc0b35b97cbf9b6283f86ec8c17f7938209c370dd10cee22c61034a2b7978ba3c35f9a6af8f8da78ed8c76c84e378006dd83b1f7e97ad6e76808c822ef88963904b74fe839da6fc8ea7794e885ac13749353335be84dd0010364c6ccfb3aa00ccbb475e0f9066b2533c2c7d82c01108eb99d1d70632df57fa98aeb1eec4219b8840895bbeb8d128893903a3bfd5a4c505e115fa7de4ac29cd678ad9569fe9327795aeb0a89b8e1f8df45f2069b9cdc4b3331097a42028f8f836a50d607a4c466873f7ea4d044bc19a7739fb494059841c44b8fb8f58f87d8f8f687af69394e2c71cbb7b0350a53db7283916a9171ccb010c8e0fa24cb95c2ccf24e58f5a3e1eaa49e29cd22c1301a04886e85352b4cc9eafa550c81afbd9baaeec6fb81adbb92ca2213ef07a5c26026749382167dd2e32e53a420fed6fea035240e0222d0de447b8b4364674ddb8b30f537b44e2f7e4ff8fbfb8e321d4058f3b86ccfbe45aa3a3dcacc9e979e5d00d6cde35853aa682e82c0f2046ad065c6c88b10cd6d688d6cc6cc3ad2428531bdcb8cf4ce9729ad2a20b0dfe0e6dfcf96486eef8822978414e08aa24a50ae980f5b4e261209d7633e632ce0796d0d1bc77bc8c52cefdf832e90847984128e58c8191800dbb7f3caca99d9c6a8af70e18acda1a6701ab9d9c520117f81c38eeb4e953d15584eac43283ad76b9075de72fba17e0ed452d78718b815b33f943b854d8b6914d98954679c21deb308277d6b803373248a8a547f352949c51b51f230c7b0f7c0ce5c3d228a4484f63fcc55749ca43222c30b6471d68e1506bf9e7405a8d17e026eee2ce35a9b01ee72c247a3a78d6fffc2ce948d056472bb18f1a0cfcdeb0b7f23700eefd971be980d7005b1d30b5b8acf81c469cad0c34e6af4f30848c5fa580658eddc38c15ec77f2f55cc08b5d694ca5c30339b71119af33307cd31045611bccebda2c599693569460491258fb19392810369655e009e1b9494d92bf376cc0a006db1b9bf79c064f36c164b829516e81ae87436ff006ab01a44adfd107632d230a4b61e8966b1b541f85884724357b0b6cb53f3bf8691ee653109da9fab0f2ca30fd3c8266ecc0930f2ece53aea59e8a195c37c1fe0c8b0ba73b846de53a9304c6149d0644c2589d1bb916972299d1c34a17193f5a5b422ee8b93371dccab1080687bba0a31ad65003b11b0f66bcdabce3246e80b436c18b986a4cfc43a5e091187f6a69738b101b0f2eeb23b711f31a439777434d2729b714c789c0c151bf4de7d7732f76ce75a4789b83d97278de59f8151ea06132a338faa743c066c9c4b6cdbbfeec227d3dd54225d5b28c6bc24bdb46a142a7de87e44fd04a0a4a23365e47d538bd66619692d3c7580aa38039bf8a0519cf2aca65623b845721160775a0e76ee772e0061b7dda8fd0f5b9efea0fb325a5d630c2845a7894c45dfb1c3a2ea7f9a213562318cbfece1a6f5c5e70af37d1124395eceb8cd842fe90acf5ddb0bde6fbe16231e61277ee1528925065c081b03950f5c22efa01963ab83379a9477cbc7188deef820c5d6ac5f8b9bc03007ee0f5bb5ba467eeebe0550396fc2a5c102844494588981d73798a5f93afcfc57e0502b8dbe5236c5ce89c07dae578cb3806e81f216b96de3c92756a2f7f9932e7a8494bdb115ef5f847da9c93a36d557b6c04d6bd890f7c7d9f2f65a4a8bf0c26b89ce11453f5d763724dac095341b561609a484638b2d6c910fe0b3a5017db5692ff7292ce6d5db6df53df7e185301bb2218e78ba83debee0c6f19db0e5728972bf08e550d9fd72d1fad33e0cdd23154dfedae608d70c05d4aa7cb5756d84a7770d0072bd974e9140ae9f1dcaf5e4c4f03b3e68668cbae5f6a39b0c3f928aeec914ecf4aacc14c53c868b01fd6100403e26abdd6bb04c473a4f5b294288f2760f971b9cbe0b91a1109e39d2d39826cb6222d45cc1e7bae794f0416ad1bcdb26779266a2c2faf403413a0093f598b7778f195401a9a514b61023fe977f568082c84424c86bba85ea04b69af3d80a7b85b9cf4c8eedbfbed6f369f66d1e8b4ea9858b10b745ac05513a944bc0de5ca43789d1be2d8b842d91741b4a2d8d5c5f03b98c3f98b318571ba5b130966d7ad352cf4c647bac736cb9fdec34078a70d9cf737926ae349d9e8bd3f692746be536701ab0164ed0897f6939d900fc9da17c6749171e62ebf5e6e1b915a5b4e65c6258492bfc0d74864aed39fc41ff034054182caa406496304fa13cb803e24617ce318911036a2cda10a46b89f36e75dd999531bfdec0708dfafe0a87681d0fb38d79e420efea165092cabedd1de9bf3edef23ea736dd97f8a940b7345d0af7d9a8507a2150351f21ef6b33cd0ce0556f18232ed4d3557ab2bc83dd9855ec180939d06bd118bb1be264846b0330f8f9aa74c559a02d316abd8f7f6783706bc70fbe4f231182c93860d160b571f92e3bcbadb71316a5c04a4c5cd37827fbace43b37f4db4e7fe00ec0921870e77d4417690ef877eba83628400ef5412cebbd347345f4161f155b70ff315ca0fd8837ac74a477e6809224b23c6ebbb83c7525c3325a48b05b56bd3606232ba94856abb7408dd9269757e89a1cb2e705741a6f7062a0fe5f6211a94117bfa968166a6008668abee67ce9f82c380ede8f4c83a57a64c1efdb59e9bb1ae727cb2a88fac3722cd5259bc58a2014fecc0d3987b0b8911ff1a9d8786eea035f4040db7706f29c88d8c366d22c81267e2a42c91a7750d013282a32f2e850949467a835e6cfc02c8d4b9c0f0a69ea81a1774abda1457a961ace72853d3c5c06d1e1d1624a4ff5f5fa069413d7df0effa3d290852d4221ea7aeb03c80394e75b51445fee31254f32addb15b92dabea9b0aa2d81ed26894e33fcdf65a846cb68966cc2bd59bcc7ddd55d16cdc61a39f22e0ebec38e48249828246162ab00531677cf95f55ab990c02b80a44629e4e78743eaa1f9f9309bb627f198d99cbf7d71bdd0c960393d6e0e9423a770585a7eb86b24aa44137dcf1c659eaa0526bed5f62dcb3506325a9ce644d7508b199fc55e50ed70ac549fab0e7a566949923f7d03a050553437a3cf2eb4f08c668eb6ecb9fe16043fa8a7cf250f17357f7325c3e9cdf102bb8d43a5e623d57c58028ae2f6c98692dc6799795aa357430e98636b57eef747740a60f6902aeb8bebafb28968cf9cee3c4e63ce8d5ca57039581ae134c2e0b916c19306f0bbbf201ad7250974bbb6336862028dd2074102a25dbc6e0e1417d603537e120cb4bc6d8c86b400e8229c91faac8a751d95163ad35f24cc97f92af5fca0515657f7b978dc1a1b30bd647598b4b939b4048266e08d0849545326027190e6bcee930071d143460a23c6bcb95d0ff9584067f9e36a2e2f7a92bdc2aaf07cf49cd9bf4b5f30fe2bc90b4783e537efe1e8f11f4d5cc0de22aa6fcb7cc9dd12891e77bf87cf1e53a38b6abf2ebf9602c6bafeeea1ff5b13c858e4676a553eb929b74c1b9fd2fcc5c91421b9ef050baf2477f4f30c1eb2d1ef824034d6db0a3203df1d4cedfc3622d7c94b16890c553bca010d11aed17e413e82929fa05785feeb07be535903c6f33c86a8b4e3bec9b37ee25e5346752465b44b174bd1be0bc70c0af247bf6e20d96908ee7e10cdc2b8b75c00f3082044becf3890e17064a0220e7ab948f75a06dbba64fe2a19ca31659b66e10409e1d18e644acc84b05a8408ac829a475f0d04648caf9ceea41fb07c680ca24e69ef0a5d9af006d2069ef222137b2dd6c44966682488fcc87ebd5bdb29ec11042df49a4a963c618f8b12ac000eb2c4a3d8686df4c6e3559edf29472f06688ccfe7abdb0d857a01f6c5b616f4eeddd60ac89435f4f67aa62cb6de3c15b3e76d5e078446c81a166798e9a8a284d6992a7d3fc02828088c60b00752c774185ca61ac990562a84f7f720c03db4e249627f55b298f5d459f4f9ce9e401e195435716c08d5daed80ddf772c5f06941a42556613eb8520b91335f528673b36e43f0d0803bd55168a11a004c6a77b9b6b3092b7fc05672f41cd94586fa9ff0cbeb08e7fd051bcdba2694acbfe68f41c04f4594a1f3fdb0ecf88284f217cda892889d0e3693fd89dcb97d995d97cedc12e6fb6df47fe3d17fb2446686a7f7aeefc1d7034d2dc76d1ac4081f773185f5267cdbcc79b4dfd144de7e9f9d12726b2fa4151122726aa171f5ff11c1de344798d1cdf76378f497a1a1fa9c8d74ee1a8437be9d934f30cc352c8a6bea5bb6c84b0f52e0743550c273f2c57c933803873b6792eb1a105d14ea7745385b87552b30d892e87442555d5f5742a6167da5aaf7625e8aaae2911659b37fe612a5ac1dec08daabdf51ee2d13474716aa9ddb52dff7e1b4024507d17271e7eb36151185b79f21f11fe5a5eb945d75146aab4e0b4331860766cf1f57fc13e5eadef75ec486b6612409655646124fb312aafd7600389497547dbe6cf2265986ac59bc8196fac7eb8d5cae100c121de66445f9efed81466ac7e425a45f4107294f5419770d0044af3648512449baa084bf6a83f2765d0404f44eb22aed27567bdd34fb08ad0e2686b6abf1ba9450efb437ff6eeebde878ace9517f9f0abacd06a7a5dba5a9bc9c296a3739f888dc67b6529f8a69039ebb477f813b6da577edcd73d7683a3141f237cc93ef728c6f68284251dc40ffa1c237c1916664e1bdb360c90886fb8df2b61abe8e4991d4f9fad8059455985f5eb6064af958af953f02e3c937366f18a84222eaa48dea6bc37f1168ee5851493ea728f8d10654db18ac26bf42a1c2c94164b3727acb852b3a1e6452418fb4d6d61c91b3e97987b069aece4c1293d72403f86bf2029612ff44249c71d0e98448d35fd486c1061b3eac299133784b59272c7ec42ce1d43ea6997424c27329356e85d43932c08ba6760e2c8e412766acf2e03b8b844d49dcc912c83de1be9b4e7fa7700ff1a83cc182e705c12026fa689514bda6d4e41b2bd6b6b40d1c501966f5c837941243216564183f8c1eee8ae859496570a1a64667aee9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hf2ecfa4143d3819ebf78105f972ebef5be362a4d04a17dfc5f91fcdc5d014be0725a9c8560817657ce55e381253d265ff5be8d5a2ce3a9f29dd4181e8469c83b236a76fde9d457b49161512a9c17e2ae8525be7200e5274b5939c32dc479d270193425d00aa7a3e5f61b49cc58b29a95a066bfd1009f8f858235a58f0e0e80a43288dc99b77ec627cae00bd3e0221f92a3fd72987b3452f714dbc8eaff02d90480d20c09cd93ef5a16ae7e457d6ee4625cfd9ec263a299a6ad209913ecc4eb0688adc271904b414916d6b988cf47aa61a05521296b1f519e40e0b68c9f33c4d0bd95f9bd7ed6b2b22788e951491118026d3f5ca9f4c76470803855b49582d76f8312c3880145d87911360b18acacc5564326fa21ab8251f0e8f3a4fbb3273e017df6bc3592f73310675aaaf30d1217d3ec945de294f9c8d9f07fc92496a204c30d6dfd2bdd547daad7b1ec7e26d773484153a55cf87e8f92f646156177038a43c7ca30816f22d9ffeb9d44009cbf2651da11540068cb12cc5ab6d73356ab2df9ef4e648f27e558b6935621a4f6382b5c9b3abbb2e26132e48d6ee550f76008d6f8997aee050770f8bc98f1188ee05ef30609f9543524a096f891f05f5f97d344b9ed5ac545ad06785a60fd2f121bda99df002fca86e1fb8a5fb9274a4b72b34d2a168299ab8acaf917bb4cc2710db56d726a6e0e33a20e678670a4c0258d0f025aeded0821a1fbb56c4eec80a41eaea9157e7bb3bfb5c48d2e346c81fb18efa90bc5a4e45c15b63b314cb0af78d318ba6f28c0bf464ee933a2ad1fa3b41dcbfd61caec74de7ad8d3e135a6ce8623f2bde6e08710ad1377658097866cbc93bd9fff09f4294981a40d04a4054f424e9989dd12ab5ec6e1f3452e8fd462497a4fee48be6c30d670091da53cf1a8506c84ca3697eabd2f190c0d4f994da499386bd4cac4467030ffde000308217d19da85e6d5bc5b83921c07a32d458fd16e6042d84e73e04fb511a7d47543848f0e70bb71d782f2531e2dd88cbbb9c88dea6fa164e3000b81174d22173700289b2dbe9fa0ac52af38b3120aad62db666ec31c657ce8bd6f54d1fd5cf685d1b962c30d8c44d925cff0461533ad811683554bf7db062d3daf4898ff8a13615f3f59a9ce7d06e4d455fd9c1082c4e4e6532d5521038ecfcd64d28ab6142dca6fa8a5a21a2acbe2946441c0874747e13773c9b07924b5da4e5dcea3bacd15a8f287809c06be687dc7e85b2f06c46c68025517405e0694c3eb9fb647a6bcdfcf47b546248c89f7c654680bf37330059e20117bfa41147209f1dc04bd0376bdd123ccdcbe37023448233d8bbb3c9fa71a0cd3b7290c5a88922ca9f8e7f8830fbdac4f3fed73cf8436943a0b3142570ef1f186250d4d2190f7e638a5267894d8856159425f40eb9a4162829159413a086fa2e9502e745aa28ae561b9454e54e352e59152a1aa46c140f6b4301ebc56d089d9b2e9d7e98f0831aec7111b50cb8578bd2d658421596db154e7f619e3d23957fed7f31bb236ef1b98eb7bef0aa317d9b48efd7108545e5e0cb599b898d0578f6f2d286aa2c0cd1f254b6326b64746c3f06d7be9416d41a8d7ab084e4f7283358ba32cbf9fdf392544d13678a46c487223d05b00186694973310f83a3a69c75545a820228c3a26de2876cfe3a4dec1f83e46d9af4ffc4e37578cb228cad7a67f36ab5b4d7153d583986dfbe38cbb472981be9e8747e6396ac19000b42050af64c1c9f51a87e720c170c055a5f6e39fd13e4e5c895b6f48c8c439efd3c65137c8c2695a0836af8192602493f371f601a2a68a05cd1a80ac0c79e5f03b632e01534db40f8c24df68e6508b3a057c91d20bdb83dd33914ddd84c2672b25d36a9a0703d6d5782223fe008f0a7ece0652293f10b183b8180f6b9fc30362935ae7cd7b0349f2acbfe7062edf5668cd75cbee95e08b995e672689b3e0d4910fb29ccf1d1a467afb486487deb543d779bb040c1f4b307027060ba82d1f2ebb1136c6bd32c7c68d6d4572125bffc1ac2ecc5d02c4c894965933d74cf8a55616c31284480ba110337f2b0eb675cba0453558ab0141250d66e21c54a6ee4908bdeec83c16203e3b70dc6c3a5609e6691e5d8e86d383f43f1ca56b64dbd95e841f98c8a75461e9d93f6ffdfdbef79584a6273c0ca9b4783139860dadba5b5b85723445630a6d3e172a4ed1955f44d5f2408f36d0c4c214258140da27e431574b6b810396837b547260a9266c80c6387872fcfd7739e09f366b8444cf8ac7735142cb0d76d8febc01620273854fc75f44bcb84e236b469e69a5824adcec52f6f47154e1fb6a477ef5997cda3fca7cfd9ea4920101afceade587f8ea34cf700500a443e4aa819a3282da23d395832df10d92930adc4a62275ce9cd4b9b4d6d6ee953b17e282a574586878fc07dc7a3e9c0ee9e763489d5ccdd6c86178731be2490e8c903c7af1f9aeb1d07340d1d5ff8e42f85cabaaab3886da507384118c0a4e0e153143082350af42fda0d84bac0fe01b6a411c6fffbe8bf514861fc97bdda642df751ce8f81f7954cee90b04401be143141cae99944c68c14aa2cce9e06bdf2eb65540aa0faaf81b28ced2335a8940fd3b1981b980ea83e91d9fe015175c02db1087285e396c94c38f7dcd8fecc84fa628f2550601f42f7cc2f64571f46db3f84440a614ba0a99e0138523e9f56b56ae51a1d119ab054576ac49e580966179eacdcc9a95ba2a687af08c3542cb7859ebd3dd494efc0aa70109616cb3683770f2eb3896355cd79ecc05370e53c5e202c45d77954a9122a626800eb98ab344624452aef636221421dee1f1d7485388355fc7d04ee8ecc6bbb47baf1708ceb576dcb3234794a7a504ebf97e53c4d40b57caceb63d121e5e7bded408bccb5a2bc99f2913ed1a228719a9e59135a5aeeadcebd479c204ed2dfa6ee9477fc2942fb76ef965d4dc5539264669bd56d5978690e50cf49e1bf9e5067b89f2a3486b02002db3faa07715f32e7736eaff232e8de319e7bd8cb7f578dc65e28eb603e58a7e51f45978ed77c1a46c9c6a3b48a7e45cebcb1ec1aa796555054e662b294fc4fd8f098128f9824e3313b1f3d0881eebd75be6d50ce3062a0b732ec5bc8f750471796c199f507de97bd06d91759eaa1b1e41433e2005fbfb4f195580ed4fa5621fe122f6e8e2b383b964d54c74e6ead26710a169a5a5ba59271211cbb699baad9c03dfb87f0daee03c3c40901fe0f2e63c8746612df0d297559920505d508f0323675a3e64bde29025c5af4092ee961506d5ea8b267c8f2fd7b0c80a8ad77ac8343836384a45dc3c16f9754775f9052bdd69e708179ac481ad08b8c107b0553c43af165c5053c721a902c45d7d9f215c885c880555f48acc0c4d3938587d1ac95d874c45d30dd801714fe0aa3749ea32b8389a37bb3507a8449884a9d8beba3b9f92022f9c931997fc11ddd23f2b79e787f89db3bb0d7726933d99d9a8ff491a7d19a77a1fcef35f01830252dcc0468e818c1899d7f4518427799806f3f4cd26abad1ddc513fb12d61fcef0b1cd781954753c6309c1a84903c60852bc4c40562673fb39139f703afc8ec73abd60d0411e4f184799062ca20d4674464ef170ce785d4333a55eb03ed62a4e373fe1e0282a6c006301d9761ad47b369da3d98673e327bc6cb528c8d0cef1ab5871fbbde184d68ba298e80fa0e4a4a16c3ea8b7b73163cd9eda2f2d79825cee3aeefe0b6c062d3bbc215b560927a2b176b19450fd35d6796bcda67dc502c30e516906577b0b51c15890dabcfb30b0d8ca334d3eebb2460a0d13087b8d8a26478d25695a0828607ed7ba76bbd1aa1769bd2979bb29a2493754e2418e9acde018cf5fe2ea0e32a2a7d464fd21e269f510153e3f86bff48a57ae10b15a104cca2fb431f63430ec88bc13d4e89708b9c32c6f577edbeead80de9dbbb243c57468646278f32f01b54b720e7099e5ae5147650197c3e5b4bb4d350e03d5a40d4f48737afa6f64e7a6a0a98591d5b4b10deb78af17bdd5f0d65c5e13ebb2eed2957ada2d7803a063dd56343d02ec105e361203c07708b556f6d50ac9621dd508d3cbffb69457c6dffcfabb45b3baccbfa92156f75397158161eddded3e547b116c1397b72cd5ec208b0db2f648c44bbcfd94659b4e4e865cf57166ee1b38a819870b13f7cf47eba561082e602e5c065a1dd422be535c846f9a870c6b8d1e9fe8c979a70f1e496067e914b8a1a1c23ce9e433dcc8ac36f49772eeba19fb3f1744edd03febef06c2a7165955ceec535b14879f19ed7c45df4b6be9e7d925cf76fcd1999e7e3f8c405621cfcdc78ec3be6815909163f91e34f78c116fabca3c007e723cba3fcf69a6c46a98509e7a4e8d07904a5a9f20087e337122b38502d41d5386844e2fa2aeb777f3e237f36cca308c56c96ed5c9e606b0b35f504942e0d545563a69d91940735162dcc837e83811a74e350bb594dcae4a937c0746d069ab8211e58f05d11076c34c8d5d8e2e3b91eddd17b682e2c478943e7ac4c5517c62521faafc871f04b9883fa41f28f8763fcd6cdb494b92e8575b1ec8b17466d97631a118c778a42b357b2fbd802204265d23590be69a71469210ae8f26fec373125c8c7406eaa43a18d6d1caefe20be6e63d66478dcb214fa43211243f6900e8c112d4c31489a2b3d04d520285062c8fa81c6768f4dbb7c59698de7f4afeb7c794ca092a49b152704219dadf10feb43448de8f94398ee5590d69d5c6bcf91b979ec935349c1671a68818f64075a4540a8d71a575b04697cf59fdbf6e72398d88536b1e55dbb6b1d36575d171068b5f15947b96f83721245e53fc0b8c3e18b06a2a259b41956b19b77c803104ed6c07ffd6603370a8b113aa8b8de6fd5095f9469eb091d29aee5a122370770a746444dab73a427bd35b5310d103b8b6cececbd9791860121910d87a6ae5c8c653451aa44228d5a06f458b64c19a914163038a9769f1ab017be7c83be1fe2d584e0677e274935b10201deab0fce8080e09e7a1841e0ba4ce2b879ec3ff02296288152b6e597575678b932fde7b299f683d5b18b3ad7e69e0f93c41d3370c52417f63e8087a26283dfec0e9082831d765443e56b77aa5ca8be68e3db97c1ccada59f44475ec69e7e6d8a3d9933077168168ea5c98b5019b99decf7ff2bc8533d8be0721c3d33f01da7fdc2c8a8eefea19d46e44ad670d8223ab6fa0764aecaf92447b14e49d6e1ca6a846707ece0e2186879fdd067c2a685663aefb96a48dc2805908e7e8fa59a10d5875d7f88dc9ed30adb1dd2608691b63dc0f20f5541db10482d78f7011d62f4b59c41e215469d40fe583b5108e4896ced3f63f178318692a0e1fdec5e299532be1f23dbc75e5e3f4d515810085e8e414b776132ccc920d0266bbb909121c795f4224f0bf27e4a55399f70b04ce8fe400b3d3015b07fb4422a1b2a0371ccac9f01ad5737c03;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'he99bb1ebc099e6a68c06335989e7b7240549b6bd235b110edf2ae0ddd3d6ab120e086d2047f4e3738088d5eb15426c239c252f01b2d205724b5ec8d799c8adee11fa2a9664902a2159610eee9069d39667830d470d3c0a9b24e4011aee90f4758cc6041ed660664a8428f3480adf0c78e9ed5171e8a5857ea9c62b0f5a6e60b1d1fabf1d21a22582c3b5821b64a6ba400d1061ece1cb8b7526b17a98fc597592e58daadd3477f8e21c3c9726e9e3e28c2f9984ce321a9e7d4dd78fd35df7bfb900e1c16b513c19c3d235dfdfcfdee74351c0182c08b1351a5df5c45fa957f362f0ea54128c981f4ad35b352714ece0f736b4c5758bd4c9ae78dd8b222fbc3e386b4e97c113a31edd7ba6fc69a15fccd0c30e78d966330f939263e74c10aa2689fc8c8e2d0a7e0c4caa60f2f9cbe508a98d30918b0b3f0f124f4a90ff0792aa406a716788e3201009f5068d674de0f5591ddcee0e220d94c5ff5bf7d98e4b871b38b7f0bc2f0aa9e4ac346fa0ac023e17603016a9e52a8db851d68e64757349efc9930475fad03891a536bdb273c7ee7e0ed4c1aacc25b2a05f2e240e59d7eab4fffe0ff94e88f74f98ca39540f61db8bb28b6c62c2131ebc41c90c4b68e881aa768ec12b12e2ef379d7dd83e8ed31ac0ad3c877752c231f429b6fc2673986c3a696d36ff5a9d4d184ed6b4f4789f0829084998e20c53bf3e10d3ed284b7aad65b15a84c9b48110c00fa7d94aee95c3ee311e1ceda011aae8567d630fa1ed2ec0c8bcddf06855d501167fe87fe4912664f74253ae05563c7b7716bdcf8d763fc1f81dc5f56215da2894dcf69c7c554bfc65563f1b0e2d08c10a380e41a4d5dbe073eb4b6b32e6784c8ec951b5ffb86581c42f8e6cc32ee1dde992d8ee8b828c2ee5ab08eb5c1b518c201485b60415dfd66a1c9f313781099178325b3a92239b99daacf13fa45fafa12e5a653fe5e88f3d17dd4f64f1cecb1929460328c061b42186000cbf809543149b09762cc01f8cf42509f9f8d0f271854e507cff41e8ebefb1baab83f273b797543ec870b25cff4ee8dd3a52eb9701128e676c0cd5505fc145f8db3eb94dc007bc4330ca4e984e54afa0160cd1611a885fee57cea208775ba7fc5095eddc9252885ae62403ea793bdffd871d73503e78ce14593d5aef9b3c2a4e200a14c9d4be00d92cd66f2a717c681787cd1f2962d508c38a7af8ea1ff3acd5c74cd3ac6494dc8770280f895516a33c361f4b1751176c7058f05e76db5e7badb06914b09c145ca60e7474f8b278bfeb760a916a463df97c726ddff7c6a0b1ecd67db262f2f58a3723586be9de05525ce70c895eac487d659945857a0d838b8f81f8532047715e8b4e41a7a2507f4586269a82beef40d752b885246aa89d90e727963b369d25ea5cece46535c17350bbf121d602c4c4f88fc8a25df4f64e017722adb9e98c9c18e0cbed0dec71ce17a7193b0d91ee4c896321a4b72b62d4c4ab1f788eb3812f60105cf2a25ed16ebefca43f22b242c0f01a62679e215495cef212a228ec8384d3e36393c3b8e865f82b85d0194e90f13fc192a32c9f7fd65510009fdedfc1edb5ef04ce2335be6c1f2910fe56daf625b0d27ca81ee5d5daedbfcdcc6ee380da5c2e6132928519ff77d8b6433b944d62ae15ea54df2b6b16b041fa8d67068395072e77e1fc75c0362a1387002349f232d2d6414172345749b139dc7a323b46794af2fb96a6e2253e7e4bffb0efb7bf80cd7772b3b1583bd210f7e5816a900affe2245ddcb9cad780d2b8b38af935b207c25ea67041cc4c59b118e0fdcf3cd90cf028638fe678e8c210c838387f13e70b1ed1f913b4c90b48963b56c1b5863ffbddb35561acc50465d7a95dafbc155eade0be23f5fd06ba673e8703f40c150bc627971ea418d3711fc0c8651f735f36b01478aa943fccfa8e88b15cf7cff2f6a0228c2d8469157114cdc85bf4705817d3b03d195994e2a201402ff07812aa48699d28c7332fcd2e92567bc9c9a71ea18254679caeadfb036bf6d6936b9f33b67ef5b04775a7c55a013b06872122a37634d17071c7025251dd2bf616033ce2037f1aef6bb3f712f1707313d3df8997bc8537f579655a26c1845f75bf7cee6f388286ec78800eb6a3e83dfa14102c8e359cff63b4875ef3b754549581ef68568a8f4ca3f6377cc79a17e483da36a6df99c1c2879f230176f590e703d866b327f49defa00565b7f478d97a7741ffd893baa059d8826d8b9aaaa4e7f1b5fa40df9b2686ac839c1c0e5dac23a54a2c15fbdd821e6f357716f5aa171f9218be05c55b8e9a16f5407082a31fe4ea2e5c81ff636ce264b16becdbad67f49d523c17a243662e32af8fe44208b67852f4c8d9e36f6824f6f5ae8d7c5f392b645d9a28c409d6b85f83066a7f7d06b535d4a1d822a0ac0b0ceb5c0057c7b9527dae4f94d2212724c4e9d46c2330061decf949738cb734c3af755c61de7bacaa39fb4304e85a4857942165b414bb712b55050f5074f65ee8b88377aab3a990ad352040b30978741e7b576aa6e4c0f8689f5a71f18835e41998a894787f4f8ba18a2183213c6226c544ad934fa5fd7fc6284c9bee201cce79a17e3040e773603a8ad7f65279ef4aac9a32b64e04180d8747fefc6c072d0f96fe3d40452aa180861c741bb9c34dd9d58afbb810303bfe2ef0708887d29788fba75965b2dedaaba89e7335fef2e88d978035bb6ee3d93746810d7457487264d18e38b8388bf9db004cc8897dbf57c481710bd28a343bb1298acbf43109a10e140db5c365024b35fdd9f6b9ec9141fdba81eb5f6d3820de3e0e45909908427b72865ec928e7b08ab9e6e7e1c72672c98741a77173e5eb621970423e51bdfe0c0a90d3d66863839246234fb2a82cb35aa3d55704b658363c17d4b2e093ab152ecdba881c6c12a24945d86f881cd87d92fcd0b4f3097ce14b88dbfb0c78367f1d1347c8ba5477773a5047d58e26bbe0bfe31fc09092fd898d08cc8b4fd1e293216e02b1976d3435c6499f64da20b5a5622fe0df81bdf51a7265130988ee15e85e60d82374abe0a821d4bf715c70eab611599e283e83131fec1da274408da45503d17d29638af37e4dbd65e8457c1bda130f31c36d7d9c9b271a3ab649acc98e15f6d7a012c3abf1360a655065cf3b6c1408f4a7cb83f81d0252650502bd9a3ada7c69db6e26b981b4dbafc7dbfb7a9d30f2a547b2c2375872094fd56d1676fe99449bf2fbcb67cbc216558c7ff4cc4fdcc00971bf02a9dc7d5967ea9e6cce68a4f57111e8204728f9330e74ef5dcdb423b985e24ed45578d001dd6a9d572fca49315c7aab692be6f2446ed0eaef7bfe5766d94dface3130c1e3e3c56f8b1caa9e8537b1db21e901c906eb73b2419b7b2cf587ab3e9d21e92ab50439d7d75855ce64d7dd3990775f4219a47552d3d40b5e5365f8a0348e7ad23eac085fd5ed964bbfca51980f5aa61b595ac953c9198bcb1ac3599ec79b5feb74eaff7462cae3705a5cb72c186c040cfa063372efc1079d1f0e3d8f58cd4a44c3b64e42fd3934280d626e2f042f8c3061908b4e4ade371b30f539623f1a17edd127787210d64d547e1940f91dcd319e85c1b11e42d00415912deb631ee74df97f9f93020a9c1da3f08aade706e40d8896e87213af810c7e5b8fac7f0748cfb34e730b53cdd48fd79e1448e9ebe878455bd12f1645f51753fc3b6f249840cffd3c05e42a6330eb30162308fe49e366e5cb5b563b8f6a354398773a37376227a1c9d6572d1309d4e30534b681d119bce54e192dab6992118460ece874eb52e28e18be2af5aecb7ad060137b811680d2200a0e0c332361ae9df6090722c47c3fe8bbceed03470d9dbf0e2a6ed7600c53093b87ede16187d96f1d057c7f4e1cf88acfa7306c193d56dd9937e5cd6cd1456dacfe9d829ba2626b5dc54b2a0fbb72e84ef581eebebd661bfb6952d569a3085f1c45f5d7e77ff95a076266556956fd3d18796478b460ae2217343d66e62cd4ccfae515aeae76bac19a5eb2e55ed1da38dc3f6d8e4ef6209886a405c53cd86b3e0969be179d7ecfbed834065db9386416e3f85c2116ae9c94f066aa92382062acfdaced2801c417ed72c4f1b073ba16b01d33c985cc458377979c0e567c096b4459c4aaa7c7e4fa67cffa8711fb604dd32adfc51b998db0dfb5559e312234f6e6f346e3a33569d452319f71c42c691a1a4870732fae593ba9d1052a577575fc20eea0a8d583706791873f592429d323198fe8491f9dfbcb3ada7b0e488a9ed2eacd152d3f57b54b94d5bbb84abdd6e21b9d70b4fc554184ca54026628009f4f3941edda0456eb273f5d57c5a405e4436dab1f0690020fae3c08badc60ad9f144e9792e1538521632bb2a7be4824855e2cecc90b18150f92f1abd2ec56afc802af3b19dd7f90321e075fc42453ad3a30b88a04d93cac9a1070924bbfaaa2b1bd4d62417bb90e6f6e40d8bb4985bf5ffbf435029319f898316429172f4ac8cf2e8106e7d1423ab70c08f18cd84e7fecb15aa9e59fac42e98881976b46e8df429474fafbefe51e6c3050d75949939efe58454cfb31f5d1f3de591174686234f07b62e536b8dc0a4a458710cac4e300ba012ae4a8d98dafe11dcee924744baf3706b98ab9a9aedba201458c93599824d9ceb9d3a01f033636fb5a7a20a6cd221818297020f974087dbf7192599887edc237c41317bf6109ecff99aac3aa314cc90dba6e668552b17a4f586b3c8f86ca47e1c86b3db3e326e87d8f72cd97ddb204e0074ab6a9e3cf352a6898809548a7cf3a28aeb27e21517a83691b2ba5e70dd6ba55620e45e9e46f04af8dd02aa8d765d65d10d502b004f751be0178a3c4ad020a7de1cbb1db47e0a7a34c33dacf4f6acf2af6c7fa57984b03e2057806657046bd2ae106526bb445059de8f4944a92aff29e74fc7c806b3d8abc8a32cbce10973f5a694037275ae3a17e25fe9fa39fe75aafdfdcce9380dd068a04773baf0144048d873515754e4d7a6629cd42938f7de13596b26278f22ecd7a9a80caf6b06df0144f7e5f9425535e6271ff4a386fb3932dd40ab1762b19656061ddac56c8cbb6b212d43bd621e75dd5d51bca72838f871e36bc3c6f1131de579747ec74f6800d203288a7cd1a6593f1998061aa672fa7288c60a06b1e7b80f53d2d3afce52538c9db03b90f673a0dba6c543d145fd8882297a2a816f9b805b7ba023934fcce873f71c6f3f559111a3019655a7bad379f1f346138395fd68ca4150a982aeb74c3a81f9415cb68be9e2070252969d07846e495c90c813f40be487b562933fc02a8b41ea35fff70b624726f1fe3073c2fd66f3dbd40da9ab6e34874ece89e0ba5677619859b5a6308df85afc73d17844e08b3c4674423fa4eb6932363fa6b65425302a8ac409b9396589e1a3cd8a3b8d244490cd40509fa1046cd9e223a5703ef6f2193cf01a59e7338da31e6f672ba7477b4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h18bfe3a0cafe032c518ffbe34c5fc079a1993cf08636ffcd2939e8362eef3ead421ded3eec7f3249d0a7cca94fa6fdc6f691051b3c7548fabd2339d252f480bb6121346aeadbaf9ee023153611b78c023b07c251d8d78b7af5d5c6239728e1c8829d96c5aa65b0a53e1ddb403e1cd747c74c511b8367780a6148234ee3e7a479975311de2fd1a16a16991cc815dd526248ed21acf23c336adfacc244d7250a258b0b89838404ba138f9ddafc9cdcb846d26f8512658ddd1d7196fd56a103cb5d09067670572f1c739307def263cc8063e8c793f79e339cd3b43812ffbc3ed457098bb946eade9b6cd41df62b7f45c21521c06ef8da7f8ec76a3df69bdd56d2bebf304269c7c8bc81c4ba765b09c0c26d4b4fa2fbdf8894bd0cab3db900e51692b8cd06af2287587400be7f959f0ff0007a564bf6633b7f6b96f4115fcc345cb40da97ca243a568adef3942cc96f04247ce0de024d7a312745da9b97b555aeded2e6469faaa822724dbacbd69c619694cd9c524581e911c057b3cb4caf476fe9515933922b45e115b43bd95aa9abeac590c29b8b5747a25e7fa08c95e4d90e469985e2a7e1192e20f58eabf4bbd259a32b13fb91916fc1f6d14f8db637c8d07b7cccf75deace2ac7a0079341ae39417e4c96330aa44d687265f48197e89bdb01b5f1b466893dfed8f7c0ea526c10acbb1013cdb906e50a1298f7702d6527504cf06ac757d39516af8f4343dde4e527a160d6665add7866b251cc83a8e2af629f461b8eb90c60c825f3f85436bd8b8cc8f47ba9682d8dc4f91882b431f0b18dbe32af88033f1a1e69fb8918e02b363d9bdec2c316e8c9536f39d824dae0ca2be63064cf2d8dadee83f810befb77fdc17df739e7ea11deb416c2f1e4afc94161f0cca872701ce86b387e8e2a02eee72cf7a06d0f0b042c99db83920a5c687ec11d5c4d4b5ef97895fbfd9e56d69a23bf84b6b9117babb03206bafafbdf5ea1b88742466ab297d5d00fe54ee9f0247de1baa03be9125b8a6a8708c29258d498acedcd90c8be16b17f5078ff07f58c1474062b32e866889ba8174866f73f43cae87cba377feba2ebadf62dfa71bbe3608728ef457b6cc9b6b1310a2c59ff00122721bdd105dd2c7345ae847a888fbe647cafdb32468e695c5c4601463370cc169770739fd839678bbfd85c1b6e360aa93e42bcb76a26737f0ac5593b1be1ef2bb965a937622ef16011723935897f6675da8281834c068fd283dd0c2181c9048902450a1cb9b891fa635101fb2f3de0b86cf06482d89d775d4d8ba9e192d7ba484b6b44795aea0f99b1a32616473ba1243cdaae3ff375bfb405a74ac766b8aa31cf1672b8da8bca5f8882c87c7d81f9e536890fcde98df0d0fb85f2087183e0b787ce58898eaac2438f5304e8388fd5cbf6eb4e97e005dce251b469f059d651ec19f1b5f87c514a6d7f66c8b7433c8914acc189c097eaaa57e9ae89eb61d9262eae5c23677ee676e03d83cc63392226d9533587194cc6f61c77d7e568e605dc43ce646c13d3a6edd26ce2867aea81877686e942f9b74db802bab06cf2464b0f5502a7c547fd543e1b7b62b783eb0fe6e3949794af28fc57d8b38cbe29bf8204a199e2d966e72bb9240f8e2c19c39ea01c8bb02e3d74d8b1ada1e8de6e269863efae547e520b596903454b2a9d30243941d725cdd55d71405a08c0613f436c04915e8b497237192e29c329121f4c52e6d1c9d9542aee8515e65f21c48e3fbcd4b870aa3158ea7f0ad879259d849dfa1676a2606dbf4e65cb48b08c7cd3d67aa2525ddc4abfb7033d110ddd7f36a0132e09b518cdb22196bc2b8c3d75c9801dab429d69acbee6d44045568881542b62ac37df39de2248c05b516a73f2468b13b154aa8c89b4a8bdf35a20c7067ebb589cbecd51c09325513af50b923a4db183f182b266c41a5181d3f6ce9fdf3b4f55f4e5f6d37cac95e6cd3e2dc7df90703a5d96905e4a3b77d1388ee51633a96ea88d32882f07bb6910a7f6c84544e3a600533fe9d1715f03ca70567c492040df87c973ab385cbaad8e71af04617de99a807b4d6407f11cfb3df09445e36cc02a419d25090fd373d1d6493702e72bd2bd6625ed241b5860e25b9c083c619db6afe2d435e8683c8d4174bd0dc1d3c6d46917364dd7f0041b2d122a3e8e5972168481e7ce931fd31d0cf7caf8ae4915802ee7cb0de9d740d8f2839f2a2d227eec0e410729f4c551fa10da23751c172ca14397240bad74fc9e5b08d7a7b795cdfe2808e2a20736ae8e047f4d6d59e43da3412d1f7ee6966b2d41fe8595905521c2c93651145e3249a7a0e0b75d9f75ca4a14676f280bf88762ab4c6ea7cd5cc6c0c8896279f175ee7c628fa3af46dd1c891b8202224dc7a8bc3d31c61d8c48034fdae05d4fb5a6189949120c0c1d80f9ab3b28766913899ebaf9d2780fd3851c4007001fad14e5b2ae8644db7f1c7926c1c7efc0a278404b1166941c807ac2f5b71ccb14bdaee9a9d3b0da29506ba1aa3241bb65a28ca0a89a481987c8f47eb1aa212096a3d73db92e1ecbcc1b0669a4370141cac585b360a1040e24112bb956d053f368fb3d77503ffe8d21a81e0a97ba8c7213a82daf2465ec49f83b5dc4675b645f203d4103592ba068ca7eb0074184759a2c36b34f13e32e14805a7f4820101895826d313e651342e656f22b3a9ebba32fd55f08683b0f489bda41607ed44db00eb30e40b9759236aec7cc33dbdaf9800dc07871035d44820f0ad55cbe54ed34fb50d65c88ea18c582dfe12ee4e07c53762cc04e982b57ff2dc408bfbd37b6d57a486e95ab9bd6dd8626da987d401379408682ecbdfde0c754a41e753a276c5c4c91bfe42290140afdb0ad83ef9f8d0d8520af46021b26b26638455b3a971b3bd6aa9a457c70bc95ae6594b27c513ebb1abed88a905f2dc3261151b1130a2c79d8d435296c41ab7c6419892b6fdcbea279cd132e25d1763b7dfc75873996aa2185366e72400d0b237697227c6a1aa2a89ff908dfdbd5253f1a7273f14ac55cfa4e5d930e4d4cc1f0fd7b405b2a0dd8efcc1006e5039d74fa0ad80afda99a8d164ba860e67c945432e27b665e5839dde17ad5e21f1869bfb07df65bc237f3aaac7e42a3e6c505352984612e94cf6409d4ae19c604ef9bca0748ca2644f70dcf6e1491fd2337c81bb1709a2f8cefc6103f98b0fa62428983a7ceef529bdc770827f6212b9ec14a2de15e539843e98c71cce980f990bb004e321f905d66d5ec3ba1d596938539c70a0d09ee5e48a2a16a49e36d85162f13a44832d04546d4f4a4ddbbcb0a43f56549f4ddcf1829452913f022eeabfbda20c9cb60b28416f8c9618e5470097c31b7879d8bfab223e426cf9cebdcd8ada5171b9f0210591821bcd8638099c6a5a818e0f431d84c61cc3177339e31e65aa918da4ecbe06de63ad06fe09fdcdaac396c99403b5d65fb9ce70fd8abb589d21b5f81aa07e2006816ba6a7ea9cbf3eb1882743e36c67b19c91765618da030e3813e3aec466a408b69c1f1fa760e81ecc934811329ca90d8e1b0035aff41dfd0eeb5e06e8656edb03fe093e84ad4f42297c652e09a9c878f61c4d5e2006d521b217d16a915b65e8742d7cc63c43fce6127c9f9dee7ea6c24fe1efcc5ecc107a81ffae49516f5ebe84acebf5fda7e94e4a86942470d7a02cc39256547c2d1b809d737c93cbc946947e0438bcfe7bdcc5c16e6c2d5835175f9963992b5c4f69316435c5cbdc51c2467b2b914bfa4ce535575f844c053fc6d53083d3047b1d9bf1b01147dcfd7c71e64507f559cb8441f2e432652a6c4c1fad57853a2fef4b48d79293bbc996245fd9dffc0a0d1995b9b63a38355bab27c47f50419ca39de44d928c5cb3743655816db7d48f20c39d505d93a6735321c51291d36ea0a3ae036e16a70b2795f84cde5d023f71cd2d0ea8e1e71cf9294126b6a480803818c2c173e2975ee25983eafbd8676aba8a5bad0d6296004036f2003433e94d016a2acb2931e9a010ce7c6a140ed95f5592a63a91626a03ca88d8fb31ad7ad5b60db14392ef0470c3811f2d1f85b00bbf171d5033de2728580e9a8f27989777d0224f67d88d03f45049b1cf34e1a3bc987705ba9121fe4224705e30b6215283899c4bba06de2ab01bca5c5a76a5234f9d861371e8b0ef85f49681790977594900e716a6830517cefdecb524212f6e993c7a73a2794b2f90739e62727d570be0a3da589a4d157e1c6d9665e020bd661656ebcb3aef19cd7f490647fecbfd3190c1b5b6016f4782a8a9ccc8d10b7ebb1c27d1a066c5abc7263e9afa20b8b826caa08befc8bd93f13e0592aecfb048929058ffa4375f0fac99ce8d9b680e322af0d71f05ace939086373c07a0f6d724fb32e6b050f67b5831c11fb52ce920c0d3c18a758a0bd7eba915955d91a5c145ccf230de8e4836900471a1e79b5d7675d491394326b5d38f48cc3b2434308d8fcc8c0aad75d386e42768457e2ab7f2247e2a241c00a6fcf7e57ce6d75c3a49821b8dd70eadf032759e60cc169381b762edb614c59728e40c5bf2eba35138629c6963354db0f80f2782a506252b467a83881df639321c69f7a1b3798a6fa069b47c3641bfb97b2bcb8fb28f0c3e2863fa67396840de112f925be2941da90bcfce7e2161e08090dfbb8c85eeba013a0a5654f01da544fbfd8b4688358017d967cb4d886c86449fac3c2cd23828ba9d1d386dfcbcfa9d2a090e50a438aabfdedf1fb184304f6d23ee85b7004b7a8fba1541be98e6354a004c4fcfdab33a63654759014f03f0dc02397271dfb11189695dc2cbde761ac9dd0107bbcbef62ddd97d1d4204af121cc6a5e3ce92641c2c8e2af78d3e66ce37768ea07964e62066b7459ddd69bba3480596e714f33727fed282531e1c4557c53278b74d3c7f8ccc1586e486311c10cf2730655a93379ddc1cf6f5343917744b18eea319eb115933e92f5b81f77f5eb9c3710e53cae89b689f1fee1f31b38deae307f96566bcaec84e9d5ddae2bba9d33fd4b40d2d5faabf45c36c381ea52576a103da7d965693ef9f741cdd880a2062da4647e59977894476577f10a063fcd2ff719be536c12119e3a64f2773c77773f320ef15a3bb4044d72d282c0710b0d8abafaf1a219156c0889772bfbe965e489f1b0084de4c47debcc4d909003befee429aad577ed52eb609e1adf49d8c56858251d56f4d8d9c27636ddfc407fe6867fc27a80d98d69a1af757cc8280bda6ab805762314dd2e842720cf739ed056d42f4ec278a681cea031c749ace5eae3a84436106c91f0c025947683920ec89ce632ebdb63eb5b04389b569e6fd1ebdaf897256cd012218bf4d23070bdc46f8fc74c5fd00534c2b571b33192ab1bdb26e6d20ce633f04c94098afc414880e01625d91fa135e29ac8b1cdc71177b5f2217b4278e1069601b060d0d132b457d0a5f1726907115c05c2a48b6338424bb8be3543ea887bb2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h720ffe123d50dca455d3d6d0e6d884838c8eaad6b626e5d65dccb116fd3b19bba3f56ff1c33c9d9c4799c5a55699bedc6e818556c53a07574dd3820f7bc0962a76e62bbd1be82ab1267ba0b14e71c960fe1764eaf3b1fab18b6e659c050c3169e0633e838571f5f1fd62ffd08f0a2248363a9487ba610be7146f044233a5637851ca23ef993228bee7bd23e9561bb83ce43ea158e6ce38273cb3c52ed876b76797ab4f22321eefd0c9f4d2e2f245f8754bfe433448f69ecb68f9b0e9883c76d9499752119d806b8e53b276a1a729780e0148002a6ff57f80409cc0fbd67a18b1b51489137ade98653e16631a3a324429a1d537697b03a5b3407cdeb18f9c9d6912c537ff4d0d4d9649932691bbff393cb2400b5880e48a223af1d50b4f8cdde9c77c3ecd048191ce90113c70436bddc9b1957a696b5136904dbb042ebbc7a498039e697883acad246bd31b958a7ec06a55a76ec026f9084740e84ed810db82cc697ce504232ce5bc6ee8348dd49cb58e043bb535a9aa49546f43214a21e9cf7939d6d8c53e3333b4492f61f8d047ff5fb92d4351fa938bfae8d43c84bacc1a75e47fc8f3bf4a67207f5e088c524e3589d1519c78b204d1df54b43d90780ab26e914612353722cba2520a291f7e823abc1cf9af299498436eed5376dd8cc20bd9e35ed236884e414c9778a8bf64264e0042386c794ea2b1c49ff46d2f68aab1f23a28227f3e8658087d46e76679595cc5fe361df2a08cb68361d4719e47578dee1277909cec0aea3d64b4c235d1500670dcda8f175a760a683da906ffc165665dce51b7183429b28c4b86a051b51adcab0012b8374627d865ce872d4eb7b172f40f5adf90a86d00e52c2dec19e70a6ca452e583cf474d1b5ece3dd5220d85f78f99b75fa8ddd4f1878f6a6d12c901084f374e79ba844f29fdc63387315639a4c1daff988543b537bef7ef97241e46a357a95cb4eeaa761f72016f5a3170595bbf335ff4fdc2e532fabb63cff40ddc5b7ac9d9369cab596bbcf39c098520671cf338ec0ff1bae76034ae6b846987ac40180d6bcd2374baac38b35c935a97c5d4fe0601c1db3a988c3369da4a54b739bc82cbf790999948e7d770b5a67a1def28ba27456fba125474b0f87f2b632e4e1c2d86386dec0766fe03971f3e91e6868577f25837cccaf3ca3f7a8aae7ec7703c2542047602f823bbca04bdea8312bbd3901ec59a1cc64788252504742c538823f591c97b137936c10ee62869c7d6ae6fbf796c42dac18668543cf6bb04a8dda30d5474876b47d59702e4829216c18f8e087a79ff49a52dab79156fa56be66c57164e105f105ec5ad10529e6d20581b3c5d89a1e39b7f64a51212211c66d88a60681eff8b0708b789b1c37671fed9d984e4692646fcb62502f7e506d9dc9ce08fd1bfb355c8d44cb29d00c095c236285bae3f202ac9e347faf96a080eaf59b1a5f25312b026e8753ade4f4816687d2f902a6c64b0fb59b6ae7d8adea1d9e3e6aca93661db1427df814977e3faeeed78e3057931912d6e4e49e7eb0e123879f122d418936016baf2a217fb631fee610415e8234a001fa4bab5b545b60f5e114ce0524f763ab50ae85a2b0b5c671eb0bfe722c1347bc9c2b780f6520a1277f1f92d86d870a5426c17c95efde0945a0662caf7cdc57a9eaf343b759f37baa07943e26357b0a8ad11651983544d2505acdc6dab01b254f37ae842761821535150992abe45e242a49f64a50e71a7dc855fc239c96822cb28ccaa71cab8f7c4fade773f79fb6cd2140857368a92bbce6c119046563278a28e4fc9fd83486d129c7a0d3e49935826f8cb11ae21c2aca635ab99ef573ce1e752df65f4b59b4a0ffbce74f94c8ca1b54a3616eceb0e692bb716bf73e95e7d51bfe1006df0918021b73ee31f0322217f54ce1be4f298142d493d6e72b8b01db1c77490d21650050e515a2b3a7a4e0e753ed9c81468ca9c9a96b6e3248bc0f01fa9aa126e34c3810307b1d43319761b122afddad37b34f36ced29565e51731f9430aefe0529e52cbb18becf1fa494a5bfc06d25a566159c349e4dc7124ed53265dca8116ae526ad6c50a192e09ffccf8e5ba59ce73ce22a8fb407b27afe21de425d1687a57bd4525713924afaedef082dd11e8c19ab381022bb09fe934443e4b18db85017f8c507ebb31cce721638907145e6f643352a4ed9a8b238aa7506c65e05f4cc0dbc8def5bf1150ea8a9cb4d6486a0b1682668bde30a6b435d0adf4513b5980a23005fb49ffb1f6480ae332fc838047a1e666a6f640576a7103747aaf926f6c411dd4969856d98ad9dfd0c08af5ca09e86aeb8b19182c884b12e8fd961ac25ee91e5965d2a2ac706311b5aa2151e25b00ba23484e5ab7b84902827b30ef80edbc2ea7c9d59267d42aaba587bbf68218ae2168509f93fda7e7de79e9a7110f0e4a0201cd83293e5e30e56fa51a8ec443f51a5497b097fa89cf8013491abc486c5ca694f6f60c958ce3422e7416cabe9b9b612e62a5c2d2af5756c586c3a9385ca30e947f16c376f67655c03ec88f2694530aadfb4be4d6352b031f50df9d02eb4ea7709ef72a9b1a3282ddfd64fbe88ff787062c57381c385eecaadfefce8a0b3688587afe29e0cd44aa0be9f937b67dcde01f1eeea2ade0f9726ff26fa3afcec617cf81bafeaecfee5c0c3048e189b05239511260894b5cf6b178a076e1be2774127d8c402ce7bc06169a6695bf2b38095673fc322048f838682a60fcad5cf6e235f5614ae77fb78d25ebfd2b902744f76ed567cddb4bb8260b2bee68c7ca74f43db345980cdb1c9359dc7d0fa6974781e5b099c35fa34495562e14a8175c87932f65d39276542e3689ee083d418bba4c240f94cd60b69153ce45fb5040f5b872a83a42898251564dfaffba4178c6409570b3a42be983c792213f466ff982ff9902e8b2539783982bc505cd1c49a55fc14c5ab95d3d36755b9571e8bcfd33b5f145e5febeebe3796fb914a3aca211d5601a7e9af16c634fab777f00186a691d4aaf4741d1424b5172437bee6d421f61bb62ab7846d4523e558f10695858d78697059b5ff12aa9b692d8172016901d5079ea9762d86e6d3a6a19abdaba1aa4da24865845b800ad0fae4ce8522f2593e82b968f05fe9b1dc8d0fcc7162b672f4e299d0aa21132271120392ec741d4440581860e4b567d6c8486bc47d49e95ef72326bba2767176086e56e17b0aff3b4f8c2838081e9dc858b74d37abd13e042812113246e791ca82bd98fa1c5b26d83ba7478c96ea90bf75bbfffe2ff7edb2827c269b23a68dc695ce71c4d2ce44f23e9cc922611307296557f9382da12b8d50d96e1775954b87f77b6318ab3197dafda098dbc49d83f2225211d7f87092c6a0045c8e45a7aa65f7818c69818bdcd865dc7b148f07451761ab56f7137a21df16e666caaade9e0ad87c971595b3d24ab48bfe922764f707f91f7231785f8269487964c52ac3500bfe6ef862fc0be93c72c729f67db54d38b0fdb37a350a0ccfc92d087f7762b2dec828c7b7d1658c5ab193d458f48a123a26825ba2174ce64efb9e01a29d93fb9edd9d773dc9fa54b984a9a559e2344b775bb69cf0067a506bf28d29d62a81669fed96f28ce623e45817cd0f137320ed34fd8672175b3d42dd5f4a9b5fa77a1a3d4e0a47cba88c505eac763f6d6066576152719f1b103140ad23f71f64172036dbaac3554e30772a705c8f82950f10176d19b3635cb6441da699013490cc6e86ffaf1da8666dab6c57379ddfa1183b34c690e40500670a947a95b71a20e15148a3681c5024524a7df2033d385291f45ac423725b728e3bc6fa74967fb8c2e406e0d0510d3668cd88ddba95c15cca34da68211aff2a2086fb2426840dee178b1da14f548a09f96309316be264747b43388cab9f6d24aa2f3947c715f38afc5e270ecb928345c3289afda94d56d9d5d9bb97f86f7087d5ec79cf2f8add9db64ef0a1eb7962ed062bf9380fd239711aa067537eadcb54d26becf914c5f9f3640745c4f8af5bb812bfb4725868b75e97ea49603ddd990246e07f94050b8d6ff29257042cc771679a57cf6fce5c823e70612fd589faed0410d32914ead2044c723bdef3b4c7fbe5669d155bb3273c41765c16737b576bf97a35cf609728fa0bcdbf5c5d3e2b54e33877718c33ee511f06625d6b1f6f1af9c721bb1fd27cf27a61babd0db8820529b27d4e6dea3d2758087eeaf309e31f59caba03a49e9556c2bad149a25ddd63137fb0e042dc7b2376dbee62aa5a474cbdb95c6b7a7b730420a5b3144498454eac7ebb05f68fd7a20e5c2e0b74331067ab70d6ebe9ebdea8a087a6ffce6f913c2725e1ccf46452b76d332cedf5505bca77bfc55cb9d3cabf548a3feb2e7d49b95a24af27d9b51f52c5b53c69776d018112733b7ce845ab5a784d0892b8dd8f40c61fef90ddc94e6f243f7dddd47ef2c81caa92caa8865da5bc5320cc8f745a2fc35a5f5d920bd2d424dd11933a2dde2c4c29c1379143a0df5345c04f567efc7dd6bd95de299dee1fe67e91419ff7ef5142e37dae7913131f238df346c6293f8131efab95f3cc758da9764752742d9f8be48910e011ca3f1c44fd580e5b651e699c7e63833b2f6276ce24c41a300138c5de4ecd72948293d6b4d6ae8a3e378619d59b327f07adda8dfb3f6feebc92122c6ceefe9d496b59883acf5ec6e667d5513e98b121fa86f051d51d91673c513fd3b66140e95c4c9b6085910431a01a08f7e2f3acf36e0471332226441d2f0d364745166efe715d31e8492ecc9006771918726d579c0f5c206ad01409a1707664272f80ac4eca6c9f1458202d59e387425c3cc0f7bbc3fcc3047f9ef0bc7280e952774b708d73f004f9221de0ffdc6f08daf8834f341ec3206e814aba2ed3a81807005a2675555fef95e83fe97713ac9c13a7119782ccccf0c0bfd826a83eff6b71f9347d2d1ef62bcc5fdbef60ae5032978d36b2b89537b17e02c67728a8219987b18d19ff18981367241e492777e53eb161769cb0d08a13223941f1586f400cd40c63162185d575bbb329adce1246922fa14d18f05e8dbdd9c002fb9a28dbacbcbc3227addc85fc3dd99e6f85bbc9e9077a40cf16c69778bd88b9ab9bbc9b5415226679116303bd0a85dc4784f13e12c33148bce91a54408675ec2623275296db08633eeff02901606fc3cfd8ea73bb077b8007a057f3ca724d3ff0cb5f4b105f01288482f4147089cba41bdf7f6c91d98f0f7a823c0fc915baf184685508ce83847cb5155c703635dbfe518c072502505c2c375963df713f5fd838ae41b06ece1f27d1ce95759cc32b8fa37727ffc2ab593f13e99d3f6ce4eedd9bb4ae84efa91c63b5a204f5a200380880cf4fa2b17c372e4fbe08d8836e2b1964718186dc60da8e04add22f74311e3c1fb0945a0f2305ee3f62ed0af0994396086592fc5ef4f19a79531b1ffc4f68d0728af03bd456bb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h34ff694ad23c86ccb4bf8647d8bdf32b55ad5775772fc679c483aa57e40c89ac92f250daf37bb1848a889209fc5ca6ba1fd07f1c24434736a45796b4a22db15135059599e097f0c9cac2ec21cb623d065447ef738bf2af085dd841759b72c72753c8408560f107be5ca37ae3255fd412663781716ac4b3664a1216e68c12d7e91aed6e7a9f72b65642863d431e3bc54bf79eb53f79b6ceabdb3d3516bc2db0403d8d079203312f75f9ecae9c0869deb49147ebfbf53813cff097103dd97580add4db584c9c90c04999418c81945d9e6f2c82ed40cc2641cdaa03e992af4dabe2081d3583b4e3a8138145d63b6cf12299ab792ad55d1149476f8e33f5821e2d1f08e38742f734650aa35713acbf7d8b10532a9f1ad4fd6df88cac83987f7574d74cd0c14e1d5f917350789a5baa21a684c320c623381ad0c60c5cf7c8529618b593f87de204f11e485cd8b4d2c5c200dab240ed902b92b99d0d13a8fcfa6245b667c78fd3a3b72b3e30e1138fd0ad84be68a2bf560d94a7732cf3a520b018b036079f42a7ce09c628fca1a5a472421340da8279e864cea21dd337145709d72384bf915c76541c4cd3c2c298070a6c8028f155a28c99c3a908ca5f04354edf47868aad913c94f5b652b572755a7d5df2f3cf0f1b19fdde348d33fe5f772db792973ff1e536dd65669e1cf7013d85feebd13d55d83202594c985eb0225fae029dcfc0d719b2fa57b646818848fc89592a216b17d80e6aca0022228277cb9322b95bf226e52b88406c24023bd719c1f03e36e48762533a71fdc562a78c111125d64475d0ec325b083e8120cc3e8acaeaf4c8f3871e2a1a80e6a1eb11f026939bc9253b5f28d286a71d96c8174d5d62b79d3b026cc28bd5acd5ac660bec7da7fad5ed99f2f1c56c3eb4e11e6b3dc5f16f3426e47a4071fa13a6ef4552c6c5c09d4f0a30be24757ed92b87167fff962fbb77589313e5cda400a3a313d481107f2f8cb8345dc9252a4cd2349a01e2a6c58487565af4ed9bf1c76f777e5f229a9bbfadf317ec4df04e3fa645e2435964927ed599682e6bbcec53368b7d04fa3786a9ceff5581c79d4b38a760746e415c85ab96a8c5c61e3e44bd33b86257beb3a5f38d6e489acafdc596600adc7be6e2e997e61cf34cbc28d14af6f8747654e39bf928405921ff6f1ecf023152c06acc28aa5e8db96564b2bc2b84725affa142c2c2b3b95584ac3df88d6a28ff07988ce50738b410a8acb9a5db379c5a5475617c0f708dc441e6b184818dcdd60bb6d2bfae229fd96edaa3abea71bf7c274190fed8f63949c8337c46e2dcb1e2e24f7214ee2f678c3765e9dc3709572b479369f9f1e80e516e7b5aea74b29dc7accdf48282bfaafad276418e826610fd4d83b42f16406331591d4c003ba59af9ab56e30730e3e9521a98cc4cedbb03db3edc1af58372845d2d4aaffe9bfb0793ca8e11f887c8d1aaf5b1464d468b7622d76d8ad55c1f07a97721feea863d99fa05e538f4122ea49f62af58c3ae0744aecfe35e836ebe08e0afb0b889ae52d4df9d980dbbb017643f592412a622d5344c0028f5aa4b11cd3d6f0770a51b07e407a35a41e7dc31a73a06b38bdc4846a8518d742fc771743bff2ab082281c33bdd75c1fb1ca75ab4487ff9d1985bb0928792e06acaacf268c463942fce28e25a7f7b14c3c98c785e194919eea50d956ee594757fffd60e518ed84ab914f1d1d9dfad8a5a350463dd31e67604be9b52c43b18f135bf18d6b229b93d343db3863d3a87ebf664a195f38dc34ec4ca0148ab4370f75fc02430b6e289ed1e8d20f2b0ec3277f8540ba6a6b2c4cde797a8043b40a0ad56e18d760e1d5d3a2b2351146f2b98ddab1c0414a1a92d2c1f8a16e57c1407b0a7b515fec09b1e499774aca3e0a7dcffb0b703cd5111e7768d55a95a726ca40757efd47746b960097ce8b254a7eb40cae898b40123bcdfc2b55986bb06df44d0049e37cab4216577f20e57778cb320565c09249ddbaae5e669e3d9a9f767796d1412a90fb91cfae35d91f93f1d53cd0ce2600cbf98eea4127349468bbdc0cb2b0de62aac0120147a0b46220b20050c04e7140b61d8fa731932355f32a828348f924727cc615300c9764b665aa0126d28b763477b89d7ce85cad3ac1fb53bcecdc7e651c979eac0e2731dea7a9d598dafbce85e5f88143340d0fa43d0c0b065be5bc728b2a68d3df1056ab1692af7b6baa8ecdd2c3c7009ef09d52753bdb76b68a5f5142251cb9ecfdf765c958a117ef1a72f859bdb1a9fe24ad1601e170b1f3642671aa993b0ce541d82a32718ae0b0dff3386e46fbe8451f38817da4b9ff12d67a0372d35fb1186b6607cddc47b98adabbc2c597c2f417c0a99a07184f324cd46feacf82bfc81ea357c9b13e0ae30a50c36aa648051ab333fc5c18da589382aaadba563a1cc89807c63266e22017e32ef40fd971e743d8567eb0ae24259faaff5e9573c520459d8694371f1b769b3dfc8797de71dc43f7448eda28660b228e69b312c0286ddcdda0435f5b5e3c67a5365ffdd2fc7865d80f9cf825c4a8fd160200fe574b65fd9440c3f76ab61b835c158a511c5f5c5b00c0508842d1ac31eb46feb15164a292dbad3db1633eaf687776f151c2d8e01afccafdf28ae2d023aee5e1239616dd9123bda733743e3003d7028ccca1d4141501fa5c8cdd5197cce22fcc7f27f379de733d9f9c0f007f561553eb2dc3630fcc6170942d707cffaff9daa1978badb3c9141301346d0d6024feb996b61083d42e798f447cdee17dc985a585ef356ee58da12b5278f9edca2b9784e53fe39bc999648d840ee4dccd317017376b14e74dae9852a121307d123f4b010674bf53a84566744e96480bf02c7f82ed51a3558481cfa68deff927c33ac0a2a9d38a7b2ee69899681a4c8067e87232ee20bd46f486609242d55400c0f935170941ff518f57862a0abd6d232119a9ea71c99c3a33f510af74aeac6861f7a1cf28c9b4c48177d566eb41d195a1b3cf7c2786d227501a4923ada6da5af7865900519a800020a8ab4e7706ec1525a017f82fca19c905b8edeae09cd72ade599888fa0744aa99520bb9f12fe39b08793ed85e0e3bac7a1afab7c80ec4ae96f06303e61deb929baaca9941c1fd174d68b3cd25759389587a391862ebd2b04e1d0890b4c7673903a9586ed3a6ad0d2393aec2e32250fa0e3e650af63150be089f149f101eaafbbee0e9092c5649d62853fea9d2eb0b2ec30bd57bc680dee86587d8a7934e37e1ead1bb936bb45288a652bdbc689189031991a23a427ce2e4532b70d9804a951b3f682eb04ed0cf07da9355376c735cb50e9d491c3092df580ec3931bf05016dcfea58886ddd208bab41cdc09b2c947dadd5d3538260e0a88b09f4acb07df3decec3c873db55d7db959d8126cfbca4385ebb3b2ffcec13348ce307bb93e250c5cbb4f7c37fee0329c1f5737a9ff7600308a8e7dcfef0f24628764fefed7d3efb09c493d715798f33f04dfe169f9f1a50c78a399cd024be0383055e93bc1ff2b3969a4e36440b6d8fb4a4bae1e32bd22a9bdbf706132ac1c24f6c511c3fca28e8c840e0f81de85550c046211f11d23afb65c5be0ecd97ea6eb79915498b50774c1c7094dd18f8192b75963561b229a307b3b142c890925bc929a8f41bf62b186f942b77576bbe9d1f8738a0df70d10e6eac9a0decd5485250b42be54f97287e9ecea5e53405e6a1511544d1668a1425994a6f31fcb34f6ed3b2b328ae7a57729252b0d595df36e43e24cb8de06038637197a68bcc9ef2de92d323dc064f851be76025e8bea6f78f216cea176647e2a01c63b643ac84cfda883d94083a96038ef0ef01c1e0d8275dff53c43fea58216ea1f7d8a734b5f1256996a31383f0d7fe618b5a5af6c1241e35816c896dd915ce73dff7241ced6069b819c077c5b88593a641889788e3e1923f2c32c59a41c7a02253c4c1e404bbc46ed9680dcaf1350a89abb0a48552e1344bb09ef9f34c88bf10d4523b248db317a17412afc52f830e7d1b87e5bdab66bbe0b5fd184890b7f1d8fdea1eaa97b6fbc6f4dcc7ad8754d61bb7301e5d23be460c7c1b373251b195bee75dfb5d65c3b266a0146ca918c41f2de72686c1c7613c34956143acf8fea69a59b6a542249fc888e3be6052794a6476d42052aa1b0a7ef879626c12ec29e045151aebed1755eebc4d598a45ad27c586c639fa6719f289d607f8ab2f52298e3ac66caee001c0ffc1b7171bea5dafd87c18e93debf325e3d5fbacbd7e9656953237b1d123064c1c110c1ce1a9364eab294aa02701fe430dd23c58a301907180e7cd8236f850282ecf135c7508e5df4470c12ee6aafd7115587b207665e5aae266e1107b656bd6cd456d10e10bd2260dfabb67d16d43d50bac02855095e87f11d82d6e6697543add1ad500f386b732a76b456a044f8177572b92b3d3160be4205c8d2da05b41679cf7fed117b92575de455e048560b4bc26d8af71cdbe443346bf02355162bbcfb72adf19947330a0f1a0ca9e3d678bacc1034935e0fee16748a7775d767779ee14be0f78073cafefa2e29f094efe8568b57f2c3a9fdf6f5530516ce7c1c8d03ffd99076cfa4d7958c22ad9da3426fccf5ed297a63d270c1a7fbce10f0b04fd35467edcfc98dc5992123522d0278c798e797b46bd342cdb492b320419470a908510de93503c78bd7fb381bf3ea212b0c71bd16f7e2c928a24ba45895f61f2664bdc06b7a2ce2ab738d6c025519e4ec56a8c7079fbd4897a3e2ae38f11eb693314c4bf2e3f580ec027b6f26cb01bd49ba0174917f20984010db0873e88fef6edad4a02cd7072618f8db7d5be82b9a5757d5208b4470c4901e870e1473eaa1933fa6a084f3fc9fb8342c40ef0b6b6e1af7ba9e5b21570cdd7d48d7dcf8d6df6bb4bac7d071a10184e236043675e864a67c83ab92b8aed5d1b2fc812c84af9aefaf4b21e8c90b262616af55c51377578c92a500a3497d895390929e7f5267fdfc3b8db77819563b5d87bbb73dbdadfa45d5dc67bbb94170627b47ce8ab736d7d9f0f8cc450f1c6221de35748a5738085de6dfba81b813aa64fc531f528c4b2ab4a0b97c8ec9d5159401af9a5339048cccb88ebb495f951d0cbbb9a64cf32f59493ed747fef53ad187e2bcde11dff05cf03c7f923700645ea8e1fa39fa1869ae34346c824a742946dec7ecd2a513b838044c6ec67ff8d20586136208ccbac913fbdf2306f5415130f4e11dbf941099afb25acf62522a1a790a00581270597ee15e2bf6403e4d2eeec380e2cfd824b1c88aa6873379f60f06289744b190b07d80e38f81264422612d306294c04a0c4d34ca1bba22901ec2c1cb765915d21860f04aa522462cc3be53f613fd55ce27847bc260cd8d49ddf121280b9294ec1ea3c84109fe722deee8e515878219c9a3196ee4900f475a34740991dc34e9a89de5bfc8bfe99a8a87d29c8eb98f34909b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h7bb490b5d3187e5a7d6d04bf1003890167f663f291987d2421da5db015ce67e50bc468198d358d82e57763fcdaed0135b96361408ca0b6d11cbfe5f4f3215575a81dc4808f7a4886af62100a812730c1335245a376884864e1810e591921e049913ce9630db94fe81d0f531b6f810a50aaadd1f32097308734945d0708b331a70f5595f39284b54ff90814405003f8ea1dd7043749c949605352ca1caad0d92f3ac6d2be02dd9ae9590dc9882d720d949c0eab3b6979e8adf3471dd36ac2b346ea5da0f143cb2982eecc076548d82498b755a4744af6026da80d87bbb769f7954ef601e4964a12ed337cffd2fe84347958acd6bba2650e5cb560595f1f5e04fdbddc45998c75c51757d6d772d753a0ccb7074de79e7fb02d0356707b53618d8895ff24fa29dfd36dde33dd8aa2708c025204e86a07a8b12eec671e90a317b8018043b31a9078b607be717b7ad74116d2b3540c5cbfef0e2f8bcd676f28caa6326bdc850395eba86538be072281a9aa334a0d49f20b1e6600c072bc8c2713a8db536ff36fe0ea03705a7477e7fe46c316e55f7b3098c9eb56152d1aa87139127ed0af5cd44c3a1a4ae20608a85eb5eda26179a68ea52f449591d7f1209b43cdc052c0820966cd466f3b8a8cf36eddca6dd54f54cd47db617e384b2f4609bf6bc4fbc70828f94c95acf28ffdd80212e77cab04c1f8780dbce89b9311fc311d0e12476711f29902b93db3a251b96b32fe890a5f44095a5196b306e881c315c782387b67e47eb788a2a7b4614edffb6cc1f4f404ff5b7e789ebca4b68b05ba237ab0175c54ddba70c4d25cf2d3a9a5a90a84e1901ec98d59f050c292d703f84557b87782f477f78c1b3738146970fe53a560877a4fe41f1da47b5df9ce2c935d4c6b8722cb4f854490a34dc1e30e9337e88842a7404a89d3c39b195d654e075a9a395c2d42eeed8cd0b6d8ff660e30ceaf4016e3692dab0120409c434fea88b6e6faddf92087dc10a5e429cad81f93034564718c4711db13fbcd66961a5202e290efe24102f8b735cd83835e523fbda8b13644ca65641d1465e0f3fbe55948647f9c22984b51567ab4718a04028e96770936e589e3205b1b24dfe9e933fbc3e7466dab53437fefd4df029080faf20dcb4bcd7f6f256b21a1f10b9e61b791be3eb9b04958df9e5dfffe02e5b38bc7be0a365b6a03bb3fd407d64147538b42bc3dbf8d62ae5a9cd9969638d8aefbba6cd34d707b96fd2ec6e2374d31ee401a8abbbde71440fa64c040c6e67003907b344fa8da8492ad75828eb0a064fd62994f85108c6b79c5078c691c06b7825985da9d1089e0efb57c4ddbcb91944fe73ff6e27ad598c84d6ed15026343cbbbc2bc08265fbd6ea8ee5393ac9121cdfb18e321828819f1f899303aefa95fc7e7759982db7bf6fb0034d050b960731d8c476c4aa9ba41677ce0a2275cf0e60bc6e63f53fe88d2bd563f89c1f70e68ddc42752695b53a7a4b02b61b3ea3fab3c0f9203cfd3643fd91e182ac6a53e114347be18857adf6f59b40a040d4937a224114eb505a0969bef85e53119ea4ec04985780cf99b11ecc0748a903b787c4ded1ad7f59a1877897359d74a5bf96406202bbd77b1f5234ca1e92e907715a5dfa35134d95bac34bf2160ba231f855d5b5aa1b94f4cf31ea0f207c63be57a3b6d701539ba8f80623baf85adf97cf925ea7ec76397ebfa32bb779895bbbae683e57146a16453967e10fc41fd88cdef594e713bb59c94c48e27eeceb579ccd042ee52195488166446a6bde1b2188ac0e64c7ef2418f2c4322aa042a503d75bd19394b4cbbcc895f4b5c9877a2878633f3c5e6d3891807be225bc716a558bd6f03ab985cfd6f8a43d2218ec3346be4b5f9ee8e5457a79e5db21f0f6ba8e7ca2c11d6fb39303b31c44839041ee5396f59d38c7caaa44d933224f327a705e54a9436163ecd5c211d5bf04587fd7206ad7e7ca0b689adb53218888fe53b89ad773a3b82f89cd92a5bd60adaf0a574fa24e7e78be59b330765b28fd77c31c546db97258bced267ad3dde4e6946d5250518ac7141e6a48b31dedb96ea0606e14162a6ea00a9ae2e70e7546e4b363734193bd32f24d0ecc740232529aff50652c9414a70ac1a60eea0143f111a4ca8f77385f851b1a6c22520083f9a5b25716a2b5d41ae352624e9d6d7d50b51d8a28ff227b5921d1b430b2025d520f749dd9568aabf2d6b24e1ff5c1b5204d915c25b10863217bf7e6a38b15127727cd6262b4acb6df353f460846a233abc06f59e5d293fd64a49f4c2d46a54da9516838ae8a812e29122b8d70d1fcb3bd1c8d94c99ed00a75c010913c4cd68c43b9b81ab05344c201e9d49a5f4018142428162078218824dcc3694ea51c40856709ab6b9b4e5c855285348770f68fa8d7179e20fa27d9ac107e99d4b42e0980238bac10254c095bce6f85a35ada1330736e9486a51b236a4dbd3bc0055bc224567abf2bb1e60a12706517378768afbf7d6d9b49636f1ae87a4352320417a627a685dfe0771f2a31614ff2d0dafab0a439b720dba62073d6bb1ac44ce0445a6d76fdc7a8f0258867ff0d17e003d8fa0471fa33278e1ced07d55088fdc37ffb7d4877fd18b0baf1693f721bc25686f6bde40cdadedfd1cde822f13da8ec83d4eed4fa7a63401c5d9567797f651312c539b8753375a02f7fa5ef348c57339cfea6b7bfce68cd369473db5f53bf294878c2e2b0a954d9aebf2ba099badb22e272b8b3412618e65922cc7fad1157c39cfb10a6b52ed45a6928bb11b5e0997de33db2e6056ec8815f985c562f558c269edb870c7467ace3f2212bd9c2bd34bc458265d1deace9095d1016495ced7ffd5f81269e86e7991aa2900f9bbda27c3f62d4fee7904bc2fe7f3fed33dda0e8aea8272a261bda9f7fb7b4bc8deb21c2a51d259b5adfb74f51bed09deea4bfb4238b028fd2a39b5412fcc62a0549a13bfe6b7711ea9199915b9c8b8f817713ab4af51da02eb3883defeca1b5e424aa0cabecd66f28bb2cfcf5da47d53a715f7691506c1549f8c97bc602f0fa86fb2eb1b110a4120cbb766266576e878c75e43c8a6216a715762b95e612d2972747937ba8c853ad36bc6426fb1b2c9182dc725a88ea22107e30045026f81d5baf9fa236b7dda7dec0034d45ce18a512db6aba3a77e24ce9175cc87ec8718a7d072e6120708a6875be1294119dc6bab42d4eb09f11b163d6dfda7df1287eb042c31e222d0bac5f5d09d97dd52fafd29223df05d0219cbb39f13d8c1416e3d50a57bdbee4e722e6b4f55b4a0915fe49667805f3089b84e9c76b40b09c4087ddb0ef10062f7f09eaccda68bbca45e95dfea03a262d6ae854973821a7fbe5f2e04b3de2d88c9de959c742295147fb38e8aff2e72faf63f54f6c7a4fd487fd856d2ad4b7566ee5f14f03af34fbcfd6c98520a1a16ceacafa21e65c3f3450caa0303b2667a0f8ef7e8c38d93fd117da9f2bcb435cc17c6c123db54fe66243da7273b87594de94e5cc180640a2a7cdede8fb554a9ad6ec9867c6c4a175d7be404b3fbf6348791e40204ca44824136fa8d85cec3225ccc41966527596e51e75db56ad61f1af41791dafc8031c3960b33b22d39b47fa59f2888c24b0a3cc23aa0edd84997aa8aa19b5084f3a32fe1ec40c7efec5200a631478b622fb1a0137215a2314471b73de2f9c1634c46a78ccf6c269f23fc75a70f7ef6c626d3e21c6428dfc8224aef2dbdab1e16e912242b2801dd0675c04a4e81b89dc803c7c38fd4190bb868bac38a218298f139793567d5df4ff2a6deba010fccc2f33a3a0490239cdecd99472c6b9202fc1e923f5da680ea41d8977fb0a9a441f1d2b069295f08a79e6a244f59d8e4bf755d9f007780fec6bb2f6e640f20d76c582a07a8a6149535be76dbbebf5dd3b42d9b3818c4264e5b8cf0885f164bbb2e3479b0f2e0eb036c58f0cae9d9306462f2d2a41e05b95ca6a0180dfe5bdc94b6aed42cbffd1b11fbeb62ee4c7bbb0862ca048d7a6bbfde36f6be30230c57787981401d841a29e7e47242355eb6c0704145c37846f280c9f05b3c297890ad36cf9534c154bbd8d4af99a38afbc73b07893829d6600b171a3be88ff0a1e88cee9712243e30c7aec0f0458d3ea42bb68a9c546f141b82bf2830c9e238eedcb5332e8142cb79a04e65a69870a89140e16d1de90323dbf5eaff15dee06c4793806ebe45b0f4577b18aaf6bf3390a57a9f95a748ec328ca182ed65f46c2f6dd4834649fdf46e887d158a7162f12aa7ea6fc0d2b923416ea69f752a45ad82766eaff3f5dc3ad7818411d8cc0ad469ce231b8dbbfc4c284ebc60281388fcb647c5bc040f3b17e09aee7a21dc17bc9933227e99cbe33bbc0cddd201d1825c77f102db3308aa5379e7a0b47fc4a7b3b2f13439f7518bcb913859e6847cd4e75c51f724b491967e23ac7f937b6dc50f9fadaa74ac54a223b13a75d9ea423dc145ab1337ae4e53a71b4d300f19ae23f1b1abe90c55694c665f6628521a631204a8a675cf18938133e74aaef595d8fdf807e9fc2b9d8782e092e49e8d83571f59bd66a20dbf0298788906e3d129e6ed5c02dd8763c8d00f63836173895a3dfe4ba85d2aa0fd4a72e4373200840ca7d3b82fb7ae709e5b4ecdf163c7a51235deb09fbb0f05bd8202d1db789494b89573532d7e7477634ac0583185d01fc402e1f56db322eb0d67ad1f7e09873447083c4d6d67548ad21cf9409f61a964a9b39e712a10ef95dffa2d2b594b76a1be5fbce71c8f13626831b3ca8b715f9bcc11de3c49af68f102c7737fd5954385cb71fa610e4984edf52f44efc0edf5466d248350cec24c007dbe52a8a9bbe78b30c19f5c4bad035013dd66ae0a245c58e3fd7022ad9c5aae17366385f5638685baffd5ba24184dadb31ccc6fb41f81d38be2b37315966e1e06983e13faf1d85113abe1d9b07ead553b3933f296b94e625cd6a314d6619f5e49b188b7c3a13d9c4717be1cc28073252f6b0904994a8dcf97dbe8dfaca0ab60a97a1c49a0b210ea437ff21fc2391328d3a22613b0930f6d1c294dc2113e023b1aca0179fc2efb71fb3eab512352be10163123ad2223e550652c35d7918a5ac52c413780913a7faa30d4c11480bdd61fec829e271b338938d1c17e412471e18ccbced3ec9206174c118b94ba3d7098e367837e093123700f6ce2435d15a096604fbcd4eb224797376da3b0fce06fabf4fc7edc7795e3df8e1827f1f97dabb502b1f254778ca95a167c168ee8371ebee9aaa85c1cc57eeb6ff1e335610950b3d6725af567b60bf8b217f44cd1903b12ef820d4769464b592128ea746fab1374ade8e202e916aeae7943ef2f12a28d6fc3e84602f0f3e1d356a4c304742059b6ee048b8366a1ac9878ea9b820fa77cd47944c4ee95758226f86f5d199c2f730016b2a99c678f7e9b6e0ed98a608da808f51a856c192105b4918ab6e2a4809867fd8c3141d7a7672ec;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'he90eb89c237321e58a53bb5a080ec762ef9a0cc693a67247547e95ee3dd51ca4fb31322cbe1b82e6d0d56a4f7db307011d1b8592d523ddfd92a4fde6d3330ff9734acbb182d6d4cfe229a61306cf4f768792dad19b230f06903d65f5dcb974a3cc2ff15f94a6b86dc7c365cfed52151f9b33ba940bb6b3ec0c3421a5f4784c67e3317905fc4098e84bff442ac3a9ed5ca51bdc7467be2420fcfe1c5613430498fb3b6d2e9176ac0194cf1756527990c2a63c21ee6c27ef7633c7c370a6d7f7aaf19d6ea39571addebcfec068ca257dd86ce28dfc64f06193e1650178562408871c622ae149d30c9bcee1c83851280413fbbf02bb2f0d131dff69045692c897157db7846d86989a91f9f48c748a31effc87d9654479762eed5471e56be3a38c1374576386d960ac0193c92df7344cbd057f673f742de4d06aee037f5abc59fb981c7e0cbab033ac44b9e2464571603d77e7b7a274bd5719974aabe760bffc429efdcb9fb780a89f78a2f2b975c112c81c5d293e1289039190b1d36cc5b34003f475aef4e527a8f5b494ce5e49c4845b97a2436154ee984b158ed199727c2eb91f47ad9c828e7fbade3caae3e28612c247dbd034107d6a66220dfd499bf8dd3ce6b4628c1107ca9d21e0f95dad01fa182499993ac0c2b25c93775434bb061f98a4b15c8cf2bad2ebe97fd69c4814b1a997054259abfebb960d5288deab783119df18505be9426238ba411147a7142202393f8e38b3282625e7c9c57ea5afbe968093bff876f6e4865760eb936b45504fb1351f7ecb144a41a257b291bc30e9a960e9dbdd374f418ae19e767e465b22eb5e3298148d734164fa23d94b40152a182e32c2803ff404723913653bdf81944c8cd69d754e1515e81dd74c56404cb8faaae352046b923d3de39caa0c89310f2962efd9994634bd780950cc65e82135e507e93c6ac7c528855e622324b11ca24551238f06274e0ed22320fa18b1be41ae4432c4fce6b7f8f246e89b83ca97ebc11173d51ad2d3b5b79f6a8cdb2eb60520f6bbe5ad41aa89ca1fb20a5001575ac39c1504199b247ee3f1075774ead3eefbca2b320da2211d1810eaf9116ad16dc24f29c9fd0bb20643af33a49098237a386ff848b573582426a7074a52b43af81541b8a25b9ddb4c7b850aec49b4f5b9c8178f6c70b607a10be603b855462a5810f79cd28f5a4455a824f2b066076f2afd25cc91e148b6e313890eb4833c8b4c96120f8cb6ba00c8860b022ea2fd01c2e45ad73f1c279f028580ec5cf0f2701deb320b4ecf14547507de5848f47a05debc84cda8399048549f30ed2fb28f07ad6d816ec127431047455c7d4cc3d63c41992a7a22842867792d6751d33c3669cd1e5c21a018c1523445bb2bbd4b15e56c482703170dc8ba63fc4c137883977f92d5ca7ac8bc4a7a9568b57d28df03491977c966d67c7294a0047a09c8b5f1e2cca289b7f2dcadb1863d838230b0eb2c8f5b4958d21068ad71628388c57a88acb6aa950009e6c5456c32b7e03f89574c8701ff47773a45eb71b8d77943004c1499a96871de9aaa52f03d5466e7f0b8ee37fefdeac0957d237913ca6d9e1f45dad59d0aaab641645e10ad8d10e1efe5516d26860ab6de925a8408a5ab93efe12e24690d3494feefcf375f59261f3cb04fee2472587d7d3e1c4d2d38415de638c774818055e3bb5171ad7c4453cb88da97e79dc03d51b25db64ac1bdd11dc83d2fd12d8569c5539d392fd13d35d443ae537ef905ff3f1545ff740aaff3b32543939934d0ddc83678a315b4068298fb6b5524b46fe24b86b86b0dbee67ceb3596d3bb871133c3abf43ddcc321397ec00b8044719911462304d06426b49d2a6a5aa8a96d80b9efc19bb31cca146c7ca4fc849824107ce3740c7d17adbf9ec1015528064e929e2cd9c993e301c982386c7975d715ebad5712c8bf7143b37f5b5482cd37e3bc67428ff1033c0790f46c02f50c20060cc01b5d8219d82ce3e3ec76949bb16c7feff504d40685f6130757f41169906dec68ab10515c5a5b6114222c2e21dd966d1cdf0a55f39739ef4c888d778536ecb0aff1069261bf6afdbd8cf6f73bf8af2e0ccc786ab17460c000c383d7cdb0d236f44c4f026c1675e8421f5f6384eb12e920563544bc7ee24ab9c8eca7fbdb8b60ab27b5a6f35898ea73f0fc2ffcb18050ad29f1aecb81e3420f67ca313bbff0c061b844ee325c15b412115fbd3f93b3045eb01330d878f951db947dcdbe5728be3ed5b7b14305cabee1a87fd355e28c3ab1e1be229b7f1f574b1da2c5bc17282b24c6b1b92b716d097248a4fe9e71c60af8facb65024c65fbf3bb518f2bf3894e639c703effab0dba0306d69c5a74f8cdfcd92706383a51deea3ca209b26d3900373defb813f218bfaef965b6119eac2ad9d2964cbf9ee48d133265eed1b69383d810b7474245707e6296d997552953d0097b5a33cd6cc07e3fa4c248d2c24b2c54931d8f03724e6d4f2ed3a6f0c51c94ecbc98296198dccd6fad33ce55b1277be143964c04c7b2f77b5910dd6088dedbc9fd1d98fdf9a9e23941f83507aaf609de9fa5bbde35601a6120866ab3a8a0407359f034489b4b54c8fc04d1d58e6ad8ed26d63ef8bc04e1b86f176d93f9a913786259e6d73767e36081d983b8d544761a3dee12931a284713c73dc714ae6df74667453cb8b97cc442a57e78012a1d5c53dc120bc777d7e7f12983743d0aa61e59a01be1b0a2bbfd4e5394819753451c2edb54a1fd377e357b0851d565cd473bebbe450a96ba0c94f5c3a577236fa42af9d6973c952f362b14dbc7645c6bbcd95aec99bcf8d40ee3be63446d1aa46d4be40e7f14323f45a5d188e5426fef69963a9e8428f922a67d5de395f65eeab318118e24e5fefce1995d65acea424b581183eb268d0c42c9df59036da4b22d2e43c80a15b777e378dc201be2b5fc5cb1aefb2744332c85ba0ed431c5c97dd42fa617cb6fa6b3497ae2dfbbb1d8b2d24b63ef0782eff234c76dacf60aac1af5b569a007c705f3dbd93eaa1aff612153035ba9fc13cf3881b6615a9c618238e2bcb73d25e8a4a61d186462f2d2708d030dd780b5c29408e1f232a12980ea02a9de208cd60a31fd84c111ea3dfa415cf852606955b6161b10bac31586b34f03a6ccccd0b824967db30057c5d88518a41c17c03421e3499a8cf23b1a6f28773eba1f38ecdfd7bad0566b259de4633dad08856aeee9d03b076ca46908ce40c0b511ab6d0308123e3c07b68a258b0c28ee0977bd706b904fa54baeb310b0e7d743f174b6158fe61a2f00263980d644538aaa8dc1dd5d81672a05c02bd889be84d654dd5a58af3ff6ec4a868da21584d46729888409030ddfb775787b52423b6a498f0b2fdb5b7c4283f959c6c80f549aa457e528177d5aa35ee824bb485a95146b44071147c705a19594f06a74574cbd6676463a9d934dad3e44eb2afb0368b5e49d69ee99221faeab7879b821b62eed1afb3052295d2010a12fec27a5eca56be04c39c7b6511ee9f4d1a2afee34fc1e755b5bf02c18e3ae5c00dc297d25ba631ef12f3a32373cab74f29052c6e750e81159a418af053df8a18d010ef4f58bc0a803c498c3bcc9dbc2a184771f2ea2b52731d4df9f394e5bc3545f1bf497742c65931083aca4ec513df583300574bccb3b40cd6d899749e97c36e2f9b8cc3a5539dea9828f1bc4871e643af78eb6e90f1f4115606f3a7f69498b161daf6b88aab8b0b18f82a3858d18ca2c20d25f3d0d6b5f77ba4b90ad39d226251cf2bb3fa8318418662373ac717997a89ad1064b73d2ba23c62537c508403f86f741df693c839e0d78f8fcf6f2a87ea08cf4a34a20599b6167ea04b1d12c15ab0600d04ff1d217478d6e84f35b580fb2b8a35878ca4ec04ec67596bbc6aa25c6b0a9bc3fc6aa5d7d8a80855b536751821267347bb1a70188698d00f574bf630f3238e8af53a62aa2a3d3bd072677c6dbf5e31c172fbb8362f418d87627a4e310c94653511bc5e0408d86f9058fab33594a27a45fc33a0564fc917da6395b7e2c65540e9613374d2b221c3f8829e0aa1d613a24c6dfffa524e3881d0c597f32c7884029c683557ca04bffc4f3b3d4e2ba8f4ec88b737796c041381e621e5cebfd87e0eb23c07f142d63153cd16d2d3628093f1c8f1c4e8403d1abcc23b775ce16718fec1706e341eb6ba12cf6b318248e5f9e6bd0b125f9aa939c706f4174dd448e7ce634c09f7f0091a703ef44e97ec86fb15bb8bc48872803aefe711425bc2b292bf1ebef65a1fc7d2fb88de54dd4b7d051164636b700c3b019bf6cc0b03d030ae0e00b2527d295572080c7e365a5127748817cd18ae121db66c4b6c7f7d3dfd0518d52f1d36b12e370bf726f8e7277295a8172d80dd07199ad967c8a67a3bd373942cf7fb5556952ba65210871b769eef069ac883ba1cfc5e28faa7d091c2b363baf918c2cc0d8f36f5df2c74662e6e6ee5b9b271e891cee963115d784ff445e7c4b7a49040b21baea8320f661d9783f8774e10f77fff5feba3fc0e92c747c3f5421e4bf46e19cf75607bfdf5b124e933fcab136e4500c56ce0784efb4c52b7db79c773f6954913a7afd8ee334f2e53418632aaed0dc7061e5fffacdc508603586098662f5773097debf8483e3f500646738b574afb754dac46d38b0d46282d8f0f49fab08ab395666665e5fb1b60b64f7bd526f678027967c548532f2296dad07c9ade54eb2dc2d4edef9cad1a5e50e3c20b552b8c6093f040193d85635e5fe9830305d266c25aa8fce78ae7ac25dc33c5f3ea403b854279ebc1e0238e67d55e75c2ff4d6a20a9a5a4ff58fb68c5d5d430546dad315d9467c0e1ee5e8ec5e3fa8753c04826ec780ec637d851513fa0e5c811438ca942d71ae4a1056b1632e3c49bfab69ae86b182b49dd0c565e2f22d56d527ca2aff9f638b0948881a08b964e4b1bd4e1c94e6811ffa0548d3e626d429b49bb27a7847bf3789821b22d1310bf4619970cb3e926631133923021ce0810ac369ddc78e978f55b521a64a4d6e626c52519e7910a6e1e82228106bf3eefa5c88c04719a804866446bdef684ff1456a9d0114714b071287e67adcf2ef9714e63bb9ff0963778e0ee33d27c8c022c635b81620c6a3a0d0404cd3f583f8f5eb7fe92ea83d01ef44ed0d6f935c8d47974fb19398093b51ff7ef38c0ddbb4f86de3d6214428c2aed7a712c6b36deef4584b12e55be31957fb674e32508cbfd5086bad96b9da4dfa620b7210b946bdd4088ac388583a384c056816c181df0b9e9ff6fc60185802139801f9bfb0c9d2af3b2e3555cbc45d29ecb52838f3bfb05bb3ba1da02ab54d375ccb94c95293230712cef153b15e753b98aefedf705f300570259809fc7f62195232e30befce14c926181a5f248d9f981389a6a01fdd804908088b4ecf01190d6f9c750c6533e90be614db25109d7b39b5e2ccbefd90191bca3ba1286db55d66d5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h45293c7dfce4f794949db2f18110285c4beb13286a8601eac8452f2a02b69a7517d1907ab1f32287cce0fead9159e44e3a2f91d16d082b4d616a1f7709fec34a1632e4df4685c125bff365112f564f5ed13d4dfda11170b6a8b68cde590df1d56de509be33c4baa9dd1af876df9d96884e2d5aa4e9af3ee694f8df5ae29e6bc7cadc35fe3f01558614254b8f07403036a98e8d723a5a36f99c315258f611ca3c80282aa16b4a7d5910fff9a798fb56638567f51f47c97e764adfb94058094206a700c60a7002a8bad63a74b7ceec28f62841660562f968455c808a549082cb5b05314ca043edc3339d18756bf35758aee750f8f926dddd60fc71ac6f7bfb78bc2fa38c22abf7831b1dfc1979cfa6eaf2b9a6a81a4264b99293ff30eaaa6e7d5b2a879d2c4b1145c92e60dc9fdd1d6be8a3929d17a8545da3d295da7d5e76beb7741a4368f75c119815bcfa09dcb588ef3d4e732ab755874a5a20a33733174c7e4e8a77a056cdeff0b0852ee152e2c55f1de4a081237b83df25631e7b7bead05c2279f0784a9a1f888ec9e33802d1b95d3a538b8155575910cc8c0d0327a2dec0ffebbdbf580607e95b9cd88d6f35f091c4719ce16844064cf2733c424a6b5d68528e063a76404cff832d25a66a3d215ac245036b2dc79c304bfff02387f3d2adde97f0a61e4765dc8105d623e0401ab288dbdb23bc3c5a939924394217f700915858d26f0c04fea5a483a4d5b3da7a8604e4786ba1e2da5759f3f0ab3dc5cc66f6ba328275d691d71bcf02f920bdbc9af4478a4c1f846821b1d58ff71389a226593baafc6570149b8282ae24a9321c8ba7aa2e0f84e6ddf7cf457648eae9ce31b8143c3df83b8ee44a3bc34435ab9f572233c02fc08dee402d5887d69ed3fa268ed5a6645f530ec2f2e665ed6c95f9d614402e9d453b687d09dba9da7ccbb55c7a5d1de28058546fc879cb1e334867c62bb9c278fcd4ddc7ad9d7e8b7858a25d09ebea8a575f75dcda5cb3111fd8d16414aa31eb8336581c66d59b2693aea27c303670fc56042df84534015f83c19621bb1b74c4323c151f6c7ff05f62ffdc9f85d83fdad8d68ef428b2f3f52fa11ff1321c78896fcab05e9b26e87f882673f9915f8d7a6d74d4008ab527392e86f4ed7382bc4715b6f128cb3318942daae992df21e37afb194c042c999d9a5a8f00977ab10924f94d318a27c681376a84db6395907b09d305faac6c1b067fad5d3c4a066b239e4a54c890b44b38447f6bd4fc01a87cf3bab109dd82195b389e1279a907672a6f6a75764cd250ff26e23d19f0358b8af6d48ca637fee6c7217c801281812d447568d77c8c39383ee57d0e9aad148e60adcf880047435c06d5c7d50225daca69ce3269c31c947312033aaa554d2cfdd9f80d3c41ff5a09c6bf429f7d2e431da473108c6b04a0e742309943aec432420d08770f608a867df57670577179d59ad3554096f457ece10ecf18e077f3921bba5571a7bd978392d69d9bdeac8cfcdfdeb2fa0def7f69d95da1106924ef7a1ba4f87921edb396f95be31e78a790da01df0f5ecf8d7eee841e16621377f18b03f33385fe22fe63037476145c6096982611bfe81593bc03fa19293db8000c38c1178b5e755d71940a7d9419fe52529fbe2ebc3c7935569f49da0022e5c9c7df36dd6a7399d14219b5196e836915eafa42c4b15205d81442372c38f71427adfc4d616cbf0de18ec3c53ca77c0bdfe4baab19d126ee39e2fb5b790046a7d32f44f9589d3da6687281c0005740b450a9157674bb03dbb13a9b543173ec5e48e2e96206bcbca41cb4daccc3053bae159eb36a712fc4612c86afbc989c49a92fea748450753186d7d66b13bf7fa2a67bf34e9599d3ffef0918060e80e20ecd80d1a8fec04c897bfd1a59c6420633749fef4dd62411607fe21860af1f3ca84642bb0d2e9cf5769c9e2fba9cfcf82ca1394ffa88383a4edd175b45963fab18e12fe69cfdf3a3f1d9b9670b68fa27544926035864e54b64c93a76114251220fa9a18ec6331c1ec8acf408e3d53a4ef7465f9f07b57f33590f58f63623143aea0b69dc02337f3811adb327897d17b32edbdcf78d3a8beea2793f084c1640adccb22bd6401e8d37af404047d0927ada13b0e68911079f7d2d772011cbc6b4cb3f7254f40c6dfb1a38696697dbf632abf964f750ba7dec310546952af2b9827206f412be0efc7352d7b21a24adf2e48c192a134c2b8632c773553df76fec404cd6aa29f7f35f832e1162d61d214ea6fd36c3bc2650f5cde97d2d721da16b7fadc02b74dbb3efe11a58cf5514e66b86e96a85dd3356b2f936a6650bb2b4bef7a2c5ae158a9014c86a13b8ce755384f22c88b55223279b7881821c68f1fc4a573495fe7d966b9cf1880b9a118f05aaea6fecb382ac586343e527fe4bd20ecbeac8c9d018e0d32e8fe9d85abab8f24a0010933aaebee3e7b675a2fdd6097dd450c54c9328503f2a7b524a47fe000142ce3fd79ec0750e6e25426b614fa1d7ef67d52469531b515d13aa795b2f8e729333f6f10025d1153de6ad26e88ede1bc7df2d718f45002c2379609b1f96acdc0ea74f100aaa84108cea44ccf60336644e485806455b2b49893638ea746efa45ba34dfd8eaffe2d12766176cddae2d0ba82b952519a70ea356b53403b07638a9cf4ae464e80108da55c640aa6d9848d920608803e19f520999f7285d7f5337e74673312f223c06f908b3ec183474a2a0b01ae37d07a3fd64f95c04780c267ab9b2b30dc0b558d4506896951db1ae3fdbaf7cb13cd5f51183775b48a2c7c34aecedc7c05c7a55ad456387af86e00e7fec4ee71464fea98367dce258c1680d7bcc75ae1d57a15486cc26bb1f936e151c0a81856ab02ff46344d91c5cc89c77400a166d759bf79df21e3357b2f35dd7116afea82fc7451e0364344146c35ed9f1ea81a2f652c3230b02485a0df2a3662ff4c97f299157f6c4665f388c5881af272bc27259fecb8952df6ecd0b0ef664bf1fa0044a328a28b2731fbc8832b4f228e01ee176749e8ac98f14507c424204dc89e558eb86010b6e4dc1e07f3f921d5b9d5795a6b51003f030ee24eafadc7a4a0485fd87e21f14857309f63c4da56d9211d05166da0555b036d0dd8b8d2e7f8e2b9b08dcb69e6fb6c48a3e316339314be5a27f044683258cfb95115e042a28031472676e16d22162f4b39b337d0ad22e4d5ace2051bc3ff9c3b0ac9bc182d411f751b31257d6b71ffa0ff29029d470148f59279dc9988ed432e14610d6259ee4e7ecdd7443486af1ad9000c133e8e7f84b99eb7b2507976efeee4cee0b5a214e6ad754a835846ed8db0188afa56e2398d703d56a9bbe471e0c710272751b3870d7b907c815d7a4e12b1cfdd773b4bb6fd2d5e6a4203212e377a484d2eb3a7b55874c2e3fb7b25acd7247732117667347e0464cc588b8b14cfcfad4e8f18f8e2c45c74216709ab77cebf0ebea5b1baca351e05655570ac55d9d340ae272feef3f034b076286ffbe199f4e197720941eb967df3422f750550f0e760230ddaee3a7d8c0b231a2cad0ff4bebe5e2cbf42fb66821c86ed102b128c5d89b7427ace8fb667467e0bfaaeaff7bd7f984d258b6d2ab9d3e5db2deb99cd1099128020468953bb24abacbce866f200986c9de9fe4085be7e235abf4f119704e87b80a27a5d360b87dae1a1110dd289383ce6457bcfd1c61fda83dc778441bbbf3170e8063e7ca611309d9ede7db23966deafb276512113ee15bbf4c96a600ef51cff547e6dbd91cbb743ca450a189c2299bc2fb77d71f5de330bee44979d37e1ddc208e27da4e383e86eb91e0ac955af438112b6362b0951cef70fc2833bcc6be7bffd797cb8a21ecb270cebb6f432360a2c7c7507e8e66238a7f1e18dd704f50d95a0d94e1e174ea5addc628184d2802012098ad0217ddbc5182a7649f2f3972ce71904c4e98e87750653bacdf28196ffcab3f0fb17d1a9c7dc1693625c965cca01b0d038b88c27b89795ad5db28105fdcd0663993ddb97aec13ad257007970fae75038daed83c50aeb51df9e04a3ee8b889e2ebc212d48b00f1b23fd4a291d81473f3c4d2a980dc4666e24314d9699b66f5eca6fb157d0b36942500a5b80fe85f2b0b2ff6148a33a9e06b104c1a31228971cf882668a5c2be49f1974e471c7b39f3e6ae51fef077a0fabed7f5ec2aa3a0e4df56aaebf44a259bbbccf9ea141b96e1f51649aadbc094a94bac03c796de88acc624c14432150824898dcf783b98f5c579e3247e7d34468839f958fdaba313a24e86ed6cdbc238597f5dd82e7e5bf633eaef6689f52c2de2729c7a3384c63cf7b51d48a7456b9da31dee6be28e015f68972f2a29578fbf23025269195a83fabf0c3bdca8ebe2a620ea47be38b620e9e33c1a475bfc06e5aa7a6bafb8412160022c52474f92003b5ce18fb65790dc58bd202493e00869bfb828f16d36664e27ef0ba9862caa49ed60edfa2cc33b62cbd637135e86ec65714142c09c300c47aea974486f1cf7e4f73032fcadd2600d6ab4251e61125df4cde162ce8db40c84579f4efaa1efc6bb49e59ca720dffba7007b9765c141ad5fa2d05b28413c893e6e42543bd8f18b1c8e6222224685d9806292f3c40281f924944d541b0f192f938af3a9e90ad46b48e41990c290601106586ca5a444006ca5fcec872737a0c79aad3f41b6569ba615e1207ca9e7f76e0ad89b135ef8d714039f0f044cad7d101dbe08b4922d9c557d60b8a45f23434b532253bdb46191859c084b8fb3e0f2dfa691b5d90e43263f77ec7760a972962421fb2922a4fa8685f0c7ef307be857017fb449a390cfc07100db78e4e3b0cfd9b6a2e2575a1e3430f5203bbf044333a0b49f74c82090aa7434c3e42088f276fc5af02d08c3d49fea219b114c832b77c4fb2885116d8b6625c58902c64c8de91084859533fb9df1fcab058b017f7fa0fdaa703eb501a0b348b0156bf4a4e367a313786937e842273819899a27e0dd2c6ebc78aa0cbed76b8458311433705db6aef3ebb6055dd94a13a019d32f8cd070bcdeb672db46103e847e32059b63925ae3d5ee848a820ea87d3f74037e5bf61684629cb10e67a1f915315214ce639c5e886e96667f73ec282e59ae28ba9c55dbded1d2d9cf00d3660e8e6b30f5232cd43872086f9da11c8a73db5e00b3a214998ed0879a782d17beaa6a7d9f1ac6278d9f727bf0cce6c595fbc26e8ce3e9065389074a17468379e4f09ca76a3bb4ca9b06777fc96d93fd53f05093b9475b4a3e7284597649fdd626270cb6b755f05717e6c3feaf14b876caa6d1372ae47e982498773f398fa7f5f4b1a10bb6ffde427402f052892b315afe371f3b32a6b1636657e596dca2dc462dcdaaa094c556ffafeaa81a8b5f931fd822d507866146a77833847328e28ac4f87d9c1e4b0a87279327e76bf13230a936e6dd9381ba032df1d2780b4b06549dab557297572c4cbd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hf6583943e81b3b6d0c8b7e86e3497dd77cdc3e4bebd34bf267cc3f0883da2adbfa35862687d75175a31c18c3d8e8873dc1453ed51290f7fb37103d925169ec1f38af5dc1e82a4991cab04401d97cd9bf5d82b64c8469972006dbc9b8bff0b889b5b4d3169225af3e252a479bb29876bd25429f650a27043469cb50ad73e9cd55d49e34580c4584fcea7cd9995da8115f88a061fd748a45fa63eca2bd6837afbc346a805e70ff6fd963ee33b1217e8873329b6cba75b14188c9b117fbb1accc4957a7370c5cc0a960f8520c2a4c7baca94d36249b4bfc67919a50ba5b4bc1d101228a638abf36469433dcac952049bc4f41670af3b9cdc9936a2e586c96d59089411ac7fb38d9d36312dc32fdd16b166c51317621b7f182ffeb04dab4e5e8fe651b4ed9fadd5dec3e5d95cbd434f0c9f766bfc41cac0cb61827989d4459a9185183dec05c92bb17f5ec43ee250055a25f1a1782b8d6cd689c369bc85debc2759938a54a37c1d4a82bd0db7f2015ac9693fa8081b81091d322ca83730067284cea51860645cbed898690cbca55cd9d5dd240604ee03a6844435772970feab1bc99d4e5b422b2cab99254fb04104115fff7fca36155fab73b9582de7f54143d5a406548a6da372371f0312f6593c62499e442ac5e4233105a109defade9efaaed4f6065170ae0b4cd00302078b8f2f2f53aeb1f117ed90a60331d90032c4db95846c7e145f3b14442e5cf5cb085900ef6d0a1ce49698cde68e0bd3075674c5c307d6b8a11b8e16fc2f00e8ac462bbc01c6652047da8f3209510a7e37ff441248b8f8286e0a2b59400103435668c39d6b48b60fcf8c4b570a6c28c1e55d72658679940623417764c6a40b4477bfd41ac3fbcfbfd84ac325cc817a3afa62f1b109b745ccf3a8b25a1110bbf790236025c66db7b7d571431e57e48c4b0d2163098773b3344553afbe63222bb04e33ac3a622c070523fd850ec1cdb4d459dadd5c3a00c01bec9a2c65961ec550e82106291b833a4116369a936e7a233fc759295738765302b464860aae432e26f332ac39b20dc024c4bf0f81a9f01d3179d379ab0140d46325e4d9a513592be36e5da4d48ed09224434043ee86e131dbabc6456ae6027af412cbfbb952127359d0b79c37032fab930cb633f24df5f59a9a84ca72cfd2b02ee5f648f23f29cacf6935c079f5faf912e5eb7241820d7439b8232c2a764f6052df1686cac44515ddf41c49cfd3f66451e819787eed45eecfe372581b6bd48978369fc9699a10dffaaaf4f617d99ef658ae93e192be1b76762638bb46104bdf31e163b948d257360a22043a2354aef7791fac0a0caea36f2fc7ac69c72df3bc12e75e5800ef83c5ab6cb4febd7323506a7fd58f1e68ac4ce04d7453c71a30b51b7f9e69a8ef5b6fd24d7013e028a1a1cf8b2f72d085371482cc250edbc7c065fe2fe7fb3f4792468d4fa6dbecd01eed5477cc5f72783923c1e36e1b5b37a7284703d31967b970d6ace15d624fc702b77584cb9e52f16f07c66ead4a42a8e2c9433a3a7484fae2eea8a01aef9e1f369c733b79db9094bf49d26e7ca9366d1cc55b6bae04026961da7c680e218e2b09a61804a2bf0af8481983112090b6d26592d26436a0ad28ef865bb988b60a8a62779cb41ae73314809bef54829946dc23cd74729d80a20fa31d1685dc2a5874296ff9462fc1d37431478f54b7acb8676b0f1d114b09af572aa819155d9fc0ad6bb1d4b162239a9624d9cf88213877251b3ffb950cedc80d8c2051bca0085e3803aab7c57c87b7ad7bcb8ccc388decfa5180356bde74ffff899b9dbfa85c39a40dc72f68857e31f11f52b3a477460a4182d259d7161dfacf2dbc8b983b3f6c96c888888c0a8ef126ab020600addee7d6747ed3b650997d289df8e7892108ea4abb74fb700c25e84c4e52ab1dfe9c0fbff6b79a07a56eed64323db61681ed3f6312ac4ad2079d90b51b493d56353e4ca7663b5fbc5ae5fbcd2d8bd1a4c36d0aaa248fb26e1980641b55c3a48d0d9bcdcc54a2b506cf1e2ebe6993be053d9acc0ad396fcca69043518045efcb5bf23652537c23af1cd521063d4560999efc6dd91246d17d6fe51b2c2fa9d3c30f55e913fc61737920cf2289f3d56741b922bfcc6bad26d0a023481bb981888035319bc2c2c51a315144483d052c6375885ac9b84338d26ac3d9164a688af2b1137ec3bd8d732ef792d73a10f4e181bd97df601f965e2f4d3d14b730e05fe50dc3255badd9ec374596d439349b5171d9b5187636e2490c906f517d5e7c3366e4974cd1e3631d0ef5ddd9432f798555d802cf9c0f78a84b9976845fde63cee9f7917b1dfd70ba710ef32c388853d1d14557ec1e69bb627044261b38e465b64d61cf2b2ae2356d16a7342d9cbb457e801c7c84acc7bf512d9708f47e2ba3a9f178947472c12c72e8461643f4f4a935a2d7b24b7f4e875601c2bfcdf1b3510ad9027d823376c1178a61beaaef06f3e1816ea50722e77db8b976884e3b0dc0d840c7e133d0e4795e2e5e104cceed79a6096861db901851f4bd45df91f82b555cc91f1618f00e3e14bdb3f8f8fd9622ff2e13705d720314a230113977a4c6da6ae2bf160153d332c1c564751a291ec65b9b8b8f1da9e8e85ab94b9276d508c55f8344d05564742f7b2007d8adbb14add42de871ca9544ea1c2379064fafac1fd5d54c1e5136b468b1f09a19b884a33cf1a72bae8c42cc208bcd38618b42077a435184d493be4c32ff5d155f6bd8fefcd73a46f6763672435bd74bc0d51bc354320c847ea0590b75e4260a93ca2c975a5448184de4145adc1fc64c6bc7724e3d7833e9fcdb27161dd9b86aa2032e4d49cab8773d4d4a859855a80a86c17e096d093c1744b5d19b48bee1f8e1032702cdc1b19549f57d4a4a4c34d162082c84a4807a980ee7fbc29e37b9745adff7c37b31c2843d785c6a2bccde0afd1529b9994ef7f7ad167ceba393b8d86d6bd477bce909f674b4bbcf5e60cdcac037faca1740a0d8a4db66633f082e1b03ee221f430de4c5ffba9d156b580046f4451394cca5f7b01e38e38ec2cc9174d152744a4ab3e1fae2d96b69ba394af7568d160cc09c94ed5c5ab463e526402b34e84c7c54aa61b00933af5177d7cc52edad2fde9335d63fd2240699e2fb691f0e5edb0c213175a7289f7d6b3dcfef23547b6cc541afbd322a760686f45f977304a365d6cdb5bdaefedba4d48be034d7a8d510afda4c8e77f3fe3b3b442b38d0218c952b1089a397aaa75672f71f0ca21cbb05e92b2dfac5c002fc97deb5c035ee9ddf8e45417de1692aa7797d32e815ab39f9dd953561bbbb5b943d5bab84beaf8eddc7f418e7b2c3d4755e02b66bc1464578c584a666f59e46fe717d662a22fc5f5ada44b77fe6b211099b3dcae986ff5535468c394c05267bc82bd5911e0453a29c33e97a9a70f79ac2b8ac56e0df61f760b092857204d1d440638ece1279e366bd77d39124d9dae9468cabb13daf9d8bab98dea4cb3df817418ffb286181490ed79dd8d4b687621e90a66c9bc1847d144e2875dcf5c21b7da63ab60f14c98a7a933aa35ceb43aead04d9cff119991a842e2651c9bb5846193159f390ffe6283ed0bda48e8a07775b8f9be183913ca2acc2d3fe9177105abe8ddcb5b587d027086302d7857569495b271690ef29068da706cf5eac8a7f51e3707703cb54cd70c1c76e5261fa3d713a4a5b13134b878999c85911af5074d2a615aeded800f24c2ea41651660833ebddaf8efc84343c11035254ee53af53b7091ca928434806e303d9be117fb36981a13573cb5ba347fe96258504c49a7c115b818b11f72ca90c9cf1bac57ff20a0721a23c7cdf0f311f4a4284c5e4dac36590850442a00a5e6d17ed64f5c6986a0fdfa7e3696cd6535980b2b3b6a6cee76d360d5ed379ec87474075aea7296f57b0cdacd699e2a7e67a54fd1b8f2cedb52df37c1d7c30fcf9b3fa3e100c325f8cfaac241ad03027f1857013cac9c03d8ecfaf5ef585843de90c69def420c72d9157f1e268507d24098ef8c1cba7feb5c21e44a1e19557ded07b1b039a3cdeab47845d33d0490c81141efb9c9da8f21e8fa361b8892fe10fbe46bb552bac6ca2aa62572b9b4dbfde2119e47635329c9f98d877a8eed7969ace6b1c20cc86994012c2d5e9f38104ceb9dfe85d13f34c2755fa922a76df948ad911484244749c694b2612dad217644c474f53c1302aa14c8d78806d2b3619ac7529564ea78507b694ac1477e7e8b6268dc354b6084e8196d212a343b4ba585e4e50826832652ff0040b2d5e18398559298f86a2518516f2957d0f142d246d59cfd3fe5c47924518a5df9fdff4a0413ea96bb4d5e90db505fbe505135b76e6bb3dd247a3e45a3cc3cde06cf038e243c5875ff16af74a73b24c857c78432e5e625485c61976773c89734873aa3711a27b3c70eb829ec9986193a83ef4e120dd36cd029894244dd9ab1e524a5fe2e67d54c3537b95f2f2bcff525571b7b8c87dc99fa2eba1f01080a08c16e755ac27fa5fff587b9b34a50af0c4b4a3467730dd4a8e3b44a60a5e1346e55fc1cbe38a2698c7b17320cb61b18a51fb3e49fc2e9f75e124f267898252897e4e0f174c43d28fe549319cbaac89427daa1372d3b1aaeb92f1426fc1d60bca6d6e022c7bc9c4dab10f24f27321520d0be66dd24be02612cdd372e6ea73264130b1d9756022a6ec1533c32a6a4f72d70114c6c4d319f1ffbe47afb15ed614579b1c50be63a777dc5b91ea8cf02cb369c947bbf308a51e08e562fc3146eb257bc85dbe74005104bb3bc40f31408ac20ca8df53e6a3c50796698fcf0099a646ed4c6acb08b2721da68be6add9e2a0a156ae6e1b3e30e9021e2054be36c62dceeee0e8a269259ce6e27665bfca33cf3591f5aa33c373d443884c7a0838b0a7d39cb5e29c48ee8103af8cf938d9fe4ce9db467e1da174c3b1f3902adc315ee070da8ea36faff9191d2c8116caf858b198be4309e315ad292d6ac3668bda6bcdc778d3650dc5ad7e6bb01a57f34a9be3de26e25ba27e6361cfd7ef102980ed15e62ad323463f87e2fa2e69f345862e9dad1587086af779ed3ff95d5b6bea64763b737a9768c6c07f178e4cb3bc4db090777e15ecb278b7fe445dc0c20239ad71f01249108b721e1aa278dffe2bd47bc5a7410a5cad38b41493316a42060e682d781adde80e419f6386e6ca37ba6ed391d2fcdcc286edee58d588093ea60a7c71019180bec8263486cccc695316dfdeaa2b10acea7123f4f706c08eb5cea10c2c4f8ca5b484bbbd181ea653dbdc20d40593f7d1c67ec3ba5a4c0f806cde0805aaca4687bb85fc893518263cc2ae275296cadd11ade1d37cfdd59fd77af40487eb0ddf594bf4b4471eac617518942bf9f002badad6eaf72175fe98ef390b66acbc9865de40ad9920d978c7f60d98b31e2e4cc92e6e009dd4a2b0a0b283d39bba65bf6af06246c409d6fe;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hf39a21e89d9d643029fc31e40f11bc242382357ffc5455d4e8beb3ed43596c9d531a25930d149b1c56a1ed563a92b1528063700fe640968855325f533012cbdd685c2bb7c70affc78163b13e78964cca678fa949e5ef3d411a234bde7e6e35cf7d60596f5b0ad406b73c2955101443ac7cf016c053bc5e3ddee233a6fcf8e27a584840b312ea404d2915903195b4841b3a93a99db73165c2b297b3eea5c590f3f67770f6c7ea39ce3696563d32b930b7e84afd8cc172899a796778edac40712e35b192d8f83c9cfc3c4447760516acaa9626cb7f5271f832520186353c31575e5dc7602cd914a3655871fd6e92ba12779cb5f731d572b2f6e9722e6b443400dde385ce50e452fdeb05cb3487375ab1f837c07f313b980abaa1f1bfe2c295da8a7b116f6450dfb82a31bc202c19176b8bf04d0c75cb8d3859c954927ed88f6e2e183f3cce9f66a7733ef82af9f0b5b14f18be2c7c81fde9a43dd48068da79b6dc1272ce2acdc081e6a944f1f0bf319868b402318eb35905492799490b0c6a614cd5776d6e506505b0a93c548bb6baad6859c65237d005ce2d52044f637d723871d9ee8fe3ae95fb3eec199ee11550174e368c00be7a6fb5fe44f05e783c8496748403c2eec0a70304f4c630bf0642e4b7771307b275e6d83f65615d5d24c02f908a35ca5c9b93baa8fdc100e8160c343a8b409fa9f64d6e71e3b3b3971117fc65912602efb20632e57ef2fee557fb25400e06d0d8bb9fce551c7f75f9be1b4e435ba64a09bf2ff130688e6b16ca6dcf5087476ec9e26249d00eeb859311875e68b3cdefdeac8582666e5f447d02f65cc7683272ddd9127732ec83867f3bedc423a53cd181687c9ac604aeab27d43c238bea49c056fb4d424eef2738ffe14fd8f6bdb311981d87f29d90b2a1f98eb3b900b2d7a3c7b00320ef7e31b3dd9b317dc087c796ff920df5a0c21155ce381fc672c8b78b3fe9561fe9838351b0a4621a1111d67abf501552d73193c2e9110f272162cabd961bfc2bdeb4c57a105ee41ba718852b23c4cb479f771cccc98b5666ec9a04a369b2283169ad3dfabae4f7318b1f6d097d9859b9f5fcd4400050ce3beb9ba7d79630564a636cf634670fa3fce5777ac621531c85fcfbd3c61a88fa9b02d8445eaa2d5b9b817705cbe5a10d1e066a2df1444e2f2533a9b0c8d940c777b1ae490e1d0551a6db68034955f13b93a261db1b122ae7d76cb6cc86962827cbd8195136800d6da9fa8636ed1e41d09f09246d9df7c805e0a96c5319ad218fe837d57c7900eb8968a61da9a90c675f69ed8bea1656e049ca6495ea9f5988360de0348abdfdf1069dd59d7a9590eaae138fb962e647e0699f9d7afbb78b63d077e3611e6f589c61297236c23f34a1ad145cf1929bee6eefd32ff4b72bd10a7e6272bdf121663c8c97102fdc85ec9caa06676bd7a6be10aee90a696e118bef3cd1166dd9802861b36aa423a441641b88408db17df934226465cc2d05ed8ce6aaacf7eb818056ec8d4d904cc7a765e60c3cb4e016225971c5a4fa725fbf4b1816e5c036fad1f0ec28e5361ddd7f5cf582b9927ab3bf02089d8aecb90451d6211338f58a7845b4292a3c48b7d34926ead0f5a3d5003bf1fd0a6051c9eedccca10c0133d4a7242567dbd71da4937fd353697d9990315491f0240f4982e2981bb05ae51a3b9c8bd53c9f063d67e07d9874578214874e22192a3d69a9772898d34c5664eab3d84429382e368b6d9685f40af034b2f490915495f7e70f384d28bf7a3bded7e493540318ce2fb46c45b1d594d2db741b370ec1d28e59f4e53a8c8010afc73b61cd0bcf88e0838981873f3c7afbf9569f97103c2651c0a484d005d6347ec381b59bc842bbd8a83c322c3053dd1b526c0090db422b8e80f1a9ac059ddc71004e489929360efee15d7b0bd2b0a9bf27f9db07efc42450abc1d52390aed98edc9d2cc60b38cfb17b89c4553599f0df16cb1a6ba73ecfd6741f33b242a3c1449f5dbba71423d041630c8420e0156576e6992da4acf21d34bb3ac92fb6b780471f08f7843c06101a3aa22ef45a90ff779280681294e4d48fbdd2ba693f872038a4e1052b511e56c304153e010b2ada683791657c269a1ec20a919068fb5fca7067272c8f589b79ecd00fe5f2962facf2f4bb1b418c386dad6be8d5cbca8baa0d6e6581066d7445bdd9582bad2ca997967645b23aca70a7eb5dfa3368700cf5628f72323f40a63ac8f3ea71ef21cc30b0b6bca9813501bcc1945ff49b71603c3f246b8807fe3ef416523abef87f9a18e331f2dc7515738e2d9dcd78d69c4d9f60a601eb3bdc7f68c429653fa1575fbd4fd0d85c22721a80dfb5f15da7b3f12ce8a1063594c239d802ee0ad2eff811db02a8a2181d2190b2ad1f3a4b9e40d5b34e7bb9d985d07252b8fdbb10a09f411343ee9d4968221d846701e34a78ba9d33c7679262a2d5956e7fe9dc41cc03a87a49fdb80c9d5b6431f181ecfaf2553d2647904573e53eef2740c169e77fd3d080d4d360629c3367879f4471a8a054a76122538ac659014f3e2b33921a5232f349066b62f775df84bb8ad52a8d14f7cd0c5d4430c6cbd8290826173042a82bc982469d5949eb8bf2d4011eac5d77c762504016060a3965a084ed1f4626a798d771f8277eb52f8b8a28511ee4710a0a0e5305b5479eaf7545079845aa3b83f2c173afbbe05b485f779524c81e0bd7abefb01d1b2c84ae908ee0b2092a15e111f5f5d3c637c701ece1aa1e1bec4aaef844acb3ac3f4fbdcf3003547aed5f6c265abeb2efa97f93f0edc84c5c7af25c6123606a1f8a8107b134d6d38c604bc1bf5b3a26de7f2572fc7ba683758c573f27ee3f79c95b0417f86d72a17869e056bc0710bf7c8d19b638921f296c78bee36b1d3d1ce212d977cabd306d62220f4d8e40503f0fb560cbfdf71362f2ddef96ca25dfd52ff26113018b7b4c87775c0bd7cff46aed332943ebddd0ee53f5be5bdf57ed354881f131097d05b98db6f33e36d40bfed648f6eca0c8c90082df17c62ed6ae70a87baa414922b02801bdc836f4455c22ee9e787e09a18dd8d1a81f1b4e05a8aa2ec51fed852c15847781b632fcfd41bc0f46399ecfe97ae15353b24b57698bcbcf29d677b72c18180bcf5e09c0763c44262c58cd311185e9f259fbd40a64c80e538620153869516d30db96d4b52da1a1e3a15a27ae3253e2d87a4f9fc2f394e4307a2e46a757a8f32be56becfb5cf926a56efc8bd9a96774e1ab91033230fbf9716bd7804b9f5312a8e661533da5e2ef548800dbda63b9f60874e00e22adf50d82321a7f106416fbcbcecab2a786bb01790c036e11fa30898e8bdb2718314f971d70077c81eccdc6fe55d9664bfde01d00505263b43820e070ad5f65a5334dd347dfd1db88845f571824f638d29ab69571b575c0724fcae73eae41fcaf4d96f4397625dffe8777f525264c1f67debda0d6b823381161b72a4b0019f8cb3a4bf4814a3aa42c99f466babdecc021ac1c51a7213c9a19b784b3ca007485df3e227eb2d53ff45aa6c09e77ce0e7fe74fecb7dd4eb0b99cb07d00c71563883a13af9f09927fe252f6859f6257f85d685dae79c6e3f7f0365aae1d1d9fd9161d12a22a4b224d9be406248fc0a7c09ae1f783f1d4da89ed61462bb91a3db8346c7aee045be3c198a747ff775622f5de63cd56c115c1e1bfae3d59717f244338d92bea55aab854aaadf3136e997564fd0fb213a98607a012ac13f83bacca1421dc13b24180c2afe7f64c66387d626cfa69e92a1d60768d34e7b65553e2e242241893ef9f8cfc7567e44a86266ff4af29465317e062201bf7e868f7049432b0fb603bb400981645dcfbd326b0bfe44cb46d711897f8a75f8aac96d34fd8ef022f8c399d009244c401fa10c776c1f37de23260c15c8a1c9a68dfc4d349c473bf57f51bed8386aeb6d64f5527f865f744fcd8852688a9deb1cd0d18b42a55052a733de87c44fe2ac630d1da1ccc766c09e4c6b6f4ab2066ed63b53a7880bbfe36ac576b828f2fbe572e456ca804cbf4081e56247484ebf52327fef03b9a229e5c1650a1a045c5cc9116adbcb4f9da1bf02d1386c856de1989111129646ef641878ebee63d3b0f33230c6b44711ca7793950230140bd01d6d257fe7df8feebf417d5e5cdc91cfd062104f34661b066dfe3c57cfc654fd59f3d3ff6c576588b6c7df1a705e04c758bcd7f95d353e8ff4a1956e298657cc3997b8f9eac8e34ed953d05cf86501854bd47be363ca543a572203618ed362eb3f8041fa73fdb4bdbe32da2d3b792c121bb489945f7dcc0f2805d3bf275478c0c670a0800361ae25126a2fe499eab9a23d3c9cd9f87741a64684892201e342da6e150d0306458eca64af0d87f8bcf90bae39c1a597e1db4d1865350726c1eb9829924af313848086b473b579d8836956680499357c74fc21141326ffabd4a4e38dbf73f0d5ae5b11b486820509f9e1ca20218122a3f335b23295dff41732b3f680184a97d714d8e81954bdcb67b0caaaf64cb7f84d398d47469c3842d3e2dd66a51e5fd0147969fbb1331a4bf75187411db6ae49ada38423576573c0480ab21f97d6d44812f06b0974006c6d646401534ad7b76bc9e88cb33b7ea91dbdaa2ed20918ead8669c8186af05854833eda5dc1faa307f9e11548517c4e0a0e1df97ef495480c879bd96b86245a4b46370062cf414346445a8f21dfc3f6ec3f72ff29ba2b8f04fc544d744ce4f98eb3df168b83213663ee5a6614a99ca3d33991b022dbc652ee424a3ae331e9ab7d3138827b51f4c5e2abd0341c0cda14569d62b367a35df33f018710142322ea91fa2a8e4eaabd6051133f8e4210c611ea0ede3cd912247ecad4f3c0c235b3f9472b02c80631bef973448b3c023369e3a0979fc28157abdd8f79169bb9501c1a54941ede0df420909b150afd2bd240cc69f0b419d570b57e54261ce8ca9d1f4e8fbf0bd24f0e3b697a4f1e6e4608dcc069e99b2f27b42a8bcdcbe7eb3772a69fe5b6c09484e34757c4ff965e6c7973952297cff2e0cf208e1de968515428c425539c1a79b0bf9dd54af864bb4ae5dcfb2a637f62991ee30811a1d08fff24c1b4ca04e64696a63441131b2cdd172a96ec82fd579cfe63e46c592f7111eeec74d4251f4ee485fddf23e91734a576f9aa419a41f2dc511f33aad074aa1eaec6a57d624dda6a814804a01beaa989e5ec36dc2c280a6e339a93e9ce05dc4a5523048a135a5fca7522cc1e233fefe8066c1de8a4a97b327640b3394d8dd3dae3d81c8369deeb40f7085fb73f8baef1d3f5532765655ec50b2816d75409c6e4279d55124da2c36f6613f32f4270ae892956b44e50db201b0cd355e83bcf1f7ec985f7ceb06b78d837373f21b0c0afcf6197affb40a6a6886857cf89be4f01dfd05318597193c8ca8d8a90dc3e5a3cba65bc6a33e054ef3b81d4ed7fea90dc301bfff900bfac0f9ccf3b6f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'he3ed3ed587e0fe62bf35bba9c26becd6acd02eddc297926d02c6ed33fe1c69b3613c7aa84f11952350779d28c70c717a93089321797be7aa4086e561526acdafa58076841f98c638a1db8ad1143d6e457f15328d01dbd1dc9681fd8804e189bd85d55e460fa3c8d778070febc626593afc54829b20cbeb549d3c6058f4955399786c564e090fe57116b973b20125b9cfdebe7dcb88b1e2d682b767c9237db04d3da14f4d04e91446aef1112bc379cf4bf72e00361a52d1884224239037d063d461156fbcadcb54d496b6c6852fea14339d6ee09755eda6bfbdbab2dbcf0eb2c33b709759389d02027932caf4ab20dd32fce3ab1b9e4a718a72fd1569175936fcaa18b1839ce068873b6810346f84bc3bc30396d9329507a5026623e24cd0b7b9a3fe72db21b60bda6d7106e3357f9ca087cf2982be1809d5543b643ef5d3d4f805a4d4e70e7ab8ca352b0c21cef882adc4c3aa0d4ea33ff013cc7e4c54a1b86629f23bd88b7dace57739221ed7c75c0be556a39ba3a2c986e1c75e95e94bb3e21558e1e095470703dc80d7152f5476975dadd44bd0cabd8df1763bde366ec3a2269dc0ffa1b8f492b3afc8c786c8f9cdcd9ad4f000c06f114f13e3e1622b1c16a65e9bb864ddc0355bc5eb11d4609934e459501d41254fdfa97be877fc9edcf9378561098f368b705b70e382d40d1fcbfa1c73b6cb054797ba20d3981ce6ea2f9b0cbb09868b0a5015a2d7ee27da23eb96cee23924a4ac0ba6243516a86e76b72e3e04d8e9325a8226f007b7571f457c9e8e88daa0cb9f61955bca5da2bbba3c7b64e1a341080bfc7f3466f93075fc0f0c09934eafb3643ac26531d1c9db520c9516633a3efc1cc73a8cdae09e2a6208d7e7ba3f3bcaaf7b376b15a80d80f9fc54625c0583b3705ef78c2a25c0dd8cbbe8b7628b6f2177a8f119a51ac0c1c42aceff90f4232ed7a5f4b65e2370c6824948401b5892f46ce3b9d7dd6f1478cf0358b355addba3a1701790e95b507bcbbaf981b72898ee684ada39321078d4c8df07d3d054bde9311dabda869468cd165c713a19a61604aa17f6f663795e412decbec6d9fe08a48727e72a9bc52b2632b249f23ad4be027f4402bcc68aae64b70f90466e2259a040d0423b28503ae0f72000f76bd12a67b4908eb8a32e63432a64d7b6c49ac0bd3aa4e084e62551c955d056a0c38b188396031c52cafb30ee5d0d47c852059b4e3debdd5ba4983b97ee23cc78fb1ee0a29cde7d508dd70721d2d5106949603586ccd5a6d563f8dce3da41b22717b1edb0a3e988c7693a404df07f0bcc45e814a964d755f8a24a6fae6d3395980d6610f6c8eacd4074bcb15650f6ea203387b6f12e1b65370c7c73fbc6434fc4b6cea94080c7e3fb52ccc0d1fbe671c6a3df7c7d4d039350db83473250025b10cc05174c87cc783e5505bb48a3fcd8cc47ca70c7556c66e1c50a11ee82564c18df3d1fa0b4fa30f4fa29073f4cd68052182d7f44e0c255647c030a872d8ff237c2d9ea7a4e3cf65d42fa8f2772b2a4264ccc9d0edd585e8ca45ae022231241eade727bb9e2d5a535488a040c84cbf22cf7a5645eb8d403b3db37b3855f3a5eac0dfeafbf2fa73098754890480ddfbe5e0baf835086c0b547868137b1fb952f6cd1a1e0ef76e652688065e4cf8871b18d1a8136acf5583ea0e1f05d31832912697aeb7b296b286b3b308282c4cca03e8a2b1fba8c1dcdf6c32e1f2a139007703fe75b4c82c0370766a7a54b88c410f965e5112659642d9628b36c96b64b9d68dd0a7b05b40b66f875ba45acc0bf40ed02c53db060e6b523c4f217afc772e504b0f30d011690f5921107319858ab2e171b57196c010700e8bf9f4be80a39291705c2a86a33f878277fc08af392bbe306a0145f71cc6ab1d418f569734e95b2394f487a79e7dfc9d64d9547ed1712a675aed42b1ed71a48d2d571e79ae76106ba73214d0788118de7628e3d9a8983ae7766e9862b8f3ca7813a44e64307dd347c7d5c30c8a3be76ff6d4c032d40791099ae0c5b8e599180ea186dd72ba0b60f5fe0dbcaf2e1bcadf72473671c12fa0eabe70270f0f3880bf751119e53e19527b2206196b27afc0fab772b6e4820ffc0ef64ef45ab3d3d6ff85a391e2f8e87f8dd7a206ce68149365296d377fd39a21f8b7ce1df5fd836a159f24a44c1dac29b3c72500f4e65b802192414df5d30fa405b7a3b09d5a5b557cebe4283571d606f9ef1bc4893310c85e3e6817305c5a1c77a9e7f0477ce5f2b493ed8593e45c70f53bb430bca7c613029d5cecddba6ebd343a36fd0c6e8a46020c908604231c0c2e7b4ae97e9a53b0a2ce0dc409654960144c337e468a7f2a50a41b90387d50b7f4b64dbfe25be6fd60ecf33d39b8b7e16463395bf471e8b0c4aab73564bd0b6266528e6fdf81e6c5358acadcc64201f6b5350e3dfafdad208ed6bfa4eae3093a3f053fd1728b59286aab39ad56617ff2cf6c443ac1d035c69b74af102f51d6d681e6504e85cad4c07748d868631ae8c38e88ed35a2e00d76c55a49a7ce4b595561aedddf7100e2235a5bd950ae27359b8c9974b997fcc60e51d64f992a0389a41f319e89ca55f19a5b2d362ecfdc2beb6734d5bea9ad6a422fd004523e7f51b3da4baf76fafd829ab95307a053269218003cde5a5ff008480fa86743af7c5bbc6212ec5beb18beea9adfa189d6b4e7fe4802697e91fe94c05355eeb7b7e4daa40751ab21ca5b386221e3e425a308d53938d6b04345a057610867d309203fd6a2c7b234fcb6224c6aa125b6ccbd4923dbafce8b936dc5ed3eb4fb3b1196a4268906d5bd7df2ccd29bdea0ac1477bd597c4c3db611ab242f4b6cb8145842a9f28ddab40dad659a9ccf539e1e7b1b524fd1d865c5f6ceed3204ed080c0b161c29717a9e72eace0f7272afec80b9e3ff6c9bfb69fa679bb441f2b3c7584f54246a520dd8dc0341e1e956b26c4b6add90f8669a815db4c181cc393e640a3d809f4a40d60c86f10f75ffc3274a6185d90168de2b70d5322a67cc277d26e36ccaba36f33b3d226171ce815fbc3673909056c37bab59cd1fc0250a9374f4186b726f23db9b07bf86993839ba1767a56992614acb0152c40c835a5b3779375ac1968899c1adf4d31321d4e46bbcca1e3fcb6bd090f69f8a7b1db4836ee5ea841a1273815ff3210cb60b5aa90a85f902c82c07555c1a6400ae4c500cc0168c4165e1be650ffbd96760914fd93f3b965d01c9dc51d54fb0abcf244f33c97979d81c90cfeae6d191d97f3528bfe4c6d17f390f2f04bf213dad304caeaf9c126f40391b0b9c7e1a0c7b85caaecf02122aea7c067bed512c17c87e6a83a14706c34a045692076bb8049a49260d111e28d4df9587a7175e05dc2c7cb958a2a0a11b36c8f5e11309c45076d75908a8f9dca3eaf7d1b51c320b5c66245121d350c142e72a8eb4efca0b06f00775398224b74869f028ac3c2c6884ae0813742147ae942de46259f6d7c82ef1ac94b5e65b4eee0b63a3fef0a55074e09058e2938da6a9ff7a85468bc03381196a246e2915573a9deea6cbe88d033a532a6e3b332ba520ccb294eedc5ba1c199df0faaed3f74f58e8cd45d8a1d70c1cabc5163625edc33729af1814322269e9a5617d0e58b9571428613ec168d85b9fac8965f02c85d4cc4bc0d8bf94fdee7666315f5b22d0b96023575ffa909cc1d2ef663a8eed2d2d4365e6fa7daaf78775935b25e2e98597982de427113f406576841eccd21edf8ca2b94a96747e1040152cb73bb0fdfbc0d6b1150098ba61a0da82f8226fc6ae8723b446b833c917111b7c000a096b7dab13a7e09b85a8dcd52669a9d84b67f2716591f08fdad139debf907da33db5ca9723ee3cbc7a8de6532a1dd2698c09050f9fa7be1242f1a7f316a501b7d91267ca60f632960b7881378834efe8ab50028f9c04922b84c132482afdd67387a1cf73834ba63c017b88db2dd559c00fec7ac451975898fb9532f9e9c05af46e1392d2d988f52ccc249a580758edfb476d7418537f507a36b9704a61dc2c6240ea11abcbfdccadee912cfd6d6c3c2f9ceb6c62abb5578ab2a69c12f3d2fd028b57367a1e11bcffed581d56aa33017dd7a957fd70370874b0cd8f73f23bd151397a01cc06aa753d1e335ace08c546f0877792e7f5bb1e748074713911f1e8350d62eb1dbfc2f695c1c3cd65e33fa0795565373f079c9ba2c7414ab9ecc6fb0a5fc43fda50fcfbe8d821c9f7b7d6c5c75a546680fed2b58ad0e0b2f55331f1511340d786872c48dfaa83180b6ac0b02e390db29755eb6df8fa69d86753fc605febfa10774adb714859ad4f94f34b6fb23d5ec5a60288505f666cd1b11633430ae8c7eb4993cd93f1c6ab2beaf11b3bb518567e1579517f4299459b4d77bcdda62199d1ca76bc4775f6f98ef2460252247ba8a4b7896b57b535ec98c283e35c587a465bb24e77ec8003ee473da41c5dad6b1dc7ed91e5127b82d40f7e8f564ae451981155529e4286c4cf1df2bd45d4a14a256143503eecf218e6e34181d8e10af3603465230c38e83db041d767bee3675bc255f83e78b37842697a87cd71772f7c4c5c09380902efa3c362c9af602ac26f0b76875caa60bd29f460c8028b7c5ce92774f952cd121599b9a43c58b51b36c331b7231677ba43b3a360fa9bcdb1dd0ddc2d442156c9f900f4f003d11fe492b882f06facc0cf9750ce415e02926ed8a5d9a5e6a8a3f43a1192277d8ae671c25820c0c361460d9ad906039135d740c3dd243a9ea5f42b8fbe03fe219ac51729fb4a9b4c47ca3a9af48a85a7b3121e3d199dee8cd43d7bc32ae9f0de601cc50fbeadf1c92da058bdc7be7c299e9429c0f741cb56b8d82e9114385ad2360ed30a6127d20c93f8ccb23cfed6de298a1b8be5f21db323e75ab15d25f70d6f55899239a42425db27be132cea341f6e17a4ea6e4a719da990fc6509bb97ed5d74d8d43f496577bd629e65e535ee14cf55cb64d0562d3ed0a79c5ba73a2e014c2f609669b2e95e8909d631612b4d56fc397141205579f4f033b208bb0fb7366b91adb651fcfb1d18fe6a990172a0df845c5c17f874ae6ad0347ebc47adb982fcc2b4147447952d9b2dc31136725ced24fd2fd71103ff9d6ea671d497b89bf0685b0a90870eaf53c422c9358b6e014d671a5fbe4a870a44fdadf9aff29dc813f1d82611484d3abcb1e34c5557526283a3023f0d670468175753746a315616b2c0eca99627cb1da50a06bfda37c3f89d8eed9c8e7028352f59831db64b03358ac9d7907e47b4df6021545a589a72fd386573395cf0374bad80bacf391a8124d4dbb110c4589958e7b88ec8d34c8a7ad1544e207ea30f7ffbe5ae12e41490d8dcef00ea288b4bbbf989e21dc92adf4ad10c3135b10434804279ba078c62f215b09b6c6af52b8c0306b88532d0736164d27f319617f9ccc7c03990846b8766ece5f1c24dfdf86151b03ba5fa11affc11;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h4a682920e5d298fc7e66f51f992575a0dfee380d2d9a98d78705f85d62623e01d6e5b95e4ca297903a8e5eaf5b946e9213eb107171eb47b0badcc93984c5ae632c85adbf07ecd2ab89585c84a8206824c3edb372256a01a6d0255324686e76887dcea45569726a01dce55450e9ba23365cada800fc33a66025797aa3aea82091469624dcd45ec20346a0053ea3bf36efb2fe8b8f066ee9ebeea61e1c5c0bec6ffd17f14b5ad1eed680e571b2ec0ef5d943d675ed86007426497c0bf78afe36e445fc32bbcab30f45cbb88871a45cd255f5c7b3cc819ed5617a0c07de877c05345f71c4962ee0e00c5d440ab8abca93c28540965406c903e8687ceca16be9d079b624bacdf5530321e720dfe4a46942ade04c6a053eabe9c88ba9adb62ac73a0b4420b6655ad235d4479d91ea56e055d7e79c457136b5e59701c21d2c124f9df181afcdb84c7c3ab27826c2ae6ee935f465468ed6a4da8fa941f119cf8f9e65d9eeea387c0a72beeb2cf2fa254050903fb9d949ceff0ae75ccefce3884c33ec65d641ce7825bceb2699bb6d2aebc4cff850907645140a2686faf8704005afa1f8ef8bb999cdd3f9fa2da114a56d4f50c17a7e884787ca8f80cce47bb256bdf3e144819dd0b83ba4d41e6d56fa736ff582d753c67b30fdb0b5dcde2fead8909989505ff391abee8a00f514a85a760cdaacc47da5d973b831b70e5b40ed4140d214cbb2fddae12e1a3cdc71344a7d813d5e3df782ebc7c959b299cdc8ede7a7fa918b5a640ae5ef2cdce2b489f6445c00c5ee8948da2fcf181860e3f1fe0f3d5ce79ced2d183e9db4102702d81cd41f4cb73a2592260a385d392f3cae90ef124db2a0f8c7da5aa57455689bfbd6a69cf9ebbc550c36e4bc95aba83ada3ea415cd4001402ac79a72b9835e0c284f69fe5553bf34648469162921d7338d71bae7373ec9f5310c8aaf7bea3ca469610d778022ff576559ac6a66c35dac11634d138a49900ea2476c6e7173034f35042a779c6ef789df031ecfa5516f4387e89ad7c24de4b56759209ddb7d32120d84588a410032ebea529c8d2d8c1bee201e09ddd85c8720149f1875fef48f29c69bccb02aaf79bee4283cfed4d2efa5556106abe6a1a75cd1690d9d7474db8e196cf7704a5563e05c485d7745632c8d719edf3019806d301388320eb63a097d878226241c36a78fb3d022ac94fa58645357f551de21bba26daa30b974df5c7922a8a4f8cb7948769bf407c50bbded7308ae444719b30089267bbf3e197ff773f84c05a25093ccdb67bddac2097e6e8711bde4569cb4817c02663c47b5d9c60212e636cea5d24087ad80866d46aa2bff8a77ca15bb8e67b2d2c8788811e6fa421c5a4a2747bac6c656ee32367a8c071bf864375df5e62a719ece466a56dcd7c51dd4ab816c4ab06e3d5b3ef0624572af8aa6ef5aa7b28a8dcc614a4faeb3f7998afc3c72d7b0e3cebb92760484a2c36f49839df982cf2915c97013f08ca84a66e1b963726f39fe4f93ced60a0c6be64016013806577fdccc6244d69c3163ca282ebbe2df54730aba341f75a5b41e246c27dd7560080e3bda829338154a33984b2fae859220313254dbdb0b4212854af7f8505d2b2b97e51bb31f6dadd47124eaff4528db4aba8c08efef3e046042c6de03e12654ed728d0c61cb82c4cfca5329c3efba5774d1e5944d8371144aa96e6608bd36a78d8101365b312cccb1e8b4fee582e0fd2424fab1d887a587b23feb27a9e55f1d62f20fef368a6f789cb9c9f6126b8aed3ac0d6537dff0f8d1d3a7b7065fd304f01f009451234c2c67b44497a1b4f670b70b743b4a57baa148992136b7a636a21b5151c150e1aaaf47e8d94b4cd0513089b27038ea6e5829a817aa703911f2429c90f7b5f74265d22d848db0f7947fba2db042797da26b29518908a13308e36f1dbb57cd718c20c570646f0a716dd01fee71e178afd39f1319776c6b7020ccb34333d7278023a3943cd69f242e961d645c87562b753b309ee0cf4169c5af37f2c9288ac164df8ba97c28d163916a41cf433247c7c2da1f2daec6d4b6ae66d5784a96aa0970f6725d57e3a91b7f65487c645ed22627bff084c52c2197d11727fa9d1942a6826eddb08bf393d643fa09a9a1c07e53149292a1c5a1d837bc6d1a4be76c99b4800655085574769a2befdeb68fe62330fc1cf9cac0f0549ecf12c453770547fa5c1dcd4715ae87145402b96e19fada052f600f21f6a1025586f698055e1e54787ccc8d0a6801c6c7dfcc308b5dab039a51337e37eb0ffb42294e32ed34d8aeadc71307ae607518da1383ec00909f69cc8aed8b9dcc93583d62d03585e8195dc149bcbd53c54b65825fcc91a284e3c2c401575cf858d06b4bde70e162ee529ffc771f1325c6a2f5d13bccf260022e3e71324640d795abad376a3aa97edd873984c0f2dcce1fbe85ce73bfe10568a6b14a42d6066b53bae9bb4e5fb4f54b24c2c2cfaaefdca72e4e888a2c6863d11fe2caf7ccb021d5034fb78cdc659956d8d1b73d219d23d287b69b9813b74329d3c2022c26dc64c2c7298ebe026abcae4a4f66d883f1f0c73e1e6a24a703e8b04422b5869dc9be4294f72fe77a528ea74f9bbfa61241d7efb9df07e3dcfdaca28c770a5e5bdc178afe6286f48adea01dbc042f0ca3444eef3c0f0fb3a69e5cc4d74ce28f75a03412e56a60ee114e6b7ab8262b591501b7f4d96a50f84bd9b25bb9b6928ca77bc9f6e13164b68794c903b1fed2fc6f043cd3d8bcb86ec999fdd7ffc6a26072dead4f60a598e556aa2e4ef860971c5f693ae208fb4330bb6f8c6462c2aa9aefaa43c01eb83ad65ed1967caa4d3d74f66869f3ca911a063545a4e2958d7be0cfccd03403ca5b527c3385619b1124a4275d5f4f31aa5177e1821faa0b5875b6c6d7da4c7fea4de368ae9eeba980ce008c13c4e214751f6614eba4262c7eb54e535f8bdf368840f8231408afaf2dfc1aa9fb1b0389e4dc3e5704abe4da873a5a9f61213e3d15b62b69a070e2aa07e82bdf731aa2686c9b8ca536a9ca3cee34cf71407c8c0ed6964b8b758a8b204553b44e3803a446012901470ce1979b3cef9c72fcca9d208e55bed938c535e06d97f44a86dd271978ab56c2cac605034bad78f70d53cb6b25abf0bd868c38a982388b7095a0fd570bb45bcc889fae51c14a328d7bfa52383c286a36def1af05b8d65d547c6f197e52550d33d049c74a54c916b5e797df8a7da40a750daeccb0b5ba9457b9d974b1a021ddf73a0c3e5a614cd392cb19576691d09ce8b65899174e3f51068a7735e3bc2ed674b0a0518ef5b2dd6ff2dfd1b64ef595b7c6b8f02fd80df247f7489bf678f9a5f4b02242a11a2066fa275a8dcbe74e3f971038742dbcb3fa71c4f4602ec88976404140c0c480a7266b7d682ef57109143ff247dea781971cc98cdd511599bcdc60c0b099a7bae44d5b424f944d018ebcb3649cd25cdfdd33ada7ba2a1a4c4d152da65ba5fd00adad7c8c5e2fbf504ea40e8d3c34261a2e5413ef7e6bc7ad3c4f61b3264e8242ff1e06ddc43c22ac35a40a92860c195e351b0748a9996cf768ef4cf6b5ec245f6adf677a720d04fb627ee38775eb01ff3afdff5f7e91cce2259f50bb54c62236a3d89524887dae41df75f025da764715e732f3427d9e7c57718b17fab10a7dbbab10862fef5f907c7c7e832759af45eb584340a497a5b27637fedfdd19e306511e1f0e1f2ae65fb4f16cade043519db961155e9a7fc9b3b59847c656086026c195856f42b6f3b9120151143cbe5cf6b2fb926ccab9186277a65359113815836a7cd5b26725f2e527e989689c7ee6dd6e042bbe4cc0490f8f711a0ecb70b6370aa90da30d63585576b7e9ba66ae77da801db7dc7bb2035057efecd7d1c851b422965a98d568f157fde37e3b3a5b019ac216d46c57487d1e38e824eb774aa3dc47dd258ebfffb7371751b866a10992f37a7cd347e92dad244920c5fd59432317b2a92a4ea18a0a893261f8ec451c21a8b819cb34c2d8b14e2c37fcc4a50921b136cb692c86777ec59b94cd931f0fe639757cae1cd074a61e6321fabe7b26b4fe3387723b97b16e15984f88b480d0ca2fefd926e74ab74a46d40825c282966fe62d5fdbf79ac172f13d6bccfa9d1cd9dd947c43ac353948ecc81fc664b2a62e355461efdefd5afe7e5bfe7fc4bab672b856a2fe9d8f159828e391d6dda0e6278661b8b7b8a4dd432e2fc6742e1e5dc8ed3c8396a4e08e6408b665089c1a6c11a09d491724da7b69e00f6d8ac80315bcbcff239882e6c0b3b90f83e76d6fa8dd245a60869d032025b00dbc1bdd2780b1aee7aef5f9a30e6e4303c9ba80f17c8f1d19277600e024cf95aa126ae57a411428ee15367f493212c9d9d3888492e95d0bd363baae847fa46c0dc7e663e910c308f2e283c2d7c16d240a568e93efb663a7942831b027eea1b3bbfdcdd0da4593bde3898b21e258833dcd73bbfcfca197cffa06c9ae8405eae7e5a8fd9938eeec709b157932a7c2274f51f3522eebb5f3c692dd738bfce1fe8a6ff876a3c0ffb2fedab1d4cb438ab80aecce856924bb3f9aae89797e73dbc99d698a94fef06a49b6b2da42de3fa1a3b6bac092e466b472d089deb6521140546f3d9c34c639c25d9b3d419b0f25b44118605333a31d9677ca83fa19afb9492cb6c0bd76f713f20dbaf3f45da31b65cdbb9c90ed58387d8fca251935c1e2ba7a0cbacb5ae9d059c5401d2e8bb9878cb362be49ec099f037598eabb59eff57ea4977ce6f67f42868ccdb062aca33b3480ea202a22ff479af7250d9a62baef58b988c53d62295dc123db6deca252571a8954b43180e2374c9f9f67327458d53cfc5f5f2097634a225532b0d2fbf6ac9133aa056443b1ab505bafe41822361fc91b3041c8cfa7d70db0d1d719789c82cde25f07830d8e4ed8ab5afbfefe7f3c5b5cbe54a7388bbf3304b6d0f2642728327e6140e95aaaad5933951f52e6cfa9340ac113da5d269f86851f425b9d28e5c9e73982967e892bdc3f8a7caa66e3c4b7c34b4630e274b45d942b11dbcb554c03b6b3605c690f5948799b91ce542709e8a88b37a09f34596e08bf788551a4cfee00a38c873357875bc1529e3462734782ccd9eb8087983eb178ef2719a5bb6d243e2d2c3695c2a4821e30740a2e25c62d1412295f2b5c74756576b687903bae4cd0ce4c174d323d9cc5b8df79eca73781da0b8c2a0f4f8d47da57b5996c96c0e45d75204d7a0065067c689655181554c7ba01f84133395e7085a60f28f6e715ad15da6f2143bbc7003058a178f8899a9f9bc723fdfe58a944fa221a91b348ee5155a235272bcef7c286d90bf600f8a67cf08d54755cbedb6bf195bbb04d7b92747ece9d53da26b08a0c5f53d45e32ce064e641a8d4968ceded735d39bdb0918aad2c64ce7cff5e29a303469e7f08c94094c811a216504521661db379932e25b7bdbd7601d8ccb5f7e1bf3d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hdb2a4ae78915cb1c7167fff10da59f171f8891099fca23d9dab7a057cd2229040b113ee974d06d825acbd8c31bf85e5cdc458c42ee0776e1f9a9b46eac404c1799c418d77b01550d9074594c30fb435283d8681b35e0ba047a44c8766a5de817a179d209b511cd5d5ae9e5658550bd695d0f7d2b4b119d22039d157b09e0a5cedbbbdb97b34a3a1de829092269518867579edd3ace4b920a11e0fd1a45994b629c26248d1806dc9cfcc0cefcd441ac690d0051f77d7ac89be53f021d656375e476cab13456439fd045cb12221112de63d61d0255aa7bfca0b737139c0312b24d2f904aeba742c4a63f89f659963cb750dc07bc3f5c1b24605a9936e18605415c8a120aa236660661f2daf20eae72d76aa8bca9f8276b77d65b2210cc0251fe50c645ba19af52ccdcf1e4c202877f85add24c6d2845bc04de0c3f76b5d78cd97780b99a1b661fc6b0ab4b6af7fe824772bbc98e687e2fad0a04e799729b215bcfac7841d34249a971f5fb035edf6f5a4c4346e500c41bf8721d59a2c43f7926faad32156345d5e596667cad9dfe4daf4a0ce8d41f916bba013b80ec9d0d99f48f58fd393599ff08f3f170b63dbb65cfd2b2649ad461559b5d74e4ba4364543d15c30df451e484c761795097183a12b49a740b6eefd31b6f8a839fc2603fb8f7251b378a4be31fd4b9fd70a7988ab898f1ed6dd889a6f10ceb5f410020e6076e29037cff3917322157f1240fb7d21ed1653fb37f62ad7ec042dcd862d31c031f799b6ec05eee57f8a84bf8bfda64f76a2c63c25d648ac106f25a3ce2b9db33a71010d5962a0d63f0709e85d5b0617be6b35c18210b97caa696b9a440d111a8b75dc26c71c30ca1a286f0386d5f5e0a8a90d6f9b82578841d61df4929da151524d034d41893e632ff8da800679069ceac3abe21a5f40b4c1d967dd3c5e8872188d47255ecfbfcf3ae349229e0bf9a7a5a2e94b401dc5bc9e033edfa631230421f923b4588bcbf6b4544a9f50fcb8b979a00980890f66f5ed28b44772ac789be1752e9c0e855c98d0cae410a1d350a1f422fb9dc009f66026a1d37d7f1bd9f67c61379743e2b53e4907f88675fcf7dc55430a771623a31e0764263c0abc25bae262722a5411f725e3a55969602d74d2534e77ae43dc339626b0532e399b5f69ebc1712da90848691dae13b928f6ee3af5cf6d8e29aa71aa93ae58fe20b06bdfe0fd1c54ee31a6813c861538fb649a411bd458c81c6215296393965f099ba981d061a43862064364945bc5dd72f03068bb0b34fe2f173925e090d5f62603533abd1d49b3931e7d37a9496d372fb38aba8f3d6e0b97d218ecb27099851d584de1d24c214177c8262c80431a49a8f5a2dbd08af45cf9314bc8568d3e0f6fa4c9c6014fc456e592fb792daefae89a99790aefb61df50274a74fe13df0d7ebc94dc8fccc045b3ec168183215d000f82d345d7b3779405b58aae9b0d9c56dc4612338d6ee01df819a344949582c93cba904b14aeb83515b10cf6bca7ecbe9cc7d38ba5e9b9001dfc870a105479847aeac4cdcfb1730e59b229cbd1df9dac4e20d7917ecbed50a2260b3458bc18a30e478433d2b764c276f59547df6ba363e9fd51cf4f3dedc759472d1ee12ecb19c8580c72fee7b7255e8019f2d58ca152104bfec1cb4e49ed0f4d9e7c4f16a6915729ea264201fdca9e5fd19f1dcb1f763eee3e72dadc9a9aa49b570ef6d97e77145ca86cc6635a35dbdafa48d8deb83da23020d0ca00135c00e11a5c6d64a77bb3e1de5f2915c6a22fe2f95d052dcc7c352ed70ecfcd851f756da3a3a86a3500b27a3be3f215ba9fc949831c1cddd33f7d6bf50cd064a4117a6857aeb018f87599bc02c59c089f559c843d0f6058ad278451d1f06a8e19e83fe8a3317cee00822766f0dacba3dcde0cdf285077bf2eca9c7b5b305b32cbd3dd2016c350af5366ff3043a137ac05dfbc5e1db933d475f0e3c2bfa1abacf9bd05113378ee8a03dcbd39dff5f532cab3e4ae12638313f1a7f2d8578eea9f601a2c2467f2a3a0ddecd03b09e4d71f4b742d4709a4324e359e8f1be3c4237f49bf20dbfad7c7d978b51cd72c7cb67a5b4bdfd4f09d9737d0bd520dbe49c88925f4b045149bcd322b498350cbffdcb1b7535760e3c602963d58482a945d1c7d828ec5fd8ec00990c5cc3dc44d22b19fe2cbc8a0786f3bf237171b5e3a62c631718cc566b4339b3435af210811900989f74d0800a7b45fd65e83b2eeeb0ef6b7f434c2465c83574a62ba2f58e299871e321ace247f8463ac17f3580faf13d1ad8262a46f22cbc5282648fc90e9d42b6f8ab04801129ac299f7f12b702fd285a33ac76534dd5a6618137a644c839ca51c73b17ab8029dae71395d9ccab5f400141545a70df1a3ee2f27eb5929de4f1b16de492c2c921ef9bc95e65315c334b322852e4636f713a43d45dff952bf4a150c67994be8388ca7738c2ad2a648820ffdaa2ea324388681bdec17d34965ffe03969d8c8cff63d8ee7fbdd8f61bf111a502c32b99e96cf6e1b36e69220233d48db45b2406e0b7a0de0f6d53a12b65e94fbd0be064dfc2eca8d0993ac1a7dd76f20a51b60cd93d6a303700278afbe982a187e83f1e3553c69798f89060a6e1e00317b02b01c5b02ecc60a72ce8837dfb8429c3268b5a1eec01c23cb146e559ebc04a2deff57ec3af7e2326714d4c1a078a70ae4c04937b91920ef50e3a546894b33992adbfe20fbec1676ab8b7f4459ed71bb6e59f67cf4b10d51500bf6a56e9c0abd3086f0ca8b20b7b0f7054af5ce01ecb51ca5fc76704f19fdec2b22869c6434d0c7e81cb9af52c351ddd15e665e9d87678d00386d25f37393248edbb98f5f6967818e6c11b3d91f181bc0ca17ff91a63532d9c830f6d786ebb86a81feb3177d193c87d0eac5381c46bcdc6e35a22ba5da1162287f19c94e54b29cbab9670ce24d983514ab8104d2f59e166f79ae4a8427b562ff924aa291280863e8895e498eeb7eba27c53633291c832429129e16d50a7f647a61044eb2e26d2ab953d90e8bf39b099df9052eb39a7b4fc1b9d5428979ed430b563d3c383e39ced650c6381d13c5c920060f8f765eae8cc97f87b0f8453bed7a1aaef9a79e4e084857d76eba22e061b01e113a753762648c2948497c2d8c68fd171f3535528c06cdc7a1b9068c4d61769238a6ee09976a31912d694b5648807c0b33ba1e5766053b8306993556a4f28a39fba9e6c5460e0b556c777634aad9117ac73e6b5c7adaaae1e06287e05c44729d632ab90853b41ec2d1613f7d6381d1b402c32ea847b0162397fa2e148d2ebec5de5a68679e5f09c5930a6c871c36f31d280f15c5d67e933f96750f0f50ced0accc759dbb9a2bafcba75be04eb5560f69f95608ac3cfc9906fcca8efeff09a6ff88afd7d553f1da434a4157513308c222270086f36611988283770460afc3d17ed479088d6738e6b8c53efc5f379560ea42fc788d8edceec6445869df0852692adac1b6ac8df71892b41b8f7e6ffcde5b4275be78259aaed2f5c6fbdbb1036bd6454bad2564b91a7e08d75917392a5cb9cd0f6c5683314429a1240976e78633ae8ee26ea5f09c2643dc334cd33c6455df45104783c124d0e16bcc65e1f325ca587780b6381708d529a616fa3ec631d303a6220be5557ea0b39acf0e24c7df2fdc12f80c7d37a82526f5425827693c35553cc55406bbae5cd42c1984baf29383afb00c96082f2296ec98dd204499b55857b756f14a2a56610e957e1603b1d9d8eff413ae4942a25ff6bedb93a92f3d64a3f83a386fef7bfb99bb609d0b94ac17026645dc2fb3635d44afcca6dee11612b957941aa9d629c8712c62628a161c973c240748fb076c5f1c6c60f4d66f84cf9ef9266b1118e9c9a323c71ba89eef048be5e9740b71b3011b67781c07ea3037e2e5203f8f7214f003d20877bfdb38ce43e07b9f6dc77e703ef61680ab2cf142d8c9ad003d6dad6dcdce2a42ef4a9480931650c2e829b5bf86c1e5c369f48ba813f7837e28326c7d0105e015b6b9e3626c965b228dad043e27cfab9f2b453bb6eb13b60b4113979e82183635f5b2e6f98fdaed3de9c298943dca94edc0ce06fdbf4631a325cd7dfaa8a1566ac96a84196841f43bb6a71a14344d272b234e6d365e9407f96d3cc869e5ace4815923b3dd241afafcbee61d28e9330ed75f3aa8eea1a13a94b49ffe764fdf2838c9678fedbaa003e711498f9b4134e33c9ac53e6e3d1db01db21de785f86db7d3c56ac29bc0b3b72f4c54f665b5dfbdcd98ebdcd01b11fe6ad7b02463ab42e535815ad3c654a5df401afcbcdb4129c86e32f8359c4066157ccdcc626b05246c6abcd2999a9f51f280bce3dc20dcff39b9fe49a521d81efa61f4c4a5e2809356d37a10ee26d62bdc5f7a0197fe4ac187dd30403eb219cdcf92a1f65fd7fd5e448b7bfa424b10df3f38d0fed16b3ef795fe41e22b5450f66358f28a9417d84ec98ac2e3af6ab1e9b404db1870a6ca70bf5a53e1ef99cc79c1768310c38b0863e4a5fd2e13252af7d8f66d116f008d5617254ec4165f1e0d163436f6470e99a241a9f7f781aac1a1e66c6fbbc0fac2de494a581a22fd3ce4a2eea1d0750aba24e7dccc044f0dc5d7d0d53bae79cf0538815eeea16a83ed69e098d954207bfa3e3845a955617d3d63dc0327d78cee937878b82ce4a99be610f50d63b1ccbfa263a84907d32d2be76a46a2671c0707eda9e2385ace1645c77800b8e5d7e1a9c2c189b9b4b96bf1931ed3fce2a760c0ec105c3ca10782258a8ed44f21befb6bed4bf6f501df26cb07f8638eb42f6364095fd9a3cafd21095d9e788ef54188e4dbad2f452f1bc4f9478af5a936381812531566e320c847216b4aa7f9a1a50424daebfc26c606d4d63471ac56bcae2be6f0f91811354d64067be9313eaa7c8d12aca31b9dd2319a9229dc4a544410f3eb94bff2a40c4f0bd315b23ba1b5a06a04c060dc5e3365723def23017463a9aae8b067a92677dc188f9e9d495c8e171839c65814a8fdd5e98c51f12a1e6d330171f9dffc43ffc4de7c4b9f19d9ea230fcc664481cbcd3c30c097cd63191d7f884d3305af805e53c596881a36965e03357eb14ae191191b8cca54980f897b222591bc2fcd85ae1aa553582875fde289dc3f7020a01a951de98c9d24fa7f860f0f7289d8269cbcbdb1a9595caa012f5e8fe413c6dc94a3c47f3c28859870047869117385cb086f86422f5287e693030f13333611dbae63ec1b5beb51b6578d493e65ad41522d8107bcf0f2ff0ba417f98be62f18d7521161e565fd802f654e9dc69a5b3e1ce1415c4c9bc4dc87e166fb00586661dbafc6a057c5fea267f28df9b3e4f5c84905f281d104d0ba6c74b2e3c92ae3680f0548ae495962d57ba892c8aba93220d0d93afd4842ea9e4cd1b3da34f6d4e4394bc1b6b7bf9da86b3e02956647e7e628e8293872f5990fe8d0ce928ee08ccd5c61e1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h5e8a9eb0c00a75d956be10d8ca1e5017b93faa32a5c47937b8634a3e6ea92876a3f023c90f3155a07f9233c8a2f9dccb511e7dcf32ad6ac25e9686b3f4c74993ba3fdb60fd9f02c97f826ce81eb134372fce3e408553116c87f15c541d6ad759917bbb8df32bf4d1ea63921cef5bbd6dcbddc37f37d77b8e92c0195bd14f46acbd7f7c74ac9755d8df90adbff37a7b4aebe8a4e35b6bc43cd6132c4042f1639ac1991330870ee0fb16d809da6887ae6269257a870f1b5e983522b20d998be124c95fdce63858c8ed08028ea6c84818a69af823e1c692803dcd04f3cef92108643ec77496c11c826fdb7f542312e1b5250dfd8078167b6fd6d0e1257000c65854274723735fe0f84c97d93ec51b86e75f46a6b3ed140b7a489ea465e490898d82c69965c5af2993bc68e2fceb527ab4b0f7c89bb894194773ec735e9fb2c0b3402a95534b55f8a60474f050a27007fb398f762e663e3c269b75d336c1c7b0c81c8a3cd1e8a0585f7c94888b4e022e9fb744628c6bde027456a474493c13efc7a9a5b6dc19f656d11b578e1a937744af368f31baaad69379585a9af232d6adb0d2fd0a0d82c8cb3f9ac12cbe9a4eb3e2d4a927e6a051e9d0ec3f4415ec539ae7150aaf2ec09a3ccb372f522b157910ff643b989e84fd79e6ed57a6208d18e1559df9cd31ae23b5b98ae8ebc365aeff622dd5fa06ffad326188e443ce51886c09f52ee8dd4deb7e3d6121701f6392b62791835cbe5eb51b6d26fc7300c7118d712d80d4573e340d838ab5455edf8430ed9ba7b438eae29619f6002c6dbbf3f444cab581b0b56671d8ec40c227cfada650de88060aa8f9a620fda74ef677590512dc451bf38cc53b4f9163b59ec5b1b73540a12c6da41f4c2b6d2666237e542bef5cecd7da6b825e1a97ad3f63266c634b5e67d974438a3e58594e6e779cbc0900c8a08a4b39d4d80a7b8f4a7d35ebe5e21ab5da4df1b614405c02284085cbe0667988172ca940dc09f9fb3a9d0b4d3b374a3d2d889b462a2911ad07353f28292f5eaf77a8681ceb2ba7442f8e11c9aa9eab247448b91c60dc5186d1b49c06ceb5456f4f8795a304fddc0016787dd852e502623743feef2b297bdbab1bad85211def7bbc658717748083f545e9bd6cfcdc17a5e9adba83caf3d379f74583c31d515320cdd7461ae0465c5ba3333d2ab14c341163d2289ce11499c227a63570a2439c18e45bd2b6c9dd7003ec0d795735ed41247e3acb9a738d79af4b23f4e72e10523ba8ebea426deef12e93dfbf0fe91cfe78750584f55767075db81f494bfec1c1900085616108c86114bea2173074cc1701b01452cafc341d224373169ccaec9a6420ad234dc0e778fc6a76825d526791cddf8ebc06932825829df222fc53735d95aada4b9c1392a821bc58ce8e011a981320e4406316f3895959ea4083d162ac1c7e347f64b22cea022d846132169e6b34b5e95924d6c55a7f9d86d3224d0abe270a0da5769c579cad731b182e32276b48e8351e73ca94846b9f00eda4c4750ce5ac9f7d5196c31369d029ce3cd0b334c7e573c625f7a84f7ca4c6a90f2119206b07afc21aee71c1f78e699db50bcb9f7a9224ba0c969ead8f3d8fd2f8172587588da81ffcbd7fab7a8a1cc8e542495b2e37e1b3481160b3bfaa59a72c604487d695405e91093664831fce319f7d5c02de583bf309682f5924126d141b0d97c93ed80434355e710a0260db28b087ad6fe11291e8b5d68565b027f893728e836ba656caf591905fc7b2f8906d487f21e30e50e3998817f5f3d6907f64dbbf3c30069c38a9498f3a1ca645d6972d518f290715e79197a0b7ced24e8d6e75e281c352ab0d2b30b31e9d8dcd35f240fcac0db741a0ddc816b1ffb05c15c917e02282d1aea1ad8326ef62a95cf3be4308a858aec328b789eb08bb1f87a1b1b3e3d4f1c4de51c0a334fbcc9d0dc0d86f351cd6eee46eca5d95187865769287dcd34629e2f91c9a55eb2d3960bdb7b355bf0155b734c0a8826cd4a303256ba9316f06ffd371a4445be901ebada951c983ddc1b9155499bc4096fd150fec8668c889777db48905320909cd8c0cdb57170c345c683a0128cbeee3ccb09068e91f3bdcf213a6adf0a63a952adb9cc7c5d070b4cc3d5145020e908f4b99d421ad9d2d805d41f5e439bc257ae8df9c66c900e946e58e9a54c9f9acf9b7b77d889d2cf3e401cb3d019c6034d7f47a2dd1a231e0061b7cfbcaa888a5a9f39a4d9d0c94be6a5d8d04adc25bc4ab8e0bdd094ce0dc548d33a9cb41cfd956349de4b2b23a5df83d254d92b575d6d2925c08f5234b4a5172ea8a085323eb38dd5d2bcd852b46cab58bd7045442bf88367f198acda53e05f29fd39718840265d358faa458d4c07e9cee9938758db7fb0d0c764369da96b5da0cb6c1f28f7d3965cf7dae36af90a73d537569f11388b5e9c734bd439e6356bf9393af66997011c4aa7f047644a70f34f750aa2d6b575f2a16ac3dc4e63f79b2ed8d3b39ca19f8ac2a7baf680df6ed810ed51f336994eee00e70e17daefbd7271fc346da8554b9c9fead127ef71e6fa293c7535cbbe1315426120a73f71895fbb02068d0026050369512ea6981798a1acae9ee60be2ab63e0f254ce33813f0b50b6c71e7681c364cd2e514e8aeeb874f66cbfdbf47f17172262c50e93255e7a174e2ac4d1496a75268e455275cfaf130c0af287f3b56706cb64e0ced0555f4f8dd63a8c5221ab774e4c03e7544ccf82273383cb64bc26a8d3464a3a4743533d11aba5bb439f3694e266909e947dd685352de83edbffbe583fa73719de97fff23cdae60f99e48c002d1a606b76abe40d76bdceb3bf1b910377f11759fd588f783c2ecdf231de5b0153399ea90deb4db335d61810a81e122cbb6ab65a58857c11f8bea83dc5ba9c07bcedee68341ffdac54737f7d6696bd90fed2c3ca05409823d1b7b59a33cb9741c76a9607afb3778a115d639ca655eef549ffdbcada6eedc95944ff2493e2e644c7fb7113e8993b8596f19d49473922bd66615ae1a9f51c598efc073c6f41f0f8f4c89d24bd9fe881ef3f4b7a35ebf59bca21a45cbab94c43cc8257ce22668b19f9c9d1906f956dd7c19af0d41ebd9079fc1641f727998d7bb81fe7f4cafe8c8af2e19cf21c8c13a940ce29216832d0d0f1af8191d6839e9a26ff2c5552f752d0c65de212e3e41809c0ed7bc695100e39409ede6614a018cfdeb2d71f494396dd60dd253dadedfd49aef985216240dd32479375e1c50d4ffc25cf5e18b25784cd7ac806813352437e7a45481bfa125acd94605420769489ee93f34a2ec585b1cbedd428448c7506524a04a2f65c61b6b6c3c2fa9eb489e493d58e9a5487f533852dacd66d5c546e59d94830c01ed81751577a6415f566c733e4df9d10801c04469c010843cdd2c2f7f96dae06d5e72c67069181987dff7f21c86e46888fbd59ed85d07b52e77c9946dcee0647f9fd754dfb2ea639b64cfebab89e09ba34ddc1a280e135dd59f98767b2242a8eeafbae152e10c09867f97b32bf81c2b4644c1c4bae92b9ca03ce4c714ce1d50d17181459cdf0c040cf43d3e081c3949e8572131bbe283870307e0367bcb20f68a654d49cc539777fd6075a3770e4c3b14bd3932fd571408c5d497e840fe640338355fb6587d78e8c260e6deed853f981e51aadff07ffcd6210c3543cfda8c6e7c1a407fef64eacb27f2a05f207fe95796d6d7278a245446f1547a7553ec3102bb6bc12f227feac9afa1ad9342914e03ad91888a41c531cf1d8b5639e27e902fed02ba798624551ea03c37d362083d97ffc31d867a9819cbf3c5c6c3f0c5fe0f1defb210c1fe4beca9fb5f05274a21a9d0032413010e2f56344a3f71f09d0f13e142530724dad59f6981fcc0dc140d0b443343845b372a2ad626da15b0ea1245ff3627e22d4b6d3cca20ce197e9479d7dd09c014d938c3a39bfaea352bcd1cd6e09947275054f932fb0800d4b4c094d5c1ddf0948e88a1f162a8aceed21e8d308d91cb505b617fc22f9a4a14f64fe1b7764ffd0f966d5f303f64ccc53b30ae2f872c1bac0d54c55a3de3547e47a55ae845c10d402d094e8dccd218abe94f7d225c11d5ae843d1d8d34aeff3dfb689d79b66c83747ae2d45518b30e2c387a4915f43bea954d37c09dadd474af45eeca6f0092a181052b9614146b42e2c33491c7fc59f59b93639e0feb13795e036fd0b2096dece0c4aef1a5460c7994b1ec973bab78298b4f6c8cadc880bdbfae35943e1fec22adf02c70670951dd97daef71553b8617ad8216bf0fde596b72ea6c6efccab83c3531f17ccf360c9e3b126f73bc0a0b74768ce02e4cb7e4976d44419d8fb1d0672e57ed215adf3cb520927d6a9c4b26a3a00a5ea571922ce4b1b7221a09cee60fdc94a94cf79331bc71308c284dc84af5897423b0cb80a33c0fce1e84ea6344e2cc29b1282b0c148cfda261192084b417f6fd41c4f5af9c4720a4e8e22c2f4b9b8a912c4964ef9efabddd3a8e6b576f28c2a2b87f755378e3a60bec4a3ba59aaf3ea971c4ee1bfe4da39f7f308e8e5b4dd2eb66a372f76f6185ca5b4d00cf467fc054084e7c5c7c80a8ba9adeacde4089fc2f1e98f0c4f93e5201026674e9f8dcc37ec8c218c8ddf97c1dde92ea71f950e6c2f066dd2c6f9197a590da6e20ca72852c8901e4ffb2f3231cbdf68caa0ea0df2940c082f71a446ea480dfc6c2b06ebad3c6cc938a9e0a071bb0f2c7aa3ddb0fab6ffe6f494f6aa3e56ab5c45e7597dd2cd1edf743f178626e5eb0ab5dc4f13d05cacb83f79df2c15013baa0f953304d6e9afcf4dfb86099325ccdf9fb9ac1e679180d6e8b2aa92699653105341d9849fbc8fe595c032df8d847ce99384d85dd856b5f441c1fc00a8b89f682afc17c535d6b4e4ac7deabd694ad9bad354c67b554bf3aabf21b1e3049f6009546deb7ac7c01e9d19949efb625ff09fcbb70a2d3e6f27472f0c40d33503e608938e69584f655d739baad5b147435cc8f020b7e78226fd02169cc095cac0f2b1e4794c0ba942fbc94fe2623007f9b7b0f0730239e955138a5436d207bbd967ac13c4206f7bb4a10e966fab75f9f3cebb1d7de743b2fde0ab9384ff581e79991e7d32a4c1facd2352377eee13f93c1eb70ee31d47321a750288d7e15442f4f142ff44d2263ff27cc2a591077996bf5306ef8114be89153e4a376463bc8863ccfaf7ebaf8692361475736c1065a0846f2a26a17e9a833547208d8169d8d26b865367f614b2e2ca6e45d016f2b4c2f2fc7ea837f6c614832d2da519563adc253fd27ce508e3443f62996873d2f42393ed9a5b265442d35f50b00e85766dbfcc34b75e8404fb9a907bc1f810c527dad749b9f8777cdd72dce05fb3f6c2abff0a3d55654fc0444799efce62711c0cb738708d49ccd14d6b4a8317f66071bf892be68540debe278bd5c90755ae8576fd4a41d6217ca74cf483b92ca44829c3a5dcf;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'ha4cd272aa602e8d25833043f4d9b14e93bdbb62e49fcd17edd905888d5caad2186c10c0ed215ca18a55b60d086cdc2e995ae9b63f6ea87331a809e33203b1cd6e8c9943dfb4b3e4b615c7d1c24f304673119d4b14d7bbc5c8f692c8ee1acbd0ebe52f4764fbd8d638dd67a45daff5453f2d0f4128357b79e7c4e3b03eab1398ef7824c9a10a83c1829a08d38f8ed7bd90f8fe05d77b5040cac0e13e4dfb1650f658447fe144e1f24a87c90c58bcd78743e91bd8f5c83b029bea904bbc70632144b36b2b4a7543bc2859e1112c2d8d63212370f3a7cb849052983cf06bc06d7d4f5f4da3ef79b0ead67721737da0000158897576420e2daf9dddb299dd06aedafa159c03df28c6ef92ed08482e6065b9fcdf1f634bae6de443b878d76b316a2025ec7e5e590f8457db70c0722d4ab9d73ef7a9949c54799479fade7ae388f86496e721acf1020fa9e19b19481bb8b535f851f54f17807c66b977f06b0a130611a8bad91a00d3db94ee1494a62fc2993e160902676ff2a8bdbf6de08c5882cf036525146bc326acaa0acfaac4cb0ebbf0870088aa4a334cdac04b92e56212a0d765921aae178fc6e973b14fb84eea503bc70750412f1bb0a78578c7b464f81cf775e1be341b0f611243deedb3c2449b5934333e38a45abb383a267c34cae6c4a1b788c4b6d15de1c13aea01c3e51bc773bde33e9a559eaa9d2673f3b0dc2dba48e4fc077078661e84635d6919d7d55b238bf7df75105080ed4c5e2a6bb22467bbd1d80e49d92d0f95006535db3b49aceaada9598694fdea4ba38d795d16b7889ea940809c7e509d919615b463f1448e45cb08caf555a6109e6c358ea0968128e8eeae6835c43dad0e08601551ede1cd572e6b6b4299681e0776a05b02037acaee4176a352abf3649d2a9e9789db0cdf3e7b6fa95ad54c65d86dc31d79d123bc0ee69abd4d17b0fd2855e2988c747ded032f3dc5c31e19f396f513cc400a235bfc26fdb795f1fcf5255506fb06d9bf0aad4123e3fe1b297947f10aa8d4722f136a7afa406185ef726cf6826d025b36c4b72e2f66661dc4e3a49828494805904b4f308c06e1bcbe123b75eb19f8543d5a7a1602fe9d386085b25bb00783297c73181d17f4b1f0bc594518d210f00442ed50b073713dc94bd65bc1185eb1634453aa3e3e695fb70cd5d6b3835349620d545992d52421b546852a7659443589c1e63adc785cc48a04f092043a4d11c3f741956f4b7158bdbe6e894c75affb98d89d6809fa292297d8ef999c64d4211e119d3cebcd9d1a22bbdcdc32b684758f4c6c967d12ad6c7f971cb52ad678545692c1a3096c35fd9e4cd27abe41cbcb97b8d52a047aad30fac2218907d74d36f707205af50957673303fd33778961999913195b7e32796d1cdab4eef83c28e0bb26f649c194217ddf19f50336ac29244971997de55566b072bba304a8e11e2c9fad09e0cc20fb044ab2b0b99faf92351f4ea21a6567636c150a44050c4e3ffb6f58f55895e7d25e35425281175d35e5bb382ca7a20be7eaca2bd7b18a513282f50374afda633977d7e4ecd82212a244b81f2751b49c72df38b998c06483be15db30aec0aa03b30cbef814110c0112ea5086b2b3b4c8e9301145611dccdc714bc271f0a056d9295c95103048ee7c8420a31dba602179c0e47956559ce3bcf54af4a5e04871e94401b9fcd2f20a2772cfc70e2dd488a05a1eb4456822d44daf0e3feb0dd4ff0739d6598aca1676ff52e3eba9ed304617532200021bb10da54cd75c757e0855a8094e1080e3f45f3714fccf096e3f8b2a8b11768e12276c8f23824fd0a24a80d6b94e2a76405cad5d3274b00cf5ed1a845a4c2599d8445ce254a2147adaf53b2b2a617dc212b91a7df4e1e5236ba004c661de5371c2926b5d82c3dbd1f39ad078ab4f2f16f672515991254b75c4598c45c4bcb3449982e4af0ace9c3de5554c347a2b3156a57e5edc124574d045ab0be68a5387795e18340de49ad69873d94c54188bc3ce7d1b6f658a1ee1170af5685395ea6e73b6f6cb4a27b80f795bd966e770e8227d513b1cb71bb668a5100cbcb9a93749294c862421d18a3104f36207bfc550c20a0382355b5a432820c1845e84cd074947b99407313911333d82d9bc0d725a920007d0db7fa6055f94f40c4a669dfd1c31d831610772c883ca1dcd146e2d464d3de25361b505afebfa6d90401fa175a68325a9cb281e757cdea5c773cc098e3f3bc33400a01abb5d99d81890bea7e3526e34ca081f880d5f39ae4e71aed7db6b83845f07f11aa63a68f36edddbb948640f1a330b9cb30b58799bc84e75f805102c22d061ba3e996d09feee82a49e41b44d8a286559ee166630d8c01e880da5799826620603d55fe6f8ca0b3edc6c66cc7b4f680a5585140e4110fe9d5b973a25c1ef1dd37c81783f15cb6abf06576da70628c6cd4c45f82615c2edc085b24759a46bd7ef2fa47138b8b0fce190a055f1cf59aed26e5ded697a878a7b036a3dddc2dec263caf8cd855e560eee548da8287812dda357a1828c5c63f035141d2c4f92ceb70dd19dbcbe55262a179042372bf182eaff296219c10752435b2e444ef2ea2e47fac7a429afe71971e71a22f796e0e6fba32eac199a2c33a1ec44dfa2976117f37ec719fd6cbbd26a5f0c7c45807ae3a92d6f0e68f6966e645d583aaf385092f30a4e7e31bd04fd32239d18a9382c11b8173db909d4d111f0bc095a43e62ddc391f0ba8b87f0e0ea02cb9741afee1f150ed722ab3bbd3d8f2552c41fed633afd58ae32b13fe176da37d36314b492948701a8f2a04749a9329a488c37081f3784f6b26250979c111f9babbc6decb47b300ff79f92d9330ae2ff31256d212118ac371835b28bdbae4f8d3c462cf63aff00adf4883179deeab2e80efe1827074ff2ba8885a264a4fc9976838682f19b21d17ee56da3ca42fe9e9f00e1332030da42084b58dbcffe20640d20366fa738a764457fd17d840098066b9d872d0a252f4785668c4c24d7d923875f39432d342d8bcf437b14cb37b180f3daf0cd9e58caed0b2ecc6a55611af362de9c66200fe08909823f3d75c8083fb320d035d571ca1caf38c3aeebb5afeb30470dd401bf252ead329cbc27caa4be4d8df869db06d066a23afaed4184cba6af2439ca4b1315fa675d8a9783382d06fc4907b3a8a747aeb3b4defb54555d9f4578982bffec3a3d544abb87ea9a0c25f9ed2e089bbbb7beec30432980bb97d25d587c65db19fdcc1844f52ee1007d208fe5a1050f2c6378b50aabc9b5ad36fc7b8211c7ac2c202ae38ff13ac00aecb70c36629c4037870f8d445ccf59a4d1312044569980f4bf17a20b65d7d1cbcbeae464a028e206818ad477f56e9bfeb177c2eafd427532c626c7eb7fc2d4ae79e1f2da85902baafd3facaaf78c2de9d569dce6c53d4a0f858f1f962c2c6b41d79fd38a05d79a8922b4d8cbdd31fdd2500caa20683c819bd1bef5ca95e8d4929d2cb5a516567dbce5b0604e2752e285ea984b4180adec30305e21a07a3504dc3024107767b5d235d1dab0ad57efd8fc3e2585cda9ca823626b9348c216d5226a9263cde1bcc4d084cbc97ca360acb4ab8a6c5f0b5d1a0fc65b8ffb8ff3b636e6cc1025b416d76b76499faa745877f054c240becdcc7a7e3a632a0c3e09f5a35fc4282c9ff79cc774bf328828f4f7d61e779fd94ff25544fe1dcfe54534f9c46edcd7e74dd32df36992d08e8da887e5b15e83c5a988db13a12a0138660bac8a9f2b21e86d26bb3c1bd0030a8d3f65ba90cbdc342b9abe3ddc19339c992c57dde9e5a8643f5893da1167d49a228bd868a16661242d9ae38c9bb22ca1b1266ac3b0bb590effd9e2a1308328628c4edd204c69c7027bbc30028ffcd4ed8698444dc3cd1772cbe4786e146a5c3a92998fd8a17aa0d30c75b59f9b04808458171101cc2a37f9aa808d3ee3a64747254f4ebc1022433dedb80fa95594c868305a9af1a34e4356b176d6a777fdeb08b0c96bcda4a69a41e4a37935a98fa4a837be4a92f54a0d855cf8d381d3625b4513d0505b8f47fb9ae100a80776ac98a80edaba0ea788984502712ff89c46157a5cd23c9d33fc27f65981d53adb043cfc6ec76c29c46ab068933da8bcf70e7d5094c02f8a0f545e6a665b00af63cf96fc60355e6b3539347f8885cda3c53f8d5591a9bff660811d9ab313ec09f9b27a7001c0be1dbd0a25776891ea55fe669a2c45d08d2e82bdd9cbd859e16d8e05177c9aac1c1ab2a4dc290bbdd4026c40960c3fcfb76ba54630851369d292e2d07df5103913fa05f22b0bde53ad4a660645fe93c7ffd522fb8745e708b5e0580bf257e2a2e29b3968817b9a35ddb8de2effbeb39b2676ad6c037d0a6762e4c900302fae73a8465a60fdd93fcdb46ee70797ca9e9a74e347b428df4ec5aaef82c9a479392ba0b7b451a3ebbfe8258a1108ad4e4e235168016b2fb3cb9ca9605dea121da79746de58bbfb3ccabe8363b39f76030be83e76f48a5910f19160213a713f9dddb2c7b60467051ef0a3f275de1e128f608a4bb4e2e023f17f687069a041027714d5efda6e2d10ccafda698886c3cb82ae294de6637815f77ffc70e41ab69b8f3968bbc705a01063230da6a4c40483d4fbfca3060f7c1f58ab5eaf4428a7414b7be031ef91b669c67573e669178595894d61eb6b95e73569e9652d3edd7091cd3ead97905142a0270c03570d94bd08866c01ca86f7bba168c151dc36a1ef7373e583e759ec74f4165b45b9668774fb730975d8c2f8c2c1757175c8b759c0a8712d48bbf5a14de54f17a307387cdb036c9b868222f3faf04ae73492c89b389e9ab02823eeabbf4f9a93678de8730a2501778048c10ba0cab82bd736a15c83a634d58f3368438d53641048f62c8840aabc4195f04af828f699323f2e4ae7b630dcf81962bef940d8e9b2fc42ccb4077493485e1d4c5624ce3dea551568006ffd74650ae37d856e2ef3f4351f11e4960cc86a8ad67d69501c9f24423db62de5606c0306ead44a2c0963e9845cfc861f80eb8a3f57824b856498f1a567f78494a33ca140cfaffe83ab492547fa21925177a952708fbcb55aaab9d2130d940409cd540e3d1b77b88fe2575ab5f574a1e0060594b4534aa3b337dd32398f84755181c5c107019480fec59d3258b757fd94deb1f6b6482e0d1b3b5088296bf222c42ced232608d9215c4e012e940da59bf2066151743c4f95af40bedd6b94121b6ae4884ba4cf5d79a3064bb42c19d6eb49d31a9a96b87220847d495ec9f0f23a050db81a29096b9737e858390b86644d383778d366791cdea7871baa80e75fce06b33d633f26feefd98eb4d7391fe2222f5bfc826efde85a7f514b8beff32c3b0b7900a387b8142f428f184de259cb61bd410bfe778b388bbc6aaf72f3fdbc000f6c0b24fa4811d6f18cd3b48f01d681a50d6212579de492520167fe7ba2163ba14c7a11f7832b67d4938;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'ha7620c64d9880cd9e9d26946d3dbbe3090806b97e027b3747ac17c6db98c8e501435d3aebf750bdd4acc8b0588b915b84175e7509987afb652d51e122317c8b864f9284a0f19eef13dc49dd688f664e10929f65651ef78469d9b5d1dd2dbfc672b88b7cb42042ac3c8cac148dd60fd9cf26f390abde6ea163ab515b59212a7d5137a74cb537076b547f1cfcf2b6f7577c766757604e7abecb9aba5ee5c78c7920c7279f559fff025e3b6d6c0cc55b9d6a0123e53d15bcb621ca85386f2c88f62d928fbbd27d5b375cf76558c8766c7177dcf58b61b1e5449a7f2aa5f9da6f81402dbe341be244cb5fa8f66177a6a73251525f30a15436288d5ad0e7e351cf1de50be016fdb4e6a7b0a4fa0be64defbc6dbc7b03cbf471c0429c7e698e7ab5a5018abb0a33950f3cc7a8d94d5aa31bc218adfb5504cbf4b8e428bc681589bd7f3f50c8f64bfc6ccf33d915b552a0de805f333fc98e20a9f9b8e4ce8011db46c4a5c1c3ac67dadf5c34ebf385e39b76c6a14cc23bb9abc0be702d9f707df6b0d3074cfa35e27f86e47b80036e75fdf35d946771f7cca298527cc72409a8167d25674df8f6261a3984b2c37d4a53951790c60f546663a9105a73de0cc6542d9010493ed151a0159413693ca3eea9d0823d93e12b30595aedc6e6a1b78e3ccf161c41e7e1da5f23176fff4cf2766d9131962e0cb5ec24d92d694601fc658c7a28108e8adbc89f76c2b2313f05e387f36a5008850bb621ac282aee14a3af9a8f3bebff5c2a609c9b0b6a875e3623c833b5a44826bc5da6c55b7182aa30308d21275e532967753953fbbd238a22e3b561789c1f170269b7059f662fec307c4935077a8b6d28e04365aeeee4300b596f0faa5683246d51e3356f37e997005801ffaeb04812556257928a7f47c96c4df5b898a9924071c4eabb77ce5a54e7681b3bf167dc23b3c52385be44e26f1745e20095ccc36a4ed72d088ec34ee9dd7d41fe1945ad4a4136288ba94b89ddd01be3ed531804d48ef937c110c85b1e18ed6cd13f6418bac9b6edf2ee81753f295ba67404cfa925dbce3d62251a569127d692a3723f5d8e22b9813f7b81fcded3576cf5582d1bad07662d59013eb077baa09aae4a4688f3049509113d06566817b5c0981d5a6ab3d384e26aa0fcbd712866253118144fab2d5eb7d521c3f17adb215cde589ae74831bb677dd7ca3aff9715d365fdbc114c9d4c51065aa9c8844bfdd21887df98f09570ff918df2d66d1edf53b0ff292655be45114fd2896c200e19ab1fe14268c85dffcbbe0a326cf3e3fdb358f6d43454b471fd1667f7ea33c2f4d4f8656079a0863897bcefa8289ee37f223561063323193181709d8e0a12aa9601d13df1fe1da44aa7393d72591659f7568fdad51ce8714ad6dc2e141bebb2c6a11bbb6050f0083b5d57c17c2d8f73a649e7e7f9eebb2af347948c8e487977769cd137d03900c202cb77cdba84c0e60546f3d0d53dbe9b5648050d7e330e71c62cf9005da111cba7d197b04c7c74c97d5850b6f10d32a9521901f91bfc88d825272d6bddbca1ef84917db53af26f1e5b2d8038a127ae6a782f9b284cb423502a97f1e2ec634e820ff1188557d4513ad28ec947b50ac48a75fc482f6815b4bffc29696b386c37328c5ec3d1eec2fb3495381902c0e1f377f1e40224fe947db83da4271749648e89a9f21a4a01300b47d82acc07e8419aee3d783716ac36457e9424addf1067def48909f8e59aa06dfeae1a2010f93d9b951139cd03bf20928243a16ad2e47219293254432c6979681d3c2e96454efbb542873be42c8d55a8c1d3707d8e63674ecee4bb6bbe5374662fb86fbf53fced8e3d872b0cf539c0ebe2d0af33c3d88fb4e09b83cd49446d22d91d2ab191b2e9a9f230c99711b4a7bc463227bb9df22e20a404f7674868562f657f4f3d8b390510b7f5d3d88412cc6bd7164423f31fd636b6c77a9b0691b57c1c8a1547fb8871cb75e80f17575c8839c2ede6f6f69f2c263f693ce3cc796302bf706f6608c118c6c7735aa60161c62d7458d35cd000d0960c92b558a20e60dc7a30dee36fb90fa13d085998fa981d32e8ebecab80b7345e5040126844f962b84f85ead0b7ada23fd0238231370b3f50c72122b369b93e0201e7e1e67c33041881cb8045caa52dd4f245aa2cf76b928ad0cb82c2e6ca5c2aab52ce20ada94248a2cb5b352d8a52b8aa2687b6d9e88d7dcb459d3650386a59056220011204f671fd6623328337ff2eca0b0a465e0d470b6e5334e4998cbfc44eb25665c05b43cff7998f2e2d9fa13f5df531d96defe981f5cff8000dc5ba4a5f63d8a501af30ce9d2befbece7ddc64f40e5d0880b95f565310384c56cec9c209e48f10db990cefa9e18370ea456ce1b5b0ea98c46e8bfe67a2ece71b917b6cc5ae421d03da814b926ce47f398d4eada6c39bbbcbc5ce7e734696d9623f0c482250692f9584178cf868768a2a74c737ece9faf34052f4f136879332dcdb8813038f922db3bc5a0db786b86490974741f6da7404ff0f452dac2a4f86ce58f2a3112c5452e9861645dde9cd904271ec47d4bd2f938f3125362106c65ee02310748526d6fb27d381b98d22e749bc3464ba936ff5bcce99e826a8740490eec3fc99fb0a0c1bcdeb0cac155cafb884f1b8acee1677add679a159ed73b3661e365fea32e3842f077e83ff4ab074d4ba15053683c5fa88bdaed0c4e623c63a66cd715280343148e2dc8a3bca86b6c94f2ad852a909bbbf5caff0249c939d0aec2cb5709d5d48103d6d01692f525a8bdbca55397b52b32ec47eac5647768942afc6b3af0e33f707e40faf599a4da4a00c05cb30cb4ed5d96a3b0115d637c39735f911dfacfbd87b2480aaf178ef87e14611b8bf54b2c17731f0596a514154262498ea64e6a4a000538ca2f3df4df47d9bd5fefe37a7455198e23454354c4a5e57943d104fad39b2e41286efbd998179b66dcffa7d3631263e39a83cec88df838155644c9d870f8c48ba342f73e6fdc1f275412c23d83efea756b35c73980c65eb2e007f14455d55fd12c90e0e49fc6ec5f7227d87a2adb0a81eb70fe4deef853f4352a4f5baf1f56c51d2fd963ed6f6c273631bc56e4fbd17706e9ce6483fbb6f3b39c3d31b273eab8152216b51b25e0d5873d1e47fdd40e11015555214895ee6560a7a9fc2db53f56ebaf40bd13560a984b8eb29911c4a12a258539ae8a28287c428cbe6d0d2c63cb233e478fa0da9cf80c3af05324bfe85ba11134e5130be817231f770b3894de4f41584909f558b7168cac9d6c549d5398dc1e155dadd8b6b7d7c858e23fad12db3fd8093417b8530af6fdbb07e5e4012deee16db92f54fefc352e3d695f1388bce6c57248c3ec3d6d513f776f4d048a1ec341ed29f45270d55b5d50cbbdf490332ccc0303493d3e58becf537869835ac3d941ed69ded78203f4a48a626e35e2425067c88965da8cad2d25450b87b320caa3761511429b86fdd1cb2f75cb534eb1b665674bfb950b1c1aac0dc5cf7ada28fc5d9dc8426ae856155acd9c5295208c3d3f7212adc450b58d8e546a835d05ccdcc4f78d10e00abf67a0bac72937dac0ef404f222f3cdc157a65be322b0e4bb0cce6b451dfcefac7dbd0a770d9c0bd7a3a36010a2b789721b24b1cb63b0c48a0cf2c10fcac8fc16b42199df79be7066b0f36749cb50a134f33819eae6ae8cd49a8c25852e1822437ef5f15ed408fb74b18df4a86eea212e2ab26c6d9711c480de89b215dd0971577dcb0cfa99ebc1ffd2f790a380077a3bec9690fd3cc2466610982c996a0f87b9a31efa6be900817131e58ff558d05c9569e9d40c323dcc00fe7c661c13e6be2278777a7db427b7b57b64b3630dfe5d3dcb2b759f6262defcee73a02670fb43d1b414d15e45a4c401e131383754d8e37850a31885f99b57e6147df9e8071a84a1ea7773c9d673fbd0f162caaeaaf25b03840b5fb2d2d4f023fb19d53876643831d6e5e67f7513b2df06340193a3a541dd34e2f9281b72fc6fab72aa9c3e1fef9f6500609dfcca076f974bd1754aadff2ada690562794a79e9089ba2b8eeabc12e2a03056dc5a3a05dcc0410e6004bf22787e8a546797035cd261289e4cb7bcc9a0c620a3deeabf3e3bcabb9e17a4a645604a71ed25b3ef9a5a743cee4a1e00c167ed37f250db6b3b8a0a6bbdee1ba5ae177a5d69d3742a1bf9d1c44726ff4935ec1cdb74b47459dff3e33ad52a869e98a622fe6a8eeeb9612ae293eae6f959295fa7b31dbca7e3beefb11f70cc387e7ed382acd1e4498dc27671c45c156937529eef80d0ac2c61b835f932be89941d754b180d75759792cfab69ddcc9104743850b0081c9372f2323f8a3487ffe964b69670a708cacdbe2097f7b2bd8fb7b71a02d3b84555d40f082a6ea50314130054e110439b33854f14881d0b2b991228c5f24ddafa2aa9a3c3967355eb5b021bb911fb212a5b65d118a614d7148b001af4b1f328a77881fc2dad643d6501b33dfd475b2e8e6c66032c9f1f69b17adac23163183c57344b0bb92616ba464b785852472936bda72cc70281919fbee7a07370cc78dee7a51c26dd41111f750c0b6f352124f1e8953e9a9ffb9ad3ffcc294ee8512ff17740c17240a93b9f179348ea860a9c614a0fadb551c0070957c898c9f64fbd43be5b33b5bcfe45d3bd144e79ec084da968cd41c88e4632a1f68fbb6c719ef8103772a4d6897fb2f9d46db09998876e97df7916773218a1e027d296cdbd432a24816137306a875631eff86f366f30ae09bc89af9eabc4d95f865956cf656a5c097a1ceae8a693aa02fe5997abdc33f97e50b6253ec9fc8cb56325858ba9ff3c4778920548652750784108499bb56e2eada8f5a0632fd5327151c316d0708f56112a85e135166bd552578f63534df6310b23f48a19453ce341ed4fcb74648a768c742fac31780461b34e748f5f4b361ec1e8c996fa2342d4f52e805ffec7c7ff2b4d440d9623daa3abd8448baae4bac4b70623826cd4feb09938f3a214858752da7ba3300e1069396a5ce95171c904f4adf7431834d3441cfcfc9c1a1b2e24efa39e249b46a7988dc0613febc7ee7104f857d94f53cb4265b9bc5d04ca812c056423c106ae7557f76739d0ce8fdf52c069c16a802903f2f63da46e8e7b61c739c0e170f520bc02886da872177b082691df68852fadf6e8f0fb8a39a910eeab97d5b52f1fb46331c3ad679a4c219e163de5bde65438a2c4a2d5242f9c291f5ea51d75903b748d15ad78cedb769b0287c7689c43f9de61388ece924da01a22060a8c84cb3dfb3f14cb4435efd0a6c9b3bc5754e3b5851e88ec74d95980933ec1679aaa739d3a1ba1df9007bb15e98a6c4afc319c3bdba768fc165a46b6f53d7ae613ae896ae689e095520c6ee87fe6249959419673ff97a399db281355fa75d4955f8b16bbd1aadce22f37cb9a0e90ea8bee2053501bedf79a39538fd26b8d6c6e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hf7fbf18162055d70c9166ac54c6ef828926629aa5b65bdd14d8dd9f026538ee47684ded960f69e0192438251c4064aa0f7766afc844335ad0ab8fd7823b7fae178a93d9ebd9179264e7d3ecf5bf210a92b77f9b076332ec45cdc921b8f58d96dff818a651550d3b8b5f33ff0d65d299eb4775561b1fecc845ae2aaf6c8ef02b2cedf307042a65f7217bdf4f43f95c458c761eba03a6fec9cb39901b31f1dd6759a0bbc3899fdcd71c84e907a21e6c1ac868469a999e5169246dc5a056fa6b979ff03395c5745ae151482aaaeddd45cd1d2f92cc1b9d4d436cc4dca0c70407fae65acbacf1685df0c7b7c34d3405b06cd179a2503625a3f4514fcb6ef68094c8dc29c6561df315562a5818b91f25c9f2722c804cc0e9ed6014cb344d72f967dc82c46e41598bcb84f4f978d056d28d193ee6548176261989b8882dce6050a84f425a60e3e8f7c37289948621f753cd49d839736d248bf28306d931d7b5c58acda77fec0dc98e4a50f33928296d07d8bac06dc1497b9c1c990adc9b170d1bd6d9dc6ebc4d8042314d296e626bad09e9074878052917f01f517a85db88a0df00261d545e4891d7483eff613b9491a289f82239249b0c31aba2d7ea05ae94ed8cccd4ccdca6ac324fcebe1910f3d065b7f218e08f91c7b0b5f2ef6ad26833be356d135b3f2e5b98d4e0f44359cdea1e32bd9fea2178087bca1c846aa51ffca2c2212265f5457fce230ded727b7581b8a1d786d14d10db4a995b8d4ea6929572f47d227e28d14483d9ac306b37ff16fca1c3cc32a4821d102b68c89d1cddc3d90a3e7e0ccd6772dc291983da4ea740fd66c788eac068237513d017bf3c5c6ecf6abd3e9e3d8caf257b97a3cd195a4097694b14521822b54d5ebf2ce5d963681598e92237766cda0060e5caac1f84dd070076d2d7d0d368c9fb764b2efb8898d765717a95b8f2477481d3850e27a80e796104d3860ff35f7757b03e4454f2bae79af93980589fc435eb92d416e67122c5e446a067461c5c836894dac4b04d7dd41b74b22d8fbd9a4f02e178e444754bc89354c5c501a7272e40a21a4a1d9c9a261eb304d0e5ec1d03cb96bad6d30ffb4434d536e91e65cb12bab7ec57b6e0854960b1efdb0255ba75e649e09b758ddff030275264de8bd62f1a8ffd9c6fa72b8379cdd9784ab1622662a3a568a14f598ca5902e13aaf3031240fa8b65ef9adf9ebce29f7326ad7fce408bfa1909deec9e6b607dd6d7c8a5bd3bef265fa252c2c9fb104f52ecf2b7e449f11a110a76e5a0cbc15a653f23ce5556598d37b2ea1d63e9d4158528d4ba80e8b54664017cd28e30f8d0feb36cfecc532f342f83a64b27b306896101d9235b4f2d281636bba4c125c9e8f0ec1cafb31a6d3cbb80a29ad5dda3001bf4de05ee816ab3aecca233e436d5c3c4c1d7d7216efa9d098c887b02b0c95897be2a14c9e088e32b710550d6e08736dc8e3d3122d7d0387b4f032a5624cf37ff076a52e64dbad6667f23df7ab7050ad1dbbe5f2370b3b45f96ea2a1a115f270be8f6894ee3503de9b9d24c32a6a9d7b9b2c800b8dc53d1a208b6da8acb9d70dbd3d26b8fabefb4598bd4d0fe74f66a9007769e28835218b71fe1f24b168d1ba2e0e87d7b184ec1fe8bbd0290c01b615ab101c46f1749658c4066e042abb74296aeccbba8626c2b1e02b38288687db21489f8c28f4eac0cc072503234846ae2fb36680cfabbc2e9dd0301dcc0c6fc33cae8c4807bedbbb87eefa96c4240e97cfb616cc040eb24beec73fb487152f90614d59492bd62b96d091e47c04885ac34fda9cfc12a2cffb576ccaaacaad2166f088a3f03ada8b3f5be022e5569b3cba2f4238c4b8d04e3bbbe92d038d47098460b9b932d2f8268d6b73c2776774102a00f983e3e49177a86be964043857a88baf0535e65f2934d29ec37b6cc91ebbcf71c429ba466066195e029582311c4a30612c2ea12474f29ccf9c9fe437dd32dd83ba2cfd6a596c40ac56381848a9910eb8d5625e25f1996f8de363d38348301f8d747df9916b70ffaa768f4d8c901941cacdab526482537c6ea763b5d6ff82d2bdc5594f8f02f906b1d82e0b8599961cddadb921a9b4af0f687322b8c22aae1fb2a6c8cc37c8a542778445ecb47a8174052d80997e40936ace9d27f47a879f88e407434a0f7f93e2234ed6ae027ec829a89a2670aaf0b2afc3d763b9cca59bbb78046addadfe4a18ec43ca8ce99766352d1b1a9887b28a242ead47d122688a0be0d16eb509a6f32039bf3e0c14a500ee16e11d7a340c93fcf3c49885753538257128593fcdce3a3a9356b0bc83927ed44f627a5d34d20166560b8d2e3ddf505d7c738a4d056d64b75bf3c3fadcf89209f224b52ff7765d5fddc1eca6f061f95f18d4d980523b9690932e4f7f48c1a998488e7e652b90c828477cd570ae6bfa84a25534b0c95e18f3eb94b71e8da0a7404eba692f8b7521d640c2f3e6aefc706b7d1a7a93e84e90c1918349239c54d54e0190f330abd8889c0492d12933edc8bf4fd5c709ad38e4846a918c2015df7ad8245a573050b220f099c09e85d0ef851254746b6b3aee0372cc71a89978310f07f594555fc0e380c2798dbc3fd6137731c4925428e9458aa16989d589f8db4b3d99a5442fcf156c57cf6834efdc9b4c6952e493ece12d61dcd0f95b427cf1aab2ebd127261c986e243213f43d0be82b79ea29eae0c038ce0e9c75ec9b1ec4a3e5d4a85e0956dec5b5c4027984809b51c817f154cfa1d8edf5344409db1e44480af56354446b5d8b7e2e8fcccc60246dd2ffa083332572f330a2ea433d5c691a6926a0941a23252bf08220caac08953904474cc7ad26b15379d54646cc6b5d0c5af9b0851f8a98fb8a57903dc250458a982aa3af78c665ebb8a667f76476b9caefc148541c047d97dac5163c8fa0fd57c5bac2729fa7ab4fad50f97d8643b758142a26feab6a5a355ccc94011fb3a2e39a12c785440a3f9bf05c11b9dacb7b5d4d5fa49badb7c3f0a0343b4f55bc1b7b5fce72ea7b27dea5ce82729269bb4b24a38fc44701b26dd9b858d29ed2cb93659cb32922e7deef62103a67cc3cec69b8483ab7a825b958cc0438df58ad41e7291eee576f25131ca967be8255987c3f4a57e5ba3338777ede53043119a06f831bef81e816a9836c324eb51b06fc8ee6a96450356159814c7acae20ba210b431e2aad3c281a66f269efbfd1b0a14818cff83a53f8d5b7dd5ec7eccd97bc27e8d9ea417b29381b598febbfde8c484ef10878732f85bc23ff6a3a2550d2e992c173609c8dc0bb406a1a2927b6d495f76dab70011dd7bd0a4ed162d44036f07a1cc3d01573b57a512496c7d6e1c37b1dcf9d4da55d4d9ddea79c7edd87ecf7247ae1e5c994f5319138d0a93dff57180c9a026793ae4272255885eae0468b60743ee8dece36a548149a51b70903fac523e0e63589ffcb45de89b1a854282183c83d4886111c5d5245154622d1a399cf816742f17c79e85218a0838bc688df4e9def1f07d58c2901093f986f60107aad900ee51d25adca51906761615675cc19e9947e2cb8170ac5dbeebf2bc52324d7a88c8e61d8a0c50d5b033a6cdbe97b679cfaba2a51bd5a5e217d4c7f97d459366a5ed447c5e09ca1fc006e26898699acef15d5bc515d86de0c81c32d5ea503056916af61dd62a7582031f2c0912b3ce5d01bc7ab16b406db60c14623066e72cefd0067b352986254f48b86affef865d4c4345be503fec50a3667969a19d20a1c8927c5dbb13cbebaa51dd4a70489f7391c67fa01a3808dcd417d9e6c4e1ba56ff7429090ce089ba3683002974cfc2dec9388a08471ae8eaa1bc126b9b9859aaa767ede0593dc5385dcbdae7d7c023c44208416ee445fb45dd6dccacd644387e42dff15bfc32adbad617954147caa75a60c2be0fd2b241e67e919922ce78c5fc87c88bd854dcf865f3b630cd88882b5c354431d6319546f96a6d82dd417c6a01e5026d19da92bf43c0273ad373fed70927db728123faf8f174faca928302c5d7748e9b9c37a8af726d2d5678768fc24e649780a02cc64b2d829523a25c03a36a74d7ba68b5be45df965539626aa772cc95ce4e2f1bbf07ad0fb1ddfb8bca93f17080a9f17f21234bb63bbe5075cb2413515635ca10a9346cd507138bd4d08e9bf5bb2e9a66e3df102be022c8dbb5fa513b5396fe8b43543fd9f8b480893c6e91cd264f4684005928ffc9f73f680613f5bf0f0e3d1885f2afe79809e294d3b5501d649ecebf75dde31befa7fb17c35b96c5c80d4690df7cbc04b771a74cf80b70b5e1fd25f28fb9388b977b4611754cd93dfa53d5fb3c6fe7cdeb8e019cb8254ac9c3c69c9a7cfb065ec0ff3e389bc0b725dccd1190a62c98f135684b8eaf5915a862a5152e830ac2487a3cedb75965ad388875cd51d2718899cc8b2fedeaf243c6c4fc74da61d9c248e73061f42e8ab19c90bbf4eb2f017abbaea5d149f00025a4466c4e62d096cf1a3ba6909d32f70e61947f4b6bb6f414dead0029bed9d969e5c7c68b91806e0ee30422c491a22872efaf7faae0b8a93a65fe299e369cf0832a54a59aa2b0140105bfb6ef658899c6e88b1dc2ad8d26e8cda804fecc67a57fc3a24e62edc02e800932c9fea3363d8e82e04d602d16f9afb3d7b41e0640769bbb863c716e223f32432ad7e4fbd1ace13db796635be0aaaaef36b251146f07c00d5c972471b6efb24162ff6e7ce4d5131570a916aab7af764f4e23bf5b4f3e4829d16259e0f9d15e93614e04f125fa73b1c5ce027f6fcc672d34d0ebcb50fdb06bc72f86dae2ec46cdafcbd58dc087fea4c5d7755cdd0e2f0bdb460b8c06c244f0e163344b126374176f65058dcdde6f5e92b94487e5eb7b88081f39f48b7a98011fce146c63f06c68f2fdcd8d2293af92882d5309f41324912d93ca504661d4f35f036a091eeb60a40b2745193a4141230194e233675272c00e7e03f9fcd4106d1c8ebdae28f103d8d87725374e4b53c28e1eac828d73798d4ec86ea8b8c96a19f97c6e3f58148acc2253b3f4d5b9634748fb1ed78797b070d2447ff4f9f7ad1a2579bb426235f85f40678e799175051e0947f0ca4fa6f604e741334c9f16d7b7bf8b08a25442f5a5572efa0fbd6e32c9ce70771597f9c5623d84313e39beb99008673c938586d26b4b1185e751e571f554c321e0d7126f55daed8e3d3cb6d3be5b6f6c90d74aff43e85ebefe9e8144e460a905464f0e9442195c48b7cab4141a9796d28214bd525ad8b3eb16c5c0a334488e1c834d9d04170027c045bbee730f680d37559b6351d6918c3f96e6782884407e502e7277ffb92f69b10ea79513586f6b67b07cc704c221c26119eb22bc01a1d2acec5e8f7902fcef4ed14c008e737d87ce474ca3d9fbfac6f3dee395d6ed9d9956753134a37c111bcc1a868051b8280ecb12037a05d0399557b912d6c4930d7f7c887b2fa860bae52639f35c22500ceb0561;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hb75f5b50b3bf3ae7ff190105aa931665f8ca17df643f5884b7588eb33b80b83624481eb5291c4fd4a063fc7992fe53e75b2a5b76bef058829a0dae7615d76c55cc47101df12a76bd582e64fc826a1f78d7ccc6afa0e74aeeff4b96f90597600b82a6794bc210cededd12ef9c9f41cb7add97d5f6f627fde1b3a97b76c5ab9857c06b89889ac6e0ae82473ca5a40ab2f45b0daf75e967123fa492e7dee7178f8688a5a4ebb269f8c4f3ddfbb6fc47cb556772f307a09ad0b92291c327e36705a6063d88c7646a586e4239d37b6950855b85daf2684b44b807d577af7a627642fe14d567487d1c93c5d4b737746fd2a2d7a6001d317563903b4ca610547855851b814b5b6686b46e137c3f0ee1c6c368f0aa069eaaa20e968c5740778a6faa04788c2c3ac28dac4146296c9c65d21951dd8c031db0c6b81ff5cfcf9bc211daec3d4494caba3239340e4c459411a80b6b24eb6737c742dc3990730a5bbb150baff42022d10d19122a5412e7a8ff0080b9377a03986561439e869b52947039a958019852606a57dde4c80effb384cccb171bc84dccee789a1f20920e03760545edc5406c63cec71458cd06c401c2283cf24cde200a52da6a9d58994a6a439c29f982495a4000f4dc165090abd39e1b2db104e3563a72e481ec957a2391237b0d69d54d26bfa9d4edef2b4bf3729354fe935110b4194d098a75e07d8626899c75278514f6a40ed78dfe46f8de0b5ba74d890bd7b2f3e75356eeb5097b8f7eb6b9ea4bc60c9df664cb15f948d8004fe7ab059522690b3dc8f7b9bd3b1b29ee637e6aa0981cb2c3af4d1d80a1d130ea10a5d27724441c55d5145809069b83d8f9c7492662c1af2796642ddb73d5f0309a53f48c656aed90d32886d129918a4071c1d34f9f2318dfc670ead0ddd21ee24861055587e1dffc75693d612a6295cf549a87e9639fa9b04b9d3e0a76663bc9a56a77bbe8e6252c9d15bc4f8e1e25018e604ddf43fa4d5c16aadbed5902dfead609ab4e3d38f9b3d25f37b49090661a89a16e14dbd1b3203c6a783cb4dbcb22a470dcb3adb306fcca3fd9bb682f77ad01838015250bb8d360a576fe5b34f18c64bd6ccf08800908a72790e80c2ede94fad519821048915c63a3a51ba07dc5ec134c2e935d0c373492397696c95b01397f27bb0e54029f4f6e994f72d276ee97bc118a2185f8a6efcc05822eee6947a08c4ae6afd693498bf3133c693f34acb5916025ad1d72654d258cf4c3ee870fe75fdfe436c7bdd7df61c76dcc4a87e75732e20b1c83bab6dcb976f760b1d88b0be4be21003bc5f04abda3b39ce61f19b0331bc4cd0222b946bf2f81e5b667d8b2079739eb7268690e1c83a5811676dbb76692ab9b0001b2be7d1e67d23a1579b0318f38034f0ec9ecd9222bb182bc67573793609f8137fe0ff67ecfbf51b35c442a62446de543a10ea965da6dcb2fda8865b7c18d863076121b1c5bb67523175e6ec65e9a998834fe7e7ba3674c3a2f5189fd34716b14c7a65adb2a18e9983291c08feaffa088b16690b5bdabc72c27b1c0ef7351e0bb384c80628c9999f23a6c4e799c7bd6b094967713c9ba7a1ce0f14e1454ebbe602dad49c3fee02a2e3399139318fdb29cb04ee29461bbb68811e4e393801fbb444a4754bdd19ee2452945f56966d0ae9b2ed9611074fc7443d5c3af01549629e39d4a6613c7de8e1b25b1de1e38cda77096d0accab939d260960a1356d9fa19ac77c7ee76a7c9b514a4adb6cbc2b2bddb493d8e210ed7b60364af03e8cf9ad0b6613e062c9807587dd409ea596beb2a66cb645eb8b57a8225e9ad129929352c39c8f299a009033d670efcaeb1dee1367debcdc0f0e99ff99e94cf4b71557597edc4fb00eca497684496db26d34f106b5f74132422ac749c61a8394eb44d719531123b1ef7b4ebb9b46f2d562e3b780bb8dcdc1508961db3653b8b5f4a75ae76f987e2e76523e14e4706da17960dcfb44f9c2be93ce29e6a71ff39f30f2fe248f56ecd7e26340cd05f75a778c97d156ea15311129b61051ed41f50b9f81c839ccc85a951feb168a627b36d548e2c3116fd6bbcf35b6e17863434701109c159b81fbc67d675b7f33b09743ef6f337e7f5094310d66c7d9935296eeeefc3835d30005308dc41f6dfd11cf78954826cd9447955a70a2f52db05cbf7f55856698c808677740e685b1687374670183c4dee1a6fa068e92b9aa6c2b2dd323b319837feb08168b822d7ef7a5658ef3a5a9b56d358a3150138a4a64b497b55261bbe7ecede0bfa6537073a5ed9a621f937f875095e2c26ad30cefc9600281a3ec09a56404bac1d6cc688247dc2e71fc212bfb4a9e432ab5a32c1369d29e4c3747114abb080c8bd3a18f2ba2c2490fa02284976b6c4e00dfd9f196e7a554210f5f94650a548d7d44355ab57d248b729eda8594b399afdbba7d7d5fa571e62c1dc68e0fe5f2e8dd509c650254e963f703c6e7f3c1ba06b16e14550ed52d6c5f467de458ca38e30b4adaf08ac1437bf8ee1a18ef39f77846a42885c5b4313c5465229f8c35f6fb4a9d49a7e862a4061fdca688e32ced219c2465961cea615687bd1bcd9107bf055cbca418af4171039dfc06b8aea3228c8ec928190db2a5ade8e0e1b03a88263e67b9fd907d5313a964b1e58636bb468909d1c9dead17787f95ad58845cbce282ddac5ebe43d46db1f25f93cce682ec77317cc7dac0b0f0b55e3054044b8c824204389260bcbcb94e8869717a72023ccd6bea03b1cad029bc228ef4c6be372f08be8f37f99106d4170406f6b1becd57733a962e3f01723e56a5af313b34d14f2d7caf4e237ccc9699eaf1975a831c6d6e2da284ff0e8e6ed054a447575ec3c2fd3c64bf609f6a02c93553390195cf2d17678203b1a6a29bc787263d8b7d63c95194c34c83a4658006aded6c8e91e9b0e88c373f0575c92d04e102b7eef4a1568112bac10776996f22e18f0f76bd99d176d6b872492cc232d48bb735e19ac122f7739e27751f239720a76038b3d8194b297acdd7bbea673a4a29a14bc67e616e41d370f7b716c9b3ca56e0a6a50b73911f9f2462acec5d74a3844703ac872d464eb46d44ff25a8385502e806e529b2285430de474700bb40af2a71fcf47713e7a970a7692c7a4f7ff29abaa3794a61110ae2dfb19eb5c2b58589f7f0669d3b6cf1a2cc1ce7149152a70331ef557c87859d622f974872ae70485a69f143d472031ef83493e218a687bee870e60e6ef598becb485ca3a8f0ba0f47a166eb8e39f72331d6d0b41f767979f4090f26c0c2f3c6abb172979c62688f1d21d9759b566bddcd580ef7b0e82eb40107ed7b744da9c6bb69ed194c3d41eb7b445c5bdda803f44a4372698c209980ed91cc74b8e498fe190bac8cfcce5526179ac41fd0452c727be2c85c9bb9b7f27864b92024b8e09af00e70dff6720b0d7b14b5c1f6a8e650e1ee84d3da88e888cf87855aaaa1a350f119aeca0dbbfb9d008eaf0f53b834fb195ee75274ecd3cf048d52f179f6ef2425ae8f50f40c97cde3465cab8f62b6627aa80f52d0c860c0ed3f9084a09a4726b346f8147ec09f1f51b6feb218d786eb14f0d6c07f3159e02e129299bad1dbb3efc4f726599587cd4b1ef28ee208808c8601602ddb6ee60e435fd252ce98bc519d296b488dc7ec3d4354d9d29ab3d8a8d0e7306980310b19fc366caa9d70d9a42f6d1d114edd9e496aa7e3fff34b107c027ef973f71f7e052d350adfdb37966b5a26914e5883beea78e3118ef48213df3ea982f60938d36f4c6a000fdd6a917d9fb2b25c73220db9589a1dcea81d1a4cb300c404623d061edb377d3a7c1257f273138e6f9b8458ec312ac5ad24651f0bde9094136041264611ac63ffd117fdc61a7a0cf598d091c036f1d6bf999885b24f62b11961364a015b9e0a0ee163c357e33bfeedf33928fe968d2a3ce4f1053f53bfcc312d629b8c65dcf67edaa76d1c4ff53c111cad2216f9516d0b81af746cb88de24c1c5444aac331f00ca0a4aaa632dd3fc95ea681a6d85701a4825f82778cd9b6315aa24c3fc2f328dd16aca6a149d1f1c0af50f87a3ea0f1fc7b418bb9807b63ce0b15209c3680bf571168e485891255c787bb008cc10673ff6a1e46db196169a5d6f384c8441cc96a031f2de14977b0916945f99f17946337a377a176919a312e1ad92f0a4344e91161dca34fa1580de07996414fd5c154e65463f81389463c963808aa151d2578163456c15a42e116850094c19b9d6dd283680c4130db61894b7304b78cf4ca7a19cf89babab480f770780a6a37f9efc3e7be4b7e3e5fe22cfe9f329f247f904a4f997ed43c0369f59e236b4c8b5e47703dbeddcc3689e8204afeb8e0a79641d0e2337f9d2dae07e024f94c2dcc19aa4f0e3c85ec5587471caaf89bccf8750e8e431254582f3419eedbc1d4a7b606d281f004c9ae280bab22868fc58b4398fd783b1ab3fd7822625e8e6070ff629cb2d5e2c6fbff51c7cb18461ae6b16d5c4450afc649583e374c554a4fcf45ab82115fe25f5b0934712929c82a87ff71da3d087455695cf1a21cdde58f45f97aff73c9489761d6261875de018d2f91841be3d203e962ab2372b3a33a2e4f5c572d6df5062fd9a3ed6b537a60b577c225a6c4e17afc4c6e125c014233bf983a7089e44fda48074407c08dfaaaa3969f3fcfe0f0e939529755d483a88270d24e889480cec3dc514388e3e494eb9deeb60eba1e5ea29d27b93b603ade9118592cd205f291a4a4103d74cc840f0da425689f937690394a146dbf728260d27aeb54bded35e6dbbbc12a7293f3670614432d6ee1727e2ee709621c90e01c880465363ecf80ecc3f4e3b85f162ed7b8aedd35a9de9228c5956be01c696c2002600a8d923514c257c0e1f4cfc65fa642b0c1d9ffdd17c3fc882ae6f665b18d67bd9aabc05fe95a298a2ff21a8c40532f4a637658f621c410efde8bd84d38f6482c97e841926fe620dfc7bfd200694d469de5dc85aaaa3c40528b4fa53e5853ce1fdf202dcbc5b9c1e5ea4816487958bbd53132b8fb51449029b0bcee4921c31d78292b7e0125010210b765208c9e7c19f26e5ae2c502141c847351d4cb381da701ee2f2934e29382cd57cea68919cff60c0557ac9d734934024529479ca01822404b45467cd60d031d232318bfd9acd8148dffb1cb165025187fc0c871040bd83d20337783a57dc254842ba2bd48efe18c8fe8bf8c579ef9995d867cceae9b3d4962c2e5b931663b41597bca847ff9e2f46545c44709cd8acb32c3e312cec4c55293b9bb577b805796e54a7904ee776daeee65b88d2a87c009c86a5b02dcaeba473bac7af9b4d93091df8bcb42014a4a7cef0ade2699ba6d8db3e315df1e26471486590c79ea6895fe72b8b357b355d8c65aade6a6d76e0fe95b3fe09abd98531d61f9c71ad1049ab05566e815f7c843f5c38a2d8134ffa498d9b161f6554404fbf7da753a385987430;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h8a3250b8d90a5aa6770953a2b50575bce4cf5d8c5166d276af39dcbbf32a9395b432b5e44040b2dbd87f9ae68554b2a2d3f0fd92ccdf610843e2a241e080f356993ea0e65ad9651fbe9fa6ed3b8ba382f8b1d403ae2e4eaa4a6027a6462c81ce67de35e26d2ff09b80822972d1fc07ea2aaa1b1fd9ef9518cee77c707988945f7cf43de14ac0e137e2a46e07a878cd8e022c47d579b5a59ac80a8bd6ee047d882216c9e64c2cfac442cae9f742723aa78b133ec5fdf617833196731df8ea75be16da295c03093e64ba3b91fd6db846112594295132e158e9daef1e9996d65b1d2327f753fb2a26a66205ed8f1eae2a519b8a4310f3b266f797959299d35205cf496f3d04072b25a4b713ca4cf1a7106923b9ba4315f3fbb7d17853d048571ba28d1e01e5b519daf9fd83d6b3d6bcb6b0dcb74437c63f4b731f4ed962d6346634c762cab0b4677280be614d7229eca379a7ec288239fc75b808738e6f6995d86ead4a5f5395a6aa1a434a91b02d2971cbd386e1eb29ea638e8f5642670f72ecc4b9ef9d16cdc9c0cd5c82d54a196ad867a703a5b216c0250ea404c1fa737f74a26b91b3db784e10352603641bffb092fceac9cc631359e775439b521ac0804f55891fb77487c6f9a70de516b28693ff2cfe6a02f8e77e234aff8e9a84def22610fc9b21203189f7abd3711a8fb2a237480220e3607a854fbbaa54c3698c9c6620d6304e73e331f665b69d50c8c6cfee8c0a5bc76ec402645613929931c38e077bdb58aa11fe4a80d6b9fe9dee384bc2f7711a5297e117ebf620672947341e010af80836fdb6ed31b1c0ddf79b532d1170e1824e95e962e88270edb77ab3f397a4463c0e914701fd8c4be5699d7bfc0e8e4d3653814e36e86c63d078e549885afeeee562e892a3c6efdeaec1dd63075f8bc19ff259effd9e39ac142ff1ec4768b61e0481bda7f691d2a474ab511af0ece9c3c277fc0b596ce79d6d021d35bd5c459cf14a2053a58932cf7b61a61025338735ed468ab35a2e577384992a08f8782b8a56258a602da37631c25a043925f5b2df8326cf63f3b57b1e0ee648754ae88e08e9a6ae146e8b7db3354114e2a6b18a44849ff1bce1c93fe83ee7d7569efddc3e5e68c77da1068e746b34f95c970b5130098ef459537d09a6ae169573b0240e8f8a960b191253f096977c817c4136294bdf283bd6238f1b680b47e27a3c368d5257518aaf2df5be1d72a13efd57ee80ee4191f6cd4989ecb7228430fc22499bfbb731ee438aed4fbfec7b5f8e78766cdb5c1cf94eb37ddd76f18dda352a29894c58017f8ffacf2c0129c3605cf0a4ce710a9d1a513fce2822b7d0c50fcad5f969bc2f0cd182ab9c276b64b97fac8e0b11fe24a508e7a3b22b5d3c482a92f08ae72f2204003eac4fcf83ec31deda72478acb14401af0d285f12e29f1f53a571966dbed7344a51b2d13c737be6e882e56ec6028fb3f2f90a68180bfdba89a48dbc45e69d1def703f2da155d8b7248e434955aa7772514d12d2848823823c27729fc41b7e01fb614d3040b56ad3b0268692e586fe8eac167dfba1780c19f05071985c7a476bf35d6e1bf81f594fef0e787fa9529fe6963eba12f58c2a4be16ef796e9a051f71b16a2efd61bdd9310e73eddbefe69878f0dca462e9b42e99024b758493d1faa5f1bc2b4ed63e4856f8a9c4a56cb207fc5033dd595ed5df0aa6b4e84b9e9e8f6e3b243bb9f03643fb178e0acd3d82e1e945af23e6a195a9ecbfbdc92bff12f48692975e88f83cde3756484b0dbc6a1f5104ec4eec5a7f304e9da1eddedbca441668ef9db2bf6d4d6a0ba2599b1bdbe8adedcfc8793230f7c8f3ec319cef19df0ba153d7569a8f8600d5905c3de9dfc0dfbb904e045cb00c70a1c41dd99d6648b4aae904fef680bdc89c331481377f6a2b12d6239c669378131e33cac5f9ac055449528615249c1e856a84fb7c7b76b407578dc20ee0f61c5508ec7e3ab58ae00e6012343b907dfd70055466fbc495d98567b1b0b4f290af8b8df46b4c5e2e1a66f45ba113ab4e7fc76b5621d75e27be26e52b2bfa799622acb9221673f027304f6d2dbf2963d1d1e296450be0488612b92d80c329904e8bb906746160d65ad45fb25ff1e83586f9caa086eb31826be967723f0664b1139b1eecad92189a6c3c7e5c57311b9933557f6d89a1e5605540d9ebcb1612887549cba9318e67f4a83f7984f6cc1e2248814d800f32983f610e14c13256a36ab2446ef4d7aa595c6b8c5f57644f6112ce38afbda9609111e95c6b08aee69d9961c5091e3cbfad0c1c62f535461ad60f8b485e2d5885c660a01f952309cb20d6687d4a2f7d9e133e9114dbc242b0688ad5ff95bca23f2e7ad5355aae17c84071404cc074811d1a629c54d142ef21dea961cd45a4f4841aa2a1a3aeb063a522e4d82e300eb62a1c4556c725c6939b47e40508620973a185f75e1917aff94110401f0d1aaf8b99570f8e61128df58d37f49dbcf730db8f11cbcb26b9bd1dcb66a4cbad6a4a94c0877f6c75dfafea18927213176a91a857989938364a1c94c0d0b98aa825135d8f2a2ae3465501ed6846b01a049217398a24fee3eebc64495aced414ca043d24b11ec0c6e8c3b221a44e1cee2d1019ba5ffdcb81c5e81ec811330d7cc871a9b27bfbd63d5992ad5ea56ef6b1e0ef23644b533fe9ee8a29622308c63ce4a40bb24a75289233bca565fe012d3e72ea27ccc68bd5a374afbaa0b10ba22502c00f75b36a2825d5d58e708b1aa927c953aded784fc81488f1edde8d39b90e45763244fe876040768d3f2b747138c8d80f2242eb82a162e7444f74c8fed2db3516549c4bcf1cb0b1213e9a8aa9f36b3886e226383865d0f0525a32463fb768647bfd424141c79cca3a0491c429e4a5a1588df0e6b6633c6d453a9658855090406dd92c92bd2a83276d1328c0b13e3d833394fc4b441282ec6569160f54e128b4e0a0660d959dc73db95266aed5b3c5c358228f6fb5c7f64d39e4aab61c4cd57590597e1fb1c7f15242213bb4de28e111373532cfb76d5ea4916724a48fd0d4d25239dd8642926f83c4702f21526f3f588a30af5fe288258bf4c216276c77a4f0aa8ceabc95a213a338914f070971bebab5cbbf4b36f907d9114ec3ccee1ac095c6f2d518ba3e0fc4da73a0d26dbd8dd0b5568eab56b0da658b27740635b5ace7389bb66648a7acdedb64ab3d488d4c346ec07b8428fce9a86636d741692f4e14df256551800c0d5975be1ec1d1fc05ab44c7e89b5d128fb9fb1904b2d24150f69795e980c3fc9fe04dd94a8550730749efe9b3025e9af11adf7d030c11987b5c1cb33a7534051a16c6fe36dad1daf8cd0e688df69424060dd088c656827b58f6606f61fbd261299414a8abc4f02775637e2e5324483640d11e3cbf40dd89d965ae5f627c0e49bdbc160a7c5fe9d32ee3135be0067eb9f3c56953d9b656990561bb763e972ca1ae639814ae12ad11ef6bb097aebb08e45dca4f0c24039128559d6305f65e63e65f6d9994f7470e67892e8486d958859ca879dd14230b21a22103745d32b1cb9105d169ba6d5243489c6dc4a0ee634bfe8447e224a3826673c4379d5ba35648cc47544af761ad1a8429cd7d21dd59c46826c6a5a361157a5a11be3acf5e68decfaf766b7f4b8882b9a462e8e54cee017e0d131efba6b64efd135b1a0763434761b11035c5dd760ce93b7f52da7cf0328018508f86404526d4d0bbb85c1c9dd925688601f788343685d883923958ac0f5149c85981ef7ea518ba1036625a1ead092560836e9f717b4620b43c8985e95b4fe67ff84cf51cb7d7bccc16ed086b494fdcaf91ad3d962d954af46c135b18d3561f914357a828a4feb79943f5a30cc72150d21cf25d1c4a9d830e0a2f253ae454b4be50afa89907df60704dd5f6c5aaabf3fe0b2ab16c1e1695ab44e9408cc2d02e8f472cb0d09e2d5194f89fe97a9f43483f72316b3d78fbf42b1c8a700fe52a365302c91fb378e6affc8bc65a4e517438c97c2004531e5059da9bb5cb7edc751d11980a63fa93e1838dec9a9e4a2360047b47c166d0b1242c5606893d4f865447a0846b9292b43710b74dfa33d270b05a8694586973ae1298927003c25a49429e5b8625feacb86d5f7012f44f2fec27c46ac644e85b3c06b3523126f3160155e50873cac9863e9406c1e5016d8fe2d09c618c6d2712d4b1a9a45af7900659100cf952fed70cd93240703be1925a9ef98e2e2074320229f10437b5fc7b9fd3a15cccd2e2a13971150ccd854befab9091d7ffcca592aeeecc2a801269815bcd3118b2cba9558dcdef1c73692f427b2965444d5d80e528da7ae436b11b477ecee7a84e7924e3e2d394933cf922d2e140d746bf8b93408b6cc8ec3f0345b49ab09774d390aa4644da9867f8ec3c6d4a21eaac560c736cbadcea7bf93194b74301e14be267c91840b427dd4616a038e6e1a9ecb775015d95c22df90e19f38bcb7004d1d5dc6c42222d0957ee676fd5fdba4daf06cb78c5754f733b952a1e6914607fb04c5a0b733bf9f56d40c59153d42603c567d760b336853525aa90958142f2b6149416132592ef30ce4f577df1c5e803b189b51c4e33b5da0f83dd849840714bcd565620315b0bb00546d77909a45158639ff52f770d5221eecf92076dadbb7533594602e9baa95ee171a7ea3d7d7a5df824e3bc9ae061953f3e7b6ce834eea8c8c814679604e4d4e9216fb30554a31cab859599ccea3ec13a80216270b1a2eeb501270709c474ec870b729ef4d5b7cbd388d0d491e01844c36bcf9dcc3ec00c656ac08eaa3e8269f6de963f3ad13169e04f9dc4e7311291243f2609a2cfc5d7df9961bcc9bda3bb3dbfd9f2791b328be627ef98979e130acf8668d22fb10e2687d4ff64b77a5d5a443114f7a637dfd2743697fa009c3cbfbaf510bbe5dbcbe0c4f964692dd3fc64fd4454e69aac38211883e99b5ac7f34a02ee04af1d9e0e8a12d5d3cf535506df7f9864e0e981578ec289390a862022f8933691f422491fcbb67e052f9069e2bcc6a34845d2b7c5ee629916f81156095a4d94086d59da189440042141134121c05348a8992ca904140f0ea46413c3d25e9ae0a440dfda403ea80affc9430e8167bd8357a4fe020ce59c44706004b721004c27c9cbfefdadb7e494ab5667e6c0c0b0c2415e60b7e30c0e3c3852e3c54671e0f1e5e62998d1ca9947694b7eb6dad7327af8b29f321311c4d67aaaf45947fd9ebe1b9c91ba5d6335e9a92efea39a051ce97b3cd95cee6bb111c801f4a8adc69512ba2716f823924da7a7da06c00dde5a767a365f4ed80c914c85ede6822bfe3693b27d84ee6d34a4aecc2e74ba20baa6f878e11e036ebcf51f3c328ff3f7a0911c44bb00016d761e98731de0fff3222bdc68d0cf04e9f64eb3cfaac867795805379cbf0ae1e0bd8f1ca013191d33ffa7d8a0c9192d1f6aaf4e5f19c06204027b6efd9e7b03;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h67b707e01bc6a1b22de87077f33bf25ebfa83e3b1b147c5b88d19b550346899fa680a1aae7f90fe9d0bf1f77bfa799024a77c8dac6cdd3ba24df66093420d04344a4e75364ba2717d52cd4bc5e92e57cea58212be58d4b559cd5b0ff9b39553ad2b865e9340316bdfc7bbe4ce114d76a50f3ee9e4e8c0778ca483485f2d7b30c4753278508abc8ded3831f458b9db20b13f04aa3231bf445271798ee16df4f66e2cd1bf0b1b161c9850652af72b1015639c30d635916a2752637918dd91752bc64081faa023cbae7f2778f16fb091953a53fb0eb2d863dd085365c251aa56b7e6a5470d5e8f66b436890a36c40ad89682e30a57b121ff9c0ce16b2f6a39cae8634578257f78eba11069e2ac6aed396bd394c52be5dc81332941478824bc393ecb43db699c016b2e81e205279ec6ee5a3662cff04efd2958c822818ac00cfe5262a62cbb8bd7bfcdaffb19073722d625e025b8360bd1fd664ce18cb984603653e95a793fc41e827159ee2207ec43a44b9fb59b89f24426910f9b35a2b24d0ef4f89334d39e0dedf26e1fb179c019af7892cf302d179f62b01cd9df6b5942783b0a6cb951b01b6be90da38cbb80b8b08fc4e6f020d2314d150a752c9dd9e6b1e7b83bec97870b607c567ba3907a90b49f30b7b745f2e5692057483905220b0b08b0a15a006e815f7617a91f85f1eb5d62365816328697841d7b8f55e6577546a968739cd9e0a5fdd6f1eeb38d7186211dfe4cfe58da3aa2978f6e47cfd5439f110084553a0795a8fe0871b4bf8032e3048280939ebef3d89a5ed25fe06a53949e94f1ed4148a44809aa1d6f06e0202bbe0da2df59b2e898ea5e18b4ae2477dc86c62b1a2819b7f953697d877e99d2f9b270cbffafcb37e488fe882d8b23fea144293c35c90bc9fe8a8c1fbb25433b6db7c4687261eb043314306396becfc4ec86d8588482a879f4b20764de265c83730e1f8a6c211f34518ca153424db4527740a0292d346940524f986bf7ecde9392724b7ad6d2d684dfaea4738a1b9b7253d7e3493c750618b5833d15331679fa4596c8e5a7b9c3e1ae1f3b6755ae16137aaf82a0ff2d869a55c65498dbf005489a34ef3a2a0666f1599b640c0d85fc2763e701b80e733085fdeff05050578265beb8c37d3a17dcd7526e6cdca297bb763c802db028ab940fdcfac2874bedf2044e809933ee685bd2a3ddca2705540f2f6b96a7a85323f00a9ebf5fd6305abe8f4a86cc1206d13fed8af34ee1b2ab5fb1973b84322df2adf9720b87956f09b4f0a8b79b93bccaafe115a88e5164ce932384f8a83ce9e40bbbd07b5becdaa8f019a581ae3e81a552cfd324e18bfdc3ec5e45c2dea428c4562c5119d48f32baf3961a4bfcac7c1ad83e5400d789f5784d1c3406d0e92668659445f1794f5c36890d9b937f9a5087434a2309962899a2a675b509b202e129a637628e52922c512918308b8c559a8149d1382cf0a9aa1918f9dad2263de67bc5a37ee642f76f5062c9462432964cb3b7c710975bc443dd9c99c0d4f17f09727361917b6c0b608056b10be604ecf1816bc5c79f64bc1b5ddabd8dd1ddb3ba070d779999590f0327e7e012f48fec46b1448cb32520655b2830be05343f0f31fbef1a03c4b3c8a65f724291b07a06d136dfb9a32c8904b11009f7ff598e79a82f6d613c47182116bd583fd2ef4726c8d4938c361b156ef935a018845c075e08ebe8950e52dd5ba22e2d26ce3dcb23d3eccbda2503bb40c8f1715004c495a8db84b41214d211765e2fc7d875997018ed0c956f0f84110b6ce8ea505229318ab03f4a4be3fbe29462e5538269bd3c1e57dfcfc0586cda7e8c5d236f9cc2a1599bc652db03484895735f66540bed8f41b8c508e3075a25067078d8d655904607d23eef6897e3fd385e2fe54bc02ac2e72a31c3362c56207a9eec30eb05dcd1a9c8f0244eca21184ccf894db462d399fafffc86ef1a5c91d898336ef0355314b09051a9eb0beb6887ecdb061d024b9bab6b1cec874bd9ee3155407239659186b74b7f27e46b1b2d561cea1e0f0e1ec6d2ec6bbcf437b9772b586de6dd75a627593555543322894fd0e77a53895daf8e663db423f167db59b4694f1c4a0bcf51e42077c0251ebd88ed857800f450e87d257cc71b5de87602210b5fcc0ddc7ec52e23a9b3e69b4708dbd7e04f3e77f9db68d438d9c87819d64c4b79e9630f1a610c9fa90047594d5cb1bba32a4084d5283dbaf385a3eb859f865153c952e4139a821007535b34c39884276c156f89c6127f5bc42debc7303a8a83f24a6397543134a94b4157a789044c3a6f7ed5abdfae536ccb54dbf2ef174e41df41c0c08697bc821e298d49c43ba8a03cf5b11c50901e66cd7570cb3f3935fcf6dc7bba913df8e4683c76c2b3a3d3c3bb23b7d39a14c4479a6f75ca4a98b26b3b6b9ea5e58a5c8af5a8c3383f43c876d76bec69b46f043b16b5c685c3a3b43e8ae67daeda87392e95b7da109d39b5de0b7c6ef11d1e7ad3562fe9098a1075953bbbb9e6cef1c85fc56027d14f8f7fe01531aec403955d3b33040003bd491f985a7375a398321c82432fa93697f5a1c81bb410e875f36bcd977b118617297cdef9691b1e985b05b1f14e9b514dc7a3d4775afd677ebd920675d506216ec889c0cae861cb66a718e58191fe8a2cde1b0583354c7a5f879fe7c2bc5530a0a30c595387edb40112a5d54b66eff55be49af981dcf5d448617cc7c38eda3b130bdcf6d312251e8d2c7f6bab3726f62c7577ef55cfd033304072417e1901d2b5706b003a97a62e282e352b6a113a41db46e72a25b4ea6f8dacfcbc0054efdb7a81c314c8c40133a097261057a47e2474cc7c4740a27db17fb5d71ba7c4e518712292636947b63d9ebd2c8c6f52d2d27bae22e24729b7d5c45cf7fef8b38f736ffea7f7a72ab6a866a70e3674364640228f617a698dcafa0512814b27646ac49c22fe0f983cc3a06339f507369c3e786a0cdc83bcb8eef9905304859b7cc51b464b219f0901c766e47db873c8cec0e7dab3859a4fdcf4d3fce45170ace85dadc6dff00d8cdb0c84153fd4a0076287662a3b6562d673cedface35287a99fbc4d1dc8ad516c72867ab8fa98c31ed196374525f1e89bf9244cfe81a64a4fd1230859f0931e090088a61482820fc55c04c0100681e5e9c87949230ec02d90198bd73891a7f71944e19500c7d007849378117dd90c735d83b66bc95408172a7ad612007a9b8d81181ecc2da2f28beedd4572f884e1a397981e33a6feb10c4551adfa23f254f4c8f2f85583e1c417cb7328b7dd7d86f7bf8a100cb137cc61c207163636c9ea3b351f6acb3a12a6d29a0725d74a7c28d6996be1066d26fe0742266cb4306e047607016f40dd59b062a9829f736628715a3fa45d130c6e69c0099c1f2ae62b45318783f35a2b443a3c18dc07098548c82bb761309dd0cb7fb051ff61307a6f04e84f73c4ed8907f5d5807cca1ea3cd71bf12f882f6cabd119619b71029efcc2c9f62d15dad98841cbdbaefa76831e3dc0221b09e0f653f38a7eabb1e0d49c5d107d21df67e5b4738dee0188efcc7a8b5a012247768fe8a6e13b130f42ddf4badf3f0742b5d30535d8552fcfb6d1793ca582df985259d5c37a0e775e9c41ac09fa6bae2a95d0a8fbdfa6258d05390605ccf93d5e18784b5a4e40862531ad0111df85a2397c32cc68116cfa922b12d616075aa5dcc52c054c97dcb51dc57567e3295a5fdb220382199a3f7adcff9ca33f4b40a530a3accc3a7628ca0e0d37620686e9823efa2034aabc63261e6da74f03ddb98f75740a42816288d4721d1dc18f1ac56d79f623ec2d5938725feb0d2b4350957ef76ee8d175aa8272f97d6c7e56597c7fd167c5c7d2e3cd3195f2a06390ffaf090a3db5db6026553b06292beffd9e016ffd090d78356a90a578517966889e4b142342841843b9b281ebec7cd71f47fb622d8ac4ac11f8a762f79c37edb997d666208e85cedcfed328d4858c4e1ff458d82b546a818e9ecebf756c11bf19da0bcc35330d7a13f815c36c782cb2f6b342d3fa7283d1a5a08f538eb7257051666056582e1c6bb2e2ac5572c2b156a17833797a21ea58cb80063706da2c14e461e39e21ba94f80df3a7b46020acb2f2e719c438c6810a23126586e45338b21b1d87f7ee41e9c29114b5aed1517376662fb89854098cd49c05ad1d5d794f5151d506538f8c339183910a55ee4ec8850209d9dbdcf8ec96e95ca0e059119d98af0e5c484892a8b1b3b22f85fca302e63d26530630fbfdfc81199958faabe04b84578474de8228dd44145da0a4d94099f3cead7175ff52f1f7ceed51d83f89d91ad854363465ba11cb5d52011bb9fd7690ef7e318643b466767b6197dcc6ac32d19945dcbc2b5888a05d2ce2182daf69e238e628da28400338221f59d5deeeda997d8db18e2896b36942cf207f0429869c37310ac5bf504c64315a1e43b692ad6cbf622fe4b82028b73930116ffc99f8641f8b305eef79d23ea0c7b46418e49aaec5386ad015e48162e0e28608bac3cec9b90c8e5c7d35bc1c9345f723645083e05fef15b00f81d071d23cad5baee5ec4673f62ca30eed6e1c0393d6f9d0fb537eaa768722039075939551c3f847110dc0a454095c84f06878dda908b892b4b927ed6da380a9b27c65b92dc9b4e44a49b91128df28c6912db59703a6b3a852bc98af2b75755b026d559972b5fbf768205133c33116278ff3612f84e7f3b1f581d8578eec06baec896f4abdb9de3f0e34efec0ade91cd56b3cad2aa95dda7a7dc0173730a8ff0dc0cb8bef4b759e8a115cc01a3702a6e724464c203a6bee7b7a95373a9ee4032ef93586992ef1ac62c63ad98e8bb2a87943704f16b5dcd77c5016df179213202b46284bce2330fdb4ade72b07628aad689f14e165720d09705b2ce8750a24f7519baf8290ab81882f521bac070d5398215e04c5190e1a944a255331528e25a87873b9c9958bfa3c61ab53707f0dfc3545d4a9d83bbe24479f989b75d7b83b4742fed89ec6950f91038efc8e0377440c04be15e57879ae80db9fcc167ce9059c4fd217e5b6183a3fbd24de6ae2e98dea4765d5f399d0b5e43d2186fda925d571da0ebee325fd14b802d3d5a2dad1ced4091600f8e2b9f748f499fe84b1cc148ae9cb4efa1675102f8ff79f529966cde4005c5b41c3c0b3ec172d3611f90a7f3e07d35fa5a706f727cc5ef57ad77ce7d223539282df7b3ca9bebdf296acdf82b7a656dfa30eef0502d6573986660cea1711cb6c72a5e0e17c7689e091659217bc04d75eda9c759bb6df3e129a63c293dc427b506e9e2ac696e469b047c89dd3e442725a1c64de663410615087136561ba4d81d95a196f1e37cc62d73a6c6c0ca7faee72774d9a922132d181690baa9e09308ed7edca79cb6fd13cdf6fa742f645ea69193734abad8c2af8a57b6027cffaf422a17478f0a04a03fcb440fd12de003ac96;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hcf7b0e223406bc1760ed03ab14194a905955f0e3a13bd3436866a5acf10663e1358e764588c83f5b42f468fec15b99b20380da077160b50fe3ba5d09a133f4f2f2dc1993140d986b3a152f90a3f407f3d32787bb00847f957c3fabaa6c12aa47e5aa38e4ba9018779b2bf36243d214846e946a00181dd1b9476adcffbc4e6947eec9ce632e7d869b2d9e277086abb9a4298adadcfa4a7775641e3390e69a3e87836c2eef861b9269f1f9d37e1da0d27216976843dd5c09c46c2bcb7eb8ff617bebba782a715e14d946e00296830e20ba362154c1fcc9047139d5ec0243dcb77058165bfc52f17b196713191752d772f7b41a33490c70aa6f2f3abecd23d87525ebdca3fdd95e56dd08e5d56373dac6d2dfc15b06c3aed02aa59171aade240a0c7f1eb4b062d0d85d52c583df02619593250be635279e1873ac28e0e7c230cc189101d4c542c89bdeef49deeea0cdd451d49602c4cc77b72b1f6e51febbc9725b03e7a74359adc7239aff62fb154f6a1695c5293bd34fa2cd7d6851238066ef2ad8cc99272b685514b3b73a24b4c0a89818cf7b9f910f4430154f971205e7d3ef4b1a8603a9215d96736bd75b5e988f6f5259a527b3e157ccd3f8e88f590733162670e3017f87bc5123911e83cf3a2d34796067a225560789f73d68deeddafa72cd66264c0426a2f1243eb021a1a2ad06581541eb16e5dbace618266fb947d5c81d8d81cdff32233f4d85448942c8e234e688bd0e750cbc1477cd925d5dbc07c264cbec55ea08d67dbe53bce8b37153499adf8f195ce319870e3373c9970aca81425c3e6339f5d42ffa59168458b37b784ab35fa8d26441ad910d049f8a8d4bb88b45035ede07e27b1998527a59794f91420f28a02e16233cc28bc03b6a98f7653ae5415f79c856764df3b991d29c2caefe3d0d5d71573ccddeb9a6ab55f4f457b9620ff292e7164fe440e28564b457261265901ff4083e6eaa244b5b56818115153924461bfd969babc3459374096dd4b77e6ad0409157c4a8ec3fe4045a241cc90ba1f6ccfde4883c846849dd5cb947fa2f1ecfb0d02582e0a834cc77a40bb8c93f58d1b9cc521ee2e3a3929e18b652d4886befba4a279dbb6cbfce3b2c9fdc6e31090ae598556a3280cad7f33af220b459898e90121d747312a639d003203bb176dccd8ad3d1a6d49cdd0e71145731c202beb7680f7b021ec3d40cae6662131216043dfdc6c799648deba26479b75f60eb6daf521036b3f612f70a997b7c2a15596e2452992d51d070ec37844265e0421a882c0cee4a9d341bcb7518151e18e4e0c1b0c0f364001923681d75d3198e331a1e0e706b6d48dc6b4a2eb35d763454e9e635e60b550c285359d2f172b269eed41a8357c80fe2bf40a3c534fc19d57d6686c1993afad8a7e3d66d2e0b2f0cee024c28bf06fb675de3bbd466b17cfd100a223fda5400909b5811fe373cf49c8f5f79fe08aed9faf7f66f39c2e4bffcc1ca58ebe3a5b9e1472b4a48b91c894ff734f5c5471b881cb5a053902f823418af961d92904e3aa620588f28ca4fc9185a276c59aeb9086ccf8a98c03d7503e4cec213b7785a65b7e32c73eace85a6ef7dcc757d2d241ef708c8693eac4c86d285bd3af487f6ec1af204102d01d04c591b8e744dc0cdbc30a7352514007e2230893a8b079a43d65a5d62f22f482152e8a84a6e14a4c4312b7eb348d6aac554f1cf9efd94e16a064f425efe82a32a78b7b4f9359a1bc504b99bdcd4b89000826d3e6e1e7e435b244ab315e1a0cfff3a4948f30161806557eb36d2eddd69502fab658d0e34f2f8a93847608f095e164958346ccd98c56e7305fd45f7d8a428dc081a95406447517860a26aa27f2f448459b9ea93c328e1bcb20f882384e3aae42285473e4f7768d086eeb5efeeafbad8f3c46170913ca8735d305c40cea604e9a9da9401db624fb8823f06d657cf2ccb8aeab5fecd15f889c0426bc3a5170d8db06ba7c8375a04513c8dc898b5e872f9a51658652cc916449434bc5aced92d93aa888753d05e49577e11c6e38b3f8aef562dee3fe7c9774aa6140e39b118e390ad9d235f3bec2b0b542b453d8104b137dec95ccc52716cd029c235113c26d2efa208ce156da15fa9277622e85343a569534bea2fd40b1d5c355c0879283be00bfe7efd160faa8d2da02d390e0c25371cb9d15b1c562ff53088809da3d5f07c66de81a7a0fd4a0f9508c6019ee5d896471904d781f680cc0664f9a75699987ec4a8b25fb60c893190ddfe7c274cac324d6c1cebf06cacd22395fb8e986080a39aedc0f18aca988515e35676713ce192b265576a58dbcb07dd5766db791ca4f47da9e5e5e02b4cf19ce9e7820ea39d68cc8cca3fa1d660de52948e0d83d4c595e06a82328f5dd7a3437a3152a89353e0a62fc58b092e91f0d77efabe8de9aa269e4d9e46a421f5987a786431e949352660cc7f96ba486e38aec5030f8aef2ec6dc83a7ece5a4233c8e9df93c723bbd984349c925beef5790e42414272538abc3d39dcf8331aa325a5829e397047e3a26e732a4b0e8e36027e7c2baa65874f70099384598793b9d22ff5ecb22ce4b5593d3cbd1ce6df87990bd8f1b1b8d369319e6db742cb29e2b55ecdc36a850f83a5ad3e0a112c00941c49166db5d893fa3d337ed921b5ad492a4c77adaa85d37b835041905cac1664372d7bfa1afc2f1138cf78d3e00972700eaf77740f9fa5b16ac3c20504a87f2d144d6f4a330afe3d04327136bf856513776dece638315aa020fe3e18f6dcf67fc8b12b9dd37ba4a0b8c48e5d24312c9ca661d044e40536072c54a4e1875d69d56a5c27efdcdba338c772d3f40ff3f8373228ff065f2ef46f9b13f25673949dcf0bdf5c819c60572bd808aa0a4619460164698cf0bc05d7d4d75fccb8060d248d24390d67ba15425cdbd3fa653f08666d56b0af3730a5bbe08510d768ea7f996871f64ef936378812909e9abf503f73081e3435b30379423fb0159085f72df49121fb1483a7d94f1b8f24ad2a1ef0354a296e67644be450ea410234b78301f76ca1d1ea1df41346fd3fc0d20d015ded15de8180acfd3b76b4cc5a193b38ca5b6aa6b35854e27ab6f1c3c0af87663bd46263ce2d83444ae2110e2c76e42e12d037c7359f81fd1bdabcaa5d5d76df551a98744c88cab51fc6d9928ebc4af2286c23417791eb20aa648e4f719be9285f8fb93947a706c8047d8a62658975aafa2f972a9adabcee842ddd342625c6c36b937722361f1eb1691d76bcf41a2a617ad706c30fc63e89fe151dd95266631566fa31909c06f3484160bfbc95be6915aa70f4481ff70d2cc0543d05efa942d0d6ddda42872056228bd4314e050707871b6677a4e695dab2aa8a36d665e39e242e5512dbfa6f4f0ebcffb34885b1ceab6a58a790eeb003a8f69b4fa932541d7f0e092af3dea8d7032c170560015eb4bcd31cf1011c6e043f72ec118b75b313c2c855646ab733935086d58195a13fc092977bc28344021fbb119c8abf9b374acf3a357e004aeece4d54bff1f3bd1198891473dda708b9de55d482fd17570f6f960009b0ebe800c609202976c0c7818d4a9ba896ebee0fc9c7e227de70a9df3696e5bf4001af78dde7089388638952c5bbdf2b7a01f2872d313187b1cd12e27480d08676644118dfb1fb7fee71ee0ae0e8de324881df447f0a7c5c2714be4c4383a6ac633a0427780121c02e546fda7f42e05768bc96eccd543cc84f87a3775f84bc9cf945971303d63ba1dc4648f25a9d4db3cdba889fa99b6af0b9ba2fce4c49c8f1aa139c285f200d225601b2074d14642d9db4dd7fe0ec778fd91a5a68672b03c7b6341b8199ec3143f6f6495d6e6b7b47d0be81332de910dc88bcf2b3c1507621a4c8c7c9116f0b2551651a235d5642ec851322757f7781d294c2ab43736480c5f43177eac1375713fea0fab6c4520ae9540ed03cbbcbb68bea73b90bf1f988be44d9ace9d11bab1b5fd7194445ca56f0e1dc6fb82cd12bbcfbcbe1824e62d2ca16eb1ad52cc330554483d33762f09c05000afccd5f3f91e293f09a55066668d915764aff7d2de0f74b9d195a95452ea70966ac0e23d6f2fae1a879a28c545469fc0ae413d1ddf5da80c5e2064408191673bec85a1df05c5e96723c95a3161712a11b5a35e011e0780efeb9a5eaa01985612668d0bd61df531a8b1a084b60e7ab3b5e8d65ab61650a6220ecd2b555e47c1ea78dab76fa7a24685df5b4a2edb59b6407d887ea1a8e236b211c48ca1a24837da1fea0363a44654860459a65ee827eec71c86daaa2c0f44fd92fa12d9e813e207497976a8ba6a1b3f883d6fa103d07c99a8ed38b73fb61654a1518d348dc065a0d9c36e08ac9839e710382fc0fb3117e5b3a5a3b906208b0a6ad951c27afb0da7275cfd2aa3daaa0a01c736d006f488b0e6f41a188d4a54fa971e9063cd50ebfc3698116fd72ff9b4aa1e87dc368174103f3d0aba6b7b7f6fd24617beda0c4bb05e2a82591a0f99f3e9b9b80bed9d8c44b37f3a6a8b67893fc13e64bff7c750099db44ea9d682a2c6a233c2473d962221be80809f92238366822081ffcc1da9b286fa55273e596a0fa349f940649de319f7acee963f269ae09a86b13bdb994a5569d954403fc83d1a5397b7db22de4816b3fdd4e9970a26ab15316e6e7ecd8d3ab3966aebe8eb15f67596b75eb7e24146a9aafc6f3bc17e030833c8b14a4f7c2ff44aa065498b3c5eeadd94734bdd5d294dae43caa95ecbfa49df62582dcce2f455b077fa72984259335ade596fdeaa879a8e268b64ef02ffb576dbb50215b62711b79c60b228821640da5f025b4beb278a4b0c522c638cd1c7c45a1819f8883456e1fd267e37fd1079c2ff26a543ae4cffe71c6315416cc80386cc298080e43a09701d05a96f16d3cbdbea6641c10635e7ed07954da9fab60be60eca7f480f2d75be0dc2c51e5856edfb45922e6dd32006c98998c7c15b1dc1dc37f3f76801aac37a1e8e51ac0b270565b6b54325aaad1f3de724e8d6a558d87b399de038ec01fb20a75f0b8240d9ca7fe3f75473acd2819fe0da59e392f72145be7f611e37e6c93095a90abfd6ce883b3eb03448ea6d71dc51774ff8c8e9640cd6f8f9ad33822b9e2ef92592d1eb395bd436ca415d8a81d97495b6c82c5237685097b2015ff2cc2a5381b95adbea9abee30b6826b170a2e404aaab49cb827d0441bd91e1b00e48b2a1b4df8beb43c178070c456e905c9c7a12f29a5893a67c9b8a3b51dc09a41babac3d01a3596d45e597a6b0a0e1b9444cc4e3f0a56ffe8b8b349d505c0b922a002a5cc076e3d8250c6211890dd718beaca0e0894fd554029cfb033b45cef62bc3a4b5ceb396bace558e70aa3fb5f9f727fe7f9c27c8f4eba8263943ac6d5ae05c5cf4d1bbc5cd3865fc1341f5ee97393d7e24d2a99accf5983a394084987d9c737ec7aabb59d320d8890806e906bbacecc5009b306a0c14ad4f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h5cdc2c5ebab2a90bb5a66e5620723500602736f8625561084732d2f222630441ceab2fd2b8032a77f3b9479ebeaa49d7aef32cf03b19dda714a1fb59d4027f067da6618a22bf6fd83d18f69a51e85c08557017892ee43b0c979f8ca1efbcf8f203f6389e4016d60499fea909dc58c1292a4d72c95cad74b4789bbcac98cc46a161567ba645831085ab9fce7410cb95e44a87693b85b97d087313d02db44cc8458afb1e19f89e9eeb47da2e3e1bdd0006f93576ac64ecbb1045bd7f885cb14d2e39a5d430d55ddb2631df56ba200b643da33ab66da8ad0ddb628533c3d3032483293b9498c9e0e42c024c04eb4fec6c7f372b4fa280db81087d362fb1976f3753e89110482ca178137ba6049dffee60700d6ad3e07b38795532d75fd3cfae087b95e26b4893ba81fde8ecda039e8625d9f221b48b57da83f564ab660f1c63e7b971bb46ccdec15c9ef582e594ec17dae3b9bf85d40d30e1ddfe8d8416309732d58df093a0206c49f1a210835316a346261e3abcc8013e4f60f740a50cf95d94ef8a398fa58cf52cb52cbaa1c1e98165e668dcfb421db425b63984c0d69f182b949379708d7fc2090dbe6cb72b518dd4cda031a5680f79f830ba3d98cef53a48cdd61c0705f1c3410aaae79b07de52b582c342c98523a944c591db2afd06f5a4f53a220da0146c864e58e8cd205c458829ec7a0909a9c27577b9844440e99428661fcee277173c86839a15c1818ca1c30f722db98d55826eb58ee9c299d4e7d43678a0cb8c14fa7f041b3d0ce779274d0d52e74e806c778fe165f94ce547aa39616b6bbf5da466a0499aa6fb66ea0180a4cfbf6ee6d79d34976f8045e1357522d2231a3374ecca64cfe8f5f48265c9eafff026d97d8899c1cb9e36536ddbcb7aa06cd00ab48595263705b4550314bc1a23f13b4ff74ea3886a945579bc5475474217b8f1e1c449247475cf00b27af58cf9ade113dc7d3be5889068e23cc8f34717e70ac41006d164d2d2179135fecff7a83bf8f71c943a72c9f85fefb8a8fd1b76ada68a83df3e552544043e8747bb84f2fbaf54acd5a59c3eac84d9cf8d7549fcb07e14f16427cd6467c095b15c4a39d508bb98fac9a426279d63b661ff4dddba65aeeb0fad7c865bb2c34b4343127fd97b1c3e0f878c5c987afb969466eb7d34415aa6b3783d669c7bef516e7b65223e8a26d8719c2057102d923c35d457923b7e998fe37a5a7d061796d9a005b77d2e77792d095b5a099d0b0d13392c0183ff0f4161df5df4416077d40a838a64e636bf317cb3ef54991c61b266684d8d3c5caff7351842c670da3f8777e42f9a3a15552bd6b0e75f94e7ea52924a4975b0f084ea3fa16b804283843463e361bd9e6fad341818bc42c263a3e6f14c211893cf9d3c5cc183d5103ad234e6b613928b8449116dcb3a890367445d4dd4116f3829130f4c01d56d4eb0edb0fc0b85a926aeec280b0bad5da4738cd0d9d7f492b1904106107babb887bfc7385bbe69b3d4810d0c2dfbcfcc8a59eead545009199f25bfeb02adda7dc407d0eb1a8599b5fd6e06aec23066d3197455b1752987687ca5399a2f3484a63b2f857dae9c02f9db9517b88598414b57495f5c128658279f7b72277738dae3b5dee18ea45a612b8a82cbdf9b68cff892f88ca1376dd9863ed7637cedcc6582fe125f813af29cdb69fbcedac576b84a365b4a23f8a004d25a350dede51936133f92bff7ab53386641b3fc7cabadd78ad4f8de8785ac4559fea69ae947ae61992856ff71e1b9f8546ccb2176c2066b840fdffb12fd07aeb53390c5efd495eb175ae049e9c70315acfc4e82af44af89843873096bf89b8259b1e3f663b25c785c17cbe25598a6d8326146d9e8044ca4aaa4e8a08fd70899526fa19b5abdc6bbefa97a1e4e770364ad1893c2e2f7f2b7c161117fbaeb72b21eddf630f45e5578d019ee5bc03f292dee91788e3b563f99962f2c99ed204982e58410660da239789cc36dc714589b701b9e89b506b88351e1b87d976854df6ba79e5a5a965d58a22f902f0edce0525cb375f757fe071a09d1fc6acb87e6faf28a5c837525a5555329c0738da5fa8fa56d3fd3030ad8ddcd99e4d97b88f893b26079f99015423970ac7395a516046818b16bc88fe85569f59724c8809ee8f5d419649dfe04c376306397e392bd1a87c81c193afb67da9cb86905485cc8bf26b9316b546ce7ce14bcc930be269c2b11522e4dd0f20097254414f504552ce10de21f563994131a54a8e875ff6eec33e6f8413701d9a0c917e4b9787ea8a369dcb8830d666a63c761abc13d6d661c1a570d4664230b2f7f8403dae09bd3ba3ab569370915eeab58651e872d57fcfe380dc64551fd0f7310afa9df59a07bfa63714fd013719798c2c869f83f0026b0b3875847f36bcdc0a1e1a8c691a048186cf842760852441fbf0da2722e956b36411e4a1157093126c39c825889f8d8b384271b2866fbeb99169a49ec672835443b98876e89f569b4ef7ef38e5327223a448c772ef490a9658d579bafc0e9fc253fdfd725d3f842f478b516d0473b1dd03990b8a291a43d7026e8e1114ca5e07284f9baa0f250b5487b2b8dd3678cf85f29ee30ef5aa490dbfb15b911d3ba6339964055cb5dd0211c082f6189180fce6c3e21687362093cd66b6fb0e6364d361a23de93ef1bf5b9038ead7581a0465191d135e0f15009862b64209fa91a30e46b910fde51179c6e09a69872f558dad1e2c0ca316b7bb7d9aaca6bea6bb7819530c5a057122158a63fd739ca00096be30fdf0ad210273168406a18fcf3ab734c3e4412e39723f4d366dbcc1be6d4a357692ae26f0f456fa825feb718efc0e05a010150274c5d21113ac725d50de1d950ce5d256bf23b7848caee4c1460d6d2c7338a4fa9e89614ad0aad8c5129974ca63626ff30c190dfe20287f73f809bcd77071046d4b942a3f5468a74607b7818d0139010cbd936c911b70f2ce2054be15568e7926ec7fa5d344112096edc1645becfe7de6dc8de8db31b4851ee10c14c1a3da7e98a2b95c364d4cbd8dfe0d7540406f5afb5e4966d1f9699b2a84927bbb5069e5073f50bb76f3cab3be5e19ab5f09a9e1ae05877e7c9d8d888c4764bdeed86eb0856257d1ee44a838deff27ed46f1ae264512c69a95d8407f6b14077fc335e41464781ff29794af3b66c7bb4151d58aed08c851f0b795f32706069500cfc84452487ea0084b54ca0016e4d061ae0749bf741ab78c62d628f0d20703899b10b95e08ed2a48f17ff1afeb6f39a395c2509402bb28db44dc0f8a509ebd2252b4e2ddd4339829b598ed67cf8d07c2b29eb9c8306d27862db870b20f57f679fed311890fda5a7f6bf90ad5ac7d26d2bcf087790a29c23aaa3f7026a843b7371bf44751984971084775eb918ff656366ce6d0d697361b0d09cb2dde23b71bdef750ccb5a641cd63b494a91673d2aa1f408ca543c6f103a43d52ba0818f7181d249fdd750fb295c67436d215a0b3cef0ab6ee6f69d8a068b7f2f82e1d54c7245c23dc96c738bda421196cb0abcffec7464de02241442f228fd089b2381789e9e32ec0d664430e5993b9ed4f0ef4c20007c097aa670ed591f225408314133e0691db783543fc3a36a5a0d966d2bcee76bbe002384cd7d8bb62c271c980e28a6d565b37bb35fc0c9f535bb899d583da10a646aa4c538d58583800d1e0ef8a81a55c5f3113b56211dc593066eca170dd045447584e897d18d2c1cd863c1b359c00314fcecb6617e84fed1f57612de2ec98d702bbb346639923c069ccaba776734314646e7b6e2a1e36ad66dfd561f5763f14f6f9823fd5eba41205e68f3d60dc7df137c0a95a775791e1ecc0c6bc9bc5dbc5c8471e736f05ca89bc1a59dcf1785ba98c271d07b3d5946c4672df9f93783f647648b21793193f2f8b42d676594a7422206b88baffb59be94bde13b4c8e61b5fa22508840eb221bc94b42187b199d6a9fe199043b6566e82a6844cb8bca93920bb3dfee54e2bd58e8e0266f10166779838afc73087b19c1a0ee474288b13aa36f98c8060893080d1726f2011fe81275a8294cab9c82ad28b9da285c4e26b5d4c9b2f9f09f54aa260e7ee3bec803d1b795457088df3f4c74dc82809f671d4bf74937ebd787feb209d798439934940507c900d208568b82a66fc3cc08195c6e6521bff0edd5cf0ed79eb3c5495557f6278be4f178721359fb09890b5ccf96cd81f03bc2fd4b9a7086c9d3e8053f58f49f3279109a019031739a0f303fe681eaa885e38f8dbb0cdb94cada6a1d71048bdec847c97b25b4119f35490ace4e4a3196cc9a3393349f3ff6213b10e612d7e6f3e54967c0e5a050dc327cfecf929e652076294bfe145b78c53619d43a82b64d56f3210a13af6625cd4f520197c3eb629880735fcabf1d3139c3eb03910ea259f638626342b2ae0467bcf42c58f17a822a07699f6e681ae4951f035020abe707f0fdd739a4b0201d5a73bf074c3ccd363f25c28dfe60e86ca346b6fb768898e68b0a717551bfba72b207afd304282dcfdc006d91e97a9893fd33fe611328ec0b4f476c1e8bfd2de5d083ef6611fd1ecff586747b2e49a24150c7b04e96feefe35017f3cf1def147d9f3a2eecd681981adee014f91c4c99806db53dc7addaeba92792dc64bb78d91b37976502965df72eb896042bf2b2dab85ba00a64f37f762e83d8552b71e10817833d2818ffacfbeb5eb70423fcda910b1131afc4baaf0915a26baea8fb9d3546c5f3ddfbefd59ca6210e272e25c9f931519ea43b4a95c67a6795420498d2b26c33c4c329f640e6114c0270697e7edd445dd506a6abff6503d6e83b066f8151dce8d9aaa518c9f75ce8e9d7edc19539a011544e62aae4fb895e833fda18b837995cceb42e291a6c1efb3b4b1170f56f21c3de008595506252521c931743d082df46c362d1546735447e7bf288717db354ecbd0aaab5abb8b28e298e5b254d3ce532bbc0e68c83ce97b584d6c93eb79e9b625857b86020959d9f21708770b6e278b010e0b32c6562a31f1a0b6a543079e2f6b0fbe31f5a5bfb1a5fab42ec80772eb20aa509b7bd797e258beebf276496f3a895b122e8cf68b310371f381879950f422ecf3ac7703b3b6daa87f5deeab45deee269aaaf63b23e8a5fc86ddc76abf63dda797879565b812adbcc694538362dcf7564a663cf947d7ebbf8ac043300ef1eeeef615ad4a0168100d8919f08f0ea6df491ec3d8a5ac00c087856d6f7713154dcaab30b06a59a98ed76959e553ea0253253795f75cca23a07826417bf22d76872eb9f47ca0edde6e30fc11741c15424db970bded20d336ceb8e0010aec5e1d7cd4325f46148e64347ae28480059c7f534568d74edf120560a0defef4792b32700a89e9890f694955fa1c56ce80e9f11a66fa2cf5f4a1991ef36235b78558d4855af97621632a884cb3c2290b79b989d0f1c2c273f62e05aa8f3f5a8f6b0fda6b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hd2777b8105a4c77756c2de12a7c58ee8bca137315eb02dfd451cccc143685ee4c87286afe005ce1897a7d1b65df960a2f51178d49b58761c0e726637087a69dc77bc4f42e92ddc137df9f349176bbb144a7c3652b5bfd3b060d8e00d7e7a907c96aa9dd150b5bab37e2e42356a42c6c06c2a2ee6104c76ebd8e3bf579fc63893c1e183ff3fe8bc9b48d979d7cb027fe4b7f37a6173b13b740f00e33b4fd70409cba115f9b075c6b5c6425a15c370fc296610d6b1196d2033b7840893bfd9655038380b4d18cf02d0e76c8bed0c13372b49fea2fc45d03c10ff15b66aba8a3e0c9bf64efbd873653b8da17a9f29d91b169ef3d838f48158dd97f987fe198e332c0e6339899ae2991df81739815f3f580e62018c40c56afc2353ca888f452e3b796491bdaa7cf436165e98f0ac578778a3968ad1b6990470fa5e5c8cc8507b8fc4008b74974141eb9204a6eda1bcb355079f1d073fd0cdabcb30c6378460cd1d0e81f9418b9e9ccebf0509c69e773e7560c9cbc1a2c088050a0f1e897791750d952697047f74139204b917ddb345b0d0e9f918649c8fef2cc182a8532ce506c5c93d1506013178f0b1927d25deb0387d9998c6e04bac11b1aafb94ea098ec8bb9fa6c9a7d238e1dec7babe50b1fb63200d1a213aecba7460105abf64e58e1d50dabbc0f86258b4a2f8c8a2d2ff7177b0a40f19353f32078b061285b44b8c2c6ce30bbf96b1bb0848f45454bf90cb8607efae1d15aa57a4c5ca9821ebd2a4e9b0d3006735bf26b09349ddc272da69134d52bac6a052b67d49fe1fc22785960ad895afa9d4ffe880793bea8180bf5d97c035ad80bca34161f857ee89d71a60e4bdfdd1aa5ec41ce9723d7e466a083f4bfc5e4674b168ae8309c2fb53245dc9906dbb57ec997b0150137cdfdf1178fbe9b7ff3ff711af6e74c1ff90a643a96e093f7185abeda671e58493ff957068c55387f036f475b978083874d922021f7912a3fc217e968cf06503bc4a68420d4b705c3e4ebe63ee327b4464e86ae2126a2896f9b924bd7f2ee38d5df241bcedeae1154130cf078d11adcc77c31b7b966fdf674b75bd57dc2244c7146db0b3667c304d775e0cdd8dcf8010a124763de405abe41f07b586382ef9fb2fa62e59952e4c6fca7dadf52d29b8ef081e392499fe05f716ac1411963806fd69bed2fa26f1558d49b1564e2f6e26c458afe213024048b8ec324a09cdf5ef993e57ce5dde67cf366445552a150c80cab91c1677ed24a7cae8a7009381e06e8cf98606347a762f8590debdc27231d49da12465c2babe4f44c34f8b8763f0010c2434c0a46797188a86eafe34c054537c163a5397bfb9a159a21795ac7e68a6b69b99a1233daed3a5aeed1e78536da2ba3c1d556012b34e6b8d3afedf39e95306b71b7196114126b88c71dff30aa6266a6ace8c49bf3b423719543232e80219f547e253f9ffc667514b296c3314ddb33048eb69c0cb4068b3d1bce877298776f123c1c2d0f76592cc051102bf7fdfe2c76bd93fe93f0ba7e0e2739354ae26c7d2ac84e6ce9c72a64beeeb3d9c92ececb6749c4ee367069e63a5bf791f4584352371dfc66e02cb26441b26b0ed2038eddb88442945fdf0b0534193399afe7cb70f694efdfead068b6f840eea1447e5589c3406bc2894f59ade21bed55ae98078b98088eb11d137b615e17f114781f67a71f299064fa91078c1750ef1e0a9b15c0a999c519b2ae7b1d49eb7bf6b4e6bcbe708451c39a00ffc2ef4b4902da85c5ac836e6f276fbd88cb5cbfb60606553fdd7e6c50dd2eada5f4157663f579604f7a9c730c3e48c6f5e397aa5d653993135d27d41bf75e025ddcd839ab792a08bb090989f9c8b269ad0d29382dcbab59a961c06ba9857e025f32c66f5bb0514ce77339dc6377e659d93021c7c5226e2d56713adac3f4a4b89787f17edac91e1563a719435df4a75849b38990c06c866f187cd4f3917f76558fc5c58a787ca618d00908b5f3fc42f937c0b97cef62a472d3be967e7d72238de7e3154272e2500fed1b4c11553ba45d79e18dbfc90bea96359ed8e617b768a8cb2cfc629daa74f91e8bb60c1ac8085296aa8e8d41caa178f784bb92ab3aab894a7359b4f3dbfb8ad8fcbe1e1918dc6bd6e34082ecb359375731cb66d9779b09bc3663a95dbb86b0fe0e3092735bf3936a92372ac8f5d4668d98bd1b1ee99dcfb5daab8a6907e2deade978e7040962874feb75201f2351ae155641b96923aa5143578c9727c8f2b2fc11d0e3c3a87001e0c1a610a6e3d97d2aca8dc3494776790f121308704b7132529a1634b70a05b6a4f9cebb65f345ce4e7f17742e4308113cddd6714451444f57fd569e33e2da2a0cba9f3d0cce926743f8401a70084f0d243d3086c990bb8136babde5643c19f970118003613acfc8069339e591f0b9d70583fea60e090fd6945b2fc7f35d180cee23055be91fe97d26e44de8d59098641406e2f83dc956826e5e2722204c635eb3ade0d62b37311815b90ad46862887adca22c8ba00137cfedcd298649850fbf0ba72b89dbe7515fb68bd6c0dcaa6815abd4d7742acede9210a89d4cdfe3e1f38533690825066c030f71d1e98bb0ef82743dc194c7e4a4e45c451f99c84f057ad36adbadcd1282712deb814c6764c448a13b5bb5ca7c448089540e5820d76ebd9850222913f49103716680abea66c0e03b57dd3153fdf2bdbae170b0f152bffd3c96764165bc0fd5178a840cb45cfd38839640d57d1361b999c9926ed6902c81bcb0364c23ba624bb5becc2fe7e83cb4ab840127f8ee3d17108bbe5e381e4d34dddc5cfb15859425e396553e538bec033327e51166649c68207d8e6bb79403dcd6e75e6ae5ad10da2e8c101b7f41e68dfc20efb53d54c99dd95e725313f85f2d6f53be32298fafb1035d5864fbcc79342bae466ed42e55e568530563bcec92b8e69df69bdc097959275c1d1078132d18bba0293dc43ac5ef5cc5a34960352e683b0ef3fc5228db00062b62c5776189798124b3cb88a7660dc6b72a526e31885097141c5d9c43b813c3b8108d14b7b8e2abec18a09de5e3d3136fa9f1ec4ddafb66374721c865a14183f18240bea792ed1b8d85eee6c1986d4f2819eab325390ab7d11f46887a996f875cd536cce8a980e9fb523c0997f57a33dbc383047828de76513436f9c4d040dfdfcab0f0f287d4b0d5652df59c027599e3183a93c1eff1e96746439e7fb3c49ad555d51cb9ee7efa49f751756a53ddafc7f22376c4daf730e665561bef02ac11dbdd6db69e01c589a23c3b2a45cacf69b611ef03d5076157b1d644c964367c53c89b1cead5a2e21ee4a8ee2143c17a1cdb45f14b7f2f5d1519083f64a9a31dfa646648fa24109c7a7fe937614a465c10561ed1f93815fbd259905cece85ee77e900f53b45e18d77c9075f20791d3d125fde32c7a3a8900dc068e42d5056ce6f90745dd1b9784ca10b755aad1548c0bf700de86b1c3a879b50cbf01683e2e8bc7fcc5e5ef8c40699c068ec26c02d36d76ef3b6422a737f7320335ae503b46100fa1ae807f926ad23f12f880b62f307ffd6bf5c42a3bec722b95509406b33b80d7508eeaf50e5fa20eee1c7abe84bf04e306acb8446f8915986c2477b7a99ed704f4da3b42bdbc6dae1ced76956fa93ec6fbd33cdf537e5e84483da14a4b711ea290a4428145c04fbcd4959ae571548a620b1833163d3b355a6ccd68218d41166bb9bb7c266467c47478531dc9be41b0eb44413291e2c4d5b04763c76cae377766d0a451a6eac0fab9bed7c0c7c9ff16be89d89f41506320601a582e97f1933f3d378d3a804613a7fb4f245473d55994a3a2994d066acb6671b5195731a81ce485a558df33b557460e16045269a6284d45af148797c29abb7d0c1fa069fd0eda615225028a10308d6dead219b13cd8afce70b747d18bc9356adefc7d191f538eae5501ad0309b45d3f744f2be1bb6c1cac862d726026418a50441a7f9081338dd6a8c632620e7fdfd47626b57ea38a3298b21fb4a92653a21da73c49e9e60443d0b62c5e76dcb33fd2492a77cf31ce45f95edfba6256b9da3913eb8f7b49b1171d40e828d1f2947959a5f3269e0bea2cd43c587b9e02e5b774bbb12f365a97132df4dee2c3be505da7e1b3d46db4aa4a3ac73be364ce3b14d5e788c4c57589aa41e55268e7e90a0b9887a2bf64270f467964317a048daa0ff073f6fca411a0c5a9ab165b13f1c5f0f1204fb9bc411e893c21da8d4142b02b643dd4f35da7fb5c62a97d4215cbda7714bd4f4200c56d30de2f30e4df2a2f8a2f306bd9c13ed35c9ffa7a185d4c387b150b41a20b33b3a7018a3647a9bd3bc9d9bd80598f0d64d050623359cf86573e583c089e3b1efb36a8c0145f925c5fbfd6627348bfcc493fe1bb3f79df55e2b45106e6694e145b170751acdc668eadecdd99e8d1ae415fd72dad356b0693a8ce75ed59523a0b86286e5262c0a8413f88e318b1f498fbb666e7a77cc7176c5b03e82dbd17d7d549f5b2a0c98815b8a84696639c3f300cb83e9267b0b3e33e177346b0e14888455efc43971fa7b3923de77ecf0bcd5ba2defcbfb16b39c72a5be01ffe49b951090e58e3e4187c96c645fd0f8fd12563b4aa25da7591214097ee5512e927201bfa92f285734b37ab38d3873f535899df1bc29aff78608e1dd8cd0749215d86b9085527c2864b72a05f519925ffe8ed42dc805473865bf6b45ffd77a6a26b1c44635f275fe5dc0d1e14b88a700b634bfa526a2f2a427b5a9732664bc34f631138951d28e45c60b2ef2986cc4528f0da9d6615961a95e924cf18ccea145f15b55968985bbf84d84ddf6c9c3e39e5e19e65fe922471ae21227d0931e52d941fc771f5b04446af3e54de9b7fc9a9125f21daa520008664a96fa842ecdcda4da710c737b77eef9d33bd8d4e1639747c25778b12e227e18507ed66c657d9590bf01f15d941011056cb86c01f021f375e9d7376e0fccca098bb0079fec55d975efc50d8edfcb5d9041427f8f1f1b9097f423eafb61ef48dcb099c88315c2279bc6026620af088c5002f7bb06a540c5ac3b79df15a564ead3b281f81a46c47858d05acecac26f4431399c10324d03ef63835759fb56419e487eef4e9c6d951cb70d70794420708938427c200126b472116bee2eaff6604f6ac242b3027efec85069593029d66e825ccdca01c2ef8b54ddbed5c475bdd8d6b960e3f7fcb377f4b4a6a15b08733c1e68198eec54a07654513835e50ca9a1b9c6acc16a58507b9ab552157d7d6aff5c43549232cba4dadf02e762c026be3d105bb6f36d4d9a6e952e792ca2598808ee4fc53c91a46f9b9662b333c91b631c7547168ae400894366c3257d40ec503cd908825c82a300a3d4f0ee30e23801ab1affec5cc2bc86b07becdbba7ba7b3bd2ff953076c89a7bdbe1836c968bd39a40a562fd56024b2fbbb1c34420b92984958a426c03948619440eeb4cd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hc9227da0cbd2504cba52815a5c166aa71a138724557d0df2e98acee9cfe19bf19e95972d970fe0bea02ff35bccebb3b83478ee26728bd92df137f9e6234794a14f94dcf60fb4105c315501b1f0dcf7d418c3cb71975d7e8b63bc5037d4d7fbef143fb819e6c2d96a3f9398e0fa34b01442d1267011d4255a8292485b9c85898bdd469fee30094eb1067a3f51600dd4f4c9cb2bf07b4f0915c39dcf9b6577647852318830d7a4f814dc9522f8600517d580f495e0cccbe33c67d10f2d703b0134bda59b78ee3fc15dc7d871025cc6954134b102945035034c7264018a67c8ecb973f744b9073c638f69312f137c7c1acd09f69bce3ebd7c351587253aa56b594e03f6f12e18bc6c0f44094463c77a643e9463ee15bd57d03553723b0ff695299340b73c84a20b1f01a7a5cb62fcd41e8ac4206530c1fff6575ceedffcefb75e38f3f5e1cade6a9875b6585c8c7aeeefffcf54cfc03bc9710897d25c27d5623d3d192dca89f2209ebb0257a5224409a29ad22eff228adacd6dbb3b76b2cebd193e867122722f7dbf332d2187c861dca5fef0c8b996bd38f98e36ed5fb66ed1b0d6750cfc0d933284f560bbabbdb36f6ef408f4f5b9c8f65673c6d0967f81704d4115fc2fa6fbcc5515394d1ea4f39f1bdd5fbe6dc985a0f07d63db5bc33dba120d333241438119abcbb6b460fa804d9de4d459c4271deb2cd5d57c92c0574b7b6e79c14f8bb7a59c6edf739b722dbd712acc4619b68d150a51b5655e96a473b56f63189768b64b2ee9c59e540408445e2119674f9479d2efd0515fea2776f210c4ebbaefd28315cf31050f3a343e3e74fe87149fa83ad010e79f2387619aae01ad6b3bd28beb135fc7cf5d56459443337a50cb56da64892c21839abdd0b35e68532bf867bf1a969aafc3dfb1413d349ca0fb2e977e361d1e5419ed73f80bd816cfafd29f573227966ddfb035e663f5a2b3dd6e1c1f4150260b7702262de2286b60143f9a77ac89de0b01e3890658beeccc9138623cc4132ff7464fd03a1e9f17313e09c5e9f563bdde50362e11a7e609f2a79488e73a0581b2f257b78b5257bd60c0d163e904784ee041cf374b669901b49530da1fab1c2bad5f5de0217ab8d067205f6900ce995201915039a9044375988a08290219e1268e3b9c8e81910b7bd131812721e360494f5a621386ff1b4bf0dc7222878d2ea5e8e9f67a02d04cfdb231e691743ff4cdbdd0223ce1f882250b2165b893c3652a6fca9e9c582cf18089ea3117c0065028190c801de858a026c00844e340e340d2ec8de15c054bd78be546e9ef495dd0a6d8001f90d134e289d09fa6ba3913bbb440be0d972328b01495c926e7845042594eca1115e57f2c6b1a34cd5daead04a135f59186569b2ae988a1617334159428e2524629594cbe354569acf1a342339a65dc11a5707642a8ca80ca4347e1667a2182390b450807a82964cec39de5d7f94cfd585bc16f273794a275b834f46278f7b7ab9961ef81848f80850da88afafea1ea63f9cb2122d6090f365a9e6ebc2a147d0d29ea58b3985dc08234d0445fef58ccfbda761e5b61db92b9da7c417c218fc5bd488b42113b99d1271417547da509cee2d724e4ff7eb51f6ae2592f60d2a2687bf5426cdee7b70915bc327a95fbba85e8d61c5adbdb75bd348093bc0ce32cb03168dddafce6c823ed31032ef23b9216f979ca37861081a41d17702482ed472ec6ff75f99bf0a9dbce43dbf401db4e860649baf18a4da3e580e12020cb8201f566739a61f0932ed2766a13555036687c00d05fea9fe8fb69802448fd45ff3916ee76e2db73b4727a8da9928053a32f64f577c2b930f4a7c7f73ccd9e92aaed6c841466c3aa845ef25a83598143ee0408da0f50e916646e4586629bc01319bafbf2869c119fa2e20af2e802809ffcdc3489a4a58915a6f643bad3fa5189fb085746c3d05251be231635358f23970077655a919232450d3c668bf8bc67f896dcec7b8e4aed80854c8d0d6460c32ab183a3eedfad8b1fe758327dfb59393d7c8001e1a79314af2c036be355f36a43d7a1307562206c5486e76096a3b0b0e3c767d72f68a98a5ff0404e05a77eea6d44293d207b45ea7bcb9b57bd2e024c64a63700ad8c51057172edea35039301a77dba4e20a3f6a94b8daba6dbe03a84fc8d2dc5737947e7bb0868716f1e5f986dca6c952278ac448739f1b7960dadd9333eae818d9f6aee493fd7c7e681c011a133a199f9f8339030354a457b727e33bb9f5ef865f90dbbf14bf0937b1753f6f551f8ed3e23b138f9ffbb3a55d0e5319c08880b0e2923db783ec35dafc5b56f770b2a77708deedb889053f0358c803f9a1deed0da69332d22534b076d8a86e358f0a3f05e48c26c6de25cdd4d996ac0acddf717554f43d753f90a8471b9072e88adaf3b72d539d4013efbf5a35b135fc304e81a38191c15105a2ceab11d0269b72648228361565b030a99f8795113e4c41ad4aa72e8a3d475403d01457dc97e42f0f89ba7f1e12ad5d59edcb5c4f5c0cdb2059fcb470bd4a7aff8883df3a4ffd69c9e38f0aed7c443bd28fda5cafbca46ea29dc27ce3eaa8ddbf77a653292d8fa9e9c22eeaee57b129aac84ca6a7b0e79e1dbcab23c3cf464bac211628e41afdad5a7e29bf3a41997b9d9213bc4c709a980fb4e546d68755e4f65cd15d9881148ce3b723ade1b05c6f6951f8898487904d3a0ab5e9b41cb63888dd2b8b962607b4c51c957c710f260076d37e305c6539c4998230477d95f2385ba4b297d30d361123a95dd9b4ac1d2749c33e2e23b9f0fbc980f8c85d8511bfd828714aaec6e5a960a7e87d86a9cc7ab61ff73ec4766c81e9d94ab50b3105cde5c7c6bb134d8b6a0e88cc600a14f2dc07f01c5c8074c53a50f8a7a3a080d04e127f6d34d4d149ff780457b6f2053e7ec231e334dfa5029423ada9d635e9ac314c8d4fe4333e16a47ce286569ffe0d70492ccf24e1ca165ee56565fa9adac1489813579cdc4a576bbc5e6995c0ae216b976b6b8c32f2f4ee50d531acb9d9a35cbed67733a7915961df6f83788d6c34d70a971f36b6065d44bae3e05f5d30ac3fb73cc5a0419facc26a85fa370c0ccb32556162763a50c8294c0022110b82a2d230755c6cefd6e7319c3c963649b30a95b9fb36ec158055f563439e8edcd1236ef1f54dd63ce3a6ddd05686c4573b207e77733cac1fac973d23b123740167c0839ba597e2418243295e497825ae53e1230ce7e7536dc6ff671b726ea6e9884bf18290e263b67f635209547ce86b7cbc87a9260c1b3e633847867dda6f8f393dcc99720e4b41823d2bc9ec46b00d729bdea38670b44db09924c4fccf649e3af929ee3451ac1b78aa7a9a4adc8c6438c90124f8615b50f768309509d76249709457ae3f4fbf2383b9e34221d737191462040a8f68e17417e06e2b500878628f78d19df68790cd715a076b41bc815f1b3b34255d53b2fc760716779f9281e8769044e8b61946bbd43aaa539cc686922bd60d158a1b1463fd1224d2d2f205576d13fd6bd02f4f593abc5602dae12013a612d739886deb96c2c16267874092cd42d65f15be1ef396dc16b5031800dc7a036e4db2e7dfeb1a6d340c8e3bf7a9ffdc710b6c2402820eb055d737b9fa6b05f8ca80e40b59e29c265d84b2dd7d265af8979bf62a522f7fc46ad243759adfd282ab77f9052f4de94b78a411d397c5d8cfa720ea3d958b09b7d1d79e06ef72260d87541292fc4d80a6edd4ab217ecfc67296726f3ec37f0363c1b40d11b39217a505c00d7ed5de592371228a18be1af1a5964b4b3060ca237e921435c649648e91f975b4486dfdc9834e6ad39caa4d9260f8b06903427b8ba262f5a482cde1eb43131a6787332047168a0634646a0b5367cddbbb87a6f66f4b83672e6386dafc668ed39876046ffe7af3faf0464c0e9a647b7b8cf349c458a18fcfffe5994c654ea90e5d5ba7cbb023d00127a861fe8f8bda9e4c2760e8b6537430a108f4e0c1e34ee129a5805d6fa20950e3346a4ab276ee259d3d7c08684b4ad0d82451d094590556695a38b154b7d2e3bbc3841dafc4edd05bb8c7807ede30ca5d9435ff99dba567fe03f31a1b25eb1ccb0bef278afc67b49c0c0e4afd04803ffea05dd528d076822f06e9622065fbd87768412666d9a54a92dfc03f990094f816cf64caa4469bfec1f35f7716389258b519cd8fe503a55772cfa119ae6cff45b06a08a14e18625ad27a7756495361435caf0c6d604012c85a9212004ff9a1747961558ea6681fe8ce19f14cfa45d6e76ec01798ed692ad37547a183be49615c7c8fd43e677c5f73639c5496fd67e00d58b26746f65f1d6caa5be17bdeab8ef65a7338c41892252eceef0237ea0e374c95fbf4410ea9be57d5a1ba89766101b25dc4e80111f8c10d98ae9b90cf339909467981250051cc3e4fa3b4f11775b080d81372c08b8fb45bd9c6689768a0c942b221b492e4623391dd9d27b06f2469f989ce2c1ebcd6d4afc289ff10ab4033012a909fd5fc4c3924f98531f9640efa1f364354009bc6a468f6ecd84cfd1f08b61667fc1c68277494226e1bd9e000999224a502f0d6ab7a8e0d722fda2f98e70571505389bc0ff59406c8815afa38bec3cafbfe69f546ef1092e414a38390176e42fb9db99ac7e3b876bf80cba98fca1635575a61cea323d2ece409d66463f44c6a76734e24de84788860ad17b695bfd28d83fd5e15b2c7c11d7a84b8da2fc65f19a2ecd30f51394baa6908f9cff9b5e3645e0bec525cb2227e1a40e985c57ec2e2fb1338fcb595146956d27ed06201c659e66a5197579f94123f75a468b805d436deb3acd2393c3cc1232f6fb6050cfa3ea3ed886e4cb86844ccb301c517e20fe7a033e4f7a36f6116d37419a396f352819bf4377aea82062b4b3ee8bfd9a4e8bc2d054e579ec9c2bfe43179ad1f359f1effed79dbf0a0390c0a7f9061730f073b574684ac042b3091a4fbb0061a713d107c1c6577ad5226b7fbb26eb621b19cb14d1ea64decbe9622b801c9dbff863e59ae4b5904ba2a95a05a494ad12fda89b922d66222d532cc619368be598323650506d578fee882272bba0c28e5edde348bb1c621f83658c7725b5e7deaa1fa0a1e6e4b5fc87a2af2572b5857de668525a63bd15d038bf8be8ab03e5b72ba1e138d493d32e011fe99e37ae17fcc355e1c160de2422b8e7eee845630a885f1c20ebed438d08d62e3222f8025e30ec9d48b3eadb50e08040fcc11b03bc5a717005704a880be5b7ea4e70d36803db2cf1a4c0488826501bd5859b1bda42be51c9ed897386ed1835cc4dd744b43e4353d5d1c2e36ac7533cab93a3f3e34f61fd0af60890f2bdf219138cf51a803ccc85a6b62b1cddc6638c093ecb29404f672fc89a072c533294e7b19a17a5580a6b0d43103db96e1b81dd54861fb150df27c2bf433f82beeee479b5aa2da0ea904a6cc634cdde59f10f9959f1237e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hc6ae87c691f3fab3c881630bc9aae9bdef208b10e57ea1a7c26981cc702320e91b6dae3ff93096acc3b6468504e6bf9c73b34f67a831c0943d694bcc23d840779441ad2778a31a7764b76dd91a4326220c68c46fbec37949086307ca24c12b70325da96001ecc84f988acb0cca6406f3f8990f4f25a448d80e4dae6bc46a8820cc90cca4fd4fa5a3fc1df70f75e3ad2f12c711ad6f617e2488d9c81e8047e50972b0faf44e91998c4d92341e1f6b92e4773fd71a1775507665d8fde988ad034eb7c149ccafc63ea613d4b41d8fdb2084faabfdfeaa270e6747ffab3a7e5f06b381085c3b9732c88d2f2aa56d4dd7a6a6d52a87bdbfbcf5a25a20333b5530ee6a7726ca81bbcf9a646a760ecc824ceb9e32dad726afcc98c08e6bb9558b31137dc7258c8de0e1e20b2912eca018f6106ad3472705b42356641c326a0fd4990bf1c0c4e67b041f4689083da8649b970118cc768c710d07cc27ea88dab2cd3b401f72fa2ad1797e2eafe6280e1877d02555c5ad52709202262fcd3cfd244ae23b891ac798e5c45cc5cafeb3b096ef38d0a1e0851a2abaa086a29b824c310c5c2914b024b5d711b1e576fc2253c967c1656e0218bc8383dfe7626bd2af8d2f6f0183d265ddf10db25753f3046316cf2fb2c264b9d7375ec8b70d637b94c64266a03efc3516f0b0cc7a4fe5a7cc090dcc248aff952d588e8c30106016f825e456d7f859fec1392848c0ba5d8c2b9703dcbe6a002934e320c6f779a4ddc4c00cc6ec63fa5dc6317c693e6113381d5f5c1246bcc44046cf2bb35c0221e42485b8665ec20fdda7c6993785da1f760d82e4b95c9858288a810922148425546df912e2290e50c695fa0b9b5bf685b4a20631ab00e98fa17313392d63b1eb62ff84545a409bbbb3d9bb39f8f83e30a3058e58df9c910fbd7dbf60577ceb0b27e97203c6f70f4226745d4f97b8cd304f0e15187eee1ab6beac4389ecd79e7fda194562c266830c0d5532f9d732606bcf05fc3317ec7e40db0aca71af24caf0ea70ebc21c7cbc9f804ffb2ab83a045575a7f1737ea8f8b5985f027bfca500ed6935c4b41f565a830ec4d4b9b9cbe0b7d688a29ed9b89b44ad7b51dc8a87ef4a52369223b097e8f26550d7e29471e3377c64e23b2cf2e72058069c1b573d738aa1618e7f8421ff0d26a054e64566caabf0d93868141d855da1ca50fd861e6d19cebb3f2ff1bfdda3de60bbb8dba2228e7a852084b59a4ba7d5c30b3fe22c10a161c167e27e7add769616c00871787ce8a38b96a7b907494170918f8eba2bab5219bf4a3970b87a27ec1c54018134e674e277bcb46ae02d8923a87ab77ccd0f67e2ca17baa01805c41602d63183ca0fb90a5ec6ba66644454a391afc7d16f304179ecf1d9345a53d1008e1f5347a2023557dd8fa05b0d90105a547dba5e12aa54a0a0fa2741b9c41dd72fb9da0f57a709e86308e1fcac1ad60e1dd0e8b952affbdb084b12ed28bff0ee736807f2604a3a5ddc7be2d6c45f775c053c13f6d8f79b87b79af6559177383dc881ed1b036353db4dae28c4893b0805852304c14bb916bba6ff4199b1239ad28ad1c9d7f59058b64664980dc6a6ec778dd618552a1d4a8f9b91d97c82aec8d8e3f39351d8ac974f455724fc01f305b018760c02298fdf1536908a59b455a6dbbcf6334663a2bb6e79d97dca9d05b7c6368c2dbd5691d7ca8b6b16623945c651fa06ac88637fb856c7a2b5fddf7a8468ec448547cd274ce79d156b9cfc0d0b845163d91c41b030863063505763c26968215c382b201d3ce397c79afc246a87e73ecb91cf81e16376076c7d60014807baf736615f5e636232856fc8b6d921797c00b12e11c575bf7a7d23b0de5567ad0fd9dd0be0be20370410665a71bcd5f3116d3f22387f3d7b07cec874ccb9a6b3c4927679708fda34d331676c06d60b07c613f14f36d44d3d0030b91db93b565c27400c94b73b960552033e55b0c316da0d6f002a0eadea9130605d58a7ad3827e5d0f5e39cf2f08520b0b60dab7ce1fabe3d7099f30def12e336a30ce24dcbfc927eb2fe557ab6728ba3008db28dd2c08cf09e3e2a75cb7b5755ed3649948fda3548f3db47ac0a33205c2ffaf58c024eae4a146360cea4beab1a340ba80201f3f3d35bd32de2a6d3074b569b5de9f2a881aaed42db602266b475729033341a90b23536a20fef80a8d3c48a6530538bd38997cf88a12a0618136b1a83896ac59ad5f45778fdccc1bfbeff205411a7dbdc9cbe338754031901fb30834d2c13ba435337729e67d9ca68e532eab14bfe7437bdbc9615cb0a8db92452a2ac1eb19b6e3e66ecb2ba9d5d4e148e04eec99143a323f1b4e6ec108696bc9322e4e5822fa08a9a68a80325b7995d5c2c328f0fc12c00626c3f35cf72bb7e2a68197ea3812273a8e634e8cfc58cef3d3b329de544d62095efb9b1ac584b5b1168f33df513cf26bf970e5bee38e09a0b34e0ef59a057ac43c44d319f11f728a5701bf36cab4557ea5d93a8b5c0dd3db9e9869c2197371ebe245e2e700af2aeaeab2205fd72348b074e6c61c8af0c216f62a201fac559c4e6e67ba209ae5fe1963e0880618a4b5efb32a52ffd579c028190060a371bfa63545eaf934b1f26b8bb8d608d5dd5dc18363b7f06a1ad963b98e7d7a09c2906a785d055fa0d38c0e1d7ce223a794a1213274fe47ab3a9cd9864ba26d29294a17b334d1c7131a5f2d00f7bc5e6389c7cbd7a22909185ea2051144916e0e27993b3d1da9081479085b519ab0b24fe1b6256bba4c25c8c32f200e090cd0ebfb2d452a7f3d21cf8b782fa2e096993ff3818d2953c83a2d5e351d09bb6b90f31ab73b7cdaebb0e4df06fe9ae095e753ea532c05b0b7a7013bdd44ceb1876eda64253314fa229604411ec59f87497adbcffb83a085e6845a42da62122e635e5c2bfdaba9e37228b60e4a27348bf1f5c8441b71ed4046cf1184858b1de1fd3e5ce23eaf734d49b5d7c8044d9c2c6e41c6ff7df049424a62ff9522715bc47eb791da8d276aa992d3da7be39b68a9787ac9ef543dcc2a0d9616db1764ef66f16ed523c822a46b6200338a76d00c69af4107de08e668723e819a5162e9676e27aaa72827064aa1bbbd1becd7ac2bbf390cccafecb1264742c1ba17314a03f1095d53e95cf87db080f6368e5705032e87f0be201df2967c0ab395c581851c678d2e32b453f8013fba028a62f80b318a51d2225c7d1bea50a67d5f509000eebc67abab379965551c40f615e466df5d05b5d60bdf52ce7fa0150362d85f53a03495af8b537e6c9d2a8eaed8648821615b9aa80459e3d56c4079974fc93527ef96be6d1d23735589a4d6727a5227944f5774c8af9243a1649f5a40b219316f0640f66c577a310759862294f14f69e50d1c637cedecef7e37dc159f28980f91347f8c8d22165063d2837f06b1a12812542f5af5fa5bdc21d6ee1193c53988465cb6cbedc495a82a8e53213d409155d62b368c5e64dfac69ccb63c6f386455e8261491a869e269eb9e20492cfdf7d65c86244e55dad39ca04983cef95e0c470b13274f0a8a48c88e3d60e9b8db31265c5ea7798e7ad66828159361b197a34e3b3aa7418b60aea100dddb3c4ac55ca401a52aec1b0eea93bf1753142b9f7acdef42b1b6addebd450049c2d183b3728db62eebbf78aa50b17ad4d024e7a313587aeba6852dfc16e64863c74ade5636b7d6bf88e9ccf2e109fe059275a499b2f2420d6e0f139d839c5ee34ee264eec60ef1cf2ccc1d52c08aeb6cf75453a7129ee4072ea3aca91cd9647f0faf57c4b8e5333f78ab4947886c3c249f5aad393660a0e79596bf498d7ac63759ec0d67d7818b37d7c975d4849a6d4b624249a922256bd80ebf3e1037175074fda97d28248b51882e595370f797c98a0c02d2358b16cef864e0f78ce390a01ca9d11c60b56dfb0cfe2e3b2effe359b961bc2e94394442cbcd8aa7fca126befdf5b709b6a8e024102b33a863f2cdaa48c72da1819da93fc29d92ae152db63c99e8ca1861a6b3619173a7e2b758412b54505b4bde04f0f4ceed34a4f529a41abf673b660d616688b1c29b6025f1cf98db3ab404378d197322e3048cb592ea53c8e47bfee755bced12b54297d0d5556703053da2c1a0c7ef6198de87dbbf63476037e5c2d5aa946d33181d50bc3778ff37d0391d62bc477c759ccf72b34d238bd964fc79fbd51b46d16af702ab5160412a5e5fe4f1b122aa1a7d1c6a35994481a954ec597bfa3c41e8c4096e1b2ee8b47c87ed619d9cf676409d9322cd2b3800a8859a07b4069d119f2f34d75401e221e94b38314b43ebad03af3c910601c10cdd6605184d67ad421edb966de755e6e9e76c0d2fee20c4dde0ba6108d26e261c0250d1774add1719f895c52e3f104e25832eb88fce2bc5c4954249fb528eef9ffaa4a2d7ad4866687aa036bec6054683bc6a8811a95fe6c5cad45a31f6532f70d67c5498e2880babe953b33acd98d3cb3e45c9651f5f88078770359a118fbd4aa514c6b8ae3c811b9fc3f0e2f48bec89e9a844afbdd7024f7db8ef28fda2c0173b15c8310fd7a9d01b51f0384c359bf0ce944315b038282136b24b8421112e19534fedc7ce14d202f90a7c8df9b955f8585224f80808128b86d5b91272769a8f3c0c5ee5bae93eefbd7e660733fce0bd817e6cd84c0d7b2caf7f253c680f229a04ef0dffb02b8ce6ac8be4bdc2b2385550f005e1ee4a51d1845701e53bb306d30edf5ebc0c5d8c183f8f304bd1e32c4679a8e1e95a05838e3ec3ddd4158fdc9c8daeb61df36f7d5bcf9f53e17593bf7283d7ca7aab9edbc06a0c10acb0cabe73960897aa3fb19f722c986081e33c3909a41190b93744dd32bb757ba7500455b86a956ec414ec0a57815a480875b3f10d6ebdd02efa0e8f800a2c3e1ebb4cd94067422f331020561b8a6da82281e8e38206ad5d13dd99983ad7cdcd9cedda007aca0b9d1ff0d0728e0415b606c762ce16453a5048b412bf7b6d669c525574bc63cd492b74d5b52cc35ebeae7af0bdf2dd0ffae6f5b0953acefbe91eed9cd01aec8b7fbec15b022b0c79e33bfbcb7681f1499c3fddebea00541f9aee4c7ea8b4086090fdd73861ecc0f87cdb27204790309ef9c015575225c4b88a61f7ac77c41db8ca7280d0f73eb1ffc111d5411fe0494749b923906bb2231054c2708f66ef8e5a359b98f979c6d51accfe202bbdd35a1dad45fe27777e08f4ff8f63a06d807756e2c8a9c3a7bace1c4a451e88b39b4e7d8ce4b180efd8e34f7ad56395437ff42b7837f8398a5b20edc477eeec7b9b8cc15e41dbd0fdf14333093bd1f21f8965e0fc7b91f0e84ca4e27bc2e71cefd9205f6edddccf6c725c53d7d028343679dd7d67671580655ec07b643d49b9dda7dfd650e2c131fa2f7c7059b360d6df3539a629425875fde7665cef96e964042299e6bcf937251a265cdf1f428c1033d2523a691688c5e3a0440b4f9954902f6;
        #1
        $finish();
    end
endmodule
